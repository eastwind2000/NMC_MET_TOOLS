netcdf gfs_r24_2018062500_f096 {
dimensions: 
 lat = 601; 
 lon = 701; 
variables:  
float lat(lat) ; 
   lat:long_name = "latitude" ;
   lat:units = "degrees_north" ;
   lat:standard_name = "latitude" ;
float lon(lon) ;
   lon:long_name = "longitude" ;
   lon:units = "degrees_east" ;
   lon:standard_name = "longitude" ;
float APCP_24(lat, lon) ;
   APCP_24:name = "APCP_24" ;
   APCP_24:long_name = "Total Precipitation" ;
   APCP_24:level = "A24" ;
   APCP_24:units = "kg/m^2" ;
   APCP_24:_FillValue = -9999.f ;
   APCP_24:init_time = "20180625_000000" ;
   APCP_24:init_time_ut = "1529884800.0" ;
   APCP_24:valid_time = "20180629_000000" ;
   APCP_24:valid_time_ut = "1530230400.0" ;
   APCP_24:accum_time = "240000" ;
   APCP_24:_FillValue = 65535 ;
   APCP_24:accum_time_sec = 86400 ;
 // global attributes: 
 :_NCProperties = "version=1|netcdflibversion=4.4.1.1" ;
	:FileOrigins = "GFS_HR_APCP24" ; 
	:MET_version = "V7.0" ;
	:Projection = "LatLon" ;
	:lat_ll = "0.0 degrees_north" ; 
	:lon_ll = "70.0 degrees_east" ; 
	:delta_lat = "0.10 degrees" ;
	:delta_lon = "0.10 degrees" ;
	:Nlat = "601 grid_points" ; 
	:Nlon = "701 grid_points" ; 
data:
lat = 0.0,0.1,0.2,0.3,0.4,0.5,0.6,0.7,0.8,0.90000004,1.0,1.1,1.2,1.3000001,1.4,1.5,1.6,1.7,1.8000001,1.9,2.0,2.1000001,2.2,2.3,2.4,2.5,2.6000001,2.7,2.8,2.9,3.0,3.1000001,3.2,3.3,3.4,3.5,3.6000001,3.7,3.8,3.9,4.0,4.1,4.2000003,4.3,4.4,4.5,4.6,4.7000003,4.8,4.9,5.0,5.1,5.2000003,5.3,5.4,5.5,5.6,5.7000003,5.8,5.9,6.0,6.1,6.2000003,6.3,6.4,6.5,6.6,6.7000003,6.8,6.9,7.0,7.1,7.2000003,7.3,7.4,7.5,7.6,7.7000003,7.8,7.9,8.0,8.1,8.2,8.3,8.400001,8.5,8.6,8.7,8.8,8.900001,9.0,9.1,9.2,9.3,9.400001,9.5,9.6,9.7,9.8,9.900001,10.0,10.1,10.2,10.3,10.400001,10.5,10.6,10.7,10.8,10.900001,11.0,11.1,11.2,11.3,11.400001,11.5,11.6,11.7,11.8,11.900001,12.0,12.1,12.2,12.3,12.400001,12.5,12.6,12.7,12.8,12.900001,13.0,13.1,13.2,13.3,13.400001,13.5,13.6,13.7,13.8,13.900001,14.0,14.1,14.2,14.3,14.400001,14.5,14.6,14.7,14.8,14.900001,15.0,15.1,15.2,15.3,15.400001,15.5,15.6,15.7,15.8,15.900001,16.0,16.1,16.2,16.300001,16.4,16.5,16.6,16.7,16.800001,16.9,17.0,17.1,17.2,17.300001,17.4,17.5,17.6,17.7,17.800001,17.9,18.0,18.1,18.2,18.300001,18.4,18.5,18.6,18.7,18.800001,18.9,19.0,19.1,19.2,19.300001,19.4,19.5,19.6,19.7,19.800001,19.9,20.0,20.1,20.2,20.300001,20.4,20.5,20.6,20.7,20.800001,20.9,21.0,21.1,21.2,21.300001,21.4,21.5,21.6,21.7,21.800001,21.9,22.0,22.1,22.2,22.300001,22.4,22.5,22.6,22.7,22.800001,22.9,23.0,23.1,23.2,23.300001,23.4,23.5,23.6,23.7,23.800001,23.9,24.0,24.1,24.2,24.300001,24.4,24.5,24.6,24.7,24.800001,24.9,25.0,25.1,25.2,25.300001,25.4,25.5,25.6,25.7,25.800001,25.9,26.0,26.1,26.2,26.300001,26.4,26.5,26.6,26.7,26.800001,26.9,27.0,27.1,27.2,27.300001,27.4,27.5,27.6,27.7,27.800001,27.9,28.0,28.1,28.2,28.300001,28.4,28.5,28.6,28.7,28.800001,28.9,29.0,29.1,29.2,29.300001,29.4,29.5,29.6,29.7,29.800001,29.9,30.0,30.1,30.2,30.300001,30.4,30.5,30.6,30.7,30.800001,30.9,31.0,31.1,31.2,31.300001,31.4,31.5,31.6,31.7,31.800001,31.9,32.0,32.100002,32.2,32.3,32.4,32.5,32.600002,32.7,32.8,32.9,33.0,33.100002,33.2,33.3,33.4,33.5,33.600002,33.7,33.8,33.9,34.0,34.100002,34.2,34.3,34.4,34.5,34.600002,34.7,34.8,34.9,35.0,35.100002,35.2,35.3,35.4,35.5,35.600002,35.7,35.8,35.9,36.0,36.100002,36.2,36.3,36.4,36.5,36.600002,36.7,36.8,36.9,37.0,37.100002,37.2,37.3,37.4,37.5,37.600002,37.7,37.8,37.9,38.0,38.100002,38.2,38.3,38.4,38.5,38.600002,38.7,38.8,38.9,39.0,39.100002,39.2,39.3,39.4,39.5,39.600002,39.7,39.8,39.9,40.0,40.100002,40.2,40.3,40.4,40.5,40.600002,40.7,40.8,40.9,41.0,41.100002,41.2,41.3,41.4,41.5,41.600002,41.7,41.8,41.9,42.0,42.100002,42.2,42.3,42.4,42.5,42.600002,42.7,42.8,42.9,43.0,43.100002,43.2,43.3,43.4,43.5,43.600002,43.7,43.8,43.9,44.0,44.100002,44.2,44.3,44.4,44.5,44.600002,44.7,44.8,44.9,45.0,45.100002,45.2,45.3,45.4,45.5,45.600002,45.7,45.8,45.9,46.0,46.100002,46.2,46.3,46.4,46.5,46.600002,46.7,46.8,46.9,47.0,47.100002,47.2,47.3,47.4,47.5,47.600002,47.7,47.8,47.9,48.0,48.100002,48.2,48.3,48.4,48.5,48.600002,48.7,48.8,48.9,49.0,49.100002,49.2,49.3,49.4,49.5,49.600002,49.7,49.8,49.9,50.0,50.100002,50.2,50.3,50.4,50.5,50.600002,50.7,50.8,50.9,51.0,51.100002,51.2,51.3,51.4,51.5,51.600002,51.7,51.8,51.9,52.0,52.100002,52.2,52.3,52.4,52.5,52.600002,52.7,52.8,52.9,53.0,53.100002,53.2,53.3,53.4,53.5,53.600002,53.7,53.8,53.9,54.0,54.100002,54.2,54.3,54.4,54.5,54.600002,54.7,54.8,54.9,55.0,55.100002,55.2,55.3,55.4,55.5,55.600002,55.7,55.8,55.9,56.0,56.100002,56.2,56.3,56.4,56.5,56.600002,56.7,56.8,56.9,57.0,57.100002,57.2,57.3,57.4,57.5,57.600002,57.7,57.8,57.9,58.0,58.100002,58.2,58.3,58.4,58.5,58.600002,58.7,58.8,58.9,59.0,59.100002,59.2,59.3,59.4,59.5,59.600002,59.7,59.8,59.9,60.0;
lon = 70.0,70.1,70.2,70.3,70.4,70.5,70.6,70.7,70.8,70.9,71.0,71.1,71.2,71.3,71.4,71.5,71.6,71.7,71.8,71.9,72.0,72.1,72.2,72.3,72.4,72.5,72.6,72.7,72.8,72.9,73.0,73.1,73.2,73.3,73.4,73.5,73.6,73.7,73.8,73.9,74.0,74.1,74.2,74.3,74.4,74.5,74.6,74.7,74.8,74.9,75.0,75.1,75.2,75.3,75.4,75.5,75.6,75.7,75.8,75.9,76.0,76.1,76.2,76.3,76.4,76.5,76.6,76.7,76.8,76.9,77.0,77.1,77.2,77.3,77.4,77.5,77.6,77.7,77.8,77.9,78.0,78.1,78.2,78.3,78.4,78.5,78.6,78.7,78.8,78.9,79.0,79.1,79.2,79.3,79.4,79.5,79.6,79.7,79.8,79.9,80.0,80.1,80.2,80.3,80.4,80.5,80.6,80.7,80.8,80.9,81.0,81.1,81.2,81.3,81.4,81.5,81.6,81.7,81.8,81.9,82.0,82.1,82.2,82.3,82.4,82.5,82.6,82.7,82.8,82.9,83.0,83.1,83.2,83.3,83.4,83.5,83.6,83.7,83.8,83.9,84.0,84.1,84.2,84.3,84.4,84.5,84.6,84.7,84.8,84.9,85.0,85.1,85.2,85.3,85.4,85.5,85.6,85.7,85.8,85.9,86.0,86.1,86.2,86.3,86.4,86.5,86.6,86.7,86.8,86.9,87.0,87.1,87.2,87.3,87.4,87.5,87.6,87.7,87.8,87.9,88.0,88.1,88.2,88.3,88.4,88.5,88.6,88.7,88.8,88.9,89.0,89.1,89.2,89.3,89.4,89.5,89.6,89.7,89.8,89.9,90.0,90.1,90.2,90.3,90.4,90.5,90.6,90.7,90.8,90.9,91.0,91.1,91.2,91.3,91.4,91.5,91.6,91.7,91.8,91.9,92.0,92.1,92.2,92.3,92.4,92.5,92.6,92.7,92.8,92.9,93.0,93.1,93.2,93.3,93.4,93.5,93.6,93.7,93.8,93.9,94.0,94.1,94.2,94.3,94.4,94.5,94.6,94.7,94.8,94.9,95.0,95.1,95.2,95.3,95.4,95.5,95.6,95.7,95.8,95.9,96.0,96.1,96.2,96.3,96.4,96.5,96.6,96.7,96.8,96.9,97.0,97.1,97.2,97.3,97.4,97.5,97.6,97.7,97.8,97.9,98.0,98.1,98.2,98.3,98.4,98.5,98.6,98.7,98.8,98.9,99.0,99.1,99.2,99.3,99.4,99.5,99.6,99.7,99.8,99.9,100.0,100.1,100.2,100.3,100.4,100.5,100.6,100.7,100.8,100.9,101.0,101.1,101.2,101.3,101.4,101.5,101.6,101.7,101.8,101.9,102.0,102.100006,102.2,102.3,102.4,102.5,102.600006,102.7,102.8,102.9,103.0,103.100006,103.2,103.3,103.4,103.5,103.600006,103.7,103.8,103.9,104.0,104.100006,104.2,104.3,104.4,104.5,104.600006,104.7,104.8,104.9,105.0,105.100006,105.2,105.3,105.4,105.5,105.600006,105.7,105.8,105.9,106.0,106.100006,106.2,106.3,106.4,106.5,106.600006,106.7,106.8,106.9,107.0,107.100006,107.2,107.3,107.4,107.5,107.600006,107.7,107.8,107.9,108.0,108.100006,108.2,108.3,108.4,108.5,108.600006,108.7,108.8,108.9,109.0,109.100006,109.2,109.3,109.4,109.5,109.600006,109.7,109.8,109.9,110.0,110.100006,110.2,110.3,110.4,110.5,110.600006,110.7,110.8,110.9,111.0,111.100006,111.2,111.3,111.4,111.5,111.600006,111.7,111.8,111.9,112.0,112.100006,112.2,112.3,112.4,112.5,112.600006,112.7,112.8,112.9,113.0,113.100006,113.2,113.3,113.4,113.5,113.600006,113.7,113.8,113.9,114.0,114.100006,114.2,114.3,114.4,114.5,114.600006,114.7,114.8,114.9,115.0,115.100006,115.2,115.3,115.4,115.5,115.600006,115.7,115.8,115.9,116.0,116.100006,116.2,116.3,116.4,116.5,116.600006,116.7,116.8,116.9,117.0,117.100006,117.2,117.3,117.4,117.5,117.600006,117.7,117.8,117.9,118.0,118.100006,118.2,118.3,118.4,118.5,118.600006,118.7,118.8,118.9,119.0,119.100006,119.2,119.3,119.4,119.5,119.600006,119.7,119.8,119.9,120.0,120.100006,120.2,120.3,120.4,120.5,120.600006,120.7,120.8,120.9,121.0,121.100006,121.2,121.3,121.4,121.5,121.600006,121.7,121.8,121.9,122.0,122.100006,122.2,122.3,122.4,122.5,122.600006,122.7,122.8,122.9,123.0,123.100006,123.2,123.3,123.4,123.5,123.600006,123.7,123.8,123.9,124.0,124.100006,124.2,124.3,124.4,124.5,124.600006,124.7,124.8,124.9,125.0,125.100006,125.2,125.3,125.4,125.5,125.600006,125.7,125.8,125.9,126.0,126.100006,126.2,126.3,126.4,126.5,126.600006,126.7,126.8,126.9,127.0,127.100006,127.2,127.3,127.4,127.5,127.600006,127.7,127.8,127.9,128.0,128.1,128.2,128.3,128.4,128.5,128.6,128.7,128.8,128.9,129.0,129.1,129.2,129.3,129.4,129.5,129.6,129.7,129.8,129.9,130.0,130.1,130.2,130.3,130.4,130.5,130.6,130.7,130.8,130.9,131.0,131.1,131.2,131.3,131.4,131.5,131.6,131.7,131.8,131.9,132.0,132.1,132.2,132.3,132.4,132.5,132.6,132.7,132.8,132.9,133.0,133.1,133.2,133.3,133.4,133.5,133.6,133.7,133.8,133.9,134.0,134.1,134.20001,134.3,134.4,134.5,134.6,134.70001,134.8,134.9,135.0,135.1,135.20001,135.3,135.4,135.5,135.6,135.70001,135.8,135.9,136.0,136.1,136.20001,136.3,136.4,136.5,136.6,136.70001,136.8,136.9,137.0,137.1,137.20001,137.3,137.4,137.5,137.6,137.70001,137.8,137.9,138.0,138.1,138.20001,138.3,138.4,138.5,138.6,138.70001,138.8,138.9,139.0,139.1,139.20001,139.3,139.4,139.5,139.6,139.70001,139.8,139.9,140.0;
APCP_24 = 0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.13778515,0.15047589,0.16316663,0.17585737,0.18673515,0.18673515,0.18673515,0.18673515,0.18673515,0.18673515,0.17585737,0.16316663,0.15047589,0.13778515,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.15047589,0.17585737,0.19942589,0.22480737,0.25018883,0.4749962,0.69980353,0.9246109,1.1494182,1.3742256,1.9996977,2.6251698,3.2506418,3.874301,4.499773,4.249584,3.9993954,3.7492065,3.5008307,3.2506418,4.361988,5.475147,6.588306,7.699652,8.812811,9.461852,10.112705,10.761745,11.4126,12.06164,12.137785,12.212116,12.28826,12.362592,12.436923,11.650098,10.863272,10.074633,9.287807,8.499168,8.399456,8.299743,8.200029,8.100317,8.000604,8.613385,9.224354,9.837135,10.449916,11.062697,11.075388,11.088079,11.10077,11.111648,11.124338,10.51337,9.900589,9.287807,8.675026,8.062244,6.9128265,5.763408,4.612177,3.4627585,2.3133402,1.8619126,1.4122978,0.96268314,0.51306844,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,1.2872034,2.4493124,3.6132345,4.7753434,5.9374523,4.749962,3.5624714,2.374981,1.1874905,0.0,1.2872034,2.5744069,3.8634233,5.1506267,6.43783,6.4994707,6.5629244,6.624565,6.688019,6.7496595,6.43783,6.1241875,5.812358,5.5005283,5.186886,4.8750563,4.5632267,4.249584,3.9377546,3.6241121,2.9369993,2.2498865,1.5627737,0.87566096,0.18673515,0.16316663,0.13778515,0.11240368,0.0870222,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,0.25018883,0.25018883,0.25018883,0.25018883,0.25018883,0.21211663,0.17585737,0.13778515,0.099712946,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.21211663,0.2374981,0.26287958,0.28826106,0.31182957,0.7124943,1.1131591,1.5120108,1.9126755,2.3133402,3.2633326,4.213325,5.163317,6.11331,7.063302,7.699652,8.337815,8.974165,9.612328,10.25049,9.686659,9.12464,8.562622,8.000604,7.4367723,7.9752226,8.511859,9.050309,9.5869465,10.125396,8.861761,7.5999393,6.338117,5.0744824,3.8126602,4.1117992,4.4127507,4.7118897,5.0128417,5.3119802,6.4759026,7.6380115,8.80012,9.96223,11.124338,12.137785,13.149418,14.162864,15.174497,16.187943,19.337059,22.487988,25.637104,28.788033,31.93715,28.586794,25.238253,21.887897,18.537542,15.187187,15.324973,15.462758,15.600543,15.738328,15.8743,15.337664,14.799213,14.262577,13.724127,13.1874895,11.961927,10.738177,9.512614,8.287052,7.063302,12.538449,18.011784,23.48693,28.962078,34.437225,31.525606,28.612175,25.700558,22.787127,19.87551,21.762802,23.650097,25.537392,27.424685,29.31198,26.300648,23.287504,20.27436,17.26303,14.249886,15.687565,17.125244,18.562923,20.000603,21.438282,18.049856,14.663241,11.274815,7.8882003,4.499773,4.8750563,5.2503395,5.6256227,6.000906,6.3743763,5.137936,3.8996825,2.663242,1.4249886,0.18673515,0.40066472,0.61278135,0.824898,1.0370146,1.2491312,2.8499773,4.4508233,6.049856,7.650702,9.249735,7.61263,5.975525,4.3366065,2.6995013,1.062396,3.8380418,6.6118746,9.38752,12.163166,14.936998,17.725336,20.511858,23.300196,26.08672,28.875055,29.86312,30.849371,31.837437,32.8255,33.811752,30.813112,27.812658,24.812206,21.811752,18.813112,21.762802,24.712494,27.662184,30.611874,33.563377,33.66309,33.762802,33.862514,33.962227,34.06194,32.374073,30.688017,29.000149,27.31228,25.624413,24.03807,22.449915,20.861761,19.275417,17.687263,17.087172,16.487082,15.8869915,15.2869005,14.68681,11.74981,8.812811,5.8758116,2.9369993,0.0,0.15047589,0.2991388,0.44961473,0.6000906,0.7505665,1.7748904,2.7992141,3.825351,4.8496747,5.8758116,6.16226,6.450521,6.736969,7.02523,7.311678,7.3370595,7.362441,7.3878226,7.413204,7.4367723,8.6877165,9.936848,11.187792,12.436923,13.687867,11.949236,10.212419,8.4756,6.736969,5.0001507,6.4632115,7.9244595,9.38752,10.850581,12.311829,10.912222,9.512614,8.113008,6.7134004,5.3119802,6.2384043,7.1630154,8.087626,9.012237,9.936848,11.537694,13.136727,14.737573,16.336605,17.937452,18.287354,18.637255,18.987158,19.337059,19.68696,17.33736,14.9877615,12.638163,10.28675,7.93715,8.113008,8.287052,8.46291,8.636953,8.812811,11.836833,14.862667,17.886688,20.912523,23.938358,20.399454,16.862366,13.325275,9.788185,6.249282,5.7869763,5.3246713,4.8623657,4.40006,3.9377546,7.9625316,11.9873085,16.012085,20.036863,24.06164,24.68711,25.312584,25.938055,26.561714,27.187187,25.637104,24.08702,22.536938,20.986855,19.436771,19.03792,18.637255,18.236591,17.837738,17.437075,17.06179,16.68832,16.313038,15.937754,15.56247,15.049402,14.538147,14.025079,13.512011,13.000754,13.125849,13.24913,13.374225,13.499319,13.6244135,13.325275,13.024323,12.725184,12.4242325,12.125093,12.763257,13.399607,14.037769,14.674119,15.312282,17.350052,19.387821,21.425592,23.461548,25.49932,22.01299,18.52485,15.036712,11.5503845,8.062244,9.461852,10.863272,12.262879,13.662486,15.062093,15.138238,15.212569,15.2869005,15.363045,15.437376,14.699501,13.961625,13.225562,12.487686,11.74981,0.05076295,0.059827764,0.07070554,0.07977036,0.09064813,0.099712946,0.11059072,0.11965553,0.13053331,0.13959812,0.15047589,0.15047589,0.15047589,0.15047589,0.15047589,0.15047589,0.13959812,0.13053331,0.11965553,0.11059072,0.099712946,0.09064813,0.07977036,0.07070554,0.059827764,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.038072214,0.06164073,0.0870222,0.11240368,0.13778515,0.21936847,0.30276474,0.38434806,0.46774435,0.5493277,0.46411842,0.38072214,0.2955129,0.21030366,0.12509441,0.15410182,0.18492219,0.21574254,0.24474995,0.2755703,0.6327239,0.9898776,1.3470312,1.7041848,2.0631514,2.7974012,3.531651,4.267714,5.0019636,5.7380266,5.8341136,5.9320135,6.0299134,6.1278133,6.2257137,6.970841,7.7141557,8.459284,9.2044115,9.949538,10.388275,10.825199,11.262123,11.700861,12.137785,12.085209,12.032633,11.980057,11.927481,11.874905,10.9774885,10.080072,9.182655,8.285239,7.3878226,7.380571,7.3733187,7.364254,7.3570023,7.3497505,7.915395,8.479226,9.04487,9.610515,10.174346,10.130835,10.085511,10.040187,9.994863,9.949538,9.47273,8.994107,8.517298,8.040489,7.5618668,6.644508,5.727149,4.8097897,3.8924308,2.9750717,2.4474995,1.9199274,1.3923552,0.86478317,0.33721104,0.27194437,0.20667773,0.14322405,0.07795739,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.07977036,0.14684997,0.21574254,0.28282216,0.34990177,0.42423326,0.50037766,0.5747091,0.6508536,0.72518504,0.6417888,0.56020546,0.47680917,0.39522585,0.31182957,0.2520018,0.19217403,0.13234627,0.072518505,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.34083697,0.67986095,1.020698,1.3597219,1.7005589,2.6233568,3.5443418,4.4671397,5.389938,6.3127356,5.4008155,4.4870825,3.5751622,2.663242,1.7495089,2.6868105,3.6241121,4.5632267,5.5005283,6.43783,6.450521,6.4632115,6.4759026,6.48678,6.4994707,6.14413,5.7906027,5.4352617,5.0799212,4.7245803,4.458075,4.1897564,3.923251,3.6549325,3.386614,2.7502642,2.1121013,1.4757515,0.8375887,0.19942589,0.17585737,0.15047589,0.12509441,0.099712946,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.014503701,0.018129626,0.01994259,0.02175555,0.025381476,0.032633327,0.03988518,0.047137026,0.054388877,0.06164073,0.09064813,0.11784257,0.14503701,0.17223145,0.19942589,0.19942589,0.19942589,0.19942589,0.19942589,0.19942589,0.17767033,0.15410182,0.13234627,0.11059072,0.0870222,0.07070554,0.052575916,0.034446288,0.018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.01994259,0.027194439,0.034446288,0.04169814,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.17223145,0.19579996,0.21755551,0.23931105,0.26287958,0.64722764,1.0333886,1.4177368,1.8020848,2.1882458,3.1944401,4.2024474,5.2104545,6.2166486,7.224656,7.855567,8.484665,9.115576,9.744674,10.375585,9.706602,9.039432,8.372261,7.705091,7.037921,7.46578,7.891826,8.319685,8.747544,9.175404,8.192778,7.210152,6.2275267,5.2449007,4.262275,4.7699046,5.277534,5.7851634,6.2927933,6.8004227,7.663393,8.52455,9.38752,10.25049,11.111648,11.671853,12.232059,12.792264,13.352469,13.912675,16.41819,18.92189,21.427404,23.932919,26.43662,24.422419,22.408218,20.392202,18.378002,16.361988,16.59586,16.827919,17.059978,17.292038,17.52591,16.537846,15.54978,14.561715,13.575464,12.5873995,13.488441,14.387671,15.2869005,16.187943,17.087172,19.819307,22.553255,25.285389,28.017523,30.749659,28.521528,26.29521,24.067078,21.84076,19.612629,20.713097,21.811752,22.912222,24.01269,25.113157,22.964798,20.818249,18.66989,16.52334,14.37498,15.787278,17.199575,18.611874,20.024172,21.438282,18.635443,15.8326025,13.029762,10.226922,7.4258947,8.033237,8.640579,9.247922,9.855265,10.462607,8.94697,7.4331465,5.91751,4.401873,2.8880494,2.7883365,2.6868105,2.5870976,2.4873846,2.3876717,3.972201,5.5567303,7.1430726,8.727602,10.312131,8.655084,6.9980354,5.3391747,3.682127,2.0250793,4.0157123,6.004532,7.995165,9.985798,11.974618,14.309713,16.64481,18.979906,21.315,23.650097,24.658104,25.664299,26.672306,27.680313,28.68832,26.396736,24.106964,21.817192,19.52742,17.237648,19.663393,22.087322,24.513067,26.936998,29.362741,29.772472,30.182201,30.59193,31.00166,31.413202,30.466837,29.522284,28.577728,27.633175,26.68681,24.371656,22.058315,19.743162,17.428009,15.112856,14.4420595,13.773077,13.102281,12.433297,11.762501,9.672155,7.5818095,5.4932766,3.4029307,1.3125849,1.1820517,1.0533313,0.922798,0.79226464,0.66173136,1.4830034,2.3024626,3.1219215,3.9431937,4.762653,5.032784,5.3029156,5.573047,5.8431783,6.11331,6.484967,6.8566246,7.230095,7.6017523,7.9752226,9.973107,11.969179,13.967064,15.964949,17.962833,15.91056,13.858286,11.804199,9.751925,7.699652,8.94697,10.194288,11.443419,12.690738,13.938056,12.857531,11.777005,10.698292,9.617766,8.537241,9.702975,10.866898,12.032633,13.196554,14.362289,15.504456,16.646622,17.790602,18.932768,20.074934,20.32331,20.569874,20.818249,21.064812,21.313189,19.070553,16.827919,14.585284,12.342649,10.100015,9.697536,9.295059,8.892582,8.490104,8.087626,11.557636,15.027647,18.497658,21.967669,25.437677,22.62396,19.812056,17.00015,14.188245,11.374527,10.667472,9.960417,9.253361,8.544493,7.837437,10.937603,14.037769,17.137936,20.238102,23.338266,23.849524,24.36259,24.87566,25.386915,25.899984,24.75419,23.610212,22.464418,21.32044,20.174648,19.415016,18.655384,17.895754,17.13431,16.374678,16.122677,15.870674,15.616859,15.364858,15.112856,14.8227825,14.532708,14.242634,13.95256,13.662486,13.492067,13.321649,13.153044,12.982625,12.812206,12.697989,12.581961,12.467744,12.351714,12.237497,12.786825,13.337966,13.887294,14.436621,14.9877615,16.905876,18.822178,20.740292,22.656593,24.574707,21.392958,18.209396,15.027647,11.845898,8.662335,10.384649,12.106964,13.829279,15.551593,17.27572,16.829731,16.385555,15.939567,15.495391,15.049402,14.235382,13.419549,12.605529,11.789696,10.975676,0.038072214,0.045324065,0.052575916,0.059827764,0.06707962,0.07433146,0.08339628,0.09064813,0.09789998,0.10515183,0.11240368,0.11240368,0.11240368,0.11240368,0.11240368,0.11240368,0.10515183,0.09789998,0.09064813,0.08339628,0.07433146,0.06707962,0.059827764,0.052575916,0.045324065,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.07433146,0.12509441,0.17585737,0.22480737,0.2755703,0.42785916,0.58014804,0.7324369,0.88472575,1.0370146,0.8557183,0.6726091,0.4894999,0.30820364,0.12509441,0.15954071,0.19579996,0.23024625,0.26469254,0.2991388,0.7904517,1.2799516,1.7694515,2.2607644,2.7502642,3.5951047,4.439945,5.2847857,6.1296263,6.9744673,7.420456,7.8646317,8.31062,8.754796,9.200785,9.577881,9.954978,10.332074,10.70917,11.088079,11.312886,11.537694,11.762501,11.9873085,12.212116,12.032633,11.853149,11.671853,11.49237,11.312886,10.304879,9.296872,8.290678,7.2826705,6.2746634,6.359873,6.445082,6.530291,6.6155005,6.70071,7.217404,7.7340984,8.252605,8.7693,9.287807,9.184468,9.082943,8.979604,8.8780775,8.774739,8.432089,8.089439,7.746789,7.404139,7.063302,6.378002,5.6927023,5.0074024,4.322103,3.636803,3.0330863,2.427557,1.8220274,1.2183108,0.61278135,0.4949388,0.3770962,0.25925365,0.14322405,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.15954071,0.2955129,0.42967212,0.5656443,0.69980353,0.85027945,1.0007553,1.1494182,1.2998942,1.4503701,1.2853905,1.1204109,0.9554313,0.7904517,0.62547207,0.5058166,0.38434806,0.26469254,0.14503701,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.6544795,1.310772,1.9652514,2.619731,3.2742105,3.9576974,4.6393714,5.3228583,6.004532,6.688019,6.049856,5.411693,4.7753434,4.137181,3.5008307,4.0882306,4.6756306,5.2630305,5.8504305,6.43783,6.399758,6.3616858,6.3254266,6.2873545,6.249282,5.8522434,5.4552045,5.0581656,4.6593137,4.262275,4.0392804,3.8180993,3.5951047,3.3721104,3.149116,2.561716,1.9743162,1.3869164,0.7995165,0.21211663,0.18673515,0.16316663,0.13778515,0.11240368,0.0870222,0.07070554,0.052575916,0.034446288,0.018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.030820364,0.034446288,0.03988518,0.045324065,0.05076295,0.065266654,0.07977036,0.09427405,0.11059072,0.12509441,0.13053331,0.13415924,0.13959812,0.14503701,0.15047589,0.15047589,0.15047589,0.15047589,0.15047589,0.15047589,0.14322405,0.13415924,0.12690738,0.11965553,0.11240368,0.09064813,0.06707962,0.045324065,0.02175555,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.018129626,0.034446288,0.052575916,0.07070554,0.0870222,0.07433146,0.06164073,0.05076295,0.038072214,0.025381476,0.03988518,0.054388877,0.07070554,0.08520924,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.13234627,0.15228885,0.17223145,0.19217403,0.21211663,0.581961,0.95180535,1.3216497,1.693307,2.0631514,3.1273603,4.1915693,5.2575917,6.3218007,7.3878226,8.009668,8.6333275,9.255174,9.87702,10.500679,9.728357,8.954222,8.1819,7.409578,6.637256,6.9545245,7.271793,7.590874,7.9081426,8.225411,7.5219817,6.8203654,6.1169357,5.4153194,4.7118897,5.42801,6.1423173,6.8566246,7.572745,8.287052,8.8508835,9.412902,9.97492,10.536939,11.10077,11.207735,11.314699,11.421664,11.530442,11.637406,13.497506,15.357606,17.217705,19.077805,20.937904,20.258043,19.578182,18.898321,18.216648,17.536787,17.864933,18.193079,18.519413,18.847559,19.175705,17.738026,16.300346,14.862667,13.424988,11.9873085,15.013144,18.037165,21.063,24.08702,27.112856,27.101978,27.092913,27.082035,27.07297,27.062092,25.51926,23.978243,22.435411,20.89258,19.34975,19.663393,19.975222,20.287052,20.600695,20.912523,19.630758,18.347181,17.065416,15.781839,14.500074,15.8869915,17.27572,18.662638,20.049553,21.438282,19.219215,17.001963,14.78471,12.567456,10.3502035,11.189605,12.03082,12.870221,13.709623,14.5508375,12.757817,10.964798,9.171778,7.380571,5.5875506,5.1741953,4.762653,4.349297,3.9377546,3.5243993,5.0944247,6.6644506,8.234476,9.804502,11.374527,9.697536,8.020547,6.341743,4.664753,2.9877625,4.1933823,5.3971896,6.60281,7.806617,9.012237,10.8959055,12.7777605,14.6596155,16.543283,18.425138,19.453089,20.479225,21.507175,22.535126,23.563074,21.982172,20.40308,18.822178,17.243088,15.662184,17.562168,19.462152,21.362139,23.262123,25.162107,25.881853,26.6016,27.323158,28.042906,28.762651,28.559599,28.35836,28.15531,27.952257,27.749205,24.707054,21.664904,18.622751,15.580601,12.536636,11.7969475,11.057259,10.31757,9.577881,8.838193,7.5945,6.352621,5.1107416,3.8670492,2.6251698,2.2154403,1.8057107,1.3941683,0.98443866,0.5747091,1.1893034,1.8057107,2.420305,3.0348995,3.6494937,3.9033084,4.15531,4.407312,4.6593137,4.9131284,5.632875,6.352621,7.072367,7.7921133,8.511859,11.258497,14.00151,16.748148,19.492973,22.237799,19.87007,17.50234,15.134612,12.766883,10.399154,11.432542,12.464118,13.497506,14.529082,15.56247,14.802839,14.043208,13.281764,12.522133,11.762501,13.167547,14.572594,15.977639,17.382685,18.787731,19.473032,20.15833,20.841818,21.527117,22.212418,22.357454,22.502491,22.647528,22.792566,22.937603,20.801933,18.668076,16.532406,14.396736,12.262879,11.282066,10.303066,9.322253,8.343254,7.362441,11.27844,15.192626,19.106813,23.022812,26.936998,24.850279,22.761745,20.675026,18.588305,16.499773,15.547967,14.594349,13.642544,12.690738,11.73712,13.912675,16.08823,18.261972,20.437527,22.613083,23.011934,23.4126,23.813263,24.212114,24.61278,23.87309,23.13159,22.391901,21.652212,20.912523,19.792112,18.671701,17.553104,16.432693,15.312282,15.181748,15.053028,14.922495,14.791962,14.663241,14.594349,14.527269,14.46019,14.39311,14.324218,13.860099,13.394168,12.930049,12.465931,11.999999,12.070704,12.139598,12.210303,12.279196,12.349901,12.812206,13.274512,13.736817,14.199123,14.663241,16.459887,18.258347,20.054993,21.851639,23.650097,20.772924,17.89394,15.016769,12.139598,9.262425,11.307447,13.352469,15.397491,17.442513,19.487535,18.523039,17.55673,16.592234,15.627737,14.663241,13.769451,12.877473,11.985496,11.091705,10.199727,0.025381476,0.030820364,0.034446288,0.03988518,0.045324065,0.05076295,0.054388877,0.059827764,0.065266654,0.07070554,0.07433146,0.07433146,0.07433146,0.07433146,0.07433146,0.07433146,0.07070554,0.065266654,0.059827764,0.054388877,0.05076295,0.045324065,0.03988518,0.034446288,0.030820364,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.11240368,0.18673515,0.26287958,0.33721104,0.41335547,0.6345369,0.8575313,1.0805258,1.3017071,1.5247015,1.2455053,0.9644961,0.6852999,0.40429065,0.12509441,0.16497959,0.20486477,0.24474995,0.28463513,0.3245203,0.9481794,1.5700256,2.1918716,2.8155308,3.437377,4.3928084,5.3482394,6.301858,7.2572894,8.212721,9.004985,9.79725,10.589515,11.381779,12.175857,12.184921,12.195799,12.2048645,12.215742,12.224807,12.237497,12.250188,12.262879,12.27557,12.28826,11.980057,11.671853,11.365462,11.057259,10.750868,9.63227,8.515485,7.3968873,6.2801023,5.163317,5.3391747,5.516845,5.6945157,5.8721857,6.049856,6.5194135,6.9907837,7.460341,7.9298983,8.399456,8.239915,8.080374,7.9208336,7.75948,7.5999393,7.3932614,7.1847706,6.978093,6.7696023,6.5629244,6.109684,5.658256,5.2050157,4.751775,4.3003473,3.6168604,2.9351864,2.2516994,1.5700256,0.8883517,0.7179332,0.5475147,0.3770962,0.20667773,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.23931105,0.44236287,0.64541465,0.8466535,1.0497054,1.2745126,1.49932,1.7241274,1.9507477,2.175555,1.9271792,1.6806163,1.4322405,1.1856775,0.93730164,0.75781834,0.57833505,0.39703882,0.21755551,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.969935,1.93987,2.909805,3.87974,4.8496747,5.292038,5.7344007,6.1767635,6.6191263,7.063302,6.70071,6.338117,5.975525,5.612932,5.2503395,5.487838,5.7253356,5.962834,6.200332,6.43783,6.350808,6.261973,6.1749506,6.0879283,6.000906,5.560356,5.1198063,4.6792564,4.2405195,3.7999697,3.6222992,3.444629,3.2669585,3.0892882,2.911618,2.374981,1.8383441,1.2998942,0.76325727,0.22480737,0.19942589,0.17585737,0.15047589,0.12509441,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.045324065,0.052575916,0.059827764,0.06707962,0.07433146,0.09789998,0.11965553,0.14322405,0.16497959,0.18673515,0.17041849,0.15228885,0.13415924,0.11784257,0.099712946,0.099712946,0.099712946,0.099712946,0.099712946,0.099712946,0.10696479,0.11421664,0.12328146,0.13053331,0.13778515,0.11059072,0.08339628,0.054388877,0.027194439,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.0870222,0.07433146,0.06164073,0.05076295,0.038072214,0.059827764,0.08339628,0.10515183,0.12690738,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.092461094,0.11059072,0.12690738,0.14503701,0.16316663,0.5166943,0.872035,1.2273756,1.5827163,1.938057,3.0602808,4.1825047,5.3047285,6.4269524,7.549176,8.165584,8.780178,9.394773,10.009366,10.625773,9.7483,8.870826,7.993352,7.115878,6.2384043,6.445082,6.6517596,6.8602505,7.066928,7.2754188,6.8529987,6.430578,6.008158,5.5857377,5.163317,6.0843024,7.0071006,7.9298983,8.852696,9.775495,10.038374,10.29944,10.56232,10.825199,11.088079,10.741803,10.397341,10.052877,9.706602,9.362139,10.576823,11.793322,13.008006,14.222692,15.437376,16.091856,16.748148,17.402628,18.057108,18.7134,19.13582,19.55824,19.980661,20.40308,20.8255,18.938208,17.050913,15.161806,13.274512,11.3872175,16.537846,21.686659,26.837286,31.987911,37.136726,34.384647,31.63257,28.880493,26.126604,23.374527,22.516994,21.659464,20.801933,19.9444,19.08687,18.611874,18.136877,17.661882,17.186886,16.71189,16.294909,15.877926,15.459132,15.0421505,14.625169,15.986704,17.350052,18.7134,20.074934,21.438282,19.804804,18.173138,16.539658,14.907991,13.274512,14.347786,15.419247,16.492521,17.565794,18.637255,16.566853,14.498261,12.427858,10.357455,8.287052,7.5618668,6.836682,6.11331,5.388125,4.6629395,6.2184615,7.7721705,9.327692,10.883214,12.436923,10.73999,9.043057,7.344311,5.6473784,3.9504454,4.36924,4.7898474,5.2104545,5.6292486,6.049856,7.4802837,8.910711,10.339326,11.769753,13.200181,14.248073,15.294152,16.342045,17.389936,18.43783,17.567608,16.697386,15.827164,14.956942,14.0867195,15.462758,16.836983,18.213022,19.587248,20.963285,21.99305,23.022812,24.052574,25.082336,26.1121,26.652363,27.192625,27.73289,28.273151,28.811602,25.042452,21.273302,17.50234,13.7331915,9.96223,9.151835,8.343254,7.5328593,6.722465,5.9120708,5.516845,5.121619,4.7282066,4.3329806,3.9377546,3.247016,2.5580902,1.8673514,1.1766127,0.48768693,0.8974165,1.3071461,1.7168756,2.126605,2.5381477,2.7720199,3.007705,3.24339,3.4772623,3.7129474,4.780782,5.846804,6.9146395,7.9824743,9.050309,12.542075,16.035654,19.52742,23.019186,26.512764,23.82958,21.148209,18.465023,15.781839,13.100468,13.918114,14.73576,15.553406,16.36924,17.186886,16.748148,16.307598,15.867048,15.428311,14.9877615,16.632118,18.278288,19.922646,21.567003,23.213173,23.439793,23.668226,23.894846,24.12328,24.349901,24.393412,24.43511,24.476809,24.520319,24.562017,22.535126,20.508232,18.479528,16.452635,14.425743,12.866595,11.30926,9.751925,8.194591,6.637256,10.997431,15.357606,19.717781,24.077955,28.438131,27.074783,25.71325,24.349901,22.988365,21.625017,20.42665,19.230095,18.031725,16.83517,15.636803,16.887747,18.136877,19.387821,20.636953,21.887897,22.174345,22.462606,22.750868,23.037315,23.325577,22.99018,22.654781,22.319382,21.985798,21.650398,20.169209,18.68983,17.210453,15.729263,14.249886,14.242634,14.235382,14.22813,14.220879,14.211814,14.367728,14.521831,14.677745,14.831847,14.9877615,14.22813,13.466686,12.707055,11.947423,11.187792,11.443419,11.697234,11.952863,12.206677,12.462305,12.837588,13.212872,13.588155,13.961625,14.336908,16.01571,17.692701,19.369692,21.046682,22.725487,20.152891,17.580297,15.007704,12.43511,9.862516,12.230246,14.597975,16.965704,19.33162,21.699348,20.214533,18.729717,17.2449,15.760084,14.275268,13.305332,12.335398,11.365462,10.395528,9.425592,0.012690738,0.014503701,0.018129626,0.01994259,0.02175555,0.025381476,0.027194439,0.030820364,0.032633327,0.034446288,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.034446288,0.032633327,0.030820364,0.027194439,0.025381476,0.02175555,0.01994259,0.018129626,0.014503701,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.15047589,0.25018883,0.34990177,0.44961473,0.5493277,0.8430276,1.1349145,1.4268016,1.7205015,2.0123885,1.6352923,1.258196,0.8792868,0.50219065,0.12509441,0.17041849,0.21574254,0.25925365,0.3045777,0.34990177,1.1040943,1.8600996,2.6142921,3.3702974,4.12449,5.1905117,6.2547207,7.320743,8.384952,9.449161,10.589515,11.729868,12.870221,14.010575,15.149116,14.791962,14.434808,14.077655,13.720501,13.363347,13.162108,12.962683,12.763257,12.562017,12.362592,11.927481,11.49237,11.057259,10.622148,10.1870365,8.9596615,7.7322855,6.5049095,5.277534,4.0501585,4.3202896,4.590421,4.860553,5.130684,5.4008155,5.823236,6.245656,6.6680765,7.0904965,7.512917,7.2953615,7.077806,6.8602505,6.642695,6.4251394,6.352621,6.2801023,6.207584,6.1350656,6.0625467,5.8431783,5.621997,5.4026284,5.18326,4.9620786,4.2024474,3.442816,2.6831846,1.9217403,1.162109,0.93911463,0.7179332,0.4949388,0.27194437,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.3208944,0.58921283,0.85934424,1.1294757,1.3996071,1.7005589,1.9996977,2.3006494,2.5997884,2.9007401,2.570781,2.2408218,1.9108626,1.5790904,1.2491312,1.0098201,0.7705091,0.5293851,0.29007402,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.2853905,2.570781,3.8543584,5.139749,6.4251394,6.628191,6.82943,7.0324817,7.2355337,7.4367723,7.3497505,7.262728,7.175706,7.0868707,6.9998484,6.887445,6.775041,6.6626377,6.550234,6.43783,6.300045,6.16226,6.0244746,5.8866897,5.750717,5.2666564,4.784408,4.3021603,3.8199122,3.3376641,3.2053177,3.0729716,2.9406252,2.808279,2.6741197,2.1882458,1.7005589,1.2128719,0.72518504,0.2374981,0.21211663,0.18673515,0.16316663,0.13778515,0.11240368,0.09064813,0.06707962,0.045324065,0.02175555,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.059827764,0.07070554,0.07977036,0.09064813,0.099712946,0.13053331,0.15954071,0.19036107,0.21936847,0.25018883,0.21030366,0.17041849,0.13053331,0.09064813,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.072518505,0.09427405,0.11784257,0.13959812,0.16316663,0.13053331,0.09789998,0.065266654,0.032633327,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.05076295,0.07977036,0.11059072,0.13959812,0.17041849,0.19942589,0.15954071,0.11965553,0.07977036,0.03988518,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.052575916,0.06707962,0.08339628,0.09789998,0.11240368,0.45324063,0.79226464,1.1331016,1.4721256,1.8129625,2.9932013,4.171627,5.351866,6.532104,7.7123427,8.319685,8.927028,9.53437,10.141713,10.750868,9.768243,8.785617,7.802991,6.8203654,5.8377395,5.9356394,6.0317264,6.1296263,6.2275267,6.3254266,6.1822023,6.0407915,5.8975673,5.754343,5.612932,6.742408,7.8718834,9.003172,10.1326475,11.262123,11.225864,11.187792,11.14972,11.111648,11.075388,10.277685,9.479981,8.682278,7.8845744,7.0868707,7.6579537,8.227224,8.798307,9.367578,9.936848,11.927481,13.918114,15.906934,17.897566,19.888199,20.404894,20.921589,21.440096,21.956789,22.475298,20.136576,17.799667,15.462758,13.125849,10.7871275,18.062546,25.337965,32.613384,39.88699,47.162407,41.66732,36.17223,30.67714,25.18205,19.68696,19.514729,19.342497,19.170267,18.998035,18.825804,17.562168,16.300346,15.036712,13.77489,12.513068,12.96087,13.406858,13.85466,14.302462,14.750263,16.08823,17.424383,18.76235,20.100317,21.438282,20.39039,19.342497,18.294605,17.246714,16.200634,17.505966,18.809486,20.11482,21.420153,22.725487,20.377699,18.029913,15.682126,13.33434,10.988366,9.949538,8.912524,7.8755093,6.836682,5.7996674,7.3406854,8.87989,10.420909,11.9601145,13.499319,11.782444,10.065568,8.34688,6.630004,4.9131284,4.5469103,4.1825047,3.8180993,3.4518807,3.0874753,4.064662,5.041849,6.0208488,6.9980354,7.9752226,9.043057,10.110892,11.176914,12.244749,13.312584,13.153044,12.99169,12.8321495,12.672608,12.513068,13.363347,14.211814,15.062093,15.912373,16.762651,18.102432,19.442211,20.78199,22.121769,23.463362,24.745127,26.026892,27.310469,28.592234,29.87581,25.37785,20.87989,16.38193,11.885782,7.3878226,6.506723,5.6274357,4.748149,3.8670492,2.9877625,3.43919,3.8924308,4.345671,4.797099,5.2503395,4.2804046,3.3104696,2.3405347,1.3705997,0.40066472,0.6055295,0.8103943,1.015259,1.2201238,1.4249886,1.6425442,1.8600996,2.077655,2.2952106,2.5127661,3.926877,5.3428006,6.7569118,8.172835,9.5869465,13.827466,18.067986,22.308504,26.54721,30.787731,27.789091,24.792263,21.795437,18.796797,15.799969,16.401873,17.005589,17.607492,18.209396,18.813112,18.691645,18.57199,18.452333,18.332678,18.213022,20.098503,21.982172,23.867653,25.753134,27.6368,27.40837,27.178122,26.947876,26.71763,26.487383,26.427555,26.367727,26.3079,26.248072,26.188244,24.266504,22.34839,20.42665,18.506721,16.586794,14.452938,12.317267,10.181598,8.047741,5.9120708,10.718235,15.522586,20.326937,25.1331,29.93745,29.299288,28.66294,28.024776,27.388426,26.750263,25.307144,23.865839,22.422722,20.979603,19.538298,19.862818,20.187338,20.511858,20.838192,21.162712,21.336756,21.512613,21.686659,21.862516,22.038374,22.107265,22.17797,22.246864,22.31757,22.388275,20.548119,18.70796,16.867804,15.027647,13.1874895,13.301706,13.417736,13.531953,13.647983,13.762199,14.139296,14.518205,14.895301,15.272397,15.649493,14.594349,13.539205,12.485873,11.430729,10.375585,10.8143215,11.254871,11.695421,12.134158,12.574709,12.862969,13.149418,13.437678,13.724127,14.012388,15.569723,17.127058,18.684393,20.241728,21.800875,19.53286,17.264843,14.996826,12.730623,10.462607,13.153044,15.84348,18.532103,21.22254,23.912977,21.90784,19.902702,17.897566,15.89243,13.887294,12.839401,11.791509,10.745429,9.697536,8.649645,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.18673515,0.31182957,0.43692398,0.5620184,0.6871128,1.0497054,1.4122978,1.7748904,2.137483,2.5000753,2.0250793,1.550083,1.0750868,0.6000906,0.12509441,0.17585737,0.22480737,0.2755703,0.3245203,0.37528324,1.261822,2.1501737,3.0367124,3.925064,4.8116026,5.9882154,7.1630154,8.337815,9.512614,10.687414,12.175857,13.662486,15.1509285,16.637558,18.124187,17.400814,16.67563,15.950445,15.22526,14.500074,14.0867195,13.675177,13.261822,12.850279,12.436923,11.874905,11.312886,10.750868,10.1870365,9.625018,8.287052,6.9508986,5.612932,4.274966,2.9369993,3.299592,3.6621845,4.024777,4.3873696,4.749962,5.125245,5.5005283,5.8758116,6.249282,6.624565,6.350808,6.0752378,5.7996674,5.524097,5.2503395,5.3119802,5.375434,5.4370747,5.5005283,5.562169,5.57486,5.5875506,5.600241,5.612932,5.6256227,4.788034,3.9504454,3.1128569,2.275268,1.4376793,1.162109,0.8883517,0.61278135,0.33721104,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.40066472,0.73787576,1.0750868,1.4122978,1.7495089,2.124792,2.5000753,2.8753586,3.2506418,3.6241121,3.2125697,2.7992141,2.3876717,1.9743162,1.5627737,1.261822,0.96268314,0.66173136,0.36259252,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.6008459,3.199879,4.800725,6.399758,8.000604,7.9625316,7.9244595,7.8882003,7.850128,7.8120556,8.000604,8.187339,8.375887,8.562622,8.749357,8.287052,7.8247466,7.362441,6.9001355,6.43783,6.249282,6.0625467,5.8758116,5.6872635,5.5005283,4.974769,4.4508233,3.925064,3.3993049,2.8753586,2.7883365,2.6995013,2.612479,2.525457,2.4366217,1.9996977,1.5627737,1.1258497,0.6871128,0.25018883,0.22480737,0.19942589,0.17585737,0.15047589,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.16316663,0.19942589,0.2374981,0.2755703,0.31182957,0.25018883,0.18673515,0.12509441,0.06164073,0.0,0.0,0.0,0.0,0.0,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.099712946,0.13778515,0.17585737,0.21211663,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.387974,0.7124943,1.0370146,1.3633479,1.6878681,2.9243085,4.162562,5.4008155,6.637256,7.8755093,8.4756,9.07569,9.675781,10.275872,10.874149,9.788185,8.700407,7.61263,6.5248523,5.4370747,5.424384,5.411693,5.4008155,5.388125,5.375434,5.5132194,5.6491914,5.7869763,5.924762,6.0625467,7.400513,8.736667,10.074633,11.4126,12.750566,12.413355,12.07433,11.73712,11.399909,11.062697,9.811753,8.562622,7.311678,6.0625467,4.8116026,4.7372713,4.6629395,4.5867953,4.512464,4.4381323,7.763106,11.088079,14.413053,17.738026,21.063,21.675781,22.286749,22.89953,23.512312,24.125093,21.336756,18.550234,15.761897,12.975373,10.1870365,19.587248,28.98746,38.38767,47.78788,57.18809,48.94999,40.711887,32.475597,24.237497,15.999394,16.512463,17.025532,17.536787,18.049856,18.562923,16.512463,14.462003,12.411542,10.362894,8.312433,9.625018,10.937603,12.250188,13.562773,14.875358,16.187943,17.500528,18.813112,20.125698,21.438282,20.974165,20.511858,20.049553,19.587248,19.124943,20.662334,22.199726,23.73712,25.274511,26.811903,24.186733,21.563377,18.938208,16.313038,13.687867,12.337211,10.988366,9.637709,8.287052,6.9382076,8.46291,9.987611,11.512312,13.037014,14.561715,12.824898,11.088079,9.349448,7.61263,5.8758116,4.7245803,3.5751622,2.4257438,1.2745126,0.12509441,0.6508536,1.1747998,1.7005589,2.2245052,2.7502642,3.8380418,4.9258194,6.011784,7.0995617,8.187339,8.736667,9.287807,9.837135,10.388275,10.937603,11.262123,11.586644,11.912977,12.237497,12.562017,14.211814,15.861609,17.513218,19.163015,20.81281,22.837889,24.862968,26.888048,28.913128,30.938206,25.711435,20.48829,15.261519,10.036561,4.8116026,3.8616104,2.913431,1.9616255,1.0116332,0.06164073,1.3633479,2.663242,3.9631362,5.2630305,6.5629244,5.3119802,4.062849,2.811905,1.5627737,0.31182957,0.31182957,0.31182957,0.31182957,0.31182957,0.31182957,0.51306844,0.7124943,0.9119202,1.1131591,1.3125849,3.0747845,4.836984,6.599184,8.363196,10.125396,15.112856,20.100317,25.087776,30.075235,35.062695,31.750414,28.438131,25.124035,21.811752,18.49947,18.887444,19.275417,19.663393,20.049553,20.437527,20.636953,20.838192,21.037619,21.237043,21.438282,23.563074,25.687866,27.812658,29.93745,32.062244,31.37513,30.688017,29.999092,29.31198,28.624866,28.4617,28.300346,28.137178,27.975826,27.812658,25.999697,24.186733,22.375584,20.562622,18.749659,16.037468,13.325275,10.613083,7.900891,5.186886,10.437225,15.687565,20.937904,26.186432,31.436771,31.525606,31.612629,31.69965,31.786673,31.875507,30.18764,28.499771,26.811903,25.125849,23.43798,22.837889,22.237799,21.637709,21.037619,20.437527,20.499168,20.562622,20.624262,20.687716,20.749357,21.224354,21.699348,22.174345,22.649342,23.124338,20.925215,18.724277,16.525154,14.326031,12.125093,12.362592,12.60009,12.837588,13.075087,13.312584,13.912675,14.512766,15.112856,15.712947,16.313038,14.96238,13.611723,12.262879,10.912222,9.563377,10.1870365,10.812509,11.437981,12.06164,12.687112,12.888351,13.087777,13.287203,13.486629,13.687867,15.125546,16.563227,18.000906,19.436771,20.87445,18.912827,16.949387,14.9877615,13.024323,11.062697,14.075842,17.087172,20.100317,23.111647,26.12479,23.599335,21.073877,18.550234,16.024776,13.499319,12.375282,11.249433,10.125396,8.999546,7.8755093,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.11059072,0.21936847,0.32995918,0.4405499,0.5493277,0.6417888,0.73424983,0.82671094,0.91917205,1.0116332,1.3633479,1.7132497,2.0631514,2.4130533,2.762955,3.1201086,3.4772623,3.834416,4.1933823,4.550536,4.0120864,3.4754493,2.9369993,2.4003625,1.8619126,2.0903459,2.3169663,2.5453994,2.7720199,3.000453,3.9848917,4.9693303,5.955582,6.9400206,7.9244595,9.1500225,10.375585,11.599335,12.824898,14.05046,14.752076,15.455506,16.157122,16.860552,17.562168,16.646622,15.732889,14.817343,13.901797,12.988064,12.618219,12.248375,11.876718,11.506873,11.137029,10.897718,10.658407,10.417283,10.177972,9.936848,8.660522,7.382384,6.104245,4.8279195,3.5497808,3.6422417,3.7347028,3.827164,3.919625,4.0120864,4.2804046,4.5469103,4.8152285,5.081734,5.3500524,5.2503395,5.1506267,5.049101,4.949388,4.8496747,4.940323,5.029158,5.1198063,5.2104545,5.2992897,5.230397,5.1596913,5.090799,5.0200934,4.949388,4.1970086,3.444629,2.6922495,1.93987,1.1874905,1.1258497,1.062396,1.0007553,0.93730164,0.87566096,0.8448406,0.81583315,0.7850128,0.7541924,0.72518504,0.99531645,1.2654479,1.5355793,1.8057107,2.0758421,2.5073273,2.9406252,3.3721104,3.8054085,4.2368937,3.9649491,3.6930048,3.4192474,3.147303,2.8753586,2.5671551,2.2607644,1.9525607,1.6443571,1.3379664,1.452183,1.5682126,1.6824293,1.7966459,1.9126755,1.8057107,1.696933,1.5899682,1.4830034,1.3742256,1.2183108,1.0605831,0.90285534,0.7451276,0.5873999,0.69255173,0.79770356,0.90285534,1.0080072,1.1131591,1.4177368,1.7223145,2.0268922,2.333283,2.6378605,4.137181,5.638314,7.137634,8.636953,10.138086,9.860703,9.583321,9.304124,9.026741,8.749357,8.664148,8.580752,8.495543,8.410334,8.325124,8.105756,7.8845744,7.665206,7.4458375,7.224656,7.3298078,7.4349594,7.5401115,7.645263,7.750415,7.413204,7.07418,6.736969,6.399758,6.0625467,5.8522434,5.6419396,5.431636,5.223145,5.0128417,4.5450974,4.077353,3.6096084,3.141864,2.6741197,2.5544643,2.4348087,2.3151531,2.1954978,2.0758421,1.6733645,1.2708868,0.8665961,0.46411842,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.072518505,0.14503701,0.21755551,0.29007402,0.36259252,0.29007402,0.21755551,0.14503701,0.072518505,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.059827764,0.07070554,0.07977036,0.09064813,0.099712946,0.13053331,0.15954071,0.19036107,0.21936847,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.054388877,0.08520924,0.11421664,0.14503701,0.17585737,0.14322405,0.11059072,0.07795739,0.045324065,0.012690738,0.014503701,0.018129626,0.01994259,0.02175555,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.099712946,0.19942589,0.2991388,0.40066472,0.50037766,0.4550536,0.40972954,0.36440548,0.3208944,0.2755703,0.37165734,0.46955732,0.56745726,0.6653573,0.76325727,0.68167394,0.60190356,0.52213323,0.44236287,0.36259252,0.29007402,0.21755551,0.14503701,0.072518505,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.37528324,0.6871128,1.0007553,1.3125849,1.6244144,2.855416,4.0846047,5.315606,6.544795,7.7757964,8.180087,8.584378,8.990481,9.394773,9.800876,8.8672,7.935337,7.0016613,6.069799,5.137936,5.2630305,5.388125,5.5132194,5.638314,5.763408,5.6927023,5.621997,5.5531044,5.482399,5.411693,6.4704633,7.5274205,8.584378,9.643148,10.700105,10.774437,10.850581,10.924912,10.999244,11.075388,9.630457,8.185526,6.740595,5.295664,3.8507326,3.7945306,3.7401419,3.6857529,3.6295512,3.5751622,6.319988,9.064813,11.809638,14.554463,17.29929,18.133251,18.9654,19.797552,20.629702,21.461851,19.43496,17.408066,15.379361,13.352469,11.325577,18.967215,26.610664,34.2523,41.895752,49.537388,42.610058,35.682728,28.7554,21.82807,14.90074,15.529838,16.160748,16.789846,17.420757,18.049856,17.304728,16.5596,15.814472,15.0693445,14.324218,14.126604,13.930804,13.7331915,13.535579,13.337966,14.904366,16.472578,18.04079,19.607191,21.175404,20.660522,20.14564,19.630758,19.115877,18.599184,19.337059,20.074934,20.81281,21.550686,22.286749,20.172834,18.057108,15.9431925,13.827466,11.711739,10.607644,9.501737,8.397643,7.2917356,6.187641,7.877322,9.567003,11.256684,12.948178,14.63786,13.274512,11.912977,10.549629,9.188094,7.8247466,6.319988,4.8152285,3.3104696,1.8057107,0.2991388,1.8329052,3.3648586,4.896812,6.430578,7.9625316,7.6833353,7.402326,7.12313,6.8421206,6.5629244,7.995165,9.427405,10.859646,12.291886,13.724127,12.989877,12.255627,11.519565,10.785315,10.049252,11.3872175,12.725184,14.06315,15.399304,16.73727,18.33993,19.942589,21.545248,23.147905,24.750565,20.575312,16.400059,12.224807,8.049554,3.874301,3.825351,3.774588,3.7256382,3.6748753,3.6241121,3.9522583,4.2804046,4.606738,4.934884,5.2630305,4.702825,4.1426196,3.5824142,3.0222087,2.4620032,2.268016,2.0722163,1.8782293,1.6824293,1.4866294,1.4195497,1.35247,1.2853905,1.2183108,1.1494182,2.9333735,4.7155156,6.497658,8.2798,10.061942,14.275268,18.48678,22.700104,26.91343,31.12494,28.197006,25.270885,22.34295,19.415016,16.487082,16.492521,16.49796,16.501585,16.507025,16.512463,17.29929,18.087927,18.874754,19.66158,20.450218,22.203352,23.954674,25.70781,27.459131,29.212267,28.361986,27.511707,26.66324,25.812962,24.962683,24.609154,24.257439,23.905725,23.552197,23.200481,22.25049,21.300497,20.350506,19.400513,18.45052,16.066475,13.684241,11.302009,8.919776,6.5375433,11.218613,15.897869,20.577126,25.256382,29.93745,30.41426,30.892883,31.369692,31.848314,32.325123,30.65901,28.99471,27.33041,25.664299,23.999998,23.069948,22.139898,21.209848,20.279799,19.34975,19.706903,20.06587,20.423023,20.780178,21.137331,21.44916,21.762802,22.074633,22.388275,22.700104,20.9651,19.230095,17.495089,15.760084,14.025079,14.075842,14.124791,14.175554,14.224504,14.275268,14.684997,15.094727,15.504456,15.914186,16.325727,15.676687,15.02946,14.382232,13.735004,13.087777,13.200181,13.312584,13.424988,13.537392,13.649796,13.716875,13.785768,13.852847,13.919927,13.987006,15.094727,16.202446,17.310167,18.417887,19.525606,18.747847,17.970085,17.192324,16.414564,15.636803,17.819609,20.002417,22.185223,24.36803,26.550837,23.978243,21.403835,18.833055,16.260462,13.687867,12.335398,10.982927,9.630457,8.2779875,6.925517,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.21936847,0.4405499,0.65991837,0.8792868,1.1004683,1.2726997,1.4449311,1.6171626,1.789394,1.9616255,2.5381477,3.1128569,3.6875658,4.262275,4.836984,5.1905117,5.542227,5.8957543,6.247469,6.599184,6.000906,5.4008155,4.800725,4.2006345,3.6005437,4.004834,4.409125,4.8152285,5.219519,5.6256227,6.7079616,7.7903004,8.872639,9.954978,11.037316,12.311829,13.588155,14.862667,16.13718,17.411694,17.330109,17.246714,17.16513,17.081734,17.00015,15.894243,14.790149,13.684241,12.580148,11.47424,11.147907,10.81976,10.491614,10.165281,9.837135,9.920531,10.002114,10.085511,10.167094,10.25049,9.03218,7.8156815,6.5973706,5.3808727,4.162562,3.9848917,3.8072214,3.6295512,3.4518807,3.2742105,3.435564,3.5951047,3.7546456,3.9141862,4.07554,4.1498713,4.2242026,4.3003473,4.3746786,4.4508233,4.5668526,4.6846952,4.802538,4.9203806,5.038223,4.8841214,4.7318325,4.5795436,4.4272547,4.274966,3.6077955,2.9406252,2.2716422,1.6044719,0.93730164,1.0877775,1.2382535,1.3869164,1.5373923,1.6878681,1.6280404,1.5682126,1.5083848,1.4467441,1.3869164,1.5899682,1.79302,1.9942589,2.1973107,2.4003625,2.8898623,3.3793623,3.870675,4.360175,4.8496747,4.7173285,4.5849824,4.4526362,4.3202896,4.1879435,3.872488,3.5570326,3.24339,2.9279346,2.612479,2.855416,3.0983531,3.339477,3.5824142,3.825351,3.6096084,3.395679,3.1799364,2.9641938,2.7502642,2.4348087,2.1193533,1.8057107,1.4902552,1.1747998,1.3851035,1.5954071,1.8057107,2.0142014,2.2245052,2.8354735,3.444629,4.0555973,4.664753,5.275721,6.6753283,8.074935,9.474543,10.874149,12.27557,11.757062,11.240368,10.721861,10.205167,9.686659,9.329506,8.972352,8.615198,8.258044,7.900891,7.9226465,7.944402,7.9679704,7.989726,8.013294,8.410334,8.807372,9.2044115,9.603263,10.000301,9.849826,9.699349,9.550687,9.400211,9.249735,8.917963,8.584378,8.252605,7.9208336,7.5872483,7.0904965,6.591932,6.09518,5.5966153,5.0998635,4.8841214,4.670192,4.454449,4.2405195,4.024777,3.245203,2.465629,1.6842422,0.90466833,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.14503701,0.29007402,0.43511102,0.58014804,0.72518504,0.58014804,0.43511102,0.29007402,0.14503701,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.045324065,0.052575916,0.059827764,0.06707962,0.07433146,0.09789998,0.11965553,0.14322405,0.16497959,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.072518505,0.09427405,0.11784257,0.13959812,0.16316663,0.13415924,0.10696479,0.07977036,0.052575916,0.025381476,0.030820364,0.034446288,0.03988518,0.045324065,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.17585737,0.34990177,0.52575916,0.69980353,0.87566096,0.79770356,0.7197462,0.6417888,0.5656443,0.48768693,0.64541465,0.8031424,0.96087015,1.1167849,1.2745126,1.1657349,1.0551442,0.9445535,0.83577573,0.72518504,0.58014804,0.43511102,0.29007402,0.14503701,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.36259252,0.66173136,0.96268314,1.261822,1.5627737,2.7847104,4.006647,5.230397,6.452334,7.6742706,7.8845744,8.094878,8.3051815,8.515485,8.725789,7.948028,7.170267,6.392506,5.614745,4.836984,5.0998635,5.3627434,5.6256227,5.8866897,6.149569,5.8721857,5.5948024,5.317419,5.040036,4.762653,5.540414,6.3181744,7.0941224,7.8718834,8.649645,9.137331,9.625018,10.112705,10.600392,11.088079,9.447348,7.8084297,6.167699,4.5269675,2.8880494,2.8517902,2.817344,2.7828975,2.7466383,2.712192,4.876869,7.041547,9.208037,11.372714,13.537392,14.590723,15.6422415,16.695572,17.747091,18.800423,17.533161,16.2659,14.996826,13.729566,12.462305,18.347181,24.232058,30.116934,36.001812,41.88669,36.27013,30.653572,25.0352,19.41683,13.800271,14.547212,15.294152,16.042906,16.789846,17.536787,18.096992,18.657198,19.217403,19.777609,20.337814,18.630003,16.922194,15.214382,13.506571,11.800573,13.622601,15.444629,17.266655,19.090496,20.912523,20.345066,19.777609,19.210152,18.642694,18.075237,18.011784,17.950142,17.886688,17.825048,17.763407,16.157122,14.55265,12.948178,11.341894,9.737422,8.8780775,8.01692,7.157576,6.298232,5.4370747,7.2917356,9.14821,11.00287,12.857531,14.712192,13.724127,12.737875,11.74981,10.761745,9.775495,7.915395,6.055295,4.195195,2.335096,0.4749962,3.0149567,5.5549173,8.094878,10.634838,13.174799,11.526816,9.880646,8.232663,6.58468,4.936697,7.25185,9.567003,11.882156,14.19731,16.512463,14.71763,12.922797,11.127964,9.333132,7.5382986,8.562622,9.5869465,10.613083,11.637406,12.661731,13.8419695,15.022208,16.202446,17.382685,18.562923,15.437376,12.311829,9.188094,6.0625467,2.9369993,3.787279,4.6375585,5.487838,6.338117,7.1883965,6.542982,5.8975673,5.2521524,4.606738,3.9631362,4.0918565,4.2223897,4.3529234,4.4816437,4.612177,4.2223897,3.832603,3.442816,3.053029,2.663242,2.327844,1.9924458,1.6570477,1.3216497,0.9880646,2.7901495,4.592234,6.394319,8.198216,10.000301,13.437678,16.875055,20.312433,23.74981,27.187187,24.645412,22.101828,19.560053,17.01828,14.474693,14.097597,13.720501,13.341592,12.964496,12.5873995,13.963438,15.337664,16.71189,18.087927,19.462152,20.841818,22.223295,23.60296,24.982624,26.36229,25.350657,24.33721,23.325577,22.31213,21.300497,20.756609,20.214533,19.672457,19.13038,18.588305,18.49947,18.412449,18.325426,18.238403,18.149569,16.097294,14.045021,11.992747,9.940474,7.8882003,11.998186,16.108173,20.218159,24.328144,28.438131,29.304728,30.173136,31.039732,31.908142,32.77474,31.132193,29.489649,27.847105,26.204561,24.562017,23.302008,22.042,20.78199,19.52198,18.261972,18.914639,19.567305,20.219973,20.872639,21.525305,21.675781,21.824444,21.97492,22.125395,22.275871,21.004984,19.734098,18.465023,17.19595,15.925063,15.787278,15.649493,15.511708,15.375735,15.23795,15.457319,15.676687,15.897869,16.117237,16.336605,16.392807,16.447197,16.503399,16.557787,16.612177,16.213324,15.812659,15.411995,15.013144,14.612478,14.547212,14.481945,14.416678,14.353225,14.287958,15.065719,15.84348,16.619429,17.397188,18.17495,18.582867,18.990784,19.396887,19.804804,20.212719,21.56519,22.91766,24.27013,25.6226,26.97507,24.35534,21.733795,19.114065,16.494333,13.874602,12.295512,10.714609,9.135518,7.554615,5.975525,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.32995918,0.65991837,0.9898776,1.3198367,1.649796,1.9017978,2.1556125,2.4076142,2.659616,2.911618,3.7129474,4.512464,5.3119802,6.11331,6.9128265,7.2591023,7.607191,7.95528,8.303369,8.649645,7.987913,7.324369,6.6626377,5.999093,5.337362,5.919323,6.5030966,7.0850577,7.667019,8.2507925,9.429218,10.609457,11.789696,12.969934,14.150173,15.475449,16.800724,18.124187,19.449463,20.774738,19.908142,19.039734,18.173138,17.304728,16.438131,15.141864,13.847408,12.552953,11.256684,9.96223,9.677594,9.39296,9.108324,8.821876,8.537241,8.943344,9.347635,9.751925,10.15803,10.56232,9.40565,8.247167,7.0904965,5.9320135,4.7753434,4.327542,3.87974,3.4319382,2.9841363,2.5381477,2.5907235,2.6432993,2.6958754,2.7466383,2.7992141,3.049403,3.299592,3.5497808,3.7999697,4.0501585,4.195195,4.3402324,4.4852695,4.6303062,4.7753434,4.539658,4.305786,4.070101,3.834416,3.6005437,3.0167696,2.4348087,1.8528478,1.2708868,0.6871128,1.0497054,1.4122978,1.7748904,2.137483,2.5000753,2.4094272,2.3205922,2.229944,2.1392958,2.0504606,2.18462,2.3205922,2.4547513,2.5907235,2.7248828,3.2723975,3.8199122,4.367427,4.914942,5.462456,5.469708,5.47696,5.484212,5.4932766,5.5005283,5.177821,4.855114,4.5324063,4.209699,3.8869917,4.256836,4.6266804,4.9983377,5.368182,5.7380266,5.4153194,5.092612,4.7699046,4.4471974,4.12449,3.6531196,3.1799364,2.7067533,2.2353828,1.7621996,2.077655,2.3931105,2.7067533,3.0222087,3.3376641,4.25321,5.1669436,6.0824895,6.9980354,7.911769,9.211663,10.51337,11.813264,13.113158,14.413053,13.655234,12.897416,12.139598,11.381779,10.625773,9.994863,9.365765,8.734854,8.105756,7.474845,7.7395372,8.00423,8.270736,8.535428,8.80012,9.490859,10.179785,10.870523,11.559449,12.250188,12.28826,12.32452,12.362592,12.400664,12.436923,11.98187,11.526816,11.071762,10.616709,10.161655,9.635896,9.108324,8.580752,8.05318,7.5256076,7.215591,6.9055743,6.5955577,6.285541,5.975525,4.8170414,3.6603715,2.5018883,1.3452182,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.21755551,0.43511102,0.6526665,0.87022203,1.0877775,0.87022203,0.6526665,0.43511102,0.21755551,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.030820364,0.034446288,0.03988518,0.045324065,0.05076295,0.065266654,0.07977036,0.09427405,0.11059072,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.09064813,0.10515183,0.11965553,0.13415924,0.15047589,0.12690738,0.10515183,0.08339628,0.059827764,0.038072214,0.045324065,0.052575916,0.059827764,0.06707962,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.25018883,0.50037766,0.7505665,1.0007553,1.2491312,1.1403534,1.0297627,0.91917205,0.8103943,0.69980353,0.91735905,1.1349145,1.35247,1.5700256,1.7875811,1.647983,1.5083848,1.3669738,1.2273756,1.0877775,0.87022203,0.6526665,0.43511102,0.21755551,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.34990177,0.63816285,0.9246109,1.2128719,1.49932,2.715818,3.930503,5.145188,6.359873,7.574558,7.590874,7.605378,7.6198816,7.6343856,7.650702,7.027043,6.4051967,5.7833505,5.1596913,4.537845,4.936697,5.337362,5.7380266,6.1368785,6.5375433,6.051669,5.567608,5.081734,4.597673,4.1117992,4.610364,5.1071157,5.6056805,6.1024323,6.599184,7.500226,8.399456,9.300498,10.199727,11.10077,9.264238,7.4295206,5.5948024,3.7600844,1.9253663,1.9108626,1.8945459,1.8800422,1.8655385,1.8492218,3.435564,5.0200934,6.604623,8.189152,9.775495,11.048194,12.31908,13.591781,14.86448,16.13718,15.62955,15.121921,14.614291,14.106662,13.600845,17.727148,21.855265,25.98338,30.109682,34.237797,29.930199,25.6226,21.315,17.007402,12.699803,13.564586,14.429369,15.294152,16.160748,17.025532,18.889257,20.754795,22.620335,24.485872,26.349598,23.13159,19.915394,16.697386,13.479377,10.263181,12.340837,14.416678,16.494333,18.57199,20.649643,20.02961,19.409578,18.789545,18.169512,17.549479,16.68832,15.825351,14.96238,14.09941,13.238253,12.143224,11.048194,9.953164,8.858135,7.763106,7.1466985,6.532104,5.91751,5.3029156,4.688321,6.7079616,8.727602,10.747242,12.766883,14.788336,14.175554,13.562773,12.949992,12.337211,11.724429,9.508988,7.2953615,5.0799212,2.864481,0.6508536,4.1970086,7.744976,11.292944,14.840912,18.387066,15.372109,12.357153,9.342196,6.3272395,3.3122826,6.510349,9.706602,12.904668,16.102734,19.3008,16.445383,13.589968,10.734551,7.8791356,5.0255322,5.7380266,6.450521,7.1630154,7.8755093,8.588004,9.345822,10.101828,10.859646,11.617464,12.375282,10.29944,8.225411,6.149569,4.07554,1.9996977,3.7492065,5.5005283,7.250037,8.999546,10.750868,9.131892,7.51473,5.8975673,4.2804046,2.663242,3.482701,4.3021603,5.123432,5.942891,6.7623506,6.1767635,5.5929894,5.0074024,4.421816,3.8380418,3.2343252,2.6324217,2.030518,1.4268016,0.824898,2.6469254,4.4707656,6.2927933,8.1148205,9.936848,12.60009,15.261519,17.92476,20.588003,23.249432,21.092007,18.934582,16.777155,14.61973,12.462305,11.702674,10.943042,10.181598,9.421967,8.662335,10.625773,12.5873995,14.5508375,16.512463,18.475903,19.482096,20.490103,21.49811,22.504305,23.512312,22.337511,21.162712,19.987913,18.813112,17.638313,16.904062,16.171627,15.439189,14.706753,13.974316,14.750263,15.524399,16.300346,17.074482,17.85043,16.128115,14.405801,12.681673,10.959359,9.237044,12.7777605,16.316664,19.85738,23.398094,26.936998,28.195194,29.451576,30.709774,31.96797,33.224354,31.605377,29.984589,28.365612,26.744823,25.125849,23.534067,21.945911,20.354132,18.765976,17.174194,18.122374,19.070553,20.01692,20.9651,21.913279,21.900587,21.887897,21.875206,21.862516,21.849825,21.04487,20.239914,19.43496,18.630003,17.825048,17.500528,17.174194,16.849674,16.525154,16.200634,16.229641,16.260462,16.289469,16.32029,16.349297,17.107115,17.864933,18.622751,19.38057,20.138388,19.224655,18.312735,17.400814,16.487082,15.575162,15.377548,15.179935,14.982323,14.78471,14.587097,15.034899,15.4827,15.930502,16.378304,16.824293,18.417887,20.009668,21.603262,23.195044,24.786825,25.31077,25.832903,26.355038,26.87717,27.399303,24.732435,22.065567,19.396887,16.730019,14.06315,12.255627,10.448103,8.640579,6.833056,5.0255322,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.4405499,0.8792868,1.3198367,1.7603867,2.1991236,2.5327086,2.864481,3.198066,3.529838,3.8616104,4.8877473,5.9120708,6.9382076,7.9625316,8.9868555,9.329506,9.672155,10.014805,10.357455,10.700105,9.97492,9.249735,8.52455,7.799365,7.07418,7.835624,8.595256,9.354887,10.114518,10.874149,12.152288,13.430427,14.706753,15.984891,17.26303,18.637255,20.013294,21.38752,22.761745,24.137783,22.484362,20.832752,19.17933,17.527721,15.8743,14.389484,12.904668,11.419851,9.935035,8.450218,8.207282,7.9643445,7.723221,7.4802837,7.2373466,7.9643445,8.693155,9.420154,10.147152,10.874149,9.7773075,8.680465,7.5818095,6.484967,5.388125,4.670192,3.9522583,3.2343252,2.518205,1.8002719,1.745883,1.6896812,1.6352923,1.5809034,1.5247015,1.9507477,2.374981,2.7992141,3.2252605,3.6494937,3.8217251,3.9957695,4.168001,4.3402324,4.512464,4.195195,3.877927,3.5606585,3.24339,2.9243085,2.427557,1.9308052,1.4322405,0.9354887,0.43692398,1.0116332,1.5881553,2.1628644,2.7375734,3.3122826,3.1926272,3.0729716,2.953316,2.8318477,2.712192,2.7792716,2.8481643,2.9152439,2.9823234,3.049403,3.6549325,4.2604623,4.8641787,5.469708,6.0752378,6.2220874,6.3707504,6.5176005,6.6644506,6.813113,6.4831543,6.153195,5.823236,5.4932766,5.163317,5.660069,6.156821,6.6553855,7.1521373,7.650702,7.219217,6.789545,6.359873,5.9302006,5.5005283,4.8696175,4.2405195,3.6096084,2.9805105,2.3495996,2.770207,3.1908143,3.6096084,4.0302157,4.4508233,5.669134,6.889258,8.109382,9.329506,10.549629,11.74981,12.949992,14.150173,15.350354,16.550535,15.553406,14.554463,13.557334,12.5602045,11.563075,10.66022,9.757364,8.854509,7.951654,7.0506115,7.558241,8.06587,8.571687,9.079316,9.5869465,10.5695715,11.552197,12.534823,13.517449,14.500074,14.724882,14.94969,15.174497,15.399304,15.624111,15.047589,14.4692545,13.892733,13.314397,12.737875,12.179482,11.622903,11.06451,10.507931,9.949538,9.545248,9.139144,8.734854,8.330563,7.9244595,6.390693,4.855114,3.3195345,1.7857682,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.29007402,0.58014804,0.87022203,1.1602961,1.4503701,1.1602961,0.87022203,0.58014804,0.29007402,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.014503701,0.018129626,0.01994259,0.02175555,0.025381476,0.032633327,0.03988518,0.047137026,0.054388877,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.10696479,0.11421664,0.12328146,0.13053331,0.13778515,0.11965553,0.10333887,0.08520924,0.06707962,0.05076295,0.059827764,0.07070554,0.07977036,0.09064813,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.3245203,0.6508536,0.97537386,1.2998942,1.6244144,1.4830034,1.3397794,1.1983683,1.0551442,0.9119202,1.1893034,1.4666867,1.745883,2.0232663,2.3006494,2.1302311,1.9598125,1.789394,1.6207886,1.4503701,1.1602961,0.87022203,0.58014804,0.29007402,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.33721104,0.61278135,0.8883517,1.162109,1.4376793,2.6451125,3.8525455,5.0599785,6.2674117,7.474845,7.2953615,7.115878,6.9345818,6.755099,6.5756154,6.107871,5.6401267,5.1723824,4.704638,4.2368937,4.7753434,5.3119802,5.8504305,6.3870673,6.925517,6.2329655,5.540414,4.847862,4.15531,3.4627585,3.680314,3.8978696,4.115425,4.3329806,4.550536,5.863121,7.175706,8.488291,9.800876,11.111648,9.082943,7.0524244,5.0219064,2.9932013,0.96268314,0.968122,0.97174793,0.97718686,0.9826257,0.9880646,1.9924458,2.9968271,4.0030212,5.0074024,6.011784,7.5056653,8.997733,10.489801,11.98187,13.475751,13.727753,13.979754,14.231756,14.485571,14.737573,17.107115,19.476658,21.848013,24.217554,26.587097,23.59027,20.593443,17.5948,14.597975,11.599335,12.581961,13.564586,14.547212,15.529838,16.512463,19.683334,22.852394,26.023266,29.192324,32.363194,27.634989,22.906782,18.18039,13.452183,8.725789,11.057259,13.390542,15.722012,18.055294,20.386765,19.714155,19.04336,18.37075,17.698141,17.025532,15.363045,13.700559,12.038072,10.375585,8.713099,8.127511,7.5419245,6.9581504,6.3725634,5.7869763,5.4171324,5.047288,4.6774435,4.307599,3.9377546,6.1223745,8.306994,10.493427,12.678047,14.862667,14.625169,14.387671,14.150173,13.912675,13.675177,11.104396,8.535428,5.964647,3.395679,0.824898,5.3808727,9.935035,14.49101,19.045172,23.599335,19.217403,14.835473,10.451729,6.069799,1.6878681,5.767034,9.848013,13.927178,18.008158,22.087322,18.173138,14.257137,10.342952,6.4269524,2.5127661,2.913431,3.3122826,3.7129474,4.1117992,4.512464,4.847862,5.18326,5.516845,5.8522434,6.187641,5.163317,4.137181,3.1128569,2.08672,1.062396,3.7129474,6.3616858,9.012237,11.662788,14.313339,11.722616,9.131892,6.542982,3.9522583,1.3633479,2.8717327,4.3819304,5.8921285,7.402326,8.912524,8.13295,7.3533764,6.5719895,5.7924156,5.0128417,4.1426196,3.2723975,2.4021754,1.5319533,0.66173136,2.5055144,4.347484,6.189454,8.033237,9.875207,11.762501,13.649796,15.537089,17.424383,19.311678,17.540413,15.767336,13.994258,12.222994,10.449916,9.30775,8.165584,7.021604,5.8794374,4.7372713,7.28811,9.837135,12.387974,14.936998,17.487837,18.122374,18.75691,19.393261,20.027798,20.662334,19.324368,17.988214,16.650248,15.312282,13.974316,13.05333,12.130532,11.207735,10.284937,9.362139,10.999244,12.638163,14.275268,15.912373,17.549479,16.157122,14.764768,13.372412,11.980057,10.587702,13.557334,16.526966,19.498413,22.468046,25.437677,27.08566,28.73183,30.379814,32.027798,33.67578,32.076748,30.479527,28.882307,27.285088,25.687866,23.767939,21.848013,19.928085,18.008158,16.08823,17.330109,18.57199,19.815681,21.05756,22.29944,22.125395,21.949537,21.775494,21.599636,21.425592,21.084755,20.745731,20.404894,20.06587,19.725033,19.211964,18.700708,18.187641,17.674572,17.163317,17.001963,16.842422,16.682882,16.52334,16.361988,17.823235,19.282671,20.742105,22.20154,23.662788,22.237799,20.81281,19.387821,17.962833,16.537846,16.207886,15.877926,15.547967,15.218008,14.888049,15.005891,15.121921,15.239763,15.357606,15.475449,18.252907,21.030367,23.807825,26.585283,29.362741,29.054539,28.748148,28.439943,28.13174,27.82535,25.109531,22.395527,19.679708,16.965704,14.249886,12.215742,10.179785,8.145641,6.109684,4.07554,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.5493277,1.1004683,1.649796,2.1991236,2.7502642,3.1618068,3.5751622,3.9867048,4.40006,4.8116026,6.0625467,7.311678,8.562622,9.811753,11.062697,11.399909,11.73712,12.07433,12.413355,12.750566,11.961927,11.175101,10.388275,9.599637,8.812811,9.750113,10.687414,11.624716,12.562017,13.499319,14.875358,16.249584,17.625622,18.999847,20.375887,21.800875,23.225864,24.650852,26.07584,27.50083,25.062395,22.625772,20.187338,17.750717,15.312282,13.637105,11.961927,10.28675,8.611572,6.9382076,6.736969,6.5375433,6.338117,6.1368785,5.9374523,6.987158,8.036863,9.088382,10.138086,11.187792,10.150778,9.11195,8.074935,7.037921,6.000906,5.0128417,4.024777,3.0367124,2.0504606,1.062396,0.89922947,0.73787576,0.5747091,0.41335547,0.25018883,0.85027945,1.4503701,2.0504606,2.6505513,3.2506418,3.4500678,3.6494937,3.8507326,4.0501585,4.249584,3.8507326,3.4500678,3.049403,2.6505513,2.2498865,1.8383441,1.4249886,1.0116332,0.6000906,0.18673515,0.97537386,1.7621996,2.5508385,3.3376641,4.12449,3.975827,3.825351,3.6748753,3.5243993,3.3757362,3.3757362,3.3757362,3.3757362,3.3757362,3.3757362,4.0374675,4.699199,5.3627434,6.0244746,6.688019,6.9744673,7.262728,7.549176,7.837437,8.125698,7.7866745,7.4494634,7.112252,6.775041,6.43783,7.063302,7.686961,8.312433,8.937905,9.563377,9.024928,8.488291,7.949841,7.413204,6.874754,6.0879283,5.2992897,4.512464,3.7256382,2.9369993,3.4627585,3.9867048,4.512464,5.038223,5.562169,7.0868707,8.611572,10.138086,11.662788,13.1874895,14.287958,15.386614,16.487082,17.58755,18.688019,17.449764,16.213324,14.975071,13.736817,12.500377,11.325577,10.150778,8.974165,7.799365,6.624565,7.3751316,8.125698,8.874452,9.625018,10.375585,11.650098,12.92461,14.200936,15.475449,16.749962,17.163317,17.57486,17.988214,18.399757,18.813112,18.11331,17.411694,16.71189,16.012085,15.312282,14.724882,14.137483,13.550082,12.962683,12.375282,11.874905,11.374527,10.874149,10.375585,9.875207,7.9625316,6.049856,4.137181,2.2245052,0.31182957,0.25018883,0.18673515,0.12509441,0.06164073,0.0,0.36259252,0.72518504,1.0877775,1.4503701,1.8129625,1.4503701,1.0877775,0.72518504,0.36259252,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.40066472,0.7995165,1.2001812,1.6008459,1.9996977,1.8256533,1.649796,1.4757515,1.2998942,1.1258497,1.4630609,1.8002719,2.137483,2.474694,2.811905,2.612479,2.4130533,2.2118144,2.0123885,1.8129625,1.4503701,1.0877775,0.72518504,0.36259252,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.3245203,0.5873999,0.85027945,1.1131591,1.3742256,2.5744069,3.774588,4.974769,6.1749506,7.3751316,6.9998484,6.624565,6.249282,5.8758116,5.5005283,5.186886,4.8750563,4.5632267,4.249584,3.9377546,4.612177,5.2865987,5.962834,6.637256,7.311678,6.412449,5.5132194,4.612177,3.7129474,2.811905,2.7502642,2.6868105,2.6251698,2.561716,2.5000753,4.2242026,5.9501433,7.6742706,9.400211,11.124338,8.899834,6.6753283,4.4508233,2.2245052,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.5493277,0.97537386,1.3996071,1.8256533,2.2498865,3.9631362,5.674573,7.3878226,9.099259,10.812509,11.825955,12.837588,13.849221,14.862667,15.8743,16.487082,17.099863,17.712645,18.325426,18.938208,17.25034,15.56247,13.874602,12.186734,10.500679,11.599335,12.699803,13.800271,14.90074,15.999394,20.4756,24.949991,29.424383,33.90059,38.374977,32.136574,25.899984,19.66158,13.424988,7.1883965,9.775495,12.362592,14.94969,17.536787,20.125698,19.400513,18.675327,17.950142,17.224958,16.499773,14.037769,11.575767,9.11195,6.6499467,4.1879435,4.1117992,4.0374675,3.9631362,3.8869917,3.8126602,3.6875658,3.5624714,3.437377,3.3122826,3.1871881,5.5367875,7.8882003,10.2378,12.5873995,14.936998,15.074784,15.212569,15.350354,15.488139,15.624111,12.699803,9.775495,6.849373,3.925064,1.0007553,6.5629244,12.125093,17.687263,23.249432,28.811602,23.062696,17.31198,11.563075,5.812358,0.06164073,5.0255322,9.987611,14.94969,19.911768,24.87566,19.899076,14.924308,9.949538,4.974769,0.0,0.0870222,0.17585737,0.26287958,0.34990177,0.43692398,0.34990177,0.26287958,0.17585737,0.0870222,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,3.6748753,7.224656,10.774437,14.324218,17.87581,14.311526,10.750868,7.1865835,3.6241121,0.06164073,2.2625773,4.461701,6.6626377,8.861761,11.062697,10.087324,9.11195,8.136576,7.1630154,6.187641,5.049101,3.9123733,2.7756457,1.6371052,0.50037766,2.3622901,4.2242026,6.0879283,7.949841,9.811753,10.924912,12.038072,13.149418,14.262577,15.375735,13.987006,12.60009,11.213174,9.824444,8.437528,6.9128265,5.388125,3.8616104,2.3369088,0.8122072,3.9504454,7.0868707,10.225109,13.361534,16.499773,16.762651,17.025532,17.288412,17.549479,17.812357,16.313038,14.811904,13.312584,11.813264,10.312131,9.200785,8.087626,6.9744673,5.863121,4.749962,7.250037,9.750113,12.250188,14.750263,17.25034,16.187943,15.125546,14.06315,13.000754,11.938358,14.336908,16.73727,19.137632,21.537996,23.938358,25.974316,28.012085,30.049854,32.087624,34.125393,32.54993,30.974466,29.400814,27.82535,26.249886,23.999998,21.750113,19.500225,17.25034,15.000452,16.537846,18.075237,19.612629,21.15002,22.687414,22.350203,22.01299,21.675781,21.336756,20.999546,21.12464,21.249735,21.374828,21.499924,21.625017,20.925215,20.22541,19.525606,18.825804,18.124187,17.774284,17.424383,17.074482,16.72458,16.374678,18.537542,20.700407,22.863272,25.024323,27.187187,25.24913,23.312885,21.374828,19.436771,17.500528,17.038223,16.574104,16.1118,15.649493,15.187187,14.975071,14.762955,14.5508375,14.336908,14.124791,18.087927,22.051064,26.012386,29.975523,33.936848,32.800117,31.66158,30.52485,29.388123,28.249582,25.486628,22.725487,19.96253,17.199575,14.436621,12.174044,9.911467,7.650702,5.388125,3.1255474,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.032633327,0.052575916,0.072518505,0.092461094,0.11240368,0.12328146,0.13234627,0.14322405,0.15228885,0.16316663,0.14322405,0.12328146,0.10333887,0.08339628,0.06164073,0.18673515,0.31182957,0.43692398,0.5620184,0.6871128,0.83940166,0.9916905,1.1457924,1.2980812,1.4503701,1.3343405,1.2201238,1.1059072,0.9898776,0.87566096,0.75781834,0.6399758,0.52213323,0.40429065,0.28826106,0.27194437,0.2574407,0.24293698,0.22662032,0.21211663,0.33177215,0.45324063,0.5728962,0.69255173,0.8122072,0.96268314,1.1131591,1.261822,1.4122978,1.5627737,1.551896,1.5428312,1.5319533,1.5228885,1.5120108,2.269829,3.0276475,3.785466,4.5432844,5.2992897,5.7053933,6.109684,6.5157876,6.9200783,7.324369,8.152893,8.979604,9.808127,10.634838,11.463363,11.650098,11.836833,12.025381,12.212116,12.400664,11.691795,10.98474,10.277685,9.570629,8.861761,9.771869,10.681975,11.592083,12.50219,13.412297,14.462003,15.511708,16.563227,17.612932,18.662638,20.207281,21.751925,23.298382,24.843027,26.38767,23.889408,21.392958,18.894695,16.398247,13.899984,12.476809,11.055446,9.63227,8.209095,6.787732,6.680767,6.5719895,6.4650245,6.35806,6.249282,7.0904965,7.9298983,8.7693,9.610515,10.449916,9.605076,8.760235,7.915395,7.0705543,6.2257137,5.3246713,4.4254417,3.5243993,2.6251698,1.7241274,1.5283275,1.3307146,1.1331016,0.9354887,0.73787576,1.260009,1.7821422,2.3042755,2.8282216,3.350355,3.5171473,3.6857529,3.8525455,4.019338,4.1879435,3.9522583,3.7183862,3.482701,3.247016,3.0131438,2.619731,2.228131,1.8347181,1.4431182,1.0497054,1.7241274,2.4003625,3.0747845,3.7492065,4.4254417,4.4127507,4.40006,4.3873696,4.3746786,4.361988,4.3873696,4.4127507,4.4381323,4.461701,4.4870825,5.243088,5.99728,6.7532854,7.507478,8.26167,8.127511,7.993352,7.85738,7.723221,7.5872483,7.3896356,7.192023,6.9944096,6.796797,6.599184,7.268167,7.935337,8.602508,9.269678,9.936848,9.590572,9.242483,8.894395,8.548119,8.200029,7.5799966,6.9599633,6.33993,5.719897,5.0998635,5.618371,6.1350656,6.6517596,7.170267,7.686961,8.9868555,10.28675,11.586644,12.888351,14.188245,14.880796,15.573349,16.2659,16.956638,17.64919,16.76084,15.870674,14.98051,14.090345,13.200181,12.322706,11.445232,10.567759,9.690285,8.812811,9.605076,10.397341,11.189605,11.98187,12.774135,14.117539,15.459132,16.802538,18.144129,19.487535,19.456715,19.427708,19.396887,19.36788,19.337059,18.655384,17.971897,17.290224,16.606737,15.925063,15.15818,14.389484,13.622601,12.855718,12.087022,11.740746,11.392657,11.044568,10.698292,10.3502035,8.7693,7.1902094,5.6093063,4.0302157,2.4493124,2.1229792,1.794833,1.4666867,1.1403534,0.8122072,0.9481794,1.0823387,1.2183108,1.35247,1.4866294,1.4830034,1.4775645,1.4721256,1.4666867,1.4630609,1.2382535,1.0116332,0.7868258,0.5620184,0.33721104,0.27013144,0.2030518,0.13415924,0.06707962,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.099712946,0.099712946,0.099712946,0.099712946,0.099712946,0.09064813,0.07977036,0.07070554,0.059827764,0.05076295,0.059827764,0.07070554,0.07977036,0.09064813,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.33177215,0.6653573,0.99712944,1.3307146,1.6624867,1.5120108,1.3633479,1.2128719,1.062396,0.9119202,1.2328146,1.551896,1.8727903,2.1918716,2.5127661,2.3532255,2.1918716,2.032331,1.8727903,1.7132497,1.3851035,1.0569572,0.7306239,0.40247768,0.07433146,0.19036107,0.3045777,0.42060733,0.53482395,0.6508536,1.0297627,1.4104849,1.789394,2.1701162,2.5508385,3.388427,4.2242026,5.0617914,5.89938,6.736969,6.506723,6.2782893,6.0480433,5.8177967,5.5875506,5.2032027,4.8170414,4.4326935,4.0483456,3.6621845,4.160749,4.6575007,5.1542525,5.6528172,6.149569,5.375434,4.599486,3.825351,3.049403,2.275268,2.220879,2.1646774,2.1102884,2.0558996,1.9996977,3.4192474,4.84061,6.26016,7.6797094,9.099259,7.5056653,5.910258,4.314851,2.7194438,1.1258497,1.3996071,1.6751775,1.9507477,2.2245052,2.5000753,2.6396735,2.7792716,2.9206827,3.0602808,3.199879,4.844236,6.490406,8.134763,9.780933,11.42529,12.15954,12.895603,13.629852,14.365915,15.100165,15.66581,16.229641,16.795286,17.359118,17.92476,16.64481,15.364858,14.084907,12.804955,11.525003,12.91192,14.300649,15.687565,17.074482,18.463211,22.283123,26.103035,29.922947,33.74286,37.56277,32.185524,26.808277,21.429218,16.051971,10.674724,12.456866,14.240821,16.022963,17.805105,19.587248,18.9654,18.341742,17.719896,17.09805,16.474392,13.947122,11.419851,8.892582,6.3653116,3.8380418,3.778214,3.7183862,3.6567454,3.5969179,3.53709,3.3702974,3.2016919,3.0348995,2.8681068,2.6995013,4.933071,7.1648283,9.398398,11.630155,13.861912,14.231756,14.601601,14.973258,15.343102,15.712947,13.017072,10.323009,7.6271334,4.933071,2.2371957,6.399758,10.56232,14.724882,18.887444,23.050007,18.867502,14.684997,10.502492,6.319988,2.137483,6.3671246,10.596766,14.828221,19.057863,23.287504,19.52742,15.767336,12.007251,8.247167,4.4870825,4.5450974,4.603112,4.6593137,4.7173285,4.7753434,4.610364,4.445384,4.2804046,4.115425,3.9504454,3.778214,3.6041696,3.4319382,3.2597067,3.0874753,5.9483304,8.807372,11.668227,14.527269,17.388124,14.703127,12.018129,9.333132,6.6481338,3.9631362,5.2032027,6.4432693,7.6833353,8.923402,10.161655,9.518054,8.872639,8.227224,7.5818095,6.9382076,6.017223,5.0980506,4.177066,3.2578938,2.3369088,3.8597972,5.382686,6.9055743,8.42665,9.949538,10.622148,11.294757,11.967366,12.639976,13.312584,12.123281,10.932164,9.742861,8.551744,7.362441,6.397945,5.431636,4.4671397,3.5026438,2.5381477,4.7771564,7.017978,9.256987,11.497808,13.736817,13.974316,14.211814,14.449312,14.68681,14.924308,13.727753,12.529385,11.332829,10.13446,8.937905,8.189152,7.4422116,6.695271,5.9483304,5.199577,7.723221,10.245051,12.766883,15.290526,17.812357,17.09805,16.38193,15.667623,14.953316,14.237195,16.233267,18.227526,20.221785,22.217857,24.212114,25.972502,27.73289,29.493275,31.251848,33.012238,31.387821,29.763407,28.137178,26.512764,24.88835,23.137028,21.38752,19.63801,17.888502,16.13718,17.384499,18.631817,19.879135,21.128265,22.375584,21.875206,21.374828,20.87445,20.375887,19.87551,19.9444,20.015106,20.085812,20.154705,20.22541,19.891825,19.560053,19.228281,18.894695,18.562923,18.394318,18.227526,18.060734,17.892128,17.725336,20.006042,22.284937,24.565643,26.844538,29.125244,26.447498,23.769753,21.092007,18.41426,15.738328,15.442815,15.147303,14.851789,14.558089,14.262577,14.262577,14.262577,14.262577,14.262577,14.262577,17.75978,21.258799,24.756004,28.251396,31.750414,30.85481,29.959208,29.065416,28.169813,27.27421,25.009819,22.745428,20.479225,18.214834,15.950445,14.132043,12.3154545,10.497053,8.680465,6.8620634,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.065266654,0.10515183,0.14503701,0.18492219,0.22480737,0.24474995,0.26469254,0.28463513,0.3045777,0.3245203,0.28463513,0.24474995,0.20486477,0.16497959,0.12509441,0.37528324,0.62547207,0.87566096,1.1258497,1.3742256,1.6806163,1.9851941,2.2897718,2.5943494,2.9007401,2.6704938,2.4402475,2.2100015,1.9797552,1.7495089,1.5156367,1.2799516,1.0442665,0.8103943,0.5747091,0.54570174,0.5148814,0.48587397,0.4550536,0.42423326,0.6653573,0.90466833,1.1457924,1.3851035,1.6244144,1.9253663,2.2245052,2.525457,2.8245957,3.1255474,3.105605,3.0856624,3.0657198,3.045777,3.0258346,3.9903307,4.954827,5.919323,6.885632,7.850128,8.247167,8.644206,9.043057,9.440096,9.837135,10.243238,10.64753,11.05182,11.457924,11.862214,11.900287,11.938358,11.974618,12.012691,12.050762,11.421664,10.794379,10.167094,9.539809,8.912524,9.795437,10.6783495,11.559449,12.442362,13.325275,14.05046,14.775645,15.50083,16.224201,16.949387,18.6155,20.279799,21.945911,23.610212,25.274511,22.718235,20.160145,17.602055,15.045776,12.487686,11.318325,10.147152,8.977791,7.806617,6.637256,6.622752,6.6082487,6.591932,6.5774283,6.5629244,7.192023,7.8229337,8.452031,9.082943,9.712041,9.059374,8.406708,7.755854,7.1031876,6.450521,5.638314,4.8242936,4.0120864,3.199879,2.3876717,2.1556125,1.9217403,1.6896812,1.4576219,1.2255627,1.6697385,2.1157274,2.5599031,3.005892,3.4500678,3.584227,3.720199,3.8543584,3.9903307,4.12449,4.0555973,3.9848917,3.9141862,3.8452935,3.774588,3.4029307,3.0294604,2.657803,2.2843328,1.9126755,2.474694,3.0367124,3.6005437,4.162562,4.7245803,4.8496747,4.974769,5.0998635,5.224958,5.3500524,5.4008155,5.4497657,5.5005283,5.5494785,5.600241,6.446895,7.2953615,8.1420145,8.990481,9.837135,9.280556,8.722163,8.165584,7.607191,7.0506115,6.9925966,6.9345818,6.87838,6.8203654,6.7623506,7.473032,8.1819,8.892582,9.603263,10.312131,10.154404,9.9966755,9.840761,9.683033,9.525306,9.072064,8.620637,8.167397,7.7141557,7.262728,7.7721705,8.281613,8.792869,9.302311,9.811753,10.88684,11.961927,13.037014,14.112101,15.187187,15.471823,15.758271,16.042906,16.327541,16.612177,16.0701,15.528025,14.984136,14.4420595,13.899984,13.319836,12.739688,12.15954,11.579392,10.999244,11.83502,12.670795,13.504758,14.340534,15.174497,16.584982,17.995466,19.404139,20.814623,22.22511,21.751925,21.280556,20.807371,20.334188,19.862818,19.19746,18.532103,17.866747,17.203201,16.537846,15.589665,14.643299,13.695119,12.74694,11.800573,11.6047735,11.410787,11.214987,11.019187,10.825199,9.577881,8.330563,7.083245,5.8341136,4.5867953,3.9957695,3.4029307,2.810092,2.2172532,1.6244144,1.5319533,1.4394923,1.3470312,1.2545701,1.162109,1.5156367,1.8673514,2.220879,2.572594,2.9243085,2.474694,2.0250793,1.5754645,1.1258497,0.6744221,0.5402629,0.40429065,0.27013144,0.13415924,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.07433146,0.07433146,0.07433146,0.07433146,0.07433146,0.06707962,0.059827764,0.052575916,0.045324065,0.038072214,0.045324065,0.052575916,0.059827764,0.06707962,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.26469254,0.5293851,0.79589057,1.0605831,1.3252757,1.2001812,1.0750868,0.9499924,0.824898,0.69980353,1.0025684,1.305333,1.6080978,1.9108626,2.2118144,2.0921588,1.9725033,1.8528478,1.7331922,1.6117238,1.3198367,1.0279498,0.73424983,0.44236287,0.15047589,0.3680314,0.5855869,0.8031424,1.020698,1.2382535,1.7350051,2.231757,2.7303216,3.2270734,3.7256382,4.2006345,4.6756306,5.1506267,5.6256227,6.1006193,6.01541,5.9302006,5.844991,5.7597823,5.674573,5.217706,4.76084,4.3021603,3.8452935,3.386614,3.7075086,4.02659,4.347484,4.668379,4.98746,4.3366065,3.6875658,3.0367124,2.3876717,1.7368182,1.6896812,1.6425442,1.5954071,1.54827,1.49932,2.6142921,3.729264,4.844236,5.959208,7.07418,6.109684,5.145188,4.1806917,3.2143826,2.2498865,2.7756457,3.299592,3.825351,4.349297,4.8750563,4.7300196,4.5849824,4.439945,4.2949085,4.1498713,5.727149,7.304426,8.881703,10.460794,12.038072,12.494938,12.951805,13.410484,13.867351,14.324218,14.842725,15.359419,15.877926,16.39462,16.913128,16.03928,15.167245,14.29521,13.423175,12.549327,14.224504,15.899682,17.57486,19.250036,20.925215,24.090647,27.254267,30.419699,33.585133,36.750565,32.232662,27.71476,23.196856,18.680767,14.162864,15.140051,16.117237,17.094423,18.071611,19.050611,18.53029,18.00997,17.48965,16.96933,16.450823,13.856473,11.26575,8.673213,6.0806766,3.48814,3.442816,3.397492,3.3521678,3.3068438,3.2633326,3.053029,2.8427253,2.6324217,2.422118,2.2118144,4.327542,6.4432693,8.557183,10.672911,12.786825,13.390542,13.992445,14.594349,15.198066,15.799969,13.33434,10.870523,8.404895,5.9392653,3.4754493,6.2384043,8.999546,11.762501,14.525456,17.288412,14.672306,12.058014,9.441909,6.827617,4.213325,7.71053,11.207735,14.70494,18.202145,21.699348,19.15395,16.610363,14.064963,11.519565,8.974165,9.003172,9.030367,9.057561,9.084756,9.11195,8.870826,8.627889,8.384952,8.1420145,7.900891,7.5292335,7.159389,6.789545,6.4197006,6.049856,8.219973,10.390089,12.5602045,14.730321,16.900436,15.092914,13.28539,11.477866,9.670342,7.8628187,8.1420145,8.423024,8.70222,8.98323,9.262425,8.94697,8.6333275,8.317872,8.002417,7.686961,6.985345,6.281915,5.580299,4.876869,4.175253,5.3573046,6.539356,7.723221,8.9052725,10.087324,10.319383,10.553255,10.785315,11.017374,11.249433,10.257742,9.264238,8.272549,7.2808576,6.2873545,5.883064,5.47696,5.0726695,4.668379,4.262275,5.6056805,6.947273,8.290678,9.63227,10.975676,11.187792,11.399909,11.612025,11.8241415,12.038072,11.142468,10.246864,9.353074,8.457471,7.5618668,7.179332,6.796797,6.414262,6.0317264,5.6491914,8.194591,10.73999,13.28539,15.828977,18.374376,18.008158,17.640125,17.272095,16.905876,16.537846,18.127813,19.717781,21.307749,22.897717,24.487686,25.97069,27.45188,28.934883,30.417887,31.90089,30.225712,28.550535,26.875357,25.20018,23.525002,22.274057,21.024927,19.775795,18.52485,17.27572,18.232965,19.190208,20.147453,21.104698,22.061941,21.40021,20.736666,20.074934,19.413204,18.749659,18.764162,18.78048,18.794983,18.809486,18.825804,18.86025,18.894695,18.929142,18.9654,18.999847,19.01435,19.030668,19.045172,19.059675,19.074179,21.472729,23.869465,26.268015,28.664751,31.063301,27.644053,24.22662,20.809185,17.393562,13.974316,13.847408,13.720501,13.591781,13.464873,13.337966,13.550082,13.762199,13.974316,14.188245,14.400362,17.433449,20.464722,23.497808,26.529081,29.562168,28.909502,28.256834,27.604168,26.953314,26.300648,24.53301,22.765371,20.997732,19.230095,17.462456,16.090042,14.71763,13.345218,11.972805,10.600392,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.09789998,0.15772775,0.21755551,0.27738327,0.33721104,0.3680314,0.39703882,0.42785916,0.45686656,0.48768693,0.42785916,0.3680314,0.30820364,0.24837588,0.18673515,0.5620184,0.93730164,1.3125849,1.6878681,2.0631514,2.520018,2.9768846,3.435564,3.8924308,4.349297,4.004834,3.6603715,3.3140955,2.9696326,2.6251698,2.2716422,1.9199274,1.5682126,1.214685,0.8629702,0.81764615,0.77232206,0.726998,0.68167394,0.63816285,0.99712944,1.357909,1.7168756,2.077655,2.4366217,2.8880494,3.3376641,3.787279,4.2368937,4.688321,4.6575007,4.6266804,4.597673,4.5668526,4.537845,5.710832,6.882006,8.054993,9.22798,10.399154,10.790753,11.18054,11.570327,11.9601145,12.349901,12.331772,12.3154545,12.297325,12.279196,12.262879,12.1504755,12.038072,11.925668,11.813264,11.700861,11.153346,10.605831,10.058316,9.510801,8.963287,9.817192,10.672911,11.526816,12.382534,13.238253,13.637105,14.037769,14.436621,14.837286,15.23795,17.021906,18.807674,20.593443,22.377398,24.163166,21.545248,18.92733,16.309412,13.693306,11.075388,10.15803,9.24067,8.323311,7.404139,6.48678,6.5647373,6.642695,6.720652,6.796797,6.874754,7.2953615,7.7141557,8.134763,8.55537,8.974165,8.515485,8.054993,7.5945,7.135821,6.6753283,5.9501433,5.224958,4.499773,3.774588,3.049403,2.7828975,2.514579,2.2480736,1.9797552,1.7132497,2.079468,2.4474995,2.8155308,3.1817493,3.5497808,3.6531196,3.7546456,3.8579843,3.9595103,4.062849,4.157123,4.25321,4.347484,4.441758,4.537845,4.1843176,3.832603,3.4808881,3.1273603,2.7756457,3.2252605,3.6748753,4.12449,4.574105,5.0255322,5.2865987,5.5494785,5.812358,6.0752378,6.338117,6.412449,6.48678,6.5629244,6.637256,6.7134004,7.652515,8.59163,9.5325575,10.471672,11.4126,10.431787,9.452786,8.471974,7.4929743,6.5121617,6.5955577,6.677141,6.7605376,6.8421206,6.925517,7.6778965,8.430276,9.182655,9.935035,10.687414,10.720048,10.752681,10.785315,10.817947,10.850581,10.564133,10.279498,9.994863,9.710228,9.425592,9.927783,10.429974,10.932164,11.434355,11.938358,12.786825,13.637105,14.487384,15.337664,16.187943,16.064661,15.9431925,15.819912,15.6966305,15.575162,15.379361,15.185374,14.989574,14.795588,14.599788,14.316965,14.034143,13.753134,13.470312,13.1874895,14.064963,14.942437,15.819912,16.697386,17.57486,19.052423,20.529987,22.007553,23.485117,24.962683,24.047136,23.133402,22.217857,21.30231,20.386765,19.739536,19.092308,18.445082,17.797853,17.150625,16.022963,14.895301,13.767638,12.639976,11.512312,11.470614,11.427103,11.385405,11.341894,11.300196,10.384649,9.470917,8.55537,7.6398244,6.7242785,5.866747,5.009216,4.1516843,3.294153,2.4366217,2.1175404,1.7966459,1.4775645,1.1566701,0.8375887,1.54827,2.2571385,2.9678197,3.6766882,4.3873696,3.7129474,3.0367124,2.3622901,1.6878681,1.0116332,0.8103943,0.6073425,0.40429065,0.2030518,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.045324065,0.03988518,0.034446288,0.030820364,0.025381476,0.030820364,0.034446288,0.03988518,0.045324065,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.19761293,0.39522585,0.59283876,0.7904517,0.9880646,0.8883517,0.7868258,0.6871128,0.5873999,0.48768693,0.77232206,1.0569572,1.3434052,1.6280404,1.9126755,1.8329052,1.7531348,1.6733645,1.5917811,1.5120108,1.2545701,0.99712944,0.73968875,0.48224804,0.22480737,0.54570174,0.86478317,1.1856775,1.504759,1.8256533,2.4402475,3.054842,3.6694362,4.2858434,4.900438,5.0128417,5.125245,5.237649,5.3500524,5.462456,5.522284,5.582112,5.6419396,5.7017674,5.7615952,5.23221,4.702825,4.171627,3.6422417,3.1128569,3.254268,3.397492,3.540716,3.682127,3.825351,3.299592,2.7756457,2.2498865,1.7241274,1.2001812,1.1602961,1.1204109,1.0805258,1.0406405,1.0007553,1.8093367,2.619731,3.4301252,4.2405195,5.049101,4.7155156,4.3801174,4.0447197,3.7093215,3.3757362,4.1498713,4.9258194,5.6999545,6.4759026,7.250037,6.8203654,6.390693,5.959208,5.529536,5.0998635,6.6100616,8.120259,9.630457,11.1406555,12.650853,12.830337,13.009819,13.189302,13.370599,13.550082,14.01964,14.489197,14.960567,15.430124,15.899682,15.435563,14.969632,14.505513,14.039582,13.575464,15.537089,17.500528,19.462152,21.425592,23.387217,25.89817,28.40731,30.918264,33.427402,35.93836,32.2798,28.623053,24.964495,21.307749,17.64919,17.823235,17.995466,18.167698,18.33993,18.512161,18.095179,17.678198,17.259403,16.842422,16.425442,13.767638,11.109835,8.452031,5.7942286,3.1382382,3.1074178,3.0765975,3.04759,3.0167696,2.9877625,2.7357605,2.4819458,2.229944,1.9779422,1.7241274,3.7220123,5.719897,7.7177815,9.715667,11.711739,12.547514,13.383289,14.217253,15.053028,15.8869915,13.651608,11.418038,9.182655,6.947273,4.7118897,6.0752378,7.4367723,8.80012,10.161655,11.525003,10.477111,9.429218,8.383139,7.3352466,6.2873545,9.052122,11.81689,14.583471,17.34824,20.113007,18.782291,17.45339,16.122677,14.791962,13.46306,13.4594345,13.457622,13.455809,13.452183,13.45037,13.129475,12.810393,12.489499,12.170418,11.849524,11.282066,10.714609,10.147152,9.579695,9.012237,10.493427,11.972805,13.452183,14.9333725,16.41275,15.4827,14.55265,13.622601,12.692551,11.762501,11.082641,10.40278,9.7229185,9.043057,8.363196,8.3777,8.392203,8.406708,8.423024,8.437528,7.951654,7.4675927,6.981719,6.497658,6.011784,6.8548117,7.6978393,8.540867,9.382081,10.225109,10.016619,9.80994,9.603263,9.394773,9.188094,8.392203,7.5981264,6.8022356,6.008158,5.2122674,5.368182,5.522284,5.678199,5.8323007,5.9882154,6.432391,6.87838,7.322556,7.7667317,8.212721,8.399456,8.588004,8.774739,8.963287,9.1500225,8.557183,7.9643445,7.3733187,6.78048,6.187641,6.169512,6.153195,6.1350656,6.1169357,6.1006193,8.667774,11.234929,13.802084,16.36924,18.938208,18.918264,18.898321,18.87838,18.856625,18.836681,20.022358,21.208036,22.391901,23.577578,24.763256,25.967064,27.172684,28.378304,29.582111,30.787731,29.06179,27.337664,25.611723,23.887594,22.161655,21.4129,20.662334,19.911768,19.163015,18.412449,19.079618,19.746788,20.415771,21.082941,21.750113,20.925215,20.100317,19.275417,18.45052,17.625622,17.585737,17.545853,17.504154,17.464268,17.424383,17.82686,18.22934,18.631817,19.034294,19.436771,19.634384,19.831997,20.02961,20.227224,20.424837,22.939415,25.455807,27.970387,30.484966,32.999546,28.842422,24.685299,20.528175,16.371052,12.212116,12.252001,12.291886,12.331772,12.371656,12.413355,12.837588,13.261822,13.687867,14.112101,14.538147,17.105303,19.672457,22.239613,24.806767,27.375734,26.964193,26.554462,26.144733,25.735004,25.325274,24.054388,22.785315,21.514427,20.245354,18.974466,18.048042,17.119806,16.193382,15.265145,14.336908,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.13053331,0.21030366,0.29007402,0.36984438,0.44961473,0.4894999,0.5293851,0.56927025,0.6091554,0.6508536,0.56927025,0.4894999,0.40972954,0.32995918,0.25018883,0.7505665,1.2491312,1.7495089,2.2498865,2.7502642,3.3594196,3.9703882,4.5795436,5.1905117,5.7996674,5.3391747,4.880495,4.420003,3.9595103,3.5008307,3.0294604,2.5599031,2.0903459,1.6207886,1.1494182,1.0895905,1.0297627,0.969935,0.9101072,0.85027945,1.3307146,1.8093367,2.2897718,2.770207,3.2506418,3.8507326,4.4508233,5.050914,5.6491914,6.249282,6.209397,6.169512,6.1296263,6.089741,6.049856,7.4295206,8.809185,10.190662,11.570327,12.949992,13.332527,13.715062,14.097597,14.480132,14.862667,14.422117,13.98338,13.54283,13.102281,12.661731,12.400664,12.137785,11.874905,11.612025,11.349146,10.883214,10.41547,9.947725,9.479981,9.012237,9.840761,10.667472,11.494183,12.322706,13.149418,13.225562,13.299893,13.374225,13.45037,13.524701,15.430124,17.335548,19.239159,21.144583,23.050007,20.372261,17.694515,15.016769,12.340837,9.663091,8.997733,8.3323765,7.667019,7.0016613,6.338117,6.506723,6.677141,6.8475595,7.017978,7.1883965,7.3968873,7.607191,7.817495,8.027799,8.238102,7.9697833,7.703278,7.4349594,7.166641,6.9001355,6.261973,5.6256227,4.98746,4.349297,3.7129474,3.4101827,3.1074178,2.8046532,2.5018883,2.1991236,2.4891977,2.7792716,3.0693457,3.3594196,3.6494937,3.720199,3.7890918,3.8597972,3.930503,3.9993954,4.2604623,4.519716,4.780782,5.040036,5.2992897,4.9675174,4.6357455,4.3021603,3.9703882,3.636803,3.975827,4.313038,4.650249,4.98746,5.3246713,5.7253356,6.1241875,6.5248523,6.925517,7.324369,7.4258947,7.5256076,7.6253204,7.7250338,7.8247466,8.858135,9.88971,10.9230995,11.954676,12.988064,11.584831,10.183411,8.780178,7.3769445,5.975525,6.1967063,6.4197006,6.642695,6.8656893,7.0868707,7.8827615,8.676839,9.47273,10.266808,11.062697,11.285692,11.506873,11.729868,11.952863,12.175857,12.058014,11.940171,11.822329,11.704487,11.586644,12.081583,12.578335,13.073273,13.568212,14.06315,14.68681,15.312282,15.937754,16.563227,17.186886,16.6575,16.128115,15.596917,15.067532,14.538147,14.690435,14.842725,14.995013,15.147303,15.299591,15.314095,15.330412,15.344915,15.359419,15.375735,16.294909,17.214079,18.135065,19.054237,19.975222,21.519865,23.06451,24.609154,26.155611,27.700254,26.342346,24.984438,23.628342,22.270432,20.912523,20.281612,19.652514,19.021603,18.392506,17.761595,16.454449,15.147303,13.840157,12.5330105,11.225864,11.334642,11.445232,11.555823,11.664601,11.775192,11.193231,10.609457,10.027496,9.445535,8.861761,7.7395372,6.6173134,5.4950895,4.3728657,3.2506418,2.7031271,2.1556125,1.6080978,1.0605831,0.51306844,1.5790904,2.6469254,3.7147603,4.782595,5.8504305,4.949388,4.0501585,3.149116,2.2498865,1.3506571,1.0805258,0.8103943,0.5402629,0.27013144,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.02175555,0.01994259,0.018129626,0.014503701,0.012690738,0.014503701,0.018129626,0.01994259,0.02175555,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13053331,0.25925365,0.38978696,0.52032024,0.6508536,0.5747091,0.50037766,0.42423326,0.34990177,0.2755703,0.5420758,0.8103943,1.0768998,1.3452182,1.6117238,1.5718386,1.5319533,1.4920682,1.452183,1.4122978,1.1893034,0.968122,0.7451276,0.52213323,0.2991388,0.72337204,1.1457924,1.5682126,1.9906329,2.4130533,3.1454902,3.877927,4.610364,5.3428006,6.0752378,5.825049,5.57486,5.3246713,5.0744824,4.8242936,5.029158,5.235836,5.4407005,5.6455655,5.8504305,5.2467136,4.64481,4.0429068,3.43919,2.8372865,2.8028402,2.7683938,2.7321346,2.6976883,2.663242,2.2625773,1.8619126,1.4630609,1.062396,0.66173136,0.629098,0.5982776,0.5656443,0.533011,0.50037766,1.0043813,1.5101979,2.0142014,2.520018,3.0258346,3.3195345,3.6150475,3.9105604,4.2042603,4.499773,5.52591,6.550234,7.574558,8.600695,9.625018,8.910711,8.194591,7.4802837,6.7641635,6.049856,7.4929743,8.934279,10.377398,11.820516,13.261822,13.165734,13.067834,12.969934,12.872034,12.774135,13.198368,13.620788,14.043208,14.465629,14.888049,14.830034,14.772019,14.715817,14.657803,14.599788,16.849674,19.099562,21.349447,23.599335,25.84922,27.705694,29.560354,31.415016,33.269676,35.124336,32.326935,29.529535,26.732134,23.934732,21.137331,20.504606,19.871883,19.239159,18.608248,17.975525,17.660069,17.344612,17.029158,16.715515,16.400059,13.67699,10.955733,8.232663,5.5095935,2.7883365,2.7720199,2.7575161,2.7430124,2.7266958,2.712192,2.4166791,2.1229792,1.8274662,1.5319533,1.2382535,3.1182957,4.9983377,6.87838,8.758422,10.636651,11.704487,12.772322,13.840157,14.907991,15.975826,13.97069,11.965553,9.960417,7.95528,5.9501433,5.9120708,5.8758116,5.8377395,5.7996674,5.763408,6.281915,6.8022356,7.322556,7.842876,8.363196,10.395528,12.427858,14.46019,16.492521,18.52485,18.410635,18.294605,18.18039,18.06436,17.950142,17.91751,17.884876,17.852243,17.819609,17.786976,17.389936,16.992899,16.59586,16.197008,15.799969,15.034899,14.269829,13.504758,12.739688,11.974618,12.76507,13.555521,14.34416,15.134612,15.925063,15.872487,15.819912,15.767336,15.71476,15.662184,14.023266,12.382534,10.741803,9.102885,7.462154,7.8084297,8.152893,8.497355,8.841819,9.188094,8.919776,8.653271,8.384952,8.116633,7.850128,8.352319,8.854509,9.3567,9.860703,10.362894,9.715667,9.066626,8.419398,7.7721705,7.124943,6.526665,5.9302006,5.331923,4.7354584,4.137181,4.853301,5.567608,6.281915,6.9980354,7.7123427,7.2591023,6.8076744,6.354434,5.903006,5.4497657,5.612932,5.774286,5.9374523,6.1006193,6.261973,5.9718986,5.6818247,5.391751,5.101677,4.8116026,5.1596913,5.5077806,5.8558693,6.202145,6.550234,9.140957,11.729868,14.320591,16.909502,19.500225,19.828371,20.154705,20.482851,20.809185,21.137331,21.916904,22.698292,23.477865,24.257439,25.037014,25.96525,26.891674,27.81991,28.748148,29.674572,27.899681,26.12479,24.349901,22.57501,20.80012,20.54993,20.299742,20.049553,19.799364,19.549175,19.928085,20.305182,20.682278,21.059374,21.438282,20.450218,19.462152,18.474089,17.487837,16.499773,16.405499,16.309412,16.215137,16.120863,16.024776,16.795286,17.565794,18.33449,19.105,19.87551,20.254417,20.63514,21.015862,21.394772,21.775494,24.407915,27.040337,29.672758,32.30518,34.937603,30.038977,25.142164,20.245354,15.348541,10.449916,10.658407,10.865085,11.071762,11.280253,11.486931,12.125093,12.763257,13.399607,14.037769,14.674119,16.777155,18.880192,20.983229,23.084452,25.187489,25.020697,24.85209,24.685299,24.516693,24.349901,23.577578,22.805256,22.032934,21.260612,20.48829,20.004229,19.52198,19.039734,18.557486,18.075237,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.16316663,0.26287958,0.36259252,0.46230546,0.5620184,0.61278135,0.66173136,0.7124943,0.76325727,0.8122072,0.7124943,0.61278135,0.51306844,0.41335547,0.31182957,0.93730164,1.5627737,2.1882458,2.811905,3.437377,4.2006345,4.9620786,5.7253356,6.48678,7.250037,6.6753283,6.1006193,5.524097,4.949388,4.3746786,3.787279,3.199879,2.612479,2.0250793,1.4376793,1.3633479,1.2872034,1.2128719,1.1367276,1.062396,1.6624867,2.2625773,2.8626678,3.4627585,4.062849,4.8116026,5.562169,6.3127356,7.063302,7.8120556,7.763106,7.7123427,7.663393,7.61263,7.5618668,9.1500225,10.738177,12.32452,13.912675,15.50083,15.8743,16.249584,16.624866,17.00015,17.375433,16.512463,15.649493,14.788336,13.925365,13.062395,12.650853,12.237497,11.8241415,11.4126,10.999244,10.613083,10.225109,9.837135,9.449161,9.063,9.862516,10.662033,11.463363,12.262879,13.062395,12.812206,12.562017,12.311829,12.06164,11.813264,13.838344,15.861609,17.886688,19.911768,21.936848,19.199274,16.4617,13.724127,10.986553,8.2507925,7.837437,7.4258947,7.0125394,6.599184,6.187641,6.450521,6.7115874,6.9744673,7.2373466,7.500226,7.500226,7.500226,7.500226,7.500226,7.500226,7.4258947,7.3497505,7.2754188,7.1992745,7.124943,6.5756154,6.0244746,5.475147,4.9258194,4.3746786,4.0374675,3.7002566,3.3630457,3.0258346,2.6868105,2.9007401,3.1128569,3.3249733,3.53709,3.7492065,3.787279,3.825351,3.8616104,3.8996825,3.9377546,4.361988,4.788034,5.2122674,5.638314,6.0625467,5.750717,5.4370747,5.125245,4.8116026,4.499773,4.7245803,4.949388,5.1741953,5.4008155,5.6256227,6.16226,6.70071,7.2373466,7.7757964,8.312433,8.437528,8.562622,8.6877165,8.812811,8.937905,10.061942,11.187792,12.311829,13.437678,14.561715,12.737875,10.912222,9.086569,7.262728,5.4370747,5.7996674,6.16226,6.5248523,6.887445,7.250037,8.087626,8.925215,9.762803,10.600392,11.437981,11.849524,12.262879,12.674421,13.087777,13.499319,13.550082,13.600845,13.649796,13.700559,13.749508,14.237195,14.724882,15.212569,15.700256,16.187943,16.586794,16.98746,17.388124,17.786976,18.187641,17.25034,16.313038,15.375735,14.436621,13.499319,13.999697,14.500074,15.000452,15.50083,15.999394,16.313038,16.624866,16.936697,17.25034,17.562168,18.52485,19.487535,20.450218,21.4129,22.375584,23.987309,25.600845,27.212568,28.824291,30.437828,28.637556,26.837286,25.037014,23.236742,21.438282,20.8255,20.212719,19.59994,18.987158,18.374376,16.887747,15.399304,13.912675,12.4242325,10.937603,11.200482,11.463363,11.724429,11.9873085,12.250188,11.999999,11.74981,11.499621,11.249433,10.999244,9.612328,8.225411,6.836682,5.4497657,4.062849,3.2869012,2.5127661,1.7368182,0.96268314,0.18673515,1.6117238,3.0367124,4.461701,5.8866897,7.311678,6.187641,5.0617914,3.9377546,2.811905,1.6878681,1.3506571,1.0116332,0.6744221,0.33721104,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06164073,0.12509441,0.18673515,0.25018883,0.31182957,0.26287958,0.21211663,0.16316663,0.11240368,0.06164073,0.31182957,0.5620184,0.8122072,1.062396,1.3125849,1.3125849,1.3125849,1.3125849,1.3125849,1.3125849,1.1258497,0.93730164,0.7505665,0.5620184,0.37528324,0.89922947,1.4249886,1.9507477,2.474694,3.000453,3.8507326,4.699199,5.5494785,6.399758,7.250037,6.637256,6.0244746,5.411693,4.800725,4.1879435,4.537845,4.8877473,5.237649,5.5875506,5.9374523,5.2630305,4.5867953,3.9123733,3.2379513,2.561716,2.3495996,2.137483,1.9253663,1.7132497,1.49932,1.2255627,0.9499924,0.6744221,0.40066472,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.19942589,0.40066472,0.6000906,0.7995165,1.0007553,1.9253663,2.8499773,3.774588,4.699199,5.6256227,6.9001355,8.174648,9.449161,10.725487,11.999999,10.999244,10.000301,8.999546,8.000604,6.9998484,8.375887,9.750113,11.124338,12.500377,13.874602,13.499319,13.125849,12.750566,12.375282,11.999999,12.375282,12.750566,13.125849,13.499319,13.874602,14.224504,14.574407,14.924308,15.27421,15.624111,18.16226,20.700407,23.236742,25.774889,28.313036,29.513218,30.711586,31.911768,33.11195,34.31213,32.374073,30.437828,28.499771,26.561714,24.625471,23.187792,21.750113,20.312433,18.874754,17.437075,17.224958,17.01284,16.800724,16.586794,16.374678,13.588155,10.799818,8.013294,5.224958,2.4366217,2.4366217,2.4366217,2.4366217,2.4366217,2.4366217,2.0994108,1.7621996,1.4249886,1.0877775,0.7505665,2.5127661,4.274966,6.037165,7.799365,9.563377,10.863272,12.163166,13.46306,14.762955,16.062849,14.287958,12.513068,10.738177,8.963287,7.1883965,5.750717,4.313038,2.8753586,1.4376793,0.0,2.088533,4.175253,6.261973,8.350506,10.437225,11.73712,13.037014,14.336908,15.636803,16.936697,18.037165,19.137632,20.238102,21.336756,22.437225,22.375584,22.31213,22.25049,22.187037,22.125395,21.650398,21.175404,20.700407,20.22541,19.750414,18.787731,17.825048,16.862366,15.899682,14.936998,15.036712,15.138238,15.23795,15.337664,15.437376,16.262274,17.087172,17.912071,18.736969,19.561867,16.962078,14.362289,11.762501,9.162713,6.5629244,7.2373466,7.911769,8.588004,9.262425,9.936848,9.8878975,9.837135,9.788185,9.737422,9.686659,9.849826,10.012992,10.174346,10.337513,10.500679,9.412902,8.325124,7.2373466,6.149569,5.0617914,4.6629395,4.262275,3.8616104,3.4627585,3.0620937,4.3384194,5.612932,6.887445,8.161958,9.438283,8.087626,6.736969,5.388125,4.0374675,2.6868105,2.8245957,2.962381,3.100166,3.2379513,3.3757362,3.386614,3.3993049,3.4119956,3.4246864,3.437377,4.1498713,4.8623657,5.57486,6.2873545,6.9998484,9.612328,12.224807,14.837286,17.449764,20.062244,20.736666,21.4129,22.087322,22.761745,23.43798,23.813263,24.186733,24.562017,24.9373,25.312584,25.963438,26.612478,27.26333,27.912373,28.563225,26.737572,24.911919,23.088078,21.262424,19.436771,19.68696,19.93715,20.187338,20.437527,20.687716,20.774738,20.861761,20.950596,21.037619,21.12464,19.975222,18.82399,17.674572,16.525154,15.375735,15.22526,15.074784,14.924308,14.775645,14.625169,15.761897,16.900436,18.037165,19.175705,20.312433,20.87445,21.438282,22.000301,22.562319,23.124338,25.874601,28.624866,31.37513,34.125393,36.87566,31.237345,25.599031,19.96253,14.326031,8.6877165,9.063,9.438283,9.811753,10.1870365,10.56232,11.4126,12.262879,13.113158,13.961625,14.811904,16.450823,18.087927,19.725033,21.362139,22.999243,23.075388,23.14972,23.225864,23.300196,23.374527,23.100769,22.8252,22.54963,22.275871,22.000301,21.962229,21.924156,21.887897,21.849825,21.811752,0.05076295,0.047137026,0.045324065,0.04169814,0.03988518,0.038072214,0.19217403,0.3480888,0.50219065,0.65810543,0.8122072,0.85027945,0.8883517,0.9246109,0.96268314,1.0007553,0.9318628,0.86478317,0.79770356,0.7306239,0.66173136,0.59283876,0.52213323,0.45324063,0.3825351,0.31182957,1.1022812,1.892733,2.6831846,3.4718235,4.262275,4.7572136,5.2521524,5.7470913,6.24203,6.736969,6.2728505,5.806919,5.3428006,4.876869,4.4127507,4.102734,3.7927177,3.482701,3.1726844,2.8626678,3.6531196,4.441758,5.23221,6.0226617,6.813113,6.8403077,6.867502,6.8946967,6.921891,6.9508986,7.12313,7.2953615,7.4675927,7.6398244,7.8120556,7.764919,7.7177815,7.6706448,7.6216946,7.574558,8.767487,9.960417,11.153346,12.344462,13.537392,13.807523,14.077655,14.347786,14.617917,14.888049,14.342347,13.796645,13.252756,12.707055,12.163166,12.067079,11.972805,11.876718,11.782444,11.6881695,11.465176,11.242181,11.019187,10.798005,10.57501,11.245807,11.91479,12.585587,13.254569,13.925365,13.318023,12.710681,12.103338,11.494183,10.88684,12.507628,14.126604,15.747393,17.368181,18.987158,16.751774,14.518205,12.282822,10.047439,7.8120556,7.5854354,7.3570023,7.130382,6.9019485,6.6753283,6.8602505,7.0451727,7.230095,7.415017,7.5999393,7.667019,7.7340984,7.802991,7.8700705,7.93715,7.9715962,8.007855,8.042302,8.076748,8.113008,8.107569,8.10213,8.096691,8.093065,8.087626,7.5274205,6.967215,6.4070096,5.846804,5.2884116,5.368182,5.4479527,5.527723,5.6074934,5.6872635,5.6655083,5.6419396,5.620184,5.5966153,5.57486,5.8522434,6.1296263,6.4070096,6.684393,6.9617763,6.495845,6.0281005,5.560356,5.092612,4.6248674,4.7554007,4.8841214,5.0146546,5.145188,5.275721,6.153195,7.0306687,7.9081426,8.785617,9.663091,9.605076,9.547061,9.490859,9.432844,9.374829,10.2378,11.10077,11.961927,12.824898,13.687867,12.186734,10.687414,9.188094,7.686961,6.187641,6.510349,6.833056,7.155763,7.476658,7.799365,8.484665,9.169965,9.855265,10.540565,11.225864,11.564888,11.9057255,12.244749,12.585587,12.92461,13.174799,13.424988,13.675177,13.925365,14.175554,14.364102,14.554463,14.744824,14.935185,15.125546,15.5878525,16.050158,16.512463,16.97477,17.437075,17.0491,16.66294,16.274965,15.8869915,15.50083,15.738328,15.975826,16.213324,16.450823,16.68832,16.875055,17.06179,17.25034,17.437075,17.625622,18.202145,18.78048,19.357002,19.935337,20.511858,22.014805,23.51775,25.020697,26.52183,28.024776,26.639671,25.254568,23.869465,22.484362,21.099258,20.404894,19.71053,19.01435,18.319986,17.625622,16.458075,15.290526,14.122978,12.955431,11.787883,11.934732,12.083396,12.230246,12.377095,12.525759,11.925668,11.325577,10.725487,10.125396,9.525306,8.482852,7.440398,6.397945,5.3554916,4.313038,3.917812,3.5225863,3.1273603,2.7321346,2.3369088,3.0874753,3.8380418,4.5867953,5.337362,6.0879283,5.139749,4.1933823,3.245203,2.2970235,1.3506571,1.0805258,0.8103943,0.5402629,0.27013144,0.0,0.034446288,0.07070554,0.10515183,0.13959812,0.17585737,0.13959812,0.10515183,0.07070554,0.034446288,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.06707962,0.072518505,0.07795739,0.08339628,0.0870222,0.07070554,0.052575916,0.034446288,0.018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.13959812,0.26831847,0.39522585,0.52213323,0.6508536,0.5293851,0.40972954,0.29007402,0.17041849,0.05076295,0.2520018,0.4550536,0.65810543,0.85934424,1.062396,1.0732739,1.0823387,1.0932164,1.1022812,1.1131591,0.9898776,0.8684091,0.7451276,0.62184614,0.50037766,1.0551442,1.6099107,2.1646774,2.7194438,3.2742105,3.9069343,4.539658,5.1723824,5.805106,6.43783,6.0679855,5.6981416,5.328297,4.95664,4.5867953,4.9167547,5.2467136,5.576673,5.906632,6.2384043,5.47696,4.7173285,3.9576974,3.198066,2.4366217,2.3876717,2.3369088,2.2879589,2.2371957,2.1882458,1.7694515,1.35247,0.9354887,0.5166943,0.099712946,0.0870222,0.07433146,0.06164073,0.05076295,0.038072214,0.19217403,0.3480888,0.50219065,0.65810543,0.8122072,1.6534219,2.4928236,3.3322253,4.171627,5.0128417,6.0480433,7.083245,8.116633,9.151835,10.1870365,9.3150015,8.442966,7.569119,6.697084,5.825049,7.037921,8.2507925,9.461852,10.674724,11.887595,12.007251,12.126906,12.248375,12.368031,12.487686,12.687112,12.888351,13.087777,13.287203,13.486629,13.595407,13.702372,13.809336,13.918114,14.025079,16.50521,18.985344,21.465477,23.94561,26.425743,26.936998,27.450066,27.963135,28.47439,28.98746,27.694817,26.402174,25.109531,23.816889,22.524246,20.963285,19.400513,17.837738,16.274965,14.712192,14.558089,14.402175,14.248073,14.092158,13.938056,11.8241415,9.712041,7.5999393,5.487838,3.3757362,3.7582715,4.1408067,4.5233417,4.9058766,5.2884116,4.8279195,4.367427,3.9069343,3.4482548,2.9877625,4.507025,6.0281005,7.5473633,9.066626,10.587702,11.853149,13.116784,14.382232,15.64768,16.913128,15.542528,14.171928,12.803142,11.432542,10.061942,9.202598,8.343254,7.4820967,6.622752,5.763408,7.1883965,8.611572,10.038374,11.463363,12.888351,13.938056,14.9877615,16.037468,17.087172,18.136877,18.869314,19.601751,20.334188,21.066626,21.800875,21.429218,21.059374,20.68953,20.319685,19.94984,19.507477,19.065115,18.622751,18.18039,17.738026,16.98746,16.236893,15.488139,14.737573,13.987006,14.157425,14.327844,14.498261,14.666867,14.837286,15.502643,16.168001,16.833357,17.496902,18.16226,15.865235,13.568212,11.269376,8.972352,6.6753283,7.170267,7.665206,8.160145,8.655084,9.1500225,9.325879,9.499924,9.675781,9.849826,10.025683,9.947725,9.869768,9.791811,9.715667,9.637709,8.669587,7.703278,6.735156,5.767034,4.800725,4.421816,4.0447197,3.6676233,3.290527,2.911618,3.972201,5.032784,6.093367,7.1521373,8.212721,7.2591023,6.3072968,5.3554916,4.401873,3.4500678,3.6023567,3.7546456,3.9069343,4.059223,4.213325,4.1933823,4.171627,4.1516843,4.1317415,4.1117992,5.029158,5.9483304,6.8656893,7.783048,8.700407,11.14972,13.599032,16.050158,18.49947,20.950596,21.563377,22.174345,22.787127,23.399908,24.01269,23.822329,23.631968,23.441607,23.253057,23.062696,23.99456,24.928236,25.860098,26.791962,27.725637,25.994257,24.26469,22.535126,20.80556,19.074179,18.941833,18.809486,18.677141,18.544794,18.412449,18.557486,18.702522,18.847559,18.992596,19.137632,18.392506,17.647377,16.90225,16.157122,15.411995,15.428311,15.442815,15.457319,15.471823,15.488139,16.49796,17.50778,18.5176,19.52742,20.537241,21.046682,21.557938,22.06738,22.576822,23.088078,25.055143,27.022207,28.989271,30.958149,32.925213,28.352922,23.778818,19.206526,14.636047,10.061942,10.455356,10.846955,11.240368,11.631968,12.025381,12.565643,13.1059065,13.644357,14.184619,14.724882,15.919624,17.114367,18.310923,19.505665,20.700407,21.15002,21.599636,22.049252,22.500679,22.950293,22.785315,22.620335,22.455355,22.290375,22.125395,22.25049,22.375584,22.500679,22.625772,22.750868,0.038072214,0.045324065,0.052575916,0.059827764,0.06707962,0.07433146,0.37165734,0.67079616,0.968122,1.2654479,1.5627737,1.5373923,1.5120108,1.4866294,1.4630609,1.4376793,1.2527572,1.067835,0.88291276,0.6979906,0.51306844,0.47318324,0.43329805,0.39159992,0.35171473,0.31182957,1.2672608,2.222692,3.1781235,4.1317415,5.087173,5.315606,5.542227,5.77066,5.99728,6.2257137,5.870373,5.5150323,5.1596913,4.804351,4.4508233,4.41819,4.3855567,4.3529234,4.3202896,4.2876563,5.942891,7.5981264,9.253361,10.906783,12.562017,12.018129,11.472427,10.926725,10.382836,9.837135,9.432844,9.026741,8.62245,8.21816,7.8120556,7.7667317,7.723221,7.6778965,7.6325727,7.5872483,8.384952,9.182655,9.980359,10.778063,11.575767,11.740746,11.9057255,12.070704,12.235684,12.400664,12.172231,11.94561,11.717177,11.490557,11.262123,11.485118,11.708113,11.929294,12.152288,12.375282,12.317267,12.259253,12.203052,12.145037,12.087022,12.627284,13.167547,13.70781,14.248073,14.788336,13.822026,12.857531,11.893035,10.926725,9.96223,11.176914,12.3916,13.608097,14.8227825,16.037468,14.304275,12.572895,10.839704,9.108324,7.3751316,7.3316207,7.2899227,7.2482243,7.2047133,7.1630154,7.26998,7.3769445,7.4857225,7.592687,7.699652,7.835624,7.9697833,8.105756,8.239915,8.375887,8.519112,8.664148,8.809185,8.954222,9.099259,9.639522,10.179785,10.720048,11.26031,11.800573,11.017374,10.234174,9.452786,8.669587,7.8882003,7.835624,7.783048,7.7304726,7.6778965,7.6253204,7.5419245,7.460341,7.3769445,7.2953615,7.211965,7.3424983,7.473032,7.6017523,7.7322855,7.8628187,7.2391596,6.6173134,5.995467,5.371808,4.749962,4.784408,4.8206677,4.855114,4.88956,4.9258194,6.1423173,7.360628,8.577126,9.795437,11.011934,10.772624,10.533313,10.292189,10.052877,9.811753,10.411844,11.011934,11.612025,12.212116,12.812206,11.637406,10.462607,9.287807,8.113008,6.9382076,7.219217,7.502039,7.7848616,8.067683,8.350506,8.881703,9.414715,9.947725,10.480737,11.011934,11.280253,11.546759,11.815077,12.083396,12.349901,12.799516,13.24913,13.700559,14.150173,14.599788,14.492823,14.385859,14.277081,14.170115,14.06315,14.587097,15.112856,15.636803,16.162561,16.68832,16.849674,17.01284,17.174194,17.33736,17.500528,17.475147,17.449764,17.424383,17.400814,17.375433,17.437075,17.500528,17.562168,17.625622,17.687263,17.879436,18.071611,18.265598,18.457771,18.649946,20.042301,21.434656,22.827011,24.219368,25.611723,24.641787,23.671852,22.701918,21.731983,20.762047,19.984287,19.208338,18.430578,17.652817,16.875055,16.028402,15.179935,14.333282,13.484816,12.638163,12.670795,12.701616,12.734249,12.766883,12.799516,11.849524,10.899531,9.949538,8.999546,8.049554,7.3533764,6.6553855,5.957395,5.2594047,4.5632267,4.5469103,4.5324063,4.517903,4.503399,4.4870825,4.5632267,4.6375585,4.7118897,4.788034,4.8623657,4.0918565,3.3231604,2.5526514,1.7821422,1.0116332,0.8103943,0.6073425,0.40429065,0.2030518,0.0,0.07070554,0.13959812,0.21030366,0.27919623,0.34990177,0.27919623,0.21030366,0.13959812,0.07070554,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.13415924,0.14503701,0.15410182,0.16497959,0.17585737,0.13959812,0.10515183,0.07070554,0.034446288,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.21755551,0.40972954,0.60190356,0.79589057,0.9880646,0.79770356,0.6073425,0.4169814,0.22662032,0.038072214,0.19217403,0.3480888,0.50219065,0.65810543,0.8122072,0.8321498,0.8520924,0.872035,0.8919776,0.9119202,0.8557183,0.79770356,0.73968875,0.68167394,0.62547207,1.209246,1.794833,2.38042,2.9641938,3.5497808,3.9649491,4.3801174,4.795286,5.2104545,5.6256227,5.4969025,5.369995,5.243088,5.1143675,4.98746,5.297477,5.6074934,5.91751,6.2275267,6.5375433,5.6927023,4.847862,4.0030212,3.1581807,2.3133402,2.4257438,2.5381477,2.6505513,2.762955,2.8753586,2.3151531,1.7549478,1.1947423,0.6345369,0.07433146,0.07433146,0.07433146,0.07433146,0.07433146,0.07433146,0.18492219,0.2955129,0.40429065,0.5148814,0.62547207,1.3796645,2.13567,2.8898623,3.6458678,4.40006,5.195951,5.9900284,6.7859187,7.5799966,8.375887,7.6307597,6.885632,6.1405044,5.3953767,4.650249,5.6999545,6.7496595,7.799365,8.8508835,9.900589,10.515183,11.129777,11.744371,12.360779,12.975373,13.000754,13.024323,13.049705,13.075087,13.100468,12.964496,12.830337,12.694364,12.5602045,12.4242325,14.848164,17.27028,19.6924,22.114517,24.536636,24.36259,24.186733,24.01269,23.836832,23.662788,23.01556,22.368332,21.719292,21.072063,20.424837,18.736969,17.050913,15.363045,13.675177,11.9873085,11.889409,11.793322,11.695421,11.597522,11.499621,10.061942,8.624263,7.1865835,5.750717,4.313038,5.0781083,5.8431783,6.6082487,7.3733187,8.138389,7.554615,6.972654,6.390693,5.806919,5.224958,6.5030966,7.7794223,9.057561,10.3357,11.612025,12.843027,14.072216,15.303217,16.532406,17.761595,16.797098,15.8326025,14.868106,13.901797,12.937301,12.654479,12.371656,12.090648,11.807825,11.525003,12.28826,13.049705,13.812962,14.574407,15.337664,16.13718,16.936697,17.738026,18.537542,19.337059,19.703278,20.067682,20.432089,20.798307,21.162712,20.484665,19.80843,19.13038,18.452333,17.774284,17.364555,16.954826,16.545097,16.135366,15.725637,15.187187,14.650551,14.112101,13.575464,13.037014,13.278138,13.517449,13.75676,13.997884,14.237195,14.743011,15.247015,15.752831,16.256836,16.762651,14.766581,12.772322,10.778063,8.781991,6.787732,7.1031876,7.41683,7.7322855,8.047741,8.363196,8.762048,9.162713,9.563377,9.96223,10.362894,10.045626,9.728357,9.409276,9.092008,8.774739,7.9280853,7.079619,6.2329655,5.384499,4.537845,4.1825047,3.827164,3.4718235,3.1182957,2.762955,3.6077955,4.4526362,5.297477,6.1423173,6.987158,6.432391,5.8776245,5.3228583,4.7680917,4.213325,4.3801174,4.5469103,4.7155156,4.882308,5.049101,4.9983377,4.945762,4.893186,4.84061,4.788034,5.910258,7.0324817,8.154706,9.27693,10.399154,12.687112,14.975071,17.26303,19.549175,21.837133,22.388275,22.937603,23.48693,24.03807,24.587399,23.833206,23.0772,22.323008,21.567003,20.81281,22.027494,23.24218,24.456865,25.67155,26.888048,25.252756,23.617464,21.982172,20.34688,18.7134,18.196705,17.681824,17.166943,16.652061,16.13718,16.34023,16.543283,16.744522,16.947575,17.150625,16.80979,16.470764,16.129929,15.790904,15.4500675,15.62955,15.810846,15.99033,16.169813,16.349297,17.23221,18.115122,18.998035,19.879135,20.762047,21.220728,21.677593,22.13446,22.59314,23.050007,24.235683,25.419548,26.605227,27.789091,28.974768,25.466686,21.960415,18.452333,14.946064,11.437981,11.847711,12.25744,12.66717,13.0769,13.486629,13.716875,13.947122,14.177367,14.407614,14.63786,15.39024,16.142618,16.894999,17.647377,18.399757,19.224655,20.049553,20.87445,21.699348,22.524246,22.469858,22.41547,22.359268,22.304878,22.25049,22.536938,22.8252,23.111647,23.399908,23.68817,0.025381476,0.04169814,0.059827764,0.07795739,0.09427405,0.11240368,0.5529536,0.9916905,1.4322405,1.8727903,2.3133402,2.2245052,2.137483,2.0504606,1.9616255,1.8746033,1.5718386,1.2708868,0.968122,0.6653573,0.36259252,0.35171473,0.34264994,0.33177215,0.32270733,0.31182957,1.4322405,2.5526514,3.673062,4.7916603,5.9120708,5.8721857,5.8323007,5.7924156,5.75253,5.712645,5.467895,5.223145,4.9783955,4.7318325,4.4870825,4.7318325,4.9783955,5.223145,5.467895,5.712645,8.232663,10.752681,13.272699,15.792717,18.312735,17.194138,16.077353,14.960567,13.8419695,12.725184,11.7425585,10.7599325,9.7773075,8.794682,7.8120556,7.7703576,7.7268467,7.6851482,7.6416373,7.5999393,8.002417,8.404895,8.807372,9.20985,9.612328,9.672155,9.731983,9.791811,9.851639,9.91328,10.002114,10.092763,10.181598,10.272246,10.362894,10.903157,11.4416065,11.98187,12.522133,13.062395,13.16936,13.278138,13.385102,13.492067,13.600845,14.010575,14.420304,14.830034,15.239763,15.649493,14.327844,13.00438,11.682731,10.359268,9.037619,9.848013,10.656594,11.466989,12.277383,13.087777,11.856775,10.627586,9.396585,8.167397,6.9382076,7.079619,7.2228427,7.364254,7.507478,7.650702,7.6797094,7.71053,7.7395372,7.7703576,7.799365,8.002417,8.205468,8.406708,8.609759,8.812811,9.066626,9.322253,9.577881,9.8316965,10.087324,11.173288,12.25744,13.343405,14.427556,15.511708,14.507326,13.502945,12.496751,11.49237,10.487988,10.303066,10.118144,9.933222,9.7483,9.563377,9.420154,9.27693,9.135518,8.992294,8.8508835,8.832754,8.814624,8.798307,8.780178,8.762048,7.9842873,7.208339,6.430578,5.6528172,4.8750563,4.8152285,4.7554007,4.695573,4.6357455,4.574105,6.1332526,7.690587,9.247922,10.805257,12.362592,11.940171,11.517752,11.095331,10.672911,10.25049,10.587702,10.924912,11.262123,11.599335,11.938358,11.088079,10.2378,9.38752,8.537241,7.686961,7.9298983,8.172835,8.415772,8.656897,8.899834,9.280556,9.659465,10.040187,10.420909,10.799818,10.995618,11.189605,11.385405,11.579392,11.775192,12.4242325,13.075087,13.724127,14.37498,15.025834,14.61973,14.21544,13.809336,13.4050455,13.000754,13.588155,14.175554,14.762955,15.350354,15.937754,16.650248,17.362743,18.075237,18.787731,19.500225,19.211964,18.925516,18.637255,18.350807,18.062546,18.000906,17.937452,17.87581,17.812357,17.750717,17.55673,17.364555,17.172382,16.980207,16.788034,18.069798,19.351562,20.63514,21.916904,23.200481,22.645716,22.089136,21.53437,20.979603,20.424837,19.565493,18.704334,17.84499,16.985647,16.124489,15.596917,15.0693445,14.541773,14.014201,13.486629,13.4050455,13.321649,13.240066,13.15667,13.075087,11.775192,10.475298,9.175404,7.8755093,6.5756154,6.2220874,5.870373,5.516845,5.1651306,4.8116026,5.177821,5.542227,5.906632,6.2728505,6.637256,6.037165,5.4370747,4.836984,4.2368937,3.636803,3.045777,2.4529383,1.8600996,1.2672608,0.6744221,0.5402629,0.40429065,0.27013144,0.13415924,0.0,0.10515183,0.21030366,0.3154555,0.42060733,0.52575916,0.42060733,0.3154555,0.21030366,0.10515183,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.2030518,0.21755551,0.23205921,0.24837588,0.26287958,0.21030366,0.15772775,0.10515183,0.052575916,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.2955129,0.5529536,0.8103943,1.067835,1.3252757,1.064209,0.80495536,0.54570174,0.28463513,0.025381476,0.13234627,0.23931105,0.3480888,0.4550536,0.5620184,0.59283876,0.62184614,0.6526665,0.68167394,0.7124943,0.7197462,0.726998,0.73424983,0.7433147,0.7505665,1.3651608,1.9797552,2.5943494,3.2107568,3.825351,4.022964,4.220577,4.41819,4.615803,4.8116026,4.9276323,5.041849,5.1578784,5.272095,5.388125,5.678199,5.9682727,6.258347,6.546608,6.836682,5.906632,4.9783955,4.0483456,3.1182957,2.1882458,2.4620032,2.7375734,3.0131438,3.2869012,3.5624714,2.8608549,2.1574254,1.455809,0.7523795,0.05076295,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.17767033,0.24293698,0.30820364,0.37165734,0.43692398,1.1077201,1.7767034,2.4474995,3.1182957,3.787279,4.3420453,4.896812,5.4533916,6.008158,6.5629244,5.9447045,5.328297,4.710077,4.0918565,3.4754493,4.361988,5.2503395,6.1368785,7.02523,7.911769,9.023115,10.1326475,11.242181,12.351714,13.46306,13.312584,13.162108,13.011633,12.862969,12.712494,12.335398,11.958302,11.579392,11.202296,10.825199,13.189302,15.555219,17.919323,20.285238,22.649342,21.788185,20.925215,20.062244,19.199274,18.338116,18.33449,18.332678,18.330864,18.327238,18.325426,16.512463,14.699501,12.8865385,11.075388,9.262425,9.222541,9.182655,9.142771,9.102885,9.063,8.299743,7.5382986,6.775041,6.011784,5.2503395,6.397945,7.5455503,8.693155,9.840761,10.988366,10.283124,9.577881,8.872639,8.167397,7.462154,8.497355,9.5325575,10.567759,11.602961,12.638163,13.832905,15.027647,16.22239,17.417131,18.611874,18.051668,17.493277,16.933071,16.372866,15.812659,16.108173,16.401873,16.697386,16.992899,17.288412,17.388124,17.487837,17.58755,17.687263,17.786976,18.338116,18.887444,19.436771,19.987913,20.537241,20.535427,20.531801,20.529987,20.528175,20.52455,19.540112,18.555672,17.56942,16.584982,15.600543,15.221634,14.844538,14.467442,14.090345,13.713249,13.386916,13.062395,12.737875,12.413355,12.087022,12.397038,12.707055,13.017072,13.327088,13.637105,13.98338,14.327844,14.672306,15.016769,15.363045,13.669738,11.978244,10.284937,8.59163,6.9001355,7.0342946,7.170267,7.304426,7.440398,7.574558,8.200029,8.825501,9.449161,10.074633,10.700105,10.141713,9.585134,9.026741,8.470161,7.911769,7.1847706,6.4577727,5.730775,5.0019636,4.274966,3.9431937,3.6096084,3.2778363,2.9442513,2.612479,3.24339,3.872488,4.503399,5.132497,5.7615952,5.6056805,5.4479527,5.290225,5.132497,4.974769,5.1578784,5.3391747,5.522284,5.7053933,5.8866897,5.803293,5.718084,5.632875,5.5476656,5.462456,6.789545,8.116633,9.445535,10.772624,12.099712,14.224504,16.349297,18.475903,20.600695,22.725487,23.213173,23.70086,24.186733,24.674421,25.162107,23.842272,22.522434,21.202597,19.882761,18.562923,20.06043,21.557938,23.055445,24.552952,26.050459,24.509441,22.970236,21.429218,19.890013,18.350807,17.451578,16.554161,15.656745,14.759329,13.861912,14.122978,14.382232,14.643299,14.902553,15.161806,15.227073,15.292339,15.357606,15.422873,15.488139,15.8326025,16.177065,16.52334,16.867804,17.212267,17.968271,18.722466,19.476658,20.232662,20.986855,21.392958,21.797249,22.203352,22.607643,23.011934,23.414412,23.816889,24.219368,24.621845,25.024323,22.582262,20.140202,17.698141,15.254267,12.812206,13.240066,13.667925,14.095784,14.521831,14.94969,14.869919,14.790149,14.710379,14.630608,14.5508375,14.860854,15.170871,15.480887,15.789091,16.099108,17.29929,18.49947,19.699652,20.899832,22.100014,22.154404,22.210604,22.264994,22.319382,22.375584,22.8252,23.274813,23.724428,24.175856,24.625471,0.012690738,0.03988518,0.06707962,0.09427405,0.12328146,0.15047589,0.7324369,1.3143979,1.8981718,2.4801328,3.0620937,2.911618,2.762955,2.612479,2.4620032,2.3133402,1.892733,1.4721256,1.0533313,0.6327239,0.21211663,0.23205921,0.2520018,0.27194437,0.291887,0.31182957,1.5972201,2.8826106,4.168001,5.4533916,6.736969,6.430578,6.1223745,5.814171,5.5077806,5.199577,5.0654173,4.9294453,4.795286,4.6593137,4.5251546,5.047288,5.569421,6.093367,6.6155005,7.137634,10.522435,13.907236,17.292038,20.676838,24.06164,22.371958,20.682278,18.992596,17.302916,15.613234,14.052273,12.493125,10.932164,9.373016,7.8120556,7.7721705,7.7322855,7.6924005,7.652515,7.61263,7.6198816,7.6271334,7.6343856,7.6416373,7.650702,7.605378,7.560054,7.51473,7.4694057,7.4258947,7.8319983,8.239915,8.647832,9.055748,9.461852,10.319383,11.176914,12.034446,12.891977,13.749508,14.023266,14.29521,14.567154,14.839099,15.112856,15.392053,15.673061,15.952258,16.233267,16.512463,14.831847,13.153044,11.472427,9.791811,8.113008,8.517298,8.921589,9.327692,9.731983,10.138086,9.409276,8.682278,7.95528,7.228282,6.4994707,6.827617,7.155763,7.4820967,7.8102427,8.138389,8.089439,8.042302,7.995165,7.948028,7.900891,8.1692095,8.439341,8.709473,8.979604,9.249735,9.6141405,9.980359,10.344765,10.70917,11.075388,12.705242,14.335095,15.964949,17.5948,19.224655,17.99728,16.769903,15.542528,14.315152,13.087777,12.770509,12.45324,12.134158,11.81689,11.499621,11.298383,11.095331,10.89228,10.689227,10.487988,10.323009,10.15803,9.99305,9.82807,9.663091,8.729415,7.797552,6.8656893,5.9320135,5.0001507,4.844236,4.690134,4.5342193,4.3801174,4.2242026,6.1223745,8.020547,9.916905,11.815077,13.713249,13.107719,12.50219,11.896661,11.292944,10.687414,10.761745,10.837891,10.912222,10.988366,11.062697,10.536939,10.012992,9.487233,8.963287,8.437528,8.640579,8.841819,9.04487,9.247922,9.449161,9.677594,9.904215,10.1326475,10.359268,10.587702,10.70917,10.832452,10.955733,11.077202,11.200482,12.050762,12.899229,13.749508,14.599788,15.4500675,14.746637,14.045021,13.341592,12.639976,11.938358,12.5873995,13.238253,13.887294,14.538147,15.187187,16.450823,17.712645,18.974466,20.238102,21.499924,20.950596,20.399454,19.850128,19.3008,18.749659,18.562923,18.374376,18.187641,17.999092,17.812357,17.235836,16.6575,16.079165,15.502643,14.924308,16.097294,17.27028,18.443268,19.614443,20.78743,20.647831,20.508232,20.366821,20.227224,20.087626,19.144884,18.202145,17.259403,16.316664,15.375735,15.167245,14.960567,14.752076,14.545399,14.336908,14.139296,13.941682,13.745882,13.548269,13.3506565,11.700861,10.049252,8.399456,6.7496595,5.0998635,5.092612,5.08536,5.0781083,5.0708566,5.0617914,5.806919,6.552047,7.2971745,8.042302,8.78743,7.512917,6.2384043,4.9620786,3.6875658,2.4130533,1.9978848,1.5827163,1.167548,0.7523795,0.33721104,0.27013144,0.2030518,0.13415924,0.06707962,0.0,0.13959812,0.27919623,0.42060733,0.56020546,0.69980353,0.56020546,0.42060733,0.27919623,0.13959812,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,0.27013144,0.29007402,0.3100166,0.32995918,0.34990177,0.27919623,0.21030366,0.13959812,0.07070554,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.37165734,0.69436467,1.017072,1.3397794,1.6624867,1.3325275,1.0025684,0.6726091,0.34264994,0.012690738,0.072518505,0.13234627,0.19217403,0.2520018,0.31182957,0.35171473,0.39159992,0.43329805,0.47318324,0.51306844,0.5855869,0.65810543,0.7306239,0.8031424,0.87566096,1.5192627,2.1646774,2.810092,3.4555066,4.099108,4.079166,4.059223,4.0392804,4.019338,3.9993954,4.358362,4.7155156,5.0726695,5.429823,5.7869763,6.057108,6.3272395,6.5973706,6.867502,7.137634,6.1223745,5.1071157,4.0918565,3.0765975,2.0631514,2.5000753,2.9369993,3.3757362,3.8126602,4.249584,3.4047437,2.5599031,1.7150626,0.87022203,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.15047589,0.17041849,0.19036107,0.21030366,0.23024625,0.25018883,0.83577573,1.4195497,2.0051367,2.5907235,3.1744974,3.489953,3.8054085,4.120864,4.4345064,4.749962,4.2604623,3.7691493,3.2796493,2.7901495,2.3006494,3.0258346,3.7492065,4.4743915,5.199577,5.924762,7.5292335,9.135518,10.73999,12.344462,13.9507475,13.6244135,13.299893,12.975373,12.650853,12.32452,11.704487,11.084454,10.46442,9.844387,9.224354,11.532255,13.840157,16.148058,18.454145,20.762047,19.211964,17.661882,16.1118,14.561715,13.011633,13.655234,14.297023,14.940624,15.582414,16.224201,14.287958,12.349901,10.411844,8.4756,6.5375433,6.5556726,6.5719895,6.590119,6.6082487,6.624565,6.5375433,6.450521,6.3616858,6.2746634,6.187641,7.7177815,9.247922,10.778063,12.308203,13.838344,13.009819,12.183108,11.354585,10.527874,9.699349,10.493427,11.285692,12.077957,12.870221,13.662486,14.8227825,15.983078,17.143373,18.301857,19.462152,19.308052,19.152136,18.998035,18.84212,18.688019,19.560053,20.432089,21.304123,22.17797,23.050007,22.487988,21.924156,21.362139,20.80012,20.238102,20.537241,20.838192,21.137331,21.438282,21.737421,21.367577,20.997732,20.627888,20.258043,19.888199,18.595556,17.302916,16.010273,14.71763,13.424988,13.080525,12.734249,12.389787,12.045323,11.700861,11.586644,11.47424,11.361836,11.249433,11.137029,11.517752,11.896661,12.277383,12.658105,13.037014,13.221936,13.406858,13.591781,13.776703,13.961625,12.572895,11.182353,9.791811,8.403082,7.0125394,6.967215,6.921891,6.87838,6.833056,6.787732,7.6380115,8.488291,9.336758,10.1870365,11.037316,10.239613,9.441909,8.644206,7.8483152,7.0506115,6.4432693,5.8359265,5.2267714,4.6194286,4.0120864,3.7020695,3.392053,3.0820365,2.7720199,2.4620032,2.8771715,3.29234,3.7075086,4.122677,4.537845,4.7771564,5.0182805,5.2575917,5.4969025,5.7380266,5.9356394,6.1332526,6.3308654,6.526665,6.7242785,6.6082487,6.490406,6.3725634,6.2547207,6.1368785,7.6706448,9.202598,10.734551,12.266505,13.800271,15.761897,17.725336,19.68696,21.650398,23.612024,24.03807,24.462305,24.88835,25.312584,25.736816,23.85315,21.967669,20.082186,18.198519,16.313038,18.093367,19.871883,21.652212,23.43254,25.212872,23.767939,22.323008,20.878077,19.433146,17.988214,16.708263,15.428311,14.14836,12.868408,11.586644,11.9057255,12.222994,12.540262,12.857531,13.174799,13.644357,14.115726,14.585284,15.054841,15.524399,16.035654,16.545097,17.054539,17.565794,18.075237,18.702522,19.329807,19.957092,20.584377,21.211662,21.56519,21.916904,22.270432,22.622147,22.975676,22.594954,22.21423,21.835321,21.4546,21.07569,19.697838,18.319986,16.942135,15.564283,14.188245,14.632421,15.07841,15.522586,15.966762,16.41275,16.022963,15.633177,15.243389,14.851789,14.462003,14.329657,14.19731,14.064963,13.932617,13.800271,15.375735,16.949387,18.52485,20.100317,21.675781,21.84076,22.00574,22.17072,22.3357,22.500679,23.111647,23.724428,24.33721,24.949991,25.562773,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.9119202,1.6371052,2.3622901,3.0874753,3.8126602,3.6005437,3.386614,3.1744974,2.962381,2.7502642,2.2118144,1.6751775,1.1367276,0.6000906,0.06164073,0.11240368,0.16316663,0.21211663,0.26287958,0.31182957,1.7621996,3.2125697,4.6629395,6.11331,7.5618668,6.987158,6.412449,5.8377395,5.2630305,4.688321,4.6629395,4.6375585,4.612177,4.5867953,4.5632267,5.3627434,6.16226,6.9617763,7.763106,8.562622,12.812206,17.06179,21.313189,25.562773,29.812357,27.54978,25.287203,23.024624,20.762047,18.49947,16.361988,14.224504,12.087022,9.949538,7.8120556,7.7757964,7.7377243,7.699652,7.663393,7.6253204,7.2373466,6.849373,6.4632115,6.0752378,5.6872635,5.5367875,5.388125,5.237649,5.087173,4.936697,5.661882,6.3870673,7.112252,7.837437,8.562622,9.737422,10.912222,12.087022,13.261822,14.436621,14.875358,15.312282,15.749206,16.187943,16.624866,16.775343,16.92582,17.074482,17.224958,17.375433,15.337664,13.299893,11.262123,9.224354,7.1883965,7.1883965,7.1883965,7.1883965,7.1883965,7.1883965,6.9617763,6.736969,6.5121617,6.2873545,6.0625467,6.5756154,7.0868707,7.5999393,8.113008,8.624263,8.499168,8.375887,8.2507925,8.125698,8.000604,8.337815,8.675026,9.012237,9.349448,9.686659,10.161655,10.636651,11.111648,11.586644,12.06164,14.237195,16.41275,18.588305,20.762047,22.937603,21.487232,20.036863,18.588305,17.137936,15.687565,15.23795,14.788336,14.336908,13.887294,13.437678,13.174799,12.91192,12.650853,12.387974,12.125093,11.813264,11.499621,11.187792,10.874149,10.56232,9.474543,8.386765,7.3008003,6.2130227,5.125245,4.8750563,4.6248674,4.3746786,4.12449,3.874301,6.11331,8.350506,10.587702,12.824898,15.062093,14.275268,13.486629,12.699803,11.912977,11.124338,10.937603,10.750868,10.56232,10.375585,10.1870365,9.987611,9.788185,9.5869465,9.38752,9.188094,9.349448,9.512614,9.675781,9.837135,10.000301,10.074633,10.150778,10.225109,10.29944,10.375585,10.424535,10.475298,10.524248,10.57501,10.625773,11.675479,12.725184,13.77489,14.824595,15.8743,14.875358,13.874602,12.87566,11.874905,10.874149,11.586644,12.299138,13.011633,13.724127,14.436621,16.249584,18.062546,19.87551,21.686659,23.49962,22.687414,21.875206,21.063,20.250792,19.436771,19.124943,18.813112,18.49947,18.187641,17.87581,16.913128,15.950445,14.9877615,14.025079,13.062395,14.124791,15.187187,16.249584,17.31198,18.374376,18.649946,18.925516,19.199274,19.474844,19.750414,18.724277,17.699953,16.67563,15.649493,14.625169,14.737573,14.849977,14.96238,15.074784,15.187187,14.875358,14.561715,14.249886,13.938056,13.6244135,11.624716,9.625018,7.6253204,5.6256227,3.6241121,3.9631362,4.3003473,4.6375585,4.974769,5.3119802,6.43783,7.5618668,8.6877165,9.811753,10.937603,8.9868555,7.037921,5.087173,3.1382382,1.1874905,0.9499924,0.7124943,0.4749962,0.2374981,0.0,0.0,0.0,0.0,0.0,0.0,0.17585737,0.34990177,0.52575916,0.69980353,0.87566096,0.69980353,0.52575916,0.34990177,0.17585737,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06164073,0.12509441,0.18673515,0.25018883,0.31182957,0.33721104,0.36259252,0.387974,0.41335547,0.43692398,0.34990177,0.26287958,0.17585737,0.0870222,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.44961473,0.8375887,1.2255627,1.6117238,1.9996977,1.6008459,1.2001812,0.7995165,0.40066472,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.11240368,0.16316663,0.21211663,0.26287958,0.31182957,0.44961473,0.5873999,0.72518504,0.8629702,1.0007553,1.6751775,2.3495996,3.0258346,3.7002566,4.3746786,4.137181,3.8996825,3.6621845,3.4246864,3.1871881,3.787279,4.3873696,4.98746,5.5875506,6.187641,6.43783,6.688019,6.9382076,7.1883965,7.4367723,6.338117,5.237649,4.137181,3.0367124,1.938057,2.5381477,3.1382382,3.738329,4.3366065,4.936697,3.9504454,2.962381,1.9743162,0.9880646,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.16316663,0.13778515,0.11240368,0.0870222,0.06164073,0.5620184,1.062396,1.5627737,2.0631514,2.561716,2.6378605,2.712192,2.7883365,2.8626678,2.9369993,2.5744069,2.2118144,1.8492218,1.4866294,1.1258497,1.6878681,2.2498865,2.811905,3.3757362,3.9377546,6.037165,8.136576,10.2378,12.337211,14.436621,13.938056,13.437678,12.937301,12.436923,11.938358,11.075388,10.212419,9.349448,8.488291,7.6253204,9.875207,12.125093,14.37498,16.624866,18.874754,16.637558,14.400362,12.163166,9.924157,7.686961,8.975978,10.263181,11.5503845,12.837588,14.124791,12.06164,10.000301,7.93715,5.8758116,3.8126602,3.8869917,3.9631362,4.0374675,4.1117992,4.1879435,4.7753434,5.3627434,5.9501433,6.5375433,7.124943,9.037619,10.950294,12.862969,14.775645,16.68832,15.738328,14.788336,13.838344,12.888351,11.938358,12.487686,13.037014,13.588155,14.137483,14.68681,15.812659,16.936697,18.062546,19.188396,20.312433,20.562622,20.81281,21.063,21.313189,21.563377,23.011934,24.462305,25.912674,27.363045,28.811602,27.587852,26.36229,25.136726,23.912977,22.687414,22.738176,22.787127,22.837889,22.886839,22.937603,22.199726,21.461851,20.725788,19.987913,19.250036,17.64919,16.050158,14.449312,12.850279,11.249433,10.937603,10.625773,10.312131,10.000301,9.686659,9.788185,9.8878975,9.987611,10.087324,10.1870365,10.636651,11.088079,11.537694,11.9873085,12.436923,12.462305,12.487686,12.513068,12.536636,12.562017,11.47424,10.388275,9.300498,8.212721,7.124943,6.9001355,6.6753283,6.450521,6.2257137,6.000906,7.07418,8.149267,9.224354,10.29944,11.374527,10.337513,9.300498,8.26167,7.224656,6.187641,5.6999545,5.2122674,4.7245803,4.2368937,3.7492065,3.4627585,3.1744974,2.8880494,2.5997884,2.3133402,2.5127661,2.712192,2.911618,3.1128569,3.3122826,3.9504454,4.5867953,5.224958,5.863121,6.4994707,6.7134004,6.925517,7.137634,7.3497505,7.5618668,7.413204,7.262728,7.112252,6.9617763,6.813113,8.549932,10.28675,12.025381,13.762199,15.50083,17.29929,19.099562,20.899832,22.700104,24.500376,24.862968,25.225561,25.588154,25.950747,26.31334,23.862213,21.4129,18.961775,16.512463,14.06315,16.124489,18.187641,20.250792,22.31213,24.375282,23.024624,21.675781,20.325123,18.974466,17.625622,15.963136,14.300649,12.638163,10.975676,9.313189,9.686659,10.061942,10.437225,10.812509,11.187792,12.063453,12.937301,13.812962,14.68681,15.56247,16.236893,16.913128,17.58755,18.261972,18.938208,19.436771,19.93715,20.437527,20.937904,21.438282,21.737421,22.038374,22.337511,22.63665,22.937603,21.775494,20.611572,19.449463,18.287354,17.125244,16.811602,16.499773,16.187943,15.8743,15.56247,16.024776,16.487082,16.949387,17.411694,17.87581,17.174194,16.474392,15.774588,15.074784,14.37498,13.800271,13.225562,12.650853,12.07433,11.499621,13.45037,15.401117,17.350052,19.298986,21.249735,21.525305,21.800875,22.074633,22.350203,22.625772,23.399908,24.175856,24.949991,25.724127,26.500074,0.012690738,0.10515183,0.19761293,0.29007402,0.3825351,0.4749962,1.167548,1.8600996,2.5526514,3.245203,3.9377546,3.7909048,3.6422417,3.4953918,3.346729,3.199879,2.9968271,2.7955883,2.5925364,2.3894846,2.1882458,2.1229792,2.0577126,1.9924458,1.9271792,1.8619126,3.0620937,4.262275,5.462456,6.6626377,7.8628187,7.360628,6.8566246,6.354434,5.8522434,5.3500524,5.105303,4.860553,4.615803,4.36924,4.12449,4.95664,5.7906027,6.622752,7.454902,8.287052,11.985496,15.682126,19.38057,23.0772,26.775644,24.882912,22.99018,21.097446,19.204712,17.31198,15.408369,13.502945,11.597522,9.692098,7.7866745,7.752228,7.7177815,7.6833353,7.647076,7.61263,7.1829576,6.7532854,6.3218007,5.8921285,5.462456,5.3808727,5.297477,5.2158933,5.132497,5.049101,5.814171,6.5792413,7.344311,8.109382,8.874452,9.902402,10.930351,11.958302,12.984438,14.012388,14.402175,14.791962,15.181748,15.573349,15.963136,15.769149,15.576975,15.384801,15.192626,15.000452,13.278138,11.555823,9.8316965,8.109382,6.3870673,6.4577727,6.526665,6.5973706,6.6680765,6.736969,6.542982,6.347182,6.153195,5.957395,5.7615952,6.285541,6.8076744,7.3298078,7.851941,8.375887,8.274362,8.174648,8.074935,7.9752226,7.8755093,8.6333275,9.389333,10.147152,10.90497,11.662788,12.179482,12.697989,13.2146845,13.7331915,14.249886,15.676687,17.105303,18.532103,19.960718,21.38752,20.04774,18.70796,17.368181,16.026588,14.68681,14.144734,13.602658,13.060582,12.516694,11.974618,11.81689,11.6591625,11.503247,11.34552,11.187792,10.899531,10.613083,10.324821,10.038374,9.750113,8.985043,8.219973,7.454902,6.6898317,5.924762,5.883064,5.8395524,5.7978544,5.754343,5.712645,7.46578,9.217102,10.970237,12.7233715,14.474693,14.039582,13.604471,13.16936,12.734249,12.299138,11.862214,11.42529,10.988366,10.549629,10.112705,9.784559,9.458226,9.130079,8.801933,8.4756,8.979604,9.48542,9.989424,10.49524,10.999244,10.872336,10.745429,10.616709,10.489801,10.362894,10.662033,10.962985,11.262123,11.563075,11.862214,12.389787,12.917358,13.44493,13.972503,14.500074,13.551895,12.605529,11.65735,10.70917,9.762803,10.40278,11.042755,11.682731,12.322706,12.962683,14.53996,16.117237,17.694515,19.271791,20.850883,20.221785,19.5945,18.967215,18.33993,17.712645,17.504154,17.297476,17.090797,16.882307,16.67563,15.80722,14.940624,14.072216,13.20562,12.337211,13.443117,14.547212,15.653119,16.757214,17.863121,17.990028,18.116936,18.245655,18.372562,18.49947,17.75253,17.005589,16.256836,15.509895,14.762955,14.654177,14.547212,14.440247,14.333282,14.224504,14.005136,13.785768,13.564586,13.345218,13.125849,11.390844,9.655839,7.9208336,6.185828,4.4508233,4.860553,5.2702823,5.6800117,6.089741,6.4994707,7.057863,7.614443,8.172835,8.729415,9.287807,7.6198816,5.9519563,4.2858434,2.617918,0.9499924,0.97718686,1.0043813,1.0333886,1.0605831,1.0877775,0.9318628,0.7777609,0.62184614,0.46774435,0.31182957,0.60190356,0.8919776,1.1820517,1.4721256,1.7621996,1.5972201,1.4322405,1.2672608,1.1022812,0.93730164,0.7505665,0.5620184,0.37528324,0.18673515,0.0,0.0,0.0,0.0,0.0,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.24837588,0.3825351,0.5166943,0.6526665,0.7868258,0.823085,0.8575313,0.8919776,0.92823684,0.96268314,0.7705091,0.57833505,0.38434806,0.19217403,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.12509441,0.21211663,0.2991388,0.387974,0.4749962,0.83940166,1.2056202,1.5700256,1.9344311,2.3006494,1.845596,1.3905423,0.9354887,0.48043507,0.025381476,0.10515183,0.18492219,0.26469254,0.3444629,0.42423326,0.49675176,0.56927025,0.6417888,0.71430725,0.7868258,1.0116332,1.2382535,1.4630609,1.6878681,1.9126755,2.465629,3.0167696,3.5697234,4.122677,4.6756306,4.4725785,4.269527,4.068288,3.8652363,3.6621845,4.157123,4.652062,5.147001,5.6419396,6.1368785,6.2873545,6.43783,6.588306,6.736969,6.887445,5.883064,4.876869,3.872488,2.8681068,1.8619126,2.3405347,2.817344,3.294153,3.7727752,4.249584,3.4047437,2.5599031,1.7150626,0.87022203,0.025381476,0.3680314,0.7106813,1.0533313,1.3941683,1.7368182,1.5718386,1.4068589,1.2418793,1.0768998,0.9119202,1.2980812,1.6824293,2.0667772,2.4529383,2.8372865,2.8245957,2.811905,2.7992141,2.7883365,2.7756457,3.0203958,3.2651455,3.5098956,3.7546456,3.9993954,3.919625,3.8398547,3.7600844,3.680314,3.6005437,6.1405044,8.680465,11.220426,13.760386,16.300346,15.584227,14.869919,14.155612,13.439491,12.725184,12.5058155,12.284635,12.065266,11.845898,11.624716,12.848466,14.070402,15.292339,16.514277,17.738026,15.950445,14.162864,12.375282,10.587702,8.80012,10.812509,12.824898,14.837286,16.849674,18.862062,15.809033,12.757817,9.704789,6.6517596,3.6005437,3.8072214,4.0157123,4.2223897,4.4308805,4.6375585,5.3391747,6.0426044,6.7442207,7.4476504,8.149267,9.764616,11.379966,12.995316,14.610665,16.224201,15.676687,15.129172,14.581658,14.034143,13.486629,13.762199,14.037769,14.313339,14.587097,14.862667,16.157122,17.451578,18.747847,20.042301,21.336756,21.74286,22.14715,22.553255,22.957544,23.361835,24.262878,25.162107,26.06315,26.96238,27.861609,27.020395,26.177366,25.33434,24.493124,23.650097,23.70086,23.74981,23.800573,23.849524,23.900286,23.044567,22.190662,21.334944,20.479225,19.62532,18.292793,16.960264,15.627737,14.29521,12.962683,12.661731,12.362592,12.06164,11.762501,11.463363,11.379966,11.298383,11.214987,11.133403,11.050007,11.381779,11.715364,12.047136,12.380721,12.712494,12.400664,12.087022,11.775192,11.463363,11.14972,10.190662,9.229793,8.270736,7.309865,6.350808,6.3145485,6.2801023,6.245656,6.209397,6.1749506,7.3570023,8.540867,9.7229185,10.90497,12.087022,11.2168,10.348391,9.4781685,8.607946,7.7377243,7.3968873,7.057863,6.717026,6.378002,6.037165,5.5458527,5.0527267,4.559601,4.068288,3.5751622,3.6077955,3.6404288,3.673062,3.7056956,3.738329,4.2894692,4.842423,5.3953767,5.9483304,6.4994707,6.7279043,6.9545245,7.1829576,7.409578,7.6380115,7.650702,7.663393,7.6742706,7.686961,7.699652,9.140957,10.58045,12.019942,13.4594345,14.90074,16.173439,17.444326,18.717026,19.989725,21.262424,21.550686,21.837133,22.125395,22.411844,22.700104,21.052122,19.404139,17.757969,16.109985,14.462003,16.13174,17.803293,19.473032,21.142769,22.812508,21.585133,20.357758,19.13038,17.903006,16.67563,15.346728,14.01964,12.692551,11.365462,10.038374,10.489801,10.943042,11.39447,11.847711,12.299138,13.16936,14.039582,14.909804,15.780026,16.650248,16.8533,17.054539,17.257591,17.460642,17.661882,18.426952,19.192022,19.957092,20.722162,21.487232,21.78456,22.081884,22.37921,22.678349,22.975676,22.098202,21.220728,20.343254,19.465778,18.588305,18.649946,18.7134,18.77504,18.836681,18.900135,18.809486,18.720652,18.630003,18.539356,18.45052,17.730774,17.009214,16.289469,15.569723,14.849977,14.168303,13.484816,12.803142,12.119655,11.437981,13.05333,14.666867,16.282217,17.897566,19.512917,20.267109,21.023113,21.777306,22.533312,23.287504,24.17767,25.067833,25.957998,26.848164,27.738327,0.025381476,0.17223145,0.3208944,0.46774435,0.61459434,0.76325727,1.4231756,2.0830941,2.7430124,3.4029307,4.062849,3.9794528,3.8978696,3.8144734,3.73289,3.6494937,3.7818398,3.9141862,4.0483456,4.1806917,4.313038,4.1317415,3.9522583,3.7727752,3.5932918,3.4119956,4.361988,5.3119802,6.261973,7.211965,8.161958,7.7322855,7.3026133,6.872941,6.4432693,6.011784,5.5476656,5.081734,4.6176157,4.1516843,3.6875658,4.552349,5.4171324,6.281915,7.1466985,8.013294,11.156972,14.302462,17.447952,20.593443,23.73712,22.21423,20.693155,19.170267,17.647377,16.124489,14.452938,12.779573,11.108022,9.434657,7.763106,7.7304726,7.6978393,7.665206,7.6325727,7.5999393,7.1267557,6.6553855,6.1822023,5.710832,5.237649,5.223145,5.2068286,5.1923246,5.177821,5.163317,5.9682727,6.773228,7.5781837,8.383139,9.188094,10.067381,10.946668,11.827768,12.707055,13.588155,13.930804,14.271642,14.614291,14.956942,15.299591,14.764768,14.229943,13.695119,13.1602955,12.625471,11.2168,9.80994,8.403082,6.9944096,5.5875506,5.727149,5.866747,6.008158,6.147756,6.2873545,6.1223745,5.957395,5.7924156,5.6274357,5.462456,5.995467,6.526665,7.059676,7.592687,8.125698,8.049554,7.9752226,7.900891,7.8247466,7.750415,8.927028,10.1054535,11.282066,12.460492,13.637105,14.19731,14.757515,15.31772,15.877926,16.438131,17.117992,17.797853,18.477715,19.157576,19.837437,18.608248,17.377247,16.148058,14.917056,13.687867,13.05333,12.416981,11.782444,11.147907,10.51337,10.460794,10.408218,10.355642,10.303066,10.25049,9.987611,9.724731,9.461852,9.200785,8.937905,8.495543,8.05318,7.610817,7.166641,6.7242785,6.889258,7.0542374,7.219217,7.3841968,7.549176,8.81825,10.085511,11.352772,12.620032,13.887294,13.80571,13.722314,13.640731,13.557334,13.475751,12.786825,12.099712,11.4126,10.725487,10.038374,9.583321,9.128266,8.673213,8.21816,7.763106,8.609759,9.458226,10.304879,11.153346,11.999999,11.67004,11.340081,11.010121,10.680162,10.3502035,10.899531,11.450671,11.999999,12.549327,13.100468,13.104094,13.109532,13.114971,13.12041,13.125849,12.230246,11.334642,10.440851,9.545248,8.649645,9.217102,9.784559,10.352016,10.919474,11.486931,12.830337,14.171928,15.515334,16.856926,18.20033,17.757969,17.315605,16.873243,16.43088,15.986704,15.885179,15.781839,15.680313,15.576975,15.475449,14.703127,13.930804,13.15667,12.384347,11.612025,12.75963,13.907236,15.054841,16.202446,17.350052,17.330109,17.310167,17.290224,17.27028,17.25034,16.78078,16.309412,15.839854,15.3702965,14.90074,14.572594,14.244447,13.918114,13.589968,13.261822,13.134913,13.008006,12.879286,12.752378,12.625471,11.155159,9.684846,8.214534,6.7442207,5.275721,5.7579694,6.240217,6.722465,7.2047133,7.686961,7.6778965,7.667019,7.6579537,7.647076,7.6380115,6.2529078,4.8678045,3.482701,2.0975976,0.7124943,1.0043813,1.2980812,1.5899682,1.8818551,2.175555,1.8655385,1.5555218,1.2455053,0.9354887,0.62547207,1.0297627,1.4358664,1.840157,2.2444477,2.6505513,2.4946365,2.3405347,2.18462,2.030518,1.8746033,1.49932,1.1258497,0.7505665,0.37528324,0.0,0.0,0.0,0.0,0.0,0.0,0.045324065,0.09064813,0.13415924,0.1794833,0.22480737,0.43329805,0.6399758,0.8466535,1.0551442,1.261822,1.3071461,1.35247,1.3977941,1.4431182,1.4866294,1.1893034,0.8919776,0.5946517,0.29732585,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.2374981,0.40066472,0.5620184,0.72518504,0.8883517,1.2291887,1.5718386,1.9144884,2.2571385,2.5997884,2.0903459,1.5809034,1.0696479,0.56020546,0.05076295,0.19761293,0.3444629,0.49312583,0.6399758,0.7868258,0.88291276,0.97718686,1.0732739,1.167548,1.261822,1.5754645,1.887294,2.1991236,2.5127661,2.8245957,3.254268,3.6857529,4.115425,4.5450974,4.974769,4.8079767,4.6393714,4.4725785,4.305786,4.137181,4.5269675,4.9167547,5.3083544,5.6981416,6.0879283,6.1368785,6.187641,6.2384043,6.2873545,6.338117,5.42801,4.517903,3.6077955,2.6976883,1.7875811,2.1429217,2.4982624,2.8517902,3.207131,3.5624714,2.8608549,2.1574254,1.455809,0.7523795,0.05076295,0.6979906,1.3452182,1.9924458,2.6396735,3.2869012,2.9823234,2.6777458,2.373168,2.0667772,1.7621996,2.032331,2.3024626,2.572594,2.8427253,3.1128569,3.0131438,2.911618,2.811905,2.712192,2.612479,3.4645715,4.3166637,5.1705694,6.0226617,6.874754,6.153195,5.429823,4.708264,3.9848917,3.2633326,6.24203,9.222541,12.203052,15.181748,18.16226,17.23221,16.30216,15.372109,14.4420595,13.512011,13.93443,14.356851,14.779271,15.201692,15.624111,15.819912,16.01571,16.209698,16.405499,16.599485,15.261519,13.925365,12.5873995,11.249433,9.91328,12.650853,15.386614,18.124187,20.861761,23.599335,19.556427,15.515334,11.472427,7.4295206,3.386614,3.727451,4.068288,4.407312,4.748149,5.087173,5.904819,6.722465,7.5401115,8.357758,9.175404,10.493427,11.809638,13.127662,14.445685,15.761897,15.616859,15.471823,15.326786,15.181748,15.036712,15.036712,15.036712,15.036712,15.036712,15.036712,16.503399,17.968271,19.433146,20.89802,22.362894,22.9231,23.483305,24.041697,24.601902,25.162107,25.512009,25.861912,26.211813,26.561714,26.911617,26.452936,25.992445,25.531952,25.073273,24.61278,24.66173,24.712494,24.763256,24.812206,24.862968,23.889408,22.91766,21.9441,20.972351,20.000603,18.934582,17.870373,16.80435,15.740141,14.674119,14.387671,14.09941,13.812962,13.524701,13.238253,12.971747,12.707055,12.442362,12.17767,11.912977,12.126906,12.342649,12.558392,12.772322,12.988064,12.337211,11.6881695,11.037316,10.388275,9.737422,8.9052725,8.073122,7.2391596,6.4070096,5.57486,5.730775,5.8848767,6.0407915,6.1948934,6.350808,7.6398244,8.930654,10.21967,11.510499,12.799516,12.097899,11.39447,10.692853,9.989424,9.287807,9.0956335,8.901647,8.709473,8.517298,8.325124,7.6271334,6.929143,6.2329655,5.5349746,4.836984,4.702825,4.5668526,4.4326935,4.2967215,4.162562,4.6303062,5.0980506,5.565795,6.0317264,6.4994707,6.742408,6.985345,7.228282,7.4694057,7.7123427,7.8882003,8.062244,8.238102,8.412147,8.588004,9.73017,10.872336,12.0145035,13.15667,14.300649,15.045776,15.789091,16.534218,17.279346,18.024473,18.238403,18.45052,18.662638,18.874754,19.08687,18.24203,17.397188,16.55235,15.707508,14.862667,16.140806,17.417131,18.69527,19.971596,21.249735,20.14564,19.039734,17.935638,16.829731,15.725637,14.732134,13.740443,12.74694,11.755249,10.761745,11.292944,11.822329,12.351714,12.882912,13.412297,14.277081,15.141864,16.006647,16.873243,17.738026,17.467894,17.197763,16.927631,16.6575,16.38737,17.417131,18.446894,19.476658,20.508232,21.537996,21.831696,22.127209,22.422722,22.718235,23.011934,22.419096,21.82807,21.235231,20.642391,20.049553,20.48829,20.925215,21.362139,21.799063,22.237799,21.594198,20.952408,20.31062,19.667019,19.025229,18.285542,17.544039,16.80435,16.064661,15.324973,14.534521,13.744069,12.955431,12.164979,11.374527,12.654479,13.93443,15.214382,16.494333,17.774284,19.010725,20.245354,21.47998,22.71461,23.949236,24.95543,25.959812,26.964193,27.970387,28.974768,0.038072214,0.23931105,0.44236287,0.64541465,0.8466535,1.0497054,1.6769904,2.3042755,2.9333735,3.5606585,4.1879435,4.169814,4.1516843,4.135368,4.117238,4.099108,4.5668526,5.034597,5.5023413,5.9700856,6.43783,6.1423173,5.846804,5.5531044,5.2575917,4.9620786,5.661882,6.3616858,7.063302,7.763106,8.46291,8.105756,7.746789,7.3896356,7.0324817,6.6753283,5.9900284,5.3047285,4.6194286,3.9341288,3.2506418,4.1480584,5.045475,5.942891,6.8403077,7.7377243,10.330261,12.922797,15.515334,18.10787,20.700407,19.547363,18.394318,17.243088,16.090042,14.936998,13.497506,12.058014,10.616709,9.177217,7.7377243,7.706904,7.6778965,7.647076,7.6180687,7.5872483,7.072367,6.5574856,6.0426044,5.527723,5.0128417,5.0654173,5.1179934,5.1705694,5.223145,5.275721,6.1205616,6.965402,7.8102427,8.655084,9.499924,10.232361,10.964798,11.697234,12.429671,13.162108,13.457622,13.753134,14.046834,14.342347,14.63786,13.760386,12.882912,12.005438,11.127964,10.25049,9.157274,8.06587,6.972654,5.8794374,4.788034,4.9983377,5.2068286,5.4171324,5.6274357,5.8377395,5.7017674,5.567608,5.431636,5.297477,5.163317,5.7053933,6.247469,6.789545,7.3316207,7.8755093,7.8247466,7.7757964,7.7250338,7.6742706,7.6253204,9.222541,10.81976,12.416981,14.014201,15.613234,16.215137,16.817041,17.420757,18.022661,18.624565,18.557486,18.490406,18.423326,18.354433,18.287354,17.166943,16.048346,14.927934,13.807523,12.687112,11.9601145,11.233116,10.504305,9.7773075,9.050309,9.102885,9.155461,9.208037,9.2606125,9.313189,9.07569,8.838193,8.600695,8.363196,8.125698,8.00423,7.8845744,7.764919,7.645263,7.5256076,7.897265,8.270736,8.642392,9.015862,9.38752,10.17072,10.952107,11.735307,12.516694,13.299893,13.5700245,13.840157,14.110288,14.380419,14.650551,13.713249,12.774135,11.836833,10.899531,9.96223,9.380268,8.798307,8.214534,7.6325727,7.0506115,8.239915,9.429218,10.620335,11.809638,13.000754,12.467744,11.934732,11.401722,10.870523,10.337513,11.137029,11.938358,12.737875,13.537392,14.336908,13.820213,13.301706,12.785012,12.268318,11.74981,10.906783,10.065568,9.222541,8.379513,7.5382986,8.033237,8.528176,9.023115,9.518054,10.012992,11.120712,12.22662,13.33434,14.4420595,15.54978,15.292339,15.034899,14.777458,14.520018,14.262577,14.26439,14.268016,14.269829,14.271642,14.275268,13.597219,12.919171,12.242936,11.564888,10.88684,12.077957,13.267261,14.458377,15.64768,16.836983,16.67019,16.503399,16.334793,16.168001,15.999394,15.80722,15.6150465,15.422873,15.230699,15.036712,14.489197,13.941682,13.394168,12.846653,12.299138,12.264692,12.230246,12.195799,12.15954,12.125093,10.919474,9.715667,8.510046,7.304426,6.1006193,6.6553855,7.210152,7.764919,8.319685,8.874452,8.29793,7.7195945,7.1430726,6.5647373,5.9882154,4.8841214,3.7818398,2.6795588,1.5772774,0.4749962,1.0333886,1.5899682,2.1483607,2.70494,3.2633326,2.7974012,2.333283,1.8673514,1.403233,0.93730164,1.4576219,1.9779422,2.4982624,3.0167696,3.53709,3.392053,3.247016,3.101979,2.956942,2.811905,2.2498865,1.6878681,1.1258497,0.5620184,0.0,0.0,0.0,0.0,0.0,0.0,0.06707962,0.13415924,0.2030518,0.27013144,0.33721104,0.61822027,0.8974165,1.1766127,1.4576219,1.7368182,1.79302,1.8474089,1.9017978,1.9579996,2.0123885,1.6099107,1.2074331,0.80495536,0.40247768,0.0,0.0,0.0,0.0,0.0,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.34990177,0.5873999,0.824898,1.062396,1.2998942,1.6207886,1.93987,2.2607644,2.5798457,2.9007401,2.335096,1.7694515,1.2056202,0.6399758,0.07433146,0.29007402,0.5058166,0.7197462,0.9354887,1.1494182,1.2672608,1.3851035,1.502946,1.6207886,1.7368182,2.137483,2.5381477,2.9369993,3.3376641,3.738329,4.0447197,4.3529234,4.6593137,4.9675174,5.275721,5.143375,5.009216,4.876869,4.744523,4.612177,4.896812,5.18326,5.467895,5.75253,6.037165,5.9882154,5.9374523,5.8866897,5.8377395,5.7869763,4.972956,4.157123,3.343103,2.5272698,1.7132497,1.9453088,2.1773682,2.4094272,2.6432993,2.8753586,2.3151531,1.7549478,1.1947423,0.6345369,0.07433146,1.0279498,1.9797552,2.9333735,3.8851788,4.836984,4.3928084,3.9468195,3.5026438,3.056655,2.612479,2.7683938,2.9224956,3.0784104,3.2325122,3.386614,3.199879,3.0131438,2.8245957,2.6378605,2.4493124,3.9105604,5.369995,6.82943,8.290678,9.750113,8.384952,7.019791,5.65463,4.2894692,2.9243085,6.345369,9.764616,13.185677,16.604925,20.024172,18.880192,17.7344,16.59042,15.444629,14.300649,15.364858,16.429068,17.495089,18.559298,19.62532,18.79317,17.959208,17.127058,16.294909,15.462758,14.574407,13.687867,12.799516,11.912977,11.024626,14.487384,17.950142,21.4129,24.87566,28.336605,23.303822,18.27285,13.240066,8.207282,3.1744974,3.6476808,4.120864,4.592234,5.0654173,5.5367875,6.4704633,7.402326,8.334189,9.267865,10.199727,11.220426,12.23931,13.260008,14.280706,15.299591,15.557032,15.814472,16.071913,16.329353,16.586794,16.313038,16.037468,15.761897,15.488139,15.212569,16.84786,18.483154,20.118446,21.751925,23.387217,24.103338,24.817644,25.531952,26.248072,26.96238,26.762953,26.561714,26.36229,26.162863,25.961624,25.885479,25.807522,25.729565,25.651608,25.575462,25.624413,25.675177,25.724127,25.774889,25.825651,24.73425,23.644657,22.555067,21.465477,20.375887,19.578182,18.78048,17.982777,17.185072,16.38737,16.1118,15.838041,15.56247,15.2869005,15.013144,14.565341,14.117539,13.669738,13.221936,12.774135,12.872034,12.969934,13.067834,13.165734,13.261822,12.27557,11.287505,10.29944,9.313189,8.325124,7.6198816,6.9146395,6.209397,5.504154,4.800725,5.145188,5.4896507,5.8341136,6.1803894,6.5248523,7.9226465,9.32044,10.718235,12.114216,13.512011,12.977186,12.442362,11.907538,11.372714,10.837891,10.792566,10.747242,10.701918,10.658407,10.613083,9.710228,8.807372,7.9045167,7.0016613,6.1006193,5.7978544,5.4950895,5.1923246,4.88956,4.5867953,4.9693303,5.351866,5.7344007,6.1169357,6.4994707,6.7569118,7.0143523,7.271793,7.5292335,7.7866745,8.125698,8.46291,8.80012,9.137331,9.474543,10.319383,11.164224,12.010877,12.855718,13.700559,13.918114,14.13567,14.353225,14.57078,14.788336,14.924308,15.062093,15.199879,15.337664,15.475449,15.431937,15.39024,15.346728,15.30503,15.263332,16.148058,17.032784,17.91751,18.802235,19.68696,18.704334,17.721708,16.739084,15.758271,14.775645,14.117539,13.4594345,12.803142,12.145037,11.486931,12.094274,12.701616,13.310771,13.918114,14.525456,15.384801,16.245958,17.105303,17.964645,18.825804,18.082489,17.339174,16.597672,15.854358,15.112856,16.40731,17.701767,18.998035,20.29249,21.586945,21.880646,22.172533,22.464418,22.75812,23.050007,22.741802,22.435411,22.127209,21.820818,21.512613,22.324821,23.137028,23.949236,24.763256,25.575462,24.38072,23.184166,21.989424,20.794682,19.59994,18.840307,18.080675,17.319231,16.5596,15.799969,14.902553,14.005136,13.107719,12.210303,11.312886,12.25744,13.201994,14.14836,15.092914,16.037468,17.75253,19.467592,21.182655,22.897717,24.61278,25.73319,26.85179,27.9722,29.092611,30.213022,0.05076295,0.30820364,0.5656443,0.823085,1.0805258,1.3379664,1.9326181,2.5272698,3.1219215,3.7183862,4.313038,4.360175,4.407312,4.454449,4.503399,4.550536,5.351866,6.155008,6.9581504,7.75948,8.562622,8.152893,7.743163,7.3316207,6.921891,6.5121617,6.9617763,7.413204,7.8628187,8.312433,8.762048,8.477413,8.192778,7.9081426,7.6216946,7.3370595,6.432391,5.527723,4.6230545,3.7183862,2.811905,3.7419548,4.6720047,5.6020546,6.532104,7.462154,9.501737,11.543133,13.582716,15.622298,17.661882,16.880495,16.097294,15.314095,14.532708,13.749508,12.542075,11.334642,10.127209,8.919776,7.7123427,7.6851482,7.6579537,7.6307597,7.6017523,7.574558,7.017978,6.4595857,5.903006,5.3446136,4.788034,4.9076896,5.027345,5.147001,5.2666564,5.388125,6.2728505,7.157576,8.042302,8.927028,9.811753,10.397341,10.982927,11.566701,12.152288,12.737875,12.984438,13.232814,13.479377,13.727753,13.974316,12.754191,11.535881,10.315757,9.0956335,7.8755093,7.0977483,6.319988,5.542227,4.764466,3.9867048,4.267714,4.5469103,4.8279195,5.1071157,5.388125,5.282973,5.177821,5.0726695,4.9675174,4.8623657,5.4153194,5.9682727,6.5194135,7.072367,7.6253204,7.5999393,7.574558,7.549176,7.5256076,7.500226,9.518054,11.534068,13.551895,15.569723,17.58755,18.232965,18.876566,19.52198,20.167397,20.81281,19.996977,19.182957,18.367125,17.553104,16.73727,15.72745,14.71763,13.70781,12.697989,11.6881695,10.866898,10.047439,9.22798,8.406708,7.5872483,7.744976,7.902704,8.0604315,8.21816,8.375887,8.161958,7.949841,7.7377243,7.5256076,7.311678,7.51473,7.7177815,7.9208336,8.122072,8.325124,8.9052725,9.48542,10.065568,10.645717,11.225864,11.5231905,11.820516,12.117842,12.415168,12.712494,13.33434,13.957999,14.579845,15.201692,15.825351,14.63786,13.45037,12.262879,11.075388,9.8878975,9.177217,8.4683485,7.757667,7.0469856,6.338117,7.8700705,9.402024,10.93579,12.467744,13.999697,13.265448,12.529385,11.795135,11.060884,10.324821,11.374527,12.4242325,13.475751,14.525456,15.575162,14.534521,13.495693,12.455053,11.4144125,10.375585,9.585134,8.794682,8.00423,7.215591,6.4251394,6.8475595,7.26998,7.6924005,8.1148205,8.537241,9.409276,10.283124,11.155159,12.027194,12.899229,12.826711,12.754191,12.681673,12.609155,12.536636,12.645414,12.752378,12.859344,12.968122,13.075087,12.493125,11.909351,11.327391,10.745429,10.161655,11.39447,12.627284,13.860099,15.092914,16.325727,16.010273,15.694818,15.379361,15.065719,14.750263,14.835473,14.920682,15.005891,15.089288,15.174497,14.407614,13.640731,12.872034,12.105151,11.338268,11.39447,11.452485,11.510499,11.566701,11.624716,10.685601,9.744674,8.805559,7.8646317,6.925517,7.552802,8.180087,8.807372,9.434657,10.061942,8.917963,7.7721705,6.628191,5.482399,4.3366065,3.5171473,2.6976883,1.8782293,1.0569572,0.2374981,1.0605831,1.8818551,2.70494,3.5280252,4.349297,3.729264,3.1092308,2.4891977,1.8691645,1.2491312,1.8854811,2.520018,3.1545548,3.7909048,4.4254417,4.2894692,4.15531,4.019338,3.8851788,3.7492065,3.000453,2.2498865,1.49932,0.7505665,0.0,0.0,0.0,0.0,0.0,0.0,0.09064813,0.1794833,0.27013144,0.36077955,0.44961473,0.8031424,1.1548572,1.5083848,1.8600996,2.2118144,2.277081,2.3423476,2.4076142,2.472881,2.5381477,2.030518,1.5228885,1.015259,0.5076295,0.0,0.0,0.0,0.0,0.0,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.46230546,0.774135,1.0877775,1.3996071,1.7132497,2.0105755,2.3079014,2.6052272,2.902553,3.199879,2.5798457,1.9598125,1.3397794,0.7197462,0.099712946,0.3825351,0.6653573,0.9481794,1.2291887,1.5120108,1.651609,1.79302,1.9326181,2.0722163,2.2118144,2.6995013,3.1871881,3.6748753,4.162562,4.650249,4.835171,5.0200934,5.2050157,5.389938,5.57486,5.47696,5.3808727,5.282973,5.185073,5.087173,5.2666564,5.4479527,5.6274357,5.806919,5.9882154,5.8377395,5.6872635,5.5367875,5.388125,5.237649,4.517903,3.7981565,3.0765975,2.3568513,1.6371052,1.7476959,1.8582866,1.9670644,2.077655,2.1882458,1.7694515,1.35247,0.9354887,0.5166943,0.099712946,1.357909,2.6142921,3.872488,5.130684,6.3870673,5.803293,5.217706,4.632119,4.0483456,3.4627585,3.5026438,3.5425289,3.5824142,3.6222992,3.6621845,3.386614,3.1128569,2.8372865,2.561716,2.2879589,4.3547363,6.4233265,8.490104,10.556881,12.625471,10.616709,8.609759,6.60281,4.59586,2.5870976,6.446895,10.306692,14.168303,18.0281,21.887897,20.528175,19.166641,17.80692,16.447197,15.087475,16.795286,18.503096,20.210907,21.916904,23.624716,21.764616,19.904516,18.044416,16.184317,14.324218,13.887294,13.45037,13.011633,12.574709,12.137785,16.325727,20.511858,24.699802,28.887745,33.07569,27.051214,21.030367,15.007704,8.985043,2.962381,3.5679104,4.171627,4.7771564,5.382686,5.9882154,7.0342946,8.082188,9.130079,10.177972,11.225864,11.947423,12.670795,13.392355,14.115726,14.837286,15.497204,16.157122,16.817041,17.47696,18.136877,17.58755,17.038223,16.487082,15.937754,15.386614,17.192324,18.998035,20.801933,22.607643,24.413355,25.281763,26.151985,27.022207,27.89243,28.762651,28.012085,27.26333,26.512764,25.762197,25.011631,25.318022,25.6226,25.927177,26.231756,26.538147,26.587097,26.63786,26.68681,26.737572,26.788336,25.579088,24.371656,23.164223,21.956789,20.749357,20.219973,19.690586,19.15939,18.630003,18.100618,17.837738,17.57486,17.31198,17.0491,16.788034,16.157122,15.528025,14.897114,14.268016,13.637105,13.617162,13.597219,13.577277,13.557334,13.537392,12.212116,10.88684,9.561564,8.238102,6.9128265,6.3344913,5.7579694,5.179634,4.603112,4.024777,4.559601,5.0944247,5.6292486,6.165886,6.70071,8.205468,9.710228,11.214987,12.719746,14.224504,13.858286,13.490254,13.122223,12.754191,12.387974,12.489499,12.592838,12.694364,12.797703,12.899229,11.793322,10.685601,9.577881,8.470161,7.362441,6.892884,6.4233265,5.9519563,5.482399,5.0128417,5.3101673,5.6074934,5.904819,6.202145,6.4994707,6.773228,7.0451727,7.317117,7.590874,7.8628187,8.363196,8.861761,9.362139,9.862516,10.362894,10.910409,11.457924,12.005438,12.552953,13.100468,12.790451,12.480434,12.170418,11.860401,11.5503845,11.612025,11.675479,11.73712,11.800573,11.862214,12.621845,13.383289,14.142921,14.902553,15.662184,16.15531,16.646622,17.139748,17.632874,18.124187,17.264843,16.405499,15.544341,14.684997,13.825653,13.502945,13.180238,12.857531,12.534823,12.212116,12.897416,13.582716,14.268016,14.953316,15.636803,16.492521,17.34824,18.202145,19.057863,19.911768,18.697083,17.482399,16.267714,15.053028,13.838344,15.397491,16.958452,18.5176,20.076748,21.637709,21.927782,22.217857,22.50793,22.798004,23.088078,23.06451,23.042755,23.019186,22.99743,22.975676,24.163166,25.350657,26.538147,27.725637,28.913128,27.165432,25.417736,23.67004,21.922344,20.174648,19.395073,18.6155,17.834112,17.054539,16.274965,15.270584,14.26439,13.260008,12.255627,11.249433,11.860401,12.469557,13.080525,13.68968,14.300649,16.494333,18.68983,20.885328,23.079014,25.274511,26.510952,27.745579,28.980207,30.214834,31.449461,0.06164073,0.37528324,0.6871128,1.0007553,1.3125849,1.6244144,2.1882458,2.7502642,3.3122826,3.874301,4.4381323,4.550536,4.6629395,4.7753434,4.8877473,5.0001507,6.1368785,7.2754188,8.412147,9.550687,10.687414,10.161655,9.637709,9.11195,8.588004,8.062244,8.26167,8.46291,8.662335,8.861761,9.063,8.8508835,8.636953,8.424837,8.212721,8.000604,6.874754,5.750717,4.6248674,3.5008307,2.374981,3.3376641,4.3003473,5.2630305,6.2257137,7.1883965,8.675026,10.161655,11.650098,13.136727,14.625169,14.211814,13.800271,13.386916,12.975373,12.562017,11.586644,10.613083,9.637709,8.662335,7.686961,7.663393,7.6380115,7.61263,7.5872483,7.5618668,6.9617763,6.3616858,5.7615952,5.163317,4.5632267,4.749962,4.936697,5.125245,5.3119802,5.5005283,6.4251394,7.3497505,8.274362,9.200785,10.125396,10.56232,10.999244,11.437981,11.874905,12.311829,12.513068,12.712494,12.91192,13.113158,13.312584,11.74981,10.1870365,8.624263,7.063302,5.5005283,5.038223,4.5759177,4.1117992,3.6494937,3.1871881,3.53709,3.8869917,4.2368937,4.5867953,4.936697,4.8623657,4.788034,4.7118897,4.6375585,4.5632267,5.125245,5.6872635,6.249282,6.813113,7.3751316,7.3751316,7.3751316,7.3751316,7.3751316,7.3751316,9.811753,12.250188,14.68681,17.125244,19.561867,20.250792,20.937904,21.625017,22.31213,22.999243,21.438282,19.87551,18.312735,16.749962,15.187187,14.287958,13.386916,12.487686,11.586644,10.687414,9.775495,8.861761,7.949841,7.037921,6.1241875,6.3870673,6.6499467,6.9128265,7.175706,7.4367723,7.250037,7.063302,6.874754,6.688019,6.4994707,7.02523,7.549176,8.074935,8.600695,9.12464,9.91328,10.700105,11.486931,12.27557,13.062395,12.87566,12.687112,12.500377,12.311829,12.125093,13.100468,14.075842,15.049402,16.024776,17.00015,15.56247,14.124791,12.687112,11.249433,9.811753,8.974165,8.138389,7.3008003,6.4632115,5.6256227,7.500226,9.374829,11.249433,13.125849,15.000452,14.06315,13.125849,12.186734,11.249433,10.312131,11.612025,12.91192,14.211814,15.511708,16.811602,15.250641,13.687867,12.125093,10.56232,8.999546,8.26167,7.5256076,6.787732,6.049856,5.3119802,5.661882,6.011784,6.3616858,6.7134004,7.063302,7.699652,8.337815,8.974165,9.612328,10.25049,10.362894,10.475298,10.587702,10.700105,10.812509,11.024626,11.236742,11.450671,11.662788,11.874905,11.3872175,10.899531,10.411844,9.924157,9.438283,10.712796,11.9873085,13.261822,14.538147,15.812659,15.350354,14.888049,14.425743,13.961625,13.499319,13.861912,14.224504,14.587097,14.94969,15.312282,14.324218,13.337966,12.349901,11.361836,10.375585,10.524248,10.674724,10.825199,10.975676,11.124338,10.449916,9.775495,9.099259,8.424837,7.750415,8.450218,9.1500225,9.849826,10.549629,11.249433,9.537996,7.8247466,6.11331,4.40006,2.6868105,2.1501737,1.6117238,1.0750868,0.53663695,0.0,1.0877775,2.175555,3.2633326,4.349297,5.4370747,4.6629395,3.8869917,3.1128569,2.3369088,1.5627737,2.3133402,3.0620937,3.8126602,4.5632267,5.3119802,5.186886,5.0617914,4.936697,4.8116026,4.688321,3.7492065,2.811905,1.8746033,0.93730164,0.0,0.0,0.0,0.0,0.0,0.0,0.11240368,0.22480737,0.33721104,0.44961473,0.5620184,0.9880646,1.4122978,1.8383441,2.2625773,2.6868105,2.762955,2.8372865,2.911618,2.9877625,3.0620937,2.4493124,1.8383441,1.2255627,0.61278135,0.0,0.0,0.0,0.0,0.0,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.5747091,0.96268314,1.3506571,1.7368182,2.124792,2.4003625,2.6741197,2.94969,3.2252605,3.5008307,2.8245957,2.1501737,1.4757515,0.7995165,0.12509441,0.4749962,0.824898,1.1747998,1.5247015,1.8746033,2.03777,2.1991236,2.3622901,2.525457,2.6868105,3.2633326,3.8380418,4.4127507,4.98746,5.562169,5.6256227,5.6872635,5.750717,5.812358,5.8758116,5.812358,5.750717,5.6872635,5.6256227,5.562169,5.638314,5.712645,5.7869763,5.863121,5.9374523,5.6872635,5.4370747,5.186886,4.936697,4.688321,4.062849,3.437377,2.811905,2.1882458,1.5627737,1.550083,1.5373923,1.5247015,1.5120108,1.49932,1.2255627,0.9499924,0.6744221,0.40066472,0.12509441,1.6878681,3.2506418,4.8134155,6.3743763,7.93715,7.211965,6.48678,5.7615952,5.038223,4.313038,4.2368937,4.162562,4.0882306,4.0120864,3.9377546,3.5751622,3.2125697,2.8499773,2.4873846,2.124792,4.800725,7.474845,10.150778,12.824898,15.50083,12.850279,10.199727,7.549176,4.900438,2.2498865,6.550234,10.850581,15.1509285,19.449463,23.74981,22.174345,20.600695,19.025229,17.449764,15.8743,18.225714,20.575312,22.924911,25.274511,27.624111,24.737875,21.849825,18.961775,16.075539,13.1874895,13.200181,13.212872,13.225562,13.238253,13.24913,18.16226,23.075388,27.988516,32.899834,37.81296,30.80042,23.787882,16.775343,9.762803,2.7502642,3.48814,4.2242026,4.9620786,5.6999545,6.43783,7.5999393,8.762048,9.924157,11.088079,12.250188,12.674421,13.100468,13.524701,13.9507475,14.37498,15.437376,16.499773,17.562168,18.624565,19.68696,18.862062,18.037165,17.212267,16.38737,15.56247,17.536787,19.512917,21.487232,23.463362,25.437677,26.462002,27.488138,28.512463,29.536787,30.562923,29.26303,27.963135,26.66324,25.363346,24.06164,24.750565,25.437677,26.12479,26.811903,27.50083,27.54978,27.600542,27.649492,27.700254,27.749205,26.425743,25.100468,23.77519,22.449915,21.12464,20.861761,20.600695,20.337814,20.074934,19.812056,19.561867,19.311678,19.063301,18.813112,18.562923,17.750717,16.936697,16.124489,15.312282,14.500074,14.362289,14.224504,14.0867195,13.9507475,13.812962,12.1504755,10.487988,8.825501,7.1630154,5.5005283,5.049101,4.599486,4.1498713,3.7002566,3.2506418,3.975827,4.699199,5.424384,6.149569,6.874754,8.488291,10.100015,11.711739,13.325275,14.936998,14.737573,14.538147,14.336908,14.137483,13.938056,14.188245,14.436621,14.68681,14.936998,15.187187,13.874602,12.562017,11.249433,9.936848,8.624263,7.987913,7.3497505,6.7115874,6.0752378,5.4370747,5.6491914,5.863121,6.0752378,6.2873545,6.4994707,6.787732,7.07418,7.362441,7.650702,7.93715,8.600695,9.262425,9.924157,10.587702,11.249433,11.499621,11.74981,11.999999,12.250188,12.500377,11.662788,10.825199,9.987611,9.1500225,8.312433,8.299743,8.287052,8.274362,8.26167,8.2507925,9.811753,11.374527,12.937301,14.500074,16.062849,16.162561,16.262274,16.361988,16.4617,16.563227,15.825351,15.087475,14.349599,13.611723,12.87566,12.888351,12.899229,12.91192,12.92461,12.937301,13.700559,14.462003,15.22526,15.986704,16.749962,17.60024,18.45052,19.3008,20.149265,20.999546,19.311678,17.625622,15.937754,14.249886,12.562017,14.387671,16.213324,18.037165,19.862818,21.686659,21.97492,22.26318,22.54963,22.837889,23.124338,23.387217,23.650097,23.912977,24.175856,24.436922,25.999697,27.56247,29.125244,30.688017,32.25079,29.950142,27.649492,25.350657,23.050007,20.749357,19.94984,19.150324,18.350807,17.549479,16.749962,15.636803,14.525456,13.412297,12.300951,11.187792,11.463363,11.73712,12.012691,12.28826,12.562017,15.23795,17.912071,20.588003,23.262123,25.938055,27.2869,28.637556,29.988214,31.337059,32.687714,0.2755703,0.5982776,0.91917205,1.2418793,1.5645868,1.887294,2.4148662,2.9424384,3.4700103,3.9975824,4.5251546,4.8152285,5.105303,5.3953767,5.6854506,5.975525,7.1992745,8.424837,9.6504,10.874149,12.099712,11.675479,11.249433,10.825199,10.399154,9.97492,9.731983,9.490859,9.247922,9.004985,8.762048,8.562622,8.363196,8.161958,7.9625316,7.763106,6.695271,5.6274357,4.559601,3.491766,2.4257438,3.2306993,4.0356545,4.84061,5.6455655,6.450521,7.5346723,8.620637,9.704789,10.790753,11.874905,11.880343,11.885782,11.889409,11.894848,11.900287,11.347333,10.794379,10.243238,9.690285,9.137331,8.861761,8.588004,8.312433,8.036863,7.763106,7.5382986,7.311678,7.0868707,6.8620634,6.637256,6.3852544,6.1332526,5.8794374,5.6274357,5.375434,6.149569,6.925517,7.699652,8.4756,9.249735,9.577881,9.904215,10.232361,10.560507,10.88684,10.995618,11.102583,11.209548,11.318325,11.42529,10.2142315,9.004985,7.795739,6.58468,5.375434,4.876869,4.3801174,3.8833659,3.3848011,2.8880494,3.529838,4.171627,4.8152285,5.4570174,6.1006193,5.8431783,5.5857377,5.328297,5.0708566,4.8116026,5.5150323,6.2166486,6.9200783,7.6216946,8.325124,8.317872,8.31062,8.303369,8.294304,8.287052,10.141713,11.998186,13.852847,15.707508,17.562168,18.301857,19.04336,19.783049,20.522736,21.262424,19.63801,18.011784,16.38737,14.762955,13.136727,12.513068,11.887595,11.262123,10.636651,10.012992,9.510801,9.006798,8.504607,8.002417,7.500226,7.5419245,7.5854354,7.6271334,7.6706448,7.7123427,7.413204,7.112252,6.813113,6.5121617,6.2130227,6.967215,7.723221,8.477413,9.233418,9.987611,10.779876,11.57214,12.364405,13.15667,13.9507475,13.753134,13.555521,13.357908,13.1602955,12.962683,13.615349,14.268016,14.920682,15.573349,16.224201,15.134612,14.045021,12.955431,11.86584,10.774437,9.933222,9.090195,8.247167,7.404139,6.5629244,8.062244,9.561564,11.062697,12.562017,14.06315,13.339779,12.618219,11.894848,11.173288,10.449916,11.684544,12.919171,14.155612,15.39024,16.624866,15.192626,13.760386,12.328146,10.894093,9.461852,8.78743,8.113008,7.4367723,6.7623506,6.0879283,6.4033837,6.717026,7.0324817,7.3479376,7.663393,8.287052,8.912524,9.537996,10.161655,10.7871275,10.846955,10.906783,10.966611,11.028252,11.088079,11.720803,12.351714,12.984438,13.617162,14.249886,14.191871,14.13567,14.077655,14.01964,13.961625,14.474693,14.9877615,15.50083,16.012085,16.525154,16.13718,15.749206,15.363045,14.975071,14.587097,14.909804,15.2325115,15.555219,15.877926,16.200634,14.947877,13.695119,12.442362,11.189605,9.936848,10.25049,10.56232,10.874149,11.187792,11.499621,11.084454,10.669285,10.254116,9.840761,9.425592,9.347635,9.269678,9.19172,9.115576,9.037619,7.6597667,6.281915,4.9040637,3.5280252,2.1501737,1.7205015,1.2908293,0.85934424,0.42967212,0.0,0.9481794,1.8945459,2.8427253,3.7909048,4.7372713,4.3003473,3.8616104,3.4246864,2.9877625,2.5508385,2.8898623,3.2306993,3.5697234,3.9105604,4.249584,4.2949085,4.3402324,4.3855567,4.4308805,4.4743915,3.83079,3.1853752,2.5399606,1.8945459,1.2491312,1.4630609,1.6751775,1.887294,2.0994108,2.3133402,1.9942589,1.6769904,1.3597219,1.0424535,0.72518504,1.0098201,1.2944553,1.5809034,1.8655385,2.1501737,2.2100015,2.269829,2.3296568,2.3894846,2.4493124,1.9598125,1.4703126,0.9808127,0.4894999,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.23205921,0.45324063,0.6726091,0.8919776,1.1131591,1.7803292,2.4474995,3.1146698,3.7818398,4.4508233,4.6593137,4.8696175,5.0799212,5.290225,5.5005283,4.7318325,3.9649491,3.198066,2.42937,1.6624867,2.0468347,2.4329958,2.817344,3.2016919,3.587853,3.8978696,4.207886,4.517903,4.8279195,5.137936,5.6274357,6.1169357,6.6082487,7.0977483,7.5872483,7.2953615,7.0016613,6.7097745,6.4178877,6.1241875,6.109684,6.09518,6.0806766,6.0643597,6.049856,5.9447045,5.8395524,5.7344007,5.6292486,5.524097,5.2648435,5.0055895,4.744523,4.4852695,4.2242026,3.8525455,3.4808881,3.1074178,2.7357605,2.3622901,2.5544643,2.7466383,2.9406252,3.1327994,3.3249733,3.002266,2.6795588,2.3568513,2.034144,1.7132497,3.1654327,4.6176157,6.069799,7.5219817,8.974165,8.334189,7.6942134,7.0542374,6.414262,5.774286,5.7017674,5.6292486,5.5567303,5.484212,5.411693,5.0581656,4.702825,4.347484,3.9921436,3.636803,5.805106,7.9715962,10.139899,12.308203,14.474693,12.219368,9.965856,7.71053,5.4552045,3.199879,6.6155005,10.029309,13.44493,16.860552,20.27436,19.08687,17.89938,16.71189,15.524399,14.336908,16.34567,18.352621,20.35957,22.368332,24.375282,22.08007,19.78486,17.48965,15.194439,12.899229,13.345218,13.789393,14.235382,14.679558,15.125546,18.247469,21.36939,24.493124,27.615046,30.736967,25.234627,19.732285,14.229943,8.727602,3.2252605,3.7618973,4.3003473,4.836984,5.375434,5.9120708,7.079619,8.247167,9.414715,10.582263,11.74981,12.308203,12.864782,13.423175,13.979754,14.538147,15.480887,16.421816,17.364555,18.307297,19.250036,18.443268,17.634687,16.827919,16.019337,15.212569,17.074482,18.938208,20.80012,22.662033,24.525759,25.113157,25.700558,26.287958,26.875357,27.462757,26.188244,24.911919,23.637405,22.362894,21.08838,21.71204,22.337511,22.962984,23.586643,24.212114,24.302763,24.391598,24.482246,24.572895,24.66173,23.532255,22.402779,21.273302,20.142014,19.012539,19.021603,19.03248,19.04336,19.052423,19.063301,18.542982,18.022661,17.50234,16.982021,16.4617,16.189756,15.917811,15.645867,15.372109,15.100165,14.889862,14.679558,14.4692545,14.260764,14.05046,12.230246,10.410031,8.589817,6.7696023,4.949388,4.710077,4.4707656,4.229642,3.9903307,3.7492065,4.4381323,5.125245,5.812358,6.4994707,7.1883965,8.500981,9.811753,11.124338,12.436923,13.749508,13.794832,13.840157,13.885481,13.930804,13.974316,14.594349,15.214382,15.834415,16.454449,17.074482,15.95951,14.844538,13.729566,12.6145935,11.499621,10.66022,9.820818,8.979604,8.140202,7.3008003,7.2427855,7.1847706,7.1267557,7.0705543,7.0125394,7.1956487,7.3769445,7.560054,7.743163,7.9244595,8.352319,8.780178,9.208037,9.634083,10.061942,10.192475,10.323009,10.451729,10.582263,10.712796,10.266808,9.822631,9.376642,8.9324665,8.488291,8.653271,8.81825,8.98323,9.14821,9.313189,10.770811,12.22662,13.684241,15.141864,16.599485,16.67019,16.740896,16.80979,16.880495,16.949387,16.334793,15.720199,15.105604,14.489197,13.874602,13.874602,13.874602,13.874602,13.874602,13.874602,14.730321,15.584227,16.439945,17.295664,18.149569,19.046986,19.9444,20.841818,21.739235,22.63665,21.392958,20.147453,18.901947,17.658255,16.41275,18.100618,19.788486,21.474543,23.16241,24.850279,24.51488,24.179482,23.845898,23.510498,23.1751,23.624716,24.07433,24.525759,24.975372,25.424988,26.980509,28.536032,30.08974,31.645262,33.200783,31.143072,29.08536,27.027647,24.969934,22.912222,22.440851,21.967669,21.494484,21.023113,20.54993,19.25185,17.955582,16.6575,15.359419,14.06315,14.567154,15.072971,15.576975,16.08279,16.586794,18.747847,20.907085,23.068136,25.227375,27.386612,28.035654,28.68288,29.330109,29.977337,30.624563,0.48768693,0.8194591,1.1530442,1.4848163,1.8184015,2.1501737,2.6432993,3.1346123,3.6277382,4.120864,4.612177,5.0799212,5.5476656,6.01541,6.4831543,6.9508986,8.26167,9.574255,10.88684,12.199425,13.512011,13.1874895,12.862969,12.536636,12.212116,11.887595,11.202296,10.516996,9.8316965,9.14821,8.46291,8.274362,8.087626,7.900891,7.7123427,7.5256076,6.5157876,5.504154,4.494334,3.484514,2.474694,3.1219215,3.7691493,4.41819,5.0654173,5.712645,6.394319,7.077806,7.75948,8.442966,9.12464,9.547061,9.969481,10.391902,10.8143215,11.236742,11.108022,10.9774885,10.846955,10.718235,10.587702,10.061942,9.537996,9.012237,8.488291,7.9625316,8.113008,8.26167,8.412147,8.562622,8.713099,8.020547,7.327995,6.635443,5.942891,5.2503395,5.8758116,6.4994707,7.124943,7.750415,8.375887,8.59163,8.809185,9.026741,9.244296,9.461852,9.4781685,9.492672,9.507175,9.52168,9.537996,8.680465,7.8229337,6.965402,6.107871,5.2503395,4.7173285,4.1843176,3.6531196,3.1201086,2.5870976,3.5225863,4.458075,5.391751,6.3272395,7.262728,6.8221784,6.3816285,5.942891,5.5023413,5.0617914,5.904819,6.7478466,7.590874,8.432089,9.275117,9.2606125,9.244296,9.229793,9.215289,9.200785,10.471672,11.744371,13.017072,14.289771,15.56247,16.354736,17.147,17.939264,18.733343,19.525606,17.837738,16.14987,14.462003,12.774135,11.088079,10.738177,10.388275,10.038374,9.686659,9.336758,9.244296,9.151835,9.059374,8.966913,8.874452,8.696781,8.519112,8.343254,8.165584,7.987913,7.574558,7.1630154,6.7496595,6.338117,5.924762,6.9092,7.895452,8.87989,9.864329,10.850581,11.648285,12.444175,13.2418785,14.039582,14.837286,14.630608,14.422117,14.21544,14.006948,13.800271,14.13023,14.46019,14.790149,15.120108,15.4500675,14.706753,13.965251,13.221936,12.480434,11.73712,10.890467,10.042,9.195346,8.34688,7.500226,8.624263,9.750113,10.874149,11.999999,13.125849,12.618219,12.11059,11.602961,11.095331,10.587702,11.757062,12.928236,14.097597,15.266958,16.438131,15.134612,13.832905,12.529385,11.227677,9.924157,9.313189,8.700407,8.087626,7.474845,6.8620634,7.1430726,7.422269,7.703278,7.9824743,8.26167,8.874452,9.487233,10.100015,10.712796,11.325577,11.332829,11.340081,11.347333,11.354585,11.361836,12.415168,13.466686,14.520018,15.573349,16.624866,16.998337,17.369995,17.741652,18.115122,18.48678,18.238403,17.988214,17.738026,17.487837,17.237648,16.92582,16.612177,16.300346,15.986704,15.674874,15.957697,16.240519,16.52334,16.80435,17.087172,15.569723,14.052273,12.534823,11.017374,9.499924,9.97492,10.449916,10.924912,11.399909,11.874905,11.720803,11.564888,11.410787,11.254871,11.10077,10.245051,9.389333,8.535428,7.6797094,6.825804,5.7833505,4.740897,3.6966307,2.6541772,1.6117238,1.2908293,0.968122,0.64541465,0.32270733,0.0,0.80676836,1.6153497,2.422118,3.2306993,4.0374675,3.9377546,3.8380418,3.738329,3.636803,3.53709,3.4681973,3.397492,3.3267863,3.2578938,3.1871881,3.4029307,3.6168604,3.832603,4.0483456,4.262275,3.9105604,3.5570326,3.2053177,2.8517902,2.5000753,2.9243085,3.350355,3.774588,4.2006345,4.6248674,3.877927,3.1291735,2.382233,1.6352923,0.8883517,1.0333886,1.1766127,1.3216497,1.4666867,1.6117238,1.6570477,1.7023718,1.7476959,1.79302,1.8383441,1.4703126,1.1022812,0.73424983,0.3680314,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.42785916,0.83033687,1.2328146,1.6352923,2.03777,2.9859493,3.9323158,4.880495,5.826862,6.775041,6.9200783,7.065115,7.210152,7.3551893,7.500226,6.639069,5.7797246,4.9203806,4.059223,3.199879,3.6204863,4.0392804,4.459888,4.880495,5.2992897,5.7579694,6.2148356,6.6717024,7.130382,7.5872483,7.993352,8.397643,8.801933,9.208037,9.612328,8.9651,8.317872,7.6706448,7.021604,6.3743763,6.4070096,6.439643,6.472276,6.5049095,6.5375433,6.2529078,5.9682727,5.6818247,5.3971896,5.1125546,4.842423,4.572292,4.3021603,4.0320287,3.7618973,3.6422417,3.5225863,3.4029307,3.2832751,3.1618068,3.5606585,3.9576974,4.3547363,4.751775,5.1506267,4.780782,4.409125,4.0392804,3.6694362,3.299592,4.6429973,5.9845896,7.327995,8.669587,10.012992,9.458226,8.901647,8.34688,7.7921133,7.2373466,7.166641,7.0977483,7.027043,6.9581504,6.887445,6.539356,6.19308,5.844991,5.4969025,5.1506267,6.8094873,8.470161,10.130835,11.789696,13.45037,11.59027,9.73017,7.8700705,6.009971,4.1498713,6.680767,9.20985,11.740746,14.269829,16.800724,15.999394,15.199879,14.400362,13.600845,12.799516,14.465629,16.129929,17.794228,19.46034,21.12464,19.422268,17.719896,16.017525,14.315152,12.612781,13.490254,14.367728,15.245202,16.122677,17.00015,18.332678,19.665205,20.997732,22.33026,23.662788,19.670645,15.6785,11.684544,7.6924005,3.7002566,4.0374675,4.3746786,4.7118897,5.049101,5.388125,6.5592985,7.7322855,8.9052725,10.078259,11.249433,11.940171,12.629097,13.319836,14.010575,14.699501,15.522586,16.34567,17.166943,17.990028,18.813112,18.022661,17.23221,16.441757,15.653119,14.862667,16.612177,18.361685,20.113007,21.862516,23.612024,23.7625,23.912977,24.06164,24.212114,24.36259,23.111647,21.862516,20.611572,19.36244,18.11331,18.675327,19.237347,19.799364,20.363195,20.925215,21.055748,21.184467,21.315,21.445534,21.574255,20.64058,19.70509,18.769602,17.834112,16.900436,17.18326,17.464268,17.747091,18.029913,18.312735,17.522284,16.731833,15.9431925,15.152741,14.362289,14.630608,14.897114,15.165432,15.431937,15.700256,15.417434,15.134612,14.851789,14.57078,14.287958,12.310016,10.332074,8.354132,6.378002,4.40006,4.36924,4.3402324,4.309412,4.2804046,4.249584,4.900438,5.5494785,6.200332,6.849373,7.500226,8.511859,9.525306,10.536939,11.5503845,12.562017,12.852092,13.142166,13.43224,13.722314,14.012388,15.002265,15.992143,16.982021,17.971897,18.961775,18.044416,17.127058,16.209698,15.292339,14.37498,13.332527,12.290073,11.24762,10.205167,9.162713,8.834567,8.508233,8.180087,7.851941,7.5256076,7.6017523,7.6797094,7.757667,7.835624,7.911769,8.105756,8.29793,8.490104,8.682278,8.874452,8.885329,8.894395,8.9052725,8.914337,8.925215,8.872639,8.820063,8.767487,8.714911,8.662335,9.004985,9.347635,9.690285,10.032935,10.375585,11.728055,13.080525,14.432995,15.785465,17.137936,17.17782,17.217705,17.257591,17.297476,17.33736,16.844234,16.352922,15.859797,15.366671,14.875358,14.862667,14.849977,14.837286,14.824595,14.811904,15.760084,16.708263,17.654629,18.60281,19.549175,20.495543,21.440096,22.38465,23.329203,24.27557,23.472427,22.669285,21.867954,21.064812,20.26167,21.811752,23.361835,24.911919,26.462002,28.012085,27.05484,26.097597,25.140352,24.183107,23.225864,23.862213,24.500376,25.136726,25.774889,26.413052,27.959509,29.507778,31.054235,32.602505,34.150776,32.334187,30.519413,28.704636,26.88986,25.075085,24.930048,24.785011,24.639975,24.494938,24.349901,22.866898,21.385706,19.902702,18.4197,16.936697,17.67276,18.40701,19.143072,19.877321,20.613384,22.257742,23.9021,25.54827,27.192625,28.836983,28.782595,28.728205,28.672003,28.617615,28.563225,0.69980353,1.0424535,1.3851035,1.7277533,2.0704033,2.4130533,2.8699198,3.3267863,3.785466,4.2423325,4.699199,5.3446136,5.9900284,6.635443,7.2808576,7.9244595,9.325879,10.725487,12.125093,13.524701,14.924308,14.699501,14.474693,14.249886,14.025079,13.800271,12.672608,11.544946,10.417283,9.28962,8.161958,7.987913,7.8120556,7.6380115,7.462154,7.28811,6.3344913,5.382686,4.4290676,3.4772623,2.525457,3.0149567,3.5044568,3.9957695,4.4852695,4.974769,5.2557783,5.5349746,5.814171,6.09518,6.3743763,7.215591,8.054993,8.894395,9.735609,10.57501,10.866898,11.160598,11.452485,11.744371,12.038072,11.262123,10.487988,9.712041,8.937905,8.161958,8.6877165,9.211663,9.737422,10.263181,10.7871275,9.655839,8.5227375,7.3896356,6.258347,5.125245,5.600241,6.0752378,6.550234,7.02523,7.500226,7.607191,7.7141557,7.8229337,7.9298983,8.036863,7.9607186,7.8827615,7.804804,7.7268467,7.650702,7.1448855,6.640882,6.1350656,5.6292486,5.125245,4.557788,3.9903307,3.4228733,2.855416,2.2879589,3.5153344,4.74271,5.9700856,7.1974616,8.424837,7.802991,7.179332,6.5574856,5.9356394,5.3119802,6.294606,7.2772317,8.259857,9.242483,10.225109,10.203354,10.179785,10.15803,10.13446,10.112705,10.801631,11.49237,12.183108,12.872034,13.562773,14.407614,15.252454,16.097294,16.942135,17.786976,16.037468,14.287958,12.536636,10.7871275,9.037619,8.963287,8.887142,8.812811,8.736667,8.662335,8.979604,9.296872,9.6141405,9.933222,10.25049,9.851639,9.4546,9.057561,8.660522,8.26167,7.7377243,7.211965,6.688019,6.16226,5.638314,6.8529987,8.067683,9.282369,10.497053,11.711739,12.514881,13.318023,14.119352,14.922495,15.725637,15.508082,15.290526,15.072971,14.855415,14.63786,14.645112,14.652364,14.6596155,14.666867,14.674119,14.280706,13.885481,13.490254,13.095029,12.699803,11.847711,10.995618,10.141713,9.28962,8.437528,9.188094,9.936848,10.687414,11.437981,12.186734,11.894848,11.602961,11.30926,11.017374,10.725487,11.829581,12.935488,14.039582,15.14549,16.249584,15.07841,13.905423,12.732436,11.559449,10.388275,9.837135,9.287807,8.736667,8.187339,7.6380115,7.8827615,8.127511,8.372261,8.617011,8.861761,9.461852,10.061942,10.662033,11.262123,11.862214,11.81689,11.773379,11.728055,11.682731,11.637406,13.109532,14.581658,16.055597,17.527721,18.999847,19.80299,20.60432,21.407463,22.210604,23.011934,22.000301,20.986855,19.975222,18.961775,17.950142,17.712645,17.475147,17.237648,17.00015,16.762651,17.005589,17.246714,17.48965,17.732588,17.975525,16.193382,14.409427,12.627284,10.845142,9.063,9.699349,10.337513,10.975676,11.612025,12.250188,12.35534,12.460492,12.565643,12.670795,12.774135,11.142468,9.510801,7.877322,6.245656,4.612177,3.9051213,3.198066,2.4891977,1.7821422,1.0750868,0.85934424,0.64541465,0.42967212,0.21574254,0.0,0.6671702,1.3343405,2.0033236,2.6704938,3.3376641,3.5751622,3.8126602,4.0501585,4.2876563,4.5251546,4.0447197,3.5642843,3.0856624,2.6052272,2.124792,2.5091403,2.8953013,3.2796493,3.6658103,4.0501585,3.9903307,3.930503,3.870675,3.8108473,3.7492065,4.3873696,5.0255322,5.661882,6.300045,6.9382076,5.7597823,4.5831695,3.4047437,2.228131,1.0497054,1.0551442,1.0605831,1.064209,1.0696479,1.0750868,1.1059072,1.1349145,1.1657349,1.1947423,1.2255627,0.9808127,0.73424983,0.4894999,0.24474995,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.62184614,1.2074331,1.79302,2.3767939,2.962381,4.1897564,5.4171324,6.644508,7.8718834,9.099259,9.180842,9.2606125,9.340384,9.420154,9.499924,8.548119,7.5945,6.642695,5.6908894,4.7372713,5.1923246,5.6473784,6.1024323,6.5574856,7.0125394,7.6180687,8.221786,8.827314,9.432844,10.038374,10.357455,10.6783495,10.997431,11.318325,11.637406,10.634838,9.63227,8.629702,7.6271334,6.624565,6.7043357,6.784106,6.8656893,6.94546,7.02523,6.5592985,6.09518,5.6292486,5.1651306,4.699199,4.420003,4.1408067,3.8597972,3.5806012,3.299592,3.4319382,3.5642843,3.6966307,3.83079,3.9631362,4.5650396,5.1669436,5.77066,6.3725634,6.9744673,6.5574856,6.1405044,5.7217097,5.3047285,4.8877473,6.1205616,7.3515635,8.584378,9.817192,11.050007,10.58045,10.110892,9.639522,9.169965,8.700407,8.6333275,8.564435,8.497355,8.430276,8.363196,8.02236,7.6833353,7.3424983,7.0016613,6.6626377,7.8156815,8.966913,10.119957,11.273002,12.4242325,10.959359,9.494485,8.029612,6.5647373,5.0998635,6.7442207,8.39039,10.034748,11.680918,13.325275,12.91192,12.500377,12.087022,11.675479,11.262123,12.585587,13.907236,15.230699,16.55235,17.87581,16.764465,15.654932,14.545399,13.435865,12.32452,13.635292,14.94425,16.255022,17.565794,18.874754,18.417887,17.959208,17.50234,17.045475,16.586794,14.104849,11.622903,9.139144,6.6571984,4.175253,4.313038,4.4508233,4.5867953,4.7245803,4.8623657,6.0407915,7.217404,8.39583,9.572442,10.750868,11.57214,12.395226,13.21831,14.039582,14.862667,15.564283,16.267714,16.96933,17.67276,18.374376,17.602055,16.829731,16.05741,15.285088,14.512766,16.14987,17.786976,19.425894,21.063,22.700104,22.411844,22.125395,21.837133,21.550686,21.262424,20.036863,18.813112,17.58755,16.361988,15.138238,15.636803,16.13718,16.637558,17.137936,17.638313,17.80692,17.977337,18.147755,18.318174,18.48678,17.747091,17.007402,16.267714,15.528025,14.788336,15.343102,15.897869,16.452635,17.007402,17.562168,16.501585,15.442815,14.382232,13.321649,12.262879,13.069647,13.878228,14.684997,15.491765,16.300346,15.945006,15.589665,15.234324,14.880796,14.525456,12.389787,10.255929,8.120259,5.9845896,3.8507326,4.0302157,4.209699,4.3891826,4.5704784,4.749962,5.3627434,5.975525,6.588306,7.1992745,7.8120556,8.52455,9.237044,9.949538,10.662033,11.374527,11.909351,12.444175,12.980812,13.515636,14.05046,15.410182,16.769903,18.129625,19.489347,20.850883,20.129324,19.409578,18.68983,17.970085,17.25034,16.004833,14.759329,13.515636,12.270131,11.024626,10.428161,9.829884,9.231606,8.63514,8.036863,8.009668,7.9824743,7.95528,7.9280853,7.900891,7.85738,7.8156815,7.7721705,7.7304726,7.686961,7.5781837,7.4675927,7.3570023,7.2482243,7.137634,7.476658,7.817495,8.158332,8.497355,8.838193,9.3567,9.87702,10.397341,10.917661,11.437981,12.685299,13.932617,15.179935,16.427254,17.674572,17.68545,17.694515,17.705393,17.714457,17.725336,17.355492,16.985647,16.615803,16.244144,15.8743,15.850732,15.825351,15.799969,15.774588,15.749206,16.789846,17.830486,18.869314,19.909956,20.950596,21.942286,22.93579,23.92748,24.91917,25.912674,25.551895,25.192928,24.832148,24.473183,24.112402,25.5247,26.936998,28.349297,29.761593,31.175705,29.5948,28.01571,26.434807,24.855717,23.274813,24.099712,24.92461,25.749508,26.574406,27.399303,28.940321,30.479527,32.020546,33.55975,35.10077,33.52712,31.955278,30.381626,28.809788,27.23795,27.419247,27.602356,27.785465,27.96676,28.14987,26.481945,24.814018,23.147905,21.47998,19.812056,20.778364,21.74286,22.707355,23.671852,24.63816,25.767637,26.897114,28.028402,29.157877,30.287354,29.529535,28.771717,28.01571,27.257893,26.500074,0.9119202,1.2654479,1.6171626,1.9706904,2.322405,2.6741197,3.0983531,3.5207734,3.9431937,4.365614,4.788034,5.6093063,6.432391,7.2554765,8.076748,8.899834,10.388275,11.874905,13.363347,14.849977,16.336605,16.213324,16.08823,15.963136,15.838041,15.712947,14.142921,12.572895,11.00287,9.432844,7.8628187,7.699652,7.5382986,7.3751316,7.211965,7.0506115,6.155008,5.2594047,4.365614,3.4700103,2.5744069,2.907992,3.2397642,3.5733492,3.9051213,4.2368937,4.115425,3.9921436,3.870675,3.7473936,3.6241121,4.882308,6.1405044,7.3968873,8.655084,9.91328,10.627586,11.341894,12.058014,12.772322,13.486629,12.462305,11.437981,10.411844,9.38752,8.363196,9.262425,10.161655,11.062697,11.961927,12.862969,11.289318,9.71748,8.145641,6.5719895,5.0001507,5.3246713,5.6491914,5.975525,6.300045,6.624565,6.622752,6.6191263,6.6173134,6.6155005,6.6118746,6.4432693,6.2728505,6.1024323,5.9320135,5.763408,5.6093063,5.4570174,5.3047285,5.1524396,5.0001507,4.3982472,3.7945306,3.1926272,2.5907235,1.987007,3.5080826,5.027345,6.548421,8.067683,9.5869465,8.781991,7.9770355,7.17208,6.3671246,5.562169,6.684393,7.806617,8.930654,10.052877,11.175101,11.144281,11.115273,11.084454,11.055446,11.024626,11.133403,11.240368,11.347333,11.454298,11.563075,12.460492,13.357908,14.255324,15.152741,16.050158,14.237195,12.4242325,10.613083,8.80012,6.987158,7.1883965,7.3878226,7.5872483,7.7866745,7.987913,8.714911,9.441909,10.17072,10.897718,11.624716,11.008308,10.390089,9.771869,9.155461,8.537241,7.900891,7.262728,6.624565,5.9882154,5.3500524,6.794984,8.239915,9.684846,11.129777,12.574709,13.383289,14.190058,14.996826,15.805408,16.612177,16.385555,16.157122,15.930502,15.702069,15.475449,15.159993,14.844538,14.530895,14.21544,13.899984,13.852847,13.80571,13.75676,13.709623,13.662486,12.804955,11.947423,11.089892,10.232361,9.374829,9.750113,10.125396,10.500679,10.874149,11.249433,11.173288,11.095331,11.017374,10.939416,10.863272,11.9021,12.9427395,13.98338,15.022208,16.062849,15.020395,13.9779415,12.935488,11.893035,10.850581,10.362894,9.875207,9.38752,8.899834,8.412147,8.62245,8.832754,9.043057,9.253361,9.461852,10.049252,10.636651,11.225864,11.813264,12.400664,12.302764,12.2048645,12.106964,12.010877,11.912977,13.80571,15.6966305,17.589363,19.482096,21.374828,22.607643,23.840458,25.073273,26.304274,27.537088,25.762197,23.987309,22.212418,20.437527,18.662638,18.49947,18.338116,18.17495,18.011784,17.85043,18.051668,18.25472,18.457771,18.660824,18.862062,16.815228,14.7683935,12.719746,10.672911,8.624263,9.425592,10.225109,11.024626,11.8241415,12.625471,12.989877,13.354282,13.720501,14.084907,14.449312,12.039885,9.630457,7.219217,4.8097897,2.4003625,2.0268922,1.6552348,1.2817645,0.9101072,0.53663695,0.42967212,0.32270733,0.21574254,0.10696479,0.0,0.5275721,1.0551442,1.5827163,2.1102884,2.6378605,3.2125697,3.787279,4.361988,4.936697,5.5132194,4.6230545,3.73289,2.8427253,1.9525607,1.062396,1.6171626,2.1719291,2.7266958,3.2832751,3.8380418,4.070101,4.3021603,4.5342193,4.7680917,5.0001507,5.8504305,6.70071,7.549176,8.399456,9.249735,7.6416373,6.035352,4.4272547,2.819157,1.2128719,1.0768998,0.94274056,0.80676836,0.6726091,0.53663695,0.5529536,0.56745726,0.581961,0.5982776,0.61278135,0.4894999,0.3680314,0.24474995,0.12328146,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.81764615,1.5845293,2.3532255,3.1201086,3.8869917,5.3953767,6.9019485,8.410334,9.916905,11.42529,11.439794,11.454298,11.470614,11.485118,11.499621,10.455356,9.409276,8.365009,7.320743,6.2746634,6.7641635,7.2554765,7.744976,8.234476,8.725789,9.4781685,10.230548,10.982927,11.735307,12.487686,12.7233715,12.957244,13.192928,13.426801,13.662486,12.304577,10.946668,9.590572,8.232663,6.874754,7.0016613,7.130382,7.2572894,7.3841968,7.512917,6.867502,6.2220874,5.576673,4.933071,4.2876563,3.9975824,3.7075086,3.4174345,3.1273603,2.8372865,3.2216346,3.6077955,3.9921436,4.3783045,4.762653,5.569421,6.378002,7.1847706,7.993352,8.80012,8.334189,7.8700705,7.404139,6.9400206,6.474089,7.5981264,8.72035,9.842574,10.964798,12.087022,11.702674,11.318325,10.932164,10.547816,10.161655,10.098202,10.032935,9.967669,9.902402,9.837135,9.5053625,9.171778,8.840006,8.508233,8.174648,8.820063,9.465478,10.110892,10.754494,11.399909,10.330261,9.2606125,8.189152,7.119504,6.049856,6.8094873,7.569119,8.330563,9.090195,9.849826,9.824444,9.800876,9.775495,9.750113,9.724731,10.705544,11.684544,12.665357,13.644357,14.625169,14.106662,13.589968,13.073273,12.554766,12.038072,13.780329,15.522586,17.264843,19.0071,20.749357,18.503096,16.255022,14.006948,11.760688,9.512614,8.540867,7.567306,6.5955577,5.621997,4.650249,4.5867953,4.5251546,4.461701,4.40006,4.3366065,5.520471,6.7025228,7.8845744,9.066626,10.25049,11.205922,12.15954,13.114971,14.070402,15.025834,15.607795,16.189756,16.771717,17.355492,17.937452,17.18326,16.427254,15.673061,14.917056,14.162864,15.687565,17.212267,18.736969,20.26167,21.788185,21.063,20.337814,19.612629,18.887444,18.16226,16.962078,15.761897,14.561715,13.363347,12.163166,12.60009,13.037014,13.475751,13.912675,14.349599,14.559902,14.770206,14.98051,15.190813,15.399304,14.855415,14.309713,13.765825,13.220123,12.674421,13.502945,14.329657,15.15818,15.984891,16.811602,15.4827,14.151986,12.823084,11.49237,10.161655,11.510499,12.857531,14.204562,15.553406,16.900436,16.472578,16.04472,15.616859,15.190813,14.762955,12.469557,10.177972,7.8845744,5.5929894,3.299592,3.6893787,4.079166,4.4707656,4.860553,5.2503395,5.825049,6.399758,6.9744673,7.549176,8.125698,8.537241,8.950596,9.362139,9.775495,10.1870365,10.968424,11.747997,12.527572,13.307145,14.0867195,15.818098,17.547665,19.277231,21.006798,22.738176,22.21423,21.692097,21.169964,20.647831,20.125698,18.677141,17.230396,15.781839,14.335095,12.888351,12.019942,11.153346,10.284937,9.418341,8.549932,8.417585,8.285239,8.152893,8.020547,7.8882003,7.610817,7.3316207,7.0542374,6.776854,6.4994707,6.2692246,6.0407915,5.810545,5.580299,5.3500524,6.0824895,6.814926,7.5473633,8.2798,9.012237,9.710228,10.408218,11.104396,11.802386,12.500377,13.642544,14.78471,15.926876,17.069042,18.213022,18.193079,18.173138,18.153194,18.133251,18.11331,17.864933,17.61837,17.369995,17.121618,16.875055,16.836983,16.800724,16.762651,16.72458,16.68832,17.819609,18.952711,20.085812,21.217102,22.350203,23.390842,24.42967,25.470312,26.509138,27.54978,27.633175,27.71476,27.798155,27.879738,27.963135,29.237648,30.51216,31.786673,33.063,34.337513,32.13476,29.932013,27.729263,25.528326,23.325577,24.33721,25.350657,26.36229,27.375734,28.387367,29.919321,31.453089,32.985043,34.516994,36.050762,34.720047,33.38933,32.06043,30.729715,29.400814,29.910257,30.419699,30.929142,31.440397,31.949839,30.096992,28.244144,26.393108,24.540262,22.687414,23.882156,25.076899,26.27164,27.468197,28.66294,29.277533,29.892128,30.506721,31.123129,31.737722,30.278288,28.81704,27.357605,25.89817,24.436922,1.1258497,1.4866294,1.8492218,2.2118144,2.5744069,2.9369993,3.3249733,3.7129474,4.099108,4.4870825,4.8750563,5.8758116,6.874754,7.8755093,8.874452,9.875207,11.450671,13.024323,14.599788,16.175253,17.750717,17.725336,17.699953,17.674572,17.64919,17.625622,15.613234,13.600845,11.586644,9.574255,7.5618668,7.413204,7.262728,7.112252,6.9617763,6.813113,5.975525,5.137936,4.3003473,3.4627585,2.6251698,2.7992141,2.9750717,3.149116,3.3249733,3.5008307,2.9750717,2.4493124,1.9253663,1.3996071,0.87566096,2.5508385,4.2242026,5.89938,7.574558,9.249735,10.388275,11.525003,12.661731,13.800271,14.936998,13.662486,12.387974,11.111648,9.837135,8.562622,9.837135,11.111648,12.387974,13.662486,14.936998,12.92461,10.912222,8.899834,6.887445,4.8750563,5.049101,5.224958,5.4008155,5.57486,5.750717,5.638314,5.52591,5.411693,5.2992897,5.186886,4.9258194,4.6629395,4.40006,4.137181,3.874301,4.07554,4.274966,4.4743915,4.6756306,4.8750563,4.2368937,3.6005437,2.962381,2.324218,1.6878681,3.5008307,5.3119802,7.124943,8.937905,10.750868,9.762803,8.774739,7.7866745,6.8004227,5.812358,7.07418,8.337815,9.599637,10.863272,12.125093,12.087022,12.050762,12.012691,11.974618,11.938358,11.463363,10.988366,10.51337,10.038374,9.563377,10.51337,11.463363,12.413355,13.363347,14.313339,12.436923,10.56232,8.6877165,6.813113,4.936697,5.411693,5.8866897,6.3616858,6.836682,7.311678,8.450218,9.5869465,10.725487,11.862214,13.000754,12.163166,11.325577,10.487988,9.6504,8.812811,8.062244,7.311678,6.5629244,5.812358,5.0617914,6.736969,8.412147,10.087324,11.762501,13.437678,14.249886,15.062093,15.8743,16.68832,17.500528,17.26303,17.025532,16.788034,16.550535,16.313038,15.674874,15.036712,14.400362,13.762199,13.125849,13.424988,13.724127,14.025079,14.324218,14.625169,13.762199,12.899229,12.038072,11.175101,10.312131,10.312131,10.312131,10.312131,10.312131,10.312131,10.449916,10.587702,10.725487,10.863272,10.999244,11.974618,12.949992,13.925365,14.90074,15.8743,14.96238,14.05046,13.136727,12.224807,11.312886,10.88684,10.462607,10.038374,9.612328,9.188094,9.362139,9.537996,9.712041,9.8878975,10.061942,10.636651,11.213174,11.787883,12.362592,12.937301,12.786825,12.638163,12.487686,12.337211,12.186734,14.500074,16.811602,19.124943,21.438282,23.74981,25.412296,27.074783,28.73727,30.399757,32.062244,29.52591,26.98776,24.449614,21.913279,19.375132,19.288109,19.199274,19.112251,19.025229,18.938208,19.099562,19.262728,19.425894,19.587248,19.750414,17.437075,15.125546,12.812206,10.500679,8.187339,9.1500225,10.112705,11.075388,12.038072,13.000754,13.6244135,14.249886,14.875358,15.50083,16.124489,12.937301,9.750113,6.5629244,3.3757362,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.0,0.0,0.0,0.0,0.0,0.387974,0.774135,1.162109,1.550083,1.938057,2.8499773,3.7618973,4.6756306,5.5875506,6.4994707,5.199577,3.8996825,2.5997884,1.2998942,0.0,0.72518504,1.4503701,2.175555,2.9007401,3.6241121,4.1498713,4.6756306,5.199577,5.7253356,6.249282,7.311678,8.374074,9.438283,10.500679,11.563075,9.525306,7.4875355,5.4497657,3.4119956,1.3742256,1.1004683,0.824898,0.5493277,0.2755703,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,1.0134461,1.9616255,2.913431,3.8616104,4.8116026,6.600997,8.386765,10.174346,11.961927,13.749508,13.700559,13.649796,13.600845,13.550082,13.499319,12.362592,11.225864,10.087324,8.950596,7.8120556,8.337815,8.861761,9.38752,9.91328,10.437225,11.338268,12.237497,13.136727,14.037769,14.936998,15.087475,15.23795,15.386614,15.537089,15.687565,13.974316,12.262879,10.549629,8.838193,7.124943,7.3008003,7.474845,7.650702,7.8247466,8.000604,7.175706,6.350808,5.524097,4.699199,3.874301,3.5751622,3.2742105,2.9750717,2.6741197,2.374981,3.0131438,3.6494937,4.2876563,4.9258194,5.562169,6.5756154,7.5872483,8.600695,9.612328,10.625773,10.112705,9.599637,9.088382,8.575313,8.062244,9.07569,10.087324,11.10077,12.112403,13.125849,12.824898,12.525759,12.224807,11.925668,11.624716,11.563075,11.499621,11.437981,11.374527,11.312886,10.988366,10.662033,10.337513,10.012992,9.686659,9.824444,9.96223,10.100015,10.2378,10.375585,9.699349,9.024928,8.350506,7.6742706,6.9998484,6.874754,6.7496595,6.624565,6.4994707,6.3743763,6.736969,7.0995617,7.462154,7.8247466,8.187339,8.825501,9.461852,10.100015,10.738177,11.374527,11.450671,11.525003,11.599335,11.675479,11.74981,13.925365,16.099108,18.274662,20.450218,22.625772,18.586493,14.5508375,10.511557,6.474089,2.4366217,2.9750717,3.5117085,4.0501585,4.5867953,5.125245,4.8623657,4.599486,4.3366065,4.07554,3.8126602,5.0001507,6.187641,7.3751316,8.562622,9.750113,10.837891,11.925668,13.011633,14.09941,15.187187,15.649493,16.1118,16.575916,17.038223,17.500528,16.762651,16.024776,15.2869005,14.5508375,13.812962,15.22526,16.637558,18.049856,19.462152,20.87445,19.712341,18.550234,17.388124,16.224201,15.062093,13.887294,12.712494,11.537694,10.362894,9.188094,9.563377,9.936848,10.312131,10.687414,11.062697,11.312886,11.563075,11.813264,12.06164,12.311829,11.961927,11.612025,11.262123,10.912222,10.56232,11.662788,12.763257,13.861912,14.96238,16.062849,14.462003,12.862969,11.262123,9.663091,8.062244,9.949538,11.836833,13.72594,15.613234,17.500528,17.00015,16.499773,15.999394,15.50083,15.000452,12.549327,10.100015,7.650702,5.199577,2.7502642,3.350355,3.9504454,4.550536,5.1506267,5.750717,6.2873545,6.825804,7.362441,7.900891,8.437528,8.549932,8.662335,8.774739,8.887142,8.999546,10.025683,11.050007,12.07433,13.100468,14.124791,16.226015,18.325426,20.424837,22.524246,24.625471,24.299137,23.974617,23.650097,23.325577,22.999243,21.349447,19.699652,18.049856,16.400059,14.750263,13.611723,12.474996,11.338268,10.199727,9.063,8.825501,8.588004,8.350506,8.113008,7.8755093,7.362441,6.849373,6.338117,5.825049,5.3119802,4.9620786,4.612177,4.262275,3.9123733,3.5624714,4.688321,5.812358,6.9382076,8.062244,9.188094,10.061942,10.937603,11.813264,12.687112,13.562773,14.599788,15.636803,16.67563,17.712645,18.749659,18.700708,18.649946,18.599184,18.550234,18.49947,18.374376,18.24928,18.124187,18.000906,17.87581,17.825048,17.774284,17.725336,17.674572,17.625622,18.849373,20.074934,21.300497,22.524246,23.74981,24.837587,25.925365,27.013142,28.099108,29.186884,29.712645,30.238403,30.762348,31.288109,31.812054,32.950596,34.087322,35.225864,36.36259,37.499317,34.67472,31.850126,29.025532,26.200935,23.374527,24.574707,25.774889,26.97507,28.175251,29.375433,30.900135,32.424835,33.94954,35.47424,37.00075,35.912975,34.8252,33.73742,32.649643,31.561865,32.399456,33.23704,34.07463,34.91222,35.74981,33.71204,31.674269,29.638311,27.600542,25.562773,26.98776,28.41275,29.837738,31.262726,32.687714,32.78743,32.887142,32.986855,33.08838,33.18809,31.025229,28.862364,26.6995,24.538448,22.375584,1.6371052,2.077655,2.518205,2.956942,3.397492,3.8380418,4.3547363,4.8732433,5.389938,5.906632,6.4251394,6.947273,7.4694057,7.993352,8.515485,9.037619,10.324821,11.612025,12.899229,14.188245,15.475449,15.616859,15.760084,15.903308,16.04472,16.187943,14.269829,12.351714,10.435412,8.517298,6.599184,6.4831543,6.3653116,6.247469,6.1296263,6.011784,5.375434,4.7372713,4.099108,3.4627585,2.8245957,2.9152439,3.005892,3.094727,3.1853752,3.2742105,3.000453,2.7248828,2.4493124,2.175555,1.8999848,3.2379513,4.574105,5.9120708,7.250037,8.588004,9.625018,10.662033,11.700861,12.737875,13.77489,12.694364,11.615651,10.535126,9.4546,8.375887,9.400211,10.424535,11.450671,12.474996,13.499319,11.7425585,9.985798,8.227224,6.4704633,4.7118897,4.9258194,5.137936,5.3500524,5.562169,5.774286,6.4251394,7.07418,7.7250338,8.375887,9.024928,8.138389,7.250037,6.3616858,5.475147,4.5867953,4.8496747,5.1125546,5.375434,5.638314,5.89938,5.6528172,5.4044414,5.1578784,4.9095025,4.6629395,5.957395,7.25185,8.548119,9.842574,11.137029,10.125396,9.11195,8.100317,7.0868707,6.0752378,7.159389,8.245354,9.329506,10.41547,11.499621,11.314699,11.129777,10.944855,10.7599325,10.57501,10.127209,9.679407,9.231606,8.785617,8.337815,9.092008,9.848013,10.602205,11.358211,12.112403,10.839704,9.567003,8.294304,7.021604,5.750717,6.01541,6.2801023,6.544795,6.8094873,7.07418,8.430276,9.784559,11.1406555,12.494938,13.849221,13.147605,12.444175,11.7425585,11.039129,10.337513,9.626831,8.917963,8.207282,7.4966,6.787732,8.537241,10.28675,12.038072,13.7875805,15.537089,16.164375,16.79166,17.420757,18.048042,18.675327,18.25472,17.834112,17.41532,16.99471,16.574104,15.903308,15.230699,14.558089,13.885481,13.212872,13.419549,13.628039,13.834718,14.043208,14.249886,13.53014,12.810393,12.090648,11.369088,10.649343,10.522435,10.395528,10.266808,10.139899,10.012992,10.087324,10.161655,10.2378,10.312131,10.388275,11.307447,12.22662,13.147605,14.066776,14.9877615,14.287958,13.588155,12.888351,12.186734,11.486931,11.019187,10.553255,10.085511,9.617766,9.1500225,9.421967,9.695724,9.967669,10.239613,10.51337,11.044568,11.5775795,12.11059,12.6417885,13.174799,13.125849,13.075087,13.024323,12.975373,12.92461,14.750263,16.574104,18.399757,20.22541,22.049252,23.398094,24.745127,26.092157,27.439188,28.788033,26.746637,24.707054,22.66747,20.627888,18.588305,18.347181,18.10787,17.866747,17.627436,17.388124,17.462456,17.536787,17.612932,17.687263,17.761595,16.050158,14.336908,12.625471,10.912222,9.200785,10.284937,11.369088,12.455053,13.539205,14.625169,14.342347,14.059525,13.776703,13.495693,13.212872,10.600392,7.987913,5.375434,2.762955,0.15047589,0.7705091,1.3905423,2.0105755,2.6306088,3.2506418,2.8282216,2.4058013,1.983381,1.5591478,1.1367276,1.3778516,1.6171626,1.8582866,2.0975976,2.3369088,3.009518,3.682127,4.3547363,5.027345,5.6999545,4.842423,3.9848917,3.1273603,2.269829,1.4122978,2.0522738,2.6922495,3.3322253,3.972201,4.612177,5.277534,5.942891,6.6082487,7.271793,7.93715,8.225411,8.511859,8.80012,9.088382,9.374829,7.7195945,6.0643597,4.409125,2.7557032,1.1004683,0.8792868,0.65991837,0.4405499,0.21936847,0.0,0.0,0.0,0.0,0.0,0.0,0.11421664,0.23024625,0.3444629,0.4604925,0.5747091,0.6979906,0.8194591,0.94274056,1.064209,1.1874905,2.0504606,2.911618,3.774588,4.6375585,5.5005283,6.892884,8.285239,9.677594,11.069949,12.462305,12.578335,12.692551,12.806767,12.922797,13.037014,12.07433,11.111648,10.150778,9.188094,8.225411,8.894395,9.56519,10.234174,10.90497,11.575767,12.444175,13.314397,14.184619,15.054841,15.925063,15.957697,15.99033,16.022963,16.055597,16.08823,14.6052265,13.122223,11.63922,10.15803,8.675026,8.537241,8.399456,8.26167,8.125698,7.987913,7.3316207,6.677141,6.0226617,5.368182,4.7118897,4.409125,4.1081734,3.8054085,3.5026438,3.199879,4.004834,4.8097897,5.614745,6.4197006,7.224656,8.01692,8.809185,9.603263,10.395528,11.187792,10.607644,10.027496,9.447348,8.8672,8.287052,9.2606125,10.232361,11.205922,12.17767,13.149418,12.66717,12.184921,11.702674,11.220426,10.738177,11.142468,11.546759,11.952863,12.357153,12.763257,13.589968,14.416678,15.245202,16.071913,16.900436,16.135366,15.3702965,14.6052265,13.840157,13.075087,11.889409,10.705544,9.519867,8.334189,7.1503243,7.0941224,7.039734,6.985345,6.929143,6.874754,7.264541,7.654328,8.044115,8.435715,8.825501,9.255174,9.684846,10.114518,10.54419,10.975676,11.222239,11.470614,11.717177,11.965553,12.212116,13.747695,15.283275,16.817041,18.352621,19.888199,16.313038,12.737875,9.162713,5.5875506,2.0123885,2.4547513,2.8971143,3.339477,3.7818398,4.2242026,4.360175,4.494334,4.6303062,4.764466,4.900438,5.89938,6.9001355,7.900891,8.899834,9.900589,11.10077,12.299138,13.499319,14.699501,15.899682,16.075539,16.249584,16.425442,16.599485,16.775343,16.017525,15.2597065,14.501887,13.745882,12.988064,14.026892,15.067532,16.108173,17.147,18.187641,17.101677,16.017525,14.93156,13.847408,12.763257,11.925668,11.088079,10.25049,9.412902,8.575313,9.015862,9.4546,9.89515,10.3357,10.774437,11.011934,11.249433,11.486931,11.724429,11.961927,11.519565,11.077202,10.634838,10.192475,9.750113,10.700105,11.650098,12.60009,13.550082,14.500074,13.410484,12.320893,11.22949,10.139899,9.050309,10.424535,11.800573,13.174799,14.5508375,15.925063,15.382988,14.840912,14.297023,13.754947,13.212872,11.234929,9.256987,7.2790446,5.3029156,3.3249733,4.220577,5.1143675,6.009971,6.9055743,7.799365,7.8102427,7.819308,7.8301854,7.83925,7.850128,7.9770355,8.105756,8.232663,8.3595705,8.488291,9.354887,10.223296,11.089892,11.958302,12.824898,14.597975,16.36924,18.142317,19.915394,21.686659,21.487232,21.287807,21.08838,20.887142,20.687716,19.342497,17.99728,16.652061,15.306843,13.961625,12.935488,11.907538,10.879588,9.853452,8.825501,8.419398,8.015107,7.610817,7.2047133,6.8004227,6.5176005,6.2347784,5.9519563,5.669134,5.388125,5.3428006,5.297477,5.2521524,5.2068286,5.163317,6.1241875,7.0868707,8.049554,9.012237,9.97492,10.845142,11.715364,12.585587,13.455809,14.324218,15.602356,16.880495,18.15682,19.43496,20.713097,20.707659,20.702219,20.696781,20.693155,20.687716,20.386765,20.087626,19.786674,19.487535,19.188396,19.308052,19.427708,19.547363,19.667019,19.786674,20.963285,22.138086,23.312885,24.487686,25.662485,26.329655,26.996826,27.66581,28.33298,29.000149,29.250338,29.500526,29.750715,29.999092,30.24928,31.645262,33.03943,34.43541,35.82958,37.22556,34.82157,32.419395,30.017221,27.615046,25.212872,25.675177,26.137482,26.599787,27.062092,27.524399,28.802536,30.080675,31.357,32.63514,33.913277,33.059372,32.20728,31.355188,30.503096,29.64919,29.92476,30.20033,30.4759,30.749659,31.025229,29.66188,28.300346,26.936998,25.575462,24.212114,26.264389,28.318476,30.370749,32.423023,34.475296,34.089134,33.70479,33.32044,32.934277,32.54993,30.793169,29.034595,27.277836,25.51926,23.7625,2.1501737,2.666868,3.1853752,3.7020695,4.220577,4.7372713,5.384499,6.0317264,6.680767,7.327995,7.9752226,8.020547,8.06587,8.109382,8.154706,8.200029,9.200785,10.199727,11.200482,12.199425,13.200181,13.510198,13.820213,14.13023,14.440247,14.750263,12.928236,11.104396,9.282369,7.460341,5.638314,5.5531044,5.467895,5.382686,5.297477,5.2122674,4.7753434,4.3384194,3.8996825,3.4627585,3.0258346,3.0294604,3.0348995,3.0403383,3.045777,3.049403,3.0258346,3.000453,2.9750717,2.94969,2.9243085,3.925064,4.9258194,5.924762,6.925517,7.9244595,8.861761,9.800876,10.738177,11.675479,12.612781,11.728055,10.843329,9.956791,9.072064,8.187339,8.963287,9.737422,10.51337,11.287505,12.06164,10.560507,9.057561,7.554615,6.051669,4.550536,4.800725,5.049101,5.2992897,5.5494785,5.7996674,7.211965,8.624263,10.038374,11.450671,12.862969,11.349146,9.837135,8.325124,6.813113,5.2992897,5.6256227,5.9501433,6.2746634,6.599184,6.925517,7.066928,7.210152,7.3533764,7.494787,7.6380115,8.415772,9.19172,9.969481,10.747242,11.525003,10.487988,9.449161,8.412147,7.3751316,6.338117,7.2445984,8.152893,9.059374,9.967669,10.874149,10.542377,10.210606,9.87702,9.545248,9.211663,8.792869,8.372261,7.951654,7.5328593,7.112252,7.6724577,8.232663,8.792869,9.353074,9.91328,9.242483,8.571687,7.902704,7.231908,6.5629244,6.6173134,6.6717024,6.7279043,6.782293,6.836682,8.410334,9.982172,11.555823,13.127662,14.699501,14.132043,13.564586,12.9971285,12.429671,11.862214,11.193231,10.522435,9.851639,9.182655,8.511859,10.337513,12.163166,13.987006,15.812659,17.638313,18.080675,18.523039,18.9654,19.407764,19.850128,19.248224,18.644506,18.042604,17.4407,16.836983,16.129929,15.422873,14.715817,14.006948,13.299893,13.41411,13.53014,13.644357,13.760386,13.874602,13.29808,12.719746,12.143224,11.564888,10.988366,10.7327385,10.477111,10.223296,9.967669,9.712041,9.724731,9.737422,9.750113,9.762803,9.775495,10.640278,11.50506,12.3698435,13.234627,14.09941,13.611723,13.125849,12.638163,12.1504755,11.662788,11.153346,10.642091,10.1326475,9.623205,9.11195,9.481794,9.851639,10.223296,10.593141,10.962985,11.452485,11.941984,12.433297,12.922797,13.412297,13.46306,13.512011,13.562773,13.611723,13.662486,15.000452,16.336605,17.674572,19.012539,20.350506,21.38208,22.41547,23.447044,24.480434,25.512009,23.96918,22.42816,20.885328,19.342497,17.799667,17.408066,17.014654,16.623055,16.229641,15.838041,15.825351,15.812659,15.799969,15.787278,15.774588,14.663241,13.550082,12.436923,11.325577,10.212419,11.419851,12.627284,13.834718,15.0421505,16.249584,15.06028,13.8691635,12.67986,11.490557,10.29944,8.26167,6.2257137,4.1879435,2.1501737,0.11240368,1.3905423,2.666868,3.9450066,5.223145,6.4994707,5.65463,4.8097897,3.9649491,3.1201086,2.275268,2.3677292,2.4601903,2.5526514,2.6451125,2.7375734,3.1708715,3.6023567,4.0356545,4.4671397,4.900438,4.4852695,4.070101,3.6549325,3.2397642,2.8245957,3.3793623,3.9341288,4.4907084,5.045475,5.600241,6.4051967,7.210152,8.015107,8.820063,9.625018,9.137331,8.649645,8.161958,7.6742706,7.1883965,5.915697,4.6429973,3.3702974,2.0975976,0.824898,0.65991837,0.4949388,0.32995918,0.16497959,0.0,0.0,0.0,0.0,0.0,0.0,0.23024625,0.4604925,0.69073874,0.91917205,1.1494182,1.3832904,1.6153497,1.8474089,2.079468,2.3133402,3.0874753,3.8616104,4.6375585,5.411693,6.187641,7.1847706,8.1819,9.180842,10.177972,11.175101,11.454298,11.735307,12.0145035,12.295512,12.574709,11.787883,10.999244,10.212419,9.425592,8.636953,9.452786,10.266808,11.082641,11.896661,12.712494,13.551895,14.39311,15.2325115,16.071913,16.913128,16.827919,16.74271,16.6575,16.57229,16.487082,15.234324,13.98338,12.730623,11.477866,10.225109,9.775495,9.325879,8.874452,8.424837,7.9752226,7.4893484,7.0052876,6.5194135,6.035352,5.5494785,5.2449007,4.940323,4.6357455,4.329355,4.024777,4.9983377,5.9700856,6.9418335,7.915395,8.887142,9.460039,10.032935,10.605831,11.176914,11.74981,11.102583,10.455356,9.808127,9.159087,8.511859,9.445535,10.377398,11.30926,12.242936,13.174799,12.509441,11.845898,11.18054,10.515183,9.849826,10.721861,11.595709,12.467744,13.339779,14.211814,16.193382,18.173138,20.152891,22.132647,24.112402,22.444477,20.778364,19.11044,17.442513,15.774588,14.079468,12.384347,10.689227,8.994107,7.3008003,7.315304,7.3298078,7.344311,7.360628,7.3751316,7.7921133,8.209095,8.627889,9.04487,9.461852,9.684846,9.907841,10.130835,10.352016,10.57501,10.995618,11.4144125,11.83502,12.255627,12.674421,13.5700245,14.465629,15.359419,16.255022,17.150625,14.037769,10.924912,7.8120556,4.699199,1.5881553,1.9344311,2.2825198,2.6306088,2.9768846,3.3249733,3.8579843,4.3891826,4.9221935,5.4552045,5.9882154,6.8004227,7.61263,8.424837,9.237044,10.049252,11.361836,12.674421,13.987006,15.299591,16.612177,16.499773,16.38737,16.274965,16.162561,16.050158,15.272397,14.494636,13.716875,12.939114,12.163166,12.830337,13.497506,14.164677,14.831847,15.50083,14.492823,13.484816,12.476809,11.470614,10.462607,9.96223,9.461852,8.963287,8.46291,7.9625316,8.4683485,8.972352,9.4781685,9.982172,10.487988,10.712796,10.937603,11.162411,11.3872175,11.612025,11.077202,10.542377,10.007553,9.47273,8.937905,9.737422,10.536939,11.338268,12.137785,12.937301,12.357153,11.777005,11.1968565,10.616709,10.038374,10.899531,11.762501,12.625471,13.486629,14.349599,13.765825,13.180238,12.594651,12.010877,11.42529,9.920531,8.415772,6.9092,5.4044414,3.8996825,5.090799,6.2801023,7.4694057,8.660522,9.849826,9.333132,8.814624,8.29793,7.7794223,7.262728,7.404139,7.5473633,7.690587,7.8319983,7.9752226,8.685904,9.394773,10.1054535,10.8143215,11.525003,12.969934,14.4148655,15.859797,17.304728,18.749659,18.675327,18.599184,18.52485,18.45052,18.374376,17.335548,16.294909,15.254267,14.21544,13.174799,12.25744,11.340081,10.422722,9.5053625,8.588004,8.015107,7.4422116,6.869315,6.298232,5.7253356,5.67276,5.620184,5.567608,5.5150323,5.462456,5.7217097,5.9827766,6.24203,6.5030966,6.7623506,7.5618668,8.363196,9.162713,9.96223,10.761745,11.628342,12.493125,13.357908,14.222692,15.087475,16.604925,18.122374,19.639824,21.157274,22.674723,22.71461,22.754494,22.794378,22.834263,22.87415,22.399153,21.924156,21.44916,20.974165,20.499168,20.789242,21.079315,21.36939,21.659464,21.949537,23.075388,24.199425,25.325274,26.44931,27.575161,27.821724,28.070099,28.316662,28.565039,28.811602,28.788033,28.762651,28.73727,28.71189,28.68832,30.33993,31.993351,33.64496,35.29657,36.94999,34.970234,32.99048,31.010725,29.03097,27.049402,26.775644,26.500074,26.224504,25.950747,25.675177,26.704939,27.734701,28.764463,29.794228,30.825802,30.207582,29.589363,28.972956,28.354734,27.738327,27.450066,27.161806,26.875357,26.587097,26.300648,25.611723,24.92461,24.237497,23.550385,22.863272,25.54283,28.22239,30.901947,33.581505,36.26288,35.392654,34.522434,33.65221,32.78199,31.911768,30.559298,29.206827,27.854357,26.501886,25.149418,2.663242,3.2578938,3.8525455,4.4471974,5.041849,5.638314,6.414262,7.192023,7.9697833,8.747544,9.525306,9.092008,8.660522,8.227224,7.795739,7.362441,8.074935,8.78743,9.499924,10.212419,10.924912,11.401722,11.880343,12.357153,12.835775,13.312584,11.584831,9.857078,8.129324,6.401571,4.6756306,4.6230545,4.5704784,4.517903,4.465327,4.4127507,4.175253,3.9377546,3.7002566,3.4627585,3.2252605,3.1454902,3.0657198,2.9841363,2.904366,2.8245957,3.049403,3.2742105,3.5008307,3.7256382,3.9504454,4.612177,5.275721,5.9374523,6.599184,7.262728,8.100317,8.937905,9.775495,10.613083,11.450671,10.7599325,10.069194,9.380268,8.689529,8.000604,8.52455,9.050309,9.574255,10.100015,10.625773,9.376642,8.129324,6.882006,5.634688,4.3873696,4.6756306,4.9620786,5.2503395,5.5367875,5.825049,8.000604,10.174346,12.349901,14.525456,16.699198,14.561715,12.4242325,10.28675,8.149267,6.011784,6.399758,6.787732,7.175706,7.5618668,7.949841,8.482852,9.015862,9.547061,10.080072,10.613083,10.872336,11.13159,11.392657,11.651911,11.912977,10.850581,9.788185,8.725789,7.66158,6.599184,7.3298078,8.0604315,8.789243,9.519867,10.25049,9.770056,9.28962,8.809185,8.330563,7.850128,7.456715,7.065115,6.6717024,6.2801023,5.8866897,6.2529078,6.6173134,6.981719,7.3479376,7.7123427,7.645263,7.5781837,7.509291,7.4422116,7.3751316,7.219217,7.065115,6.9092,6.755099,6.599184,8.39039,10.179785,11.969179,13.760386,15.54978,15.118295,14.684997,14.2516985,13.820213,13.386916,12.757817,12.126906,11.497808,10.866898,10.2378,12.137785,14.037769,15.937754,17.837738,19.737724,19.995165,20.252605,20.510046,20.767487,21.024927,20.239914,19.4549,18.66989,17.884876,17.099863,16.358362,15.6150465,14.871732,14.13023,13.386916,13.410484,13.43224,13.455809,13.477564,13.499319,13.064208,12.63091,12.195799,11.760688,11.325577,10.943042,10.560507,10.177972,9.795437,9.412902,9.362139,9.313189,9.262425,9.211663,9.162713,9.973107,10.781689,11.592083,12.402477,13.212872,12.937301,12.661731,12.387974,12.112403,11.836833,11.285692,10.7327385,10.179785,9.626831,9.07569,9.541622,10.009366,10.477111,10.944855,11.4126,11.860401,12.308203,12.754191,13.201994,13.649796,13.800271,13.9507475,14.09941,14.249886,14.400362,15.250641,16.099108,16.949387,17.799667,18.649946,19.36788,20.085812,20.801933,21.519865,22.237799,21.19172,20.147453,19.103188,18.057108,17.01284,16.467138,15.92325,15.377548,14.831847,14.287958,14.188245,14.0867195,13.987006,13.887294,13.7875805,13.274512,12.763257,12.250188,11.73712,11.225864,12.554766,13.885481,15.214382,16.545097,17.87581,15.7782135,13.680615,11.583018,9.48542,7.3878226,5.924762,4.461701,3.000453,1.5373923,0.07433146,2.0105755,3.9450066,5.8794374,7.8156815,9.750113,8.482852,7.215591,5.9483304,4.6792564,3.4119956,3.3576066,3.303218,3.247016,3.1926272,3.1382382,3.3304121,3.5225863,3.7147603,3.9069343,4.099108,4.1281157,4.15531,4.1825047,4.209699,4.2368937,4.708264,5.177821,5.6473784,6.1169357,6.588306,7.5328593,8.477413,9.421967,10.368333,11.312886,10.049252,8.78743,7.5256076,6.261973,5.0001507,4.1099863,3.2198215,2.3296568,1.4394923,0.5493277,0.4405499,0.32995918,0.21936847,0.11059072,0.0,0.0,0.0,0.0,0.0,0.0,0.3444629,0.69073874,1.0352017,1.3796645,1.7241274,2.0667772,2.4094272,2.752077,3.094727,3.437377,4.12449,4.8116026,5.5005283,6.187641,6.874754,7.476658,8.080374,8.682278,9.284182,9.8878975,10.332074,10.778063,11.222239,11.668227,12.112403,11.499621,10.88684,10.275872,9.663091,9.050309,10.009366,10.970237,11.929294,12.890164,13.849221,14.6596155,15.47001,16.280403,17.090797,17.89938,17.698141,17.495089,17.292038,17.090797,16.887747,15.865235,14.842725,13.820213,12.797703,11.775192,11.011934,10.25049,9.487233,8.725789,7.9625316,7.647076,7.3316207,7.017978,6.7025228,6.3870673,6.0806766,5.772473,5.464269,5.1578784,4.8496747,5.9900284,7.130382,8.270736,9.409276,10.549629,10.903157,11.254871,11.608399,11.9601145,12.311829,11.597522,10.883214,10.167094,9.452786,8.736667,9.630457,10.522435,11.4144125,12.308203,13.200181,12.351714,11.50506,10.656594,9.80994,8.963287,10.303066,11.642846,12.982625,14.322405,15.662184,18.794983,21.927782,25.060581,28.19338,31.324368,28.7554,26.184618,23.61565,21.04487,18.475903,16.269526,14.064963,11.860401,9.655839,7.4494634,7.5346723,7.6198816,7.705091,7.7903004,7.8755093,8.319685,8.765674,9.20985,9.655839,10.100015,10.114518,10.130835,10.145339,10.1598425,10.174346,10.767185,11.3600235,11.952863,12.545701,13.136727,13.392355,13.647983,13.901797,14.157425,14.413053,11.762501,9.11195,6.4632115,3.8126602,1.162109,1.4141108,1.6679256,1.9199274,2.1719291,2.4257438,3.3557937,4.2858434,5.2158933,6.14413,7.07418,7.699652,8.325124,8.950596,9.574255,10.199727,11.624716,13.049705,14.474693,15.899682,17.32467,16.92582,16.525154,16.124489,15.725637,15.324973,14.527269,13.729566,12.931862,12.134158,11.338268,11.631968,11.927481,12.222994,12.516694,12.812206,11.882156,10.952107,10.022058,9.092008,8.161958,8.000604,7.837437,7.6742706,7.512917,7.3497505,7.9208336,8.490104,9.059374,9.630457,10.199727,10.411844,10.625773,10.837891,11.050007,11.262123,10.634838,10.007553,9.380268,8.752983,8.125698,8.774739,9.425592,10.074633,10.725487,11.374527,11.3056345,11.234929,11.164224,11.095331,11.024626,11.374527,11.724429,12.07433,12.4242325,12.774135,12.14685,11.519565,10.89228,10.264994,9.637709,8.604321,7.572745,6.539356,5.5077806,4.4743915,5.959208,7.4458375,8.930654,10.41547,11.900287,10.854207,9.80994,8.765674,7.7195945,6.6753283,6.833056,6.9907837,7.1466985,7.304426,7.462154,8.015107,8.568061,9.119202,9.672155,10.225109,11.341894,12.460492,13.577277,14.695875,15.812659,15.861609,15.912373,15.963136,16.012085,16.062849,15.326786,14.592536,13.858286,13.122223,12.387974,11.579392,10.772624,9.965856,9.157274,8.350506,7.610817,6.869315,6.1296263,5.389938,4.650249,4.8279195,5.0055895,5.18326,5.3591175,5.5367875,6.1024323,6.6680765,7.231908,7.797552,8.363196,8.999546,9.637709,10.275872,10.912222,11.5503845,12.409729,13.2690735,14.13023,14.989574,15.850732,17.607492,19.364254,21.122828,22.879587,24.63816,24.723372,24.806767,24.891975,24.977186,25.062395,24.413355,23.7625,23.111647,22.462606,21.811752,22.272245,22.732738,23.19323,23.65191,24.112402,25.187489,26.262575,27.337664,28.41275,29.487837,29.315605,29.143373,28.96933,28.797098,28.624866,28.325727,28.024776,27.725637,27.424685,27.125546,29.034595,30.945457,32.854507,34.76537,36.67442,35.117085,33.55975,32.002415,30.44508,28.887745,27.8743,26.862667,25.84922,24.837587,23.82414,24.607342,25.390541,26.171928,26.955128,27.738327,27.355793,26.973257,26.590723,26.208187,25.825651,24.975372,24.125093,23.274813,22.424534,21.574255,21.563377,21.550686,21.537996,21.525305,21.512613,24.819458,28.128115,31.434958,34.741802,38.050457,36.694363,35.34008,33.985798,32.6297,31.275417,30.327238,29.379059,28.432692,27.484512,26.538147,3.1744974,3.8471067,4.519716,5.1923246,5.864934,6.5375433,7.4458375,8.352319,9.2606125,10.167094,11.075388,10.165281,9.255174,8.345067,7.4349594,6.5248523,6.9508986,7.3751316,7.799365,8.225411,8.649645,9.295059,9.940474,10.585889,11.22949,11.874905,10.243238,8.609759,6.978093,5.3446136,3.7129474,3.6930048,3.673062,3.6531196,3.633177,3.6132345,3.5751622,3.53709,3.5008307,3.4627585,3.4246864,3.2597067,3.094727,2.9297476,2.764768,2.5997884,3.0747845,3.5497808,4.024777,4.499773,4.974769,5.2992897,5.6256227,5.9501433,6.2746634,6.599184,7.3370595,8.074935,8.812811,9.550687,10.28675,9.791811,9.296872,8.801933,8.306994,7.8120556,8.087626,8.363196,8.636953,8.912524,9.188094,8.194591,7.2029004,6.209397,5.217706,4.2242026,4.550536,4.8750563,5.199577,5.52591,5.8504305,8.78743,11.724429,14.663241,17.60024,20.537241,17.774284,15.013144,12.250188,9.487233,6.7242785,7.175706,7.6253204,8.074935,8.52455,8.974165,9.896963,10.81976,11.7425585,12.665357,13.588155,13.330714,13.073273,12.815832,12.558392,12.299138,11.213174,10.125396,9.037619,7.949841,6.8620634,7.415017,7.9679704,8.520925,9.072064,9.625018,8.997733,8.370448,7.743163,7.115878,6.48678,6.1223745,5.7579694,5.391751,5.027345,4.6629395,4.8333583,5.0019636,5.1723824,5.3428006,5.5132194,6.0480433,6.582867,7.117691,7.652515,8.187339,7.8229337,7.456715,7.0923095,6.7279043,6.3616858,8.370448,10.377398,12.384347,14.39311,16.400059,16.102734,15.805408,15.508082,15.210756,14.911617,14.322405,13.7331915,13.142166,12.552953,11.961927,13.938056,15.912373,17.886688,19.862818,21.837133,21.909653,21.982172,22.05469,22.127209,22.199726,21.233418,20.265295,19.297174,18.330864,17.362743,16.584982,15.80722,15.02946,14.2516985,13.475751,13.4050455,13.33434,13.265448,13.194741,13.125849,12.8321495,12.540262,12.248375,11.954676,11.662788,11.153346,10.642091,10.1326475,9.623205,9.11195,8.999546,8.887142,8.774739,8.662335,8.549932,9.304124,10.060129,10.8143215,11.570327,12.32452,12.262879,12.199425,12.137785,12.07433,12.012691,11.418038,10.823386,10.226922,9.63227,9.037619,9.603263,10.167094,10.7327385,11.298383,11.862214,12.268318,12.672608,13.0769,13.483003,13.887294,14.137483,14.387671,14.63786,14.888049,15.138238,15.50083,15.861609,16.224201,16.586794,16.949387,17.351866,17.754343,18.15682,18.559298,18.961775,18.41426,17.866747,17.319231,16.771717,16.224201,15.528025,14.830034,14.132043,13.435865,12.737875,12.549327,12.362592,12.175857,11.9873085,11.800573,11.887595,11.974618,12.06164,12.1504755,12.237497,13.68968,15.141864,16.59586,18.048042,19.500225,16.494333,13.490254,10.484363,7.4802837,4.4743915,3.587853,2.6995013,1.8129625,0.9246109,0.038072214,2.6306088,5.223145,7.8156815,10.408218,13.000754,11.30926,9.619579,7.9298983,6.240217,4.550536,4.347484,4.1444325,3.9431937,3.7401419,3.53709,3.489953,3.442816,3.395679,3.346729,3.299592,3.7691493,4.2405195,4.710077,5.179634,5.6491914,6.035352,6.4197006,6.8058615,7.1902094,7.574558,8.660522,9.744674,10.830639,11.91479,13.000754,10.962985,8.925215,6.887445,4.8496747,2.811905,2.3042755,1.7966459,1.2908293,0.78319985,0.2755703,0.21936847,0.16497959,0.11059072,0.054388877,0.0,0.0,0.0,0.0,0.0,0.0,0.4604925,0.91917205,1.3796645,1.840157,2.3006494,2.752077,3.2053177,3.6567454,4.1099863,4.5632267,5.163317,5.7615952,6.3616858,6.9617763,7.5618668,7.7703576,7.9770355,8.185526,8.392203,8.600695,9.20985,9.820818,10.429974,11.039129,11.650098,11.213174,10.774437,10.337513,9.900589,9.461852,10.567759,11.671853,12.7777605,13.881854,14.9877615,15.767336,16.54691,17.328297,18.10787,18.887444,18.568363,18.247469,17.928387,17.607492,17.286598,16.494333,15.702069,14.909804,14.117539,13.325275,12.250188,11.175101,10.100015,9.024928,7.949841,7.804804,7.6597667,7.51473,7.369693,7.224656,6.9146395,6.604623,6.294606,5.9845896,5.674573,6.981719,8.290678,9.597824,10.90497,12.212116,12.344462,12.476809,12.609155,12.743314,12.87566,12.092461,11.30926,10.527874,9.744674,8.963287,9.815379,10.667472,11.519565,12.371656,13.225562,12.195799,11.164224,10.13446,9.104698,8.074935,9.882459,11.689982,13.497506,15.30503,17.112555,21.398397,25.682428,29.968271,34.2523,38.538147,35.06451,31.592686,28.11905,24.647226,21.175404,18.459585,15.74558,13.029762,10.315757,7.5999393,7.755854,7.909956,8.06587,8.219973,8.375887,8.847258,9.32044,9.791811,10.264994,10.738177,10.54419,10.352016,10.1598425,9.967669,9.775495,10.540565,11.3056345,12.070704,12.835775,13.600845,13.2146845,12.830337,12.444175,12.059827,11.675479,9.487233,7.3008003,5.1125546,2.9243085,0.73787576,0.89560354,1.0533313,1.209246,1.3669738,1.5247015,2.8517902,4.1806917,5.5077806,6.834869,8.161958,8.600695,9.037619,9.474543,9.91328,10.3502035,11.887595,13.424988,14.96238,16.499773,18.037165,17.350052,16.66294,15.975826,15.2869005,14.599788,13.782142,12.964496,12.14685,11.329204,10.51337,10.435412,10.357455,10.279498,10.203354,10.125396,9.273304,8.419398,7.567306,6.7152133,5.863121,6.037165,6.2130227,6.3870673,6.5629244,6.736969,7.3733187,8.007855,8.642392,9.27693,9.91328,10.112705,10.312131,10.51337,10.712796,10.912222,10.192475,9.47273,8.752983,8.033237,7.311678,7.8120556,8.312433,8.812811,9.313189,9.811753,10.252303,10.692853,11.133403,11.57214,12.012691,11.849524,11.6881695,11.525003,11.361836,11.200482,10.529687,9.860703,9.189907,8.519112,7.850128,7.2899227,6.7297173,6.169512,5.6093063,5.049101,6.82943,8.609759,10.390089,12.170418,13.9507475,12.377095,10.805257,9.231606,7.6597667,6.0879283,6.26016,6.432391,6.604623,6.776854,6.9508986,7.344311,7.7395372,8.134763,8.529989,8.925215,9.715667,10.504305,11.294757,12.085209,12.87566,13.049705,13.225562,13.399607,13.575464,13.749508,13.319836,12.890164,12.460492,12.03082,11.599335,10.903157,10.205167,9.507175,8.809185,8.113008,7.2047133,6.298232,5.389938,4.4834566,3.5751622,3.9830787,4.3891826,4.797099,5.2050157,5.612932,6.4831543,7.3533764,8.221786,9.092008,9.96223,10.437225,10.912222,11.3872175,11.862214,12.337211,13.192928,14.046834,14.902553,15.758271,16.612177,18.610062,20.607946,22.605831,24.601902,26.599787,26.73032,26.860853,26.989574,27.120108,27.25064,26.425743,25.600845,24.774134,23.949236,23.124338,23.755249,24.384346,25.015257,25.644356,26.275267,27.299591,28.325727,29.350052,30.374374,31.400513,30.807673,30.214834,29.621996,29.029158,28.438131,27.861609,27.2869,26.71219,26.137482,25.562773,27.729263,29.897566,32.06587,34.23236,36.40066,35.265747,34.12902,32.994106,31.859192,30.724277,28.974768,27.22526,25.47575,23.724428,21.97492,22.509743,23.044567,23.579391,24.114216,24.650852,24.50219,24.35534,24.206676,24.059826,23.912977,22.500679,21.086567,19.67427,18.261972,16.849674,17.513218,18.17495,18.836681,19.500225,20.161957,24.097898,28.03384,31.96797,35.9021,39.83804,37.997883,36.157726,34.31757,32.477413,30.637255,30.095179,29.553102,29.009214,28.467138,27.925062,3.6875658,4.4381323,5.186886,5.9374523,6.688019,7.4367723,8.4756,9.512614,10.549629,11.586644,12.625471,11.236742,9.849826,8.46291,7.07418,5.6872635,5.825049,5.962834,6.1006193,6.2384043,6.3743763,7.1865835,8.000604,8.812811,9.625018,10.437225,8.899834,7.362441,5.825049,4.2876563,2.7502642,2.762955,2.7756457,2.7883365,2.7992141,2.811905,2.9750717,3.1382382,3.299592,3.4627585,3.6241121,3.3757362,3.1255474,2.8753586,2.6251698,2.374981,3.100166,3.825351,4.550536,5.275721,6.000906,5.9882154,5.975525,5.962834,5.9501433,5.9374523,6.5756154,7.211965,7.850128,8.488291,9.12464,8.825501,8.52455,8.225411,7.9244595,7.6253204,7.650702,7.6742706,7.699652,7.7250338,7.750415,7.0125394,6.2746634,5.5367875,4.800725,4.062849,4.4254417,4.788034,5.1506267,5.5132194,5.8758116,9.574255,13.274512,16.97477,20.675026,24.375282,20.986855,17.60024,14.211814,10.825199,7.4367723,7.949841,8.46291,8.974165,9.487233,10.000301,11.312886,12.625471,13.938056,15.250641,16.563227,15.787278,15.013144,14.237195,13.46306,12.687112,11.575767,10.462607,9.349448,8.238102,7.124943,7.500226,7.8755093,8.2507925,8.624263,8.999546,8.225411,7.4494634,6.6753283,5.89938,5.125245,4.788034,4.4508233,4.1117992,3.774588,3.437377,3.4119956,3.386614,3.3630457,3.3376641,3.3122826,4.4508233,5.5875506,6.7242785,7.8628187,8.999546,8.424837,7.850128,7.2754188,6.70071,6.1241875,8.350506,10.57501,12.799516,15.025834,17.25034,17.087172,16.92582,16.762651,16.599485,16.438131,15.8869915,15.337664,14.788336,14.237195,13.687867,15.738328,17.786976,19.837437,21.887897,23.938358,23.82414,23.711737,23.599335,23.48693,23.374527,22.22511,21.07569,19.92446,18.77504,17.625622,16.813416,15.999394,15.187187,14.37498,13.562773,13.399607,13.238253,13.075087,12.91192,12.750566,12.60009,12.449615,12.299138,12.1504755,11.999999,11.361836,10.725487,10.087324,9.449161,8.812811,8.636953,8.46291,8.287052,8.113008,7.93715,8.636953,9.336758,10.038374,10.738177,11.437981,11.586644,11.73712,11.887595,12.038072,12.186734,11.5503845,10.912222,10.275872,9.637709,8.999546,9.663091,10.324821,10.988366,11.650098,12.311829,12.674421,13.037014,13.399607,13.762199,14.124791,14.474693,14.824595,15.174497,15.524399,15.8743,15.749206,15.624111,15.50083,15.375735,15.250641,15.337664,15.4246855,15.511708,15.600543,15.687565,15.636803,15.5878525,15.537089,15.488139,15.437376,14.587097,13.736817,12.888351,12.038072,11.187792,10.912222,10.636651,10.362894,10.087324,9.811753,10.500679,11.187792,11.874905,12.562017,13.24913,14.824595,16.400059,17.975525,19.549175,21.12464,17.212267,13.299893,9.38752,5.475147,1.5627737,1.2491312,0.93730164,0.62547207,0.31182957,0.0,3.2506418,6.4994707,9.750113,13.000754,16.249584,14.137483,12.025381,9.91328,7.799365,5.6872635,5.337362,4.98746,4.6375585,4.2876563,3.9377546,3.6494937,3.3630457,3.0747845,2.7883365,2.5000753,3.4119956,4.325729,5.237649,6.149569,7.063302,7.362441,7.663393,7.9625316,8.26167,8.562622,9.788185,11.011934,12.237497,13.46306,14.68681,11.874905,9.063,6.249282,3.437377,0.62547207,0.50037766,0.37528324,0.25018883,0.12509441,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.5747091,1.1494182,1.7241274,2.3006494,2.8753586,3.437377,3.9993954,4.5632267,5.125245,5.6872635,6.200332,6.7115874,7.224656,7.7377243,8.2507925,8.062244,7.8755093,7.686961,7.500226,7.311678,8.087626,8.861761,9.637709,10.411844,11.187792,10.924912,10.662033,10.399154,10.138086,9.875207,11.124338,12.375282,13.6244135,14.875358,16.124489,16.875055,17.625622,18.374376,19.124943,19.87551,19.436771,18.999847,18.562923,18.124187,17.687263,17.125244,16.563227,15.999394,15.437376,14.875358,13.486629,12.099712,10.712796,9.325879,7.93715,7.9625316,7.987913,8.013294,8.036863,8.062244,7.750415,7.4367723,7.124943,6.813113,6.4994707,7.9752226,9.449161,10.924912,12.400664,13.874602,13.7875805,13.700559,13.611723,13.524701,13.437678,12.5873995,11.73712,10.88684,10.038374,9.188094,10.000301,10.812509,11.624716,12.436923,13.24913,12.038072,10.825199,9.612328,8.399456,7.1883965,9.461852,11.73712,14.012388,16.287657,18.562923,23.999998,29.437073,34.87596,40.313038,45.75011,41.37543,37.00075,32.62426,28.249582,23.874905,20.649643,17.424383,14.199123,10.975676,7.750415,7.9752226,8.200029,8.424837,8.649645,8.874452,9.374829,9.875207,10.375585,10.874149,11.374527,10.975676,10.57501,10.174346,9.775495,9.374829,10.312131,11.249433,12.186734,13.125849,14.06315,13.037014,12.012691,10.988366,9.96223,8.937905,7.211965,5.487838,3.7618973,2.03777,0.31182957,0.37528324,0.43692398,0.50037766,0.5620184,0.62547207,2.3495996,4.07554,5.7996674,7.5256076,9.249735,9.499924,9.750113,10.000301,10.25049,10.500679,12.1504755,13.800271,15.4500675,17.099863,18.749659,17.774284,16.800724,15.825351,14.849977,13.874602,13.037014,12.199425,11.361836,10.524248,9.686659,9.237044,8.78743,8.337815,7.8882003,7.4367723,6.6626377,5.8866897,5.1125546,4.3366065,3.5624714,4.07554,4.5867953,5.0998635,5.612932,6.1241875,6.825804,7.5256076,8.225411,8.925215,9.625018,9.811753,10.000301,10.1870365,10.375585,10.56232,9.750113,8.937905,8.125698,7.311678,6.4994707,6.849373,7.1992745,7.549176,7.900891,8.2507925,9.200785,10.150778,11.10077,12.050762,13.000754,12.32452,11.650098,10.975676,10.29944,9.625018,8.912524,8.200029,7.4875355,6.775041,6.0625467,5.975525,5.8866897,5.7996674,5.712645,5.6256227,7.699652,9.775495,11.849524,13.925365,15.999394,13.899984,11.800573,9.699349,7.5999393,5.5005283,5.6872635,5.8758116,6.0625467,6.249282,6.43783,6.6753283,6.9128265,7.1503243,7.3878226,7.6253204,8.087626,8.549932,9.012237,9.474543,9.936848,10.2378,10.536939,10.837891,11.137029,11.437981,11.312886,11.187792,11.062697,10.937603,10.812509,10.225109,9.637709,9.050309,8.46291,7.8755093,6.8004227,5.7253356,4.650249,3.5751622,2.5000753,3.1382382,3.774588,4.4127507,5.049101,5.6872635,6.8620634,8.036863,9.211663,10.388275,11.563075,11.874905,12.186734,12.500377,12.812206,13.125849,13.974316,14.824595,15.674874,16.525154,17.375433,19.612629,21.849825,24.08702,26.324217,28.563225,28.73727,28.913128,29.087172,29.26303,29.437073,28.438131,27.437376,26.43662,25.437677,24.436922,25.238253,26.03777,26.837286,27.6368,28.438131,29.411692,30.387066,31.36244,32.337814,33.313187,32.29974,31.288109,30.274662,29.26303,28.249582,27.399303,26.549025,25.700558,24.850279,23.999998,26.425743,28.849674,31.275417,33.69935,36.12509,35.412598,34.700104,33.98761,33.275116,32.562622,30.075235,27.587852,25.100468,22.613083,20.125698,20.412146,20.700407,20.986855,21.275116,21.563377,21.650398,21.737421,21.824444,21.913279,22.000301,20.024172,18.049856,16.075539,14.09941,12.125093,13.46306,14.801026,16.13718,17.475147,18.813112,23.374527,27.937754,32.50098,37.062393,41.62562,39.29959,36.975372,34.64934,32.325123,30.000904,29.86312,29.725334,29.58755,29.449764,29.31198,3.5117085,4.213325,4.9131284,5.612932,6.3127356,7.0125394,7.9770355,8.943344,9.907841,10.872336,11.836833,10.556881,9.27693,7.996978,6.717026,5.4370747,5.774286,6.11331,6.450521,6.787732,7.124943,7.5219817,7.9208336,8.317872,8.714911,9.11195,7.842876,6.5719895,5.3029156,4.0320287,2.762955,2.9243085,3.0874753,3.2506418,3.4119956,3.5751622,3.8180993,4.059223,4.3021603,4.5450974,4.788034,4.365614,3.9431937,3.5207734,3.0983531,2.6741197,3.3376641,3.9993954,4.6629395,5.3246713,5.9882154,6.2365913,6.48678,6.736969,6.987158,7.2373466,7.5056653,7.7721705,8.040489,8.306994,8.575313,8.412147,8.2507925,8.087626,7.9244595,7.763106,7.7848616,7.806617,7.8301854,7.851941,7.8755093,7.324369,6.775041,6.2257137,5.674573,5.125245,5.522284,5.919323,6.3181744,6.7152133,7.112252,10.199727,13.287203,16.374678,19.462152,22.54963,19.518354,16.48527,13.452183,10.419096,7.3878226,7.8319983,8.2779875,8.722163,9.168152,9.612328,10.502492,11.392657,12.282822,13.172986,14.06315,13.515636,12.968122,12.420607,11.873092,11.325577,10.567759,9.80994,9.052122,8.294304,7.5382986,7.7177815,7.897265,8.076748,8.258044,8.437528,7.6851482,6.932769,6.1803894,5.42801,4.6756306,4.3891826,4.1045475,3.8199122,3.5352771,3.2506418,3.2125697,3.1744974,3.1382382,3.100166,3.0620937,3.972201,4.882308,5.7924156,6.7025228,7.61263,7.3370595,7.063302,6.787732,6.5121617,6.2384043,8.140202,10.042,11.94561,13.847408,15.749206,16.090042,16.43088,16.769903,17.11074,17.449764,16.875055,16.300346,15.725637,15.149116,14.574407,17.072668,19.569118,22.06738,24.565643,27.062092,26.19731,25.332525,24.467743,23.60296,22.738176,21.677593,20.61701,19.55824,18.497658,17.437075,16.599485,15.761897,14.924308,14.0867195,13.24913,13.022511,12.79589,12.567456,12.340837,12.112403,12.0416975,11.972805,11.9021,11.833207,11.762501,11.213174,10.662033,10.112705,9.563377,9.012237,8.72035,8.42665,8.134763,7.842876,7.549176,8.185526,8.820063,9.4546,10.089137,10.725487,10.990179,11.254871,11.519565,11.784257,12.050762,11.782444,11.514126,11.24762,10.979301,10.712796,11.124338,11.537694,11.949236,12.362592,12.774135,13.035201,13.294455,13.555521,13.8147745,14.075842,14.4148655,14.755702,15.094727,15.435563,15.774588,15.600543,15.4246855,15.250641,15.074784,14.90074,15.283275,15.66581,16.048346,16.43088,16.811602,16.361988,15.912373,15.462758,15.013144,14.561715,14.01964,13.477564,12.935488,12.3916,11.849524,11.418038,10.98474,10.553255,10.119957,9.686659,10.234174,10.781689,11.329204,11.876718,12.4242325,13.735004,15.045776,16.354736,17.665508,18.974466,15.430124,11.885782,8.339628,4.795286,1.2491312,1.0007553,0.7505665,0.50037766,0.25018883,0.0,2.8608549,5.719897,8.580752,11.439794,14.300649,12.397038,10.49524,8.59163,6.6898317,4.788034,4.7227674,4.6575007,4.592234,4.5269675,4.461701,4.3202896,4.177066,4.0356545,3.8924308,3.7492065,4.3873696,5.0255322,5.661882,6.300045,6.9382076,7.5382986,8.138389,8.736667,9.336758,9.936848,10.587702,11.236742,11.887595,12.536636,13.1874895,10.658407,8.127511,5.5966153,3.0675328,0.53663695,0.9808127,1.4231756,1.8655385,2.3079014,2.7502642,2.6741197,2.5997884,2.525457,2.4493124,2.374981,2.030518,1.6842422,1.3397794,0.99531645,0.6508536,1.2745126,1.8999848,2.525457,3.149116,3.774588,4.494334,5.2140803,5.9356394,6.6553855,7.3751316,7.51473,7.654328,7.795739,7.935337,8.074935,7.9824743,7.890013,7.797552,7.705091,7.61263,8.274362,8.937905,9.599637,10.263181,10.924912,10.903157,10.879588,10.857833,10.834265,10.812509,12.230246,13.647983,15.065719,16.481644,17.89938,18.397943,18.894695,19.393261,19.890013,20.386765,20.343254,20.29793,20.252605,20.207281,20.161957,19.079618,17.99728,16.914942,15.8326025,14.750263,13.602658,12.455053,11.307447,10.1598425,9.012237,9.155461,9.296872,9.440096,9.583321,9.724731,9.211663,8.700407,8.187339,7.6742706,7.1630154,8.180087,9.197159,10.2142315,11.233116,12.250188,12.344462,12.440549,12.534823,12.629097,12.725184,12.1504755,11.575767,10.999244,10.424535,9.849826,10.774437,11.700861,12.625471,13.550082,14.474693,13.780329,13.084151,12.389787,11.695421,10.999244,13.029762,15.06028,17.090797,19.119503,21.15002,26.599787,32.049553,37.499317,42.950897,48.40066,44.174644,39.950443,35.724426,31.500225,27.27421,23.236742,19.199274,15.161806,11.124338,7.0868707,7.440398,7.7921133,8.145641,8.497355,8.8508835,9.139144,9.429218,9.719293,10.009366,10.29944,10.529687,10.7599325,10.990179,11.220426,11.450671,11.635593,11.820516,12.005438,12.19036,12.375282,11.836833,11.300196,10.761745,10.225109,9.686659,8.073122,6.4577727,4.842423,3.2270734,1.6117238,1.3905423,1.167548,0.9445535,0.72337204,0.50037766,2.1628644,3.825351,5.487838,7.1503243,8.812811,9.345822,9.87702,10.410031,10.943042,11.47424,12.687112,13.899984,15.112856,16.325727,17.536787,16.39462,15.252454,14.110288,12.968122,11.8241415,11.044568,10.264994,9.48542,8.705847,7.9244595,7.6742706,7.4258947,7.175706,6.925517,6.6753283,5.910258,5.145188,4.3801174,3.6150475,2.8499773,3.2597067,3.6694362,4.079166,4.4907084,4.900438,5.467895,6.035352,6.60281,7.170267,7.7377243,8.1420145,8.548119,8.952409,9.3567,9.762803,9.367578,8.972352,8.577126,8.1819,7.7866745,7.877322,7.9679704,8.056806,8.147454,8.238102,8.890768,9.541622,10.194288,10.846955,11.499621,10.872336,10.245051,9.617766,8.990481,8.363196,7.8682575,7.3733187,6.87838,6.3816285,5.8866897,5.857682,5.826862,5.7978544,5.767034,5.7380266,7.4802837,9.222541,10.964798,12.707055,14.449312,13.009819,11.570327,10.130835,8.689529,7.250037,7.3352466,7.420456,7.5056653,7.590874,7.6742706,7.690587,7.705091,7.7195945,7.7340984,7.750415,8.161958,8.575313,8.9868555,9.400211,9.811753,10.225109,10.636651,11.050007,11.463363,11.874905,11.845898,11.815077,11.784257,11.755249,11.724429,11.095331,10.46442,9.835322,9.2044115,8.575313,7.723221,6.869315,6.017223,5.1651306,4.313038,4.8623657,5.411693,5.962834,6.5121617,7.063302,8.241728,9.421967,10.602205,11.782444,12.962683,13.247317,13.531953,13.8184,14.103036,14.387671,15.392053,16.398247,17.402628,18.40701,19.413204,21.574255,23.73712,25.899984,28.062847,30.225712,29.906631,29.589363,29.272095,28.954826,28.637556,27.729263,26.82278,25.914488,25.008005,24.099712,25.044266,25.990631,26.935184,27.879738,28.824291,29.645565,30.465023,31.284483,32.105755,32.925213,31.93715,30.949083,29.962833,28.974768,27.986704,27.025833,26.06315,25.100468,24.137783,23.1751,25.497505,27.81991,30.142317,32.46472,34.787125,34.254116,33.722916,33.189907,32.656895,32.125698,30.082489,28.03928,25.997883,23.954674,21.913279,22.217857,22.522434,22.827011,23.13159,23.43798,23.360023,23.282066,23.204107,23.127964,23.050007,21.521679,19.995165,18.466837,16.940323,15.411995,16.483456,17.553104,18.622751,19.6924,20.762047,25.047892,29.333735,33.617764,37.901794,42.18764,39.596916,37.008007,34.417282,31.828371,29.237648,28.800724,28.361986,27.925062,27.488138,27.049402,3.3376641,3.9867048,4.6375585,5.2884116,5.9374523,6.588306,7.4802837,8.372261,9.264238,10.15803,11.050007,9.87702,8.705847,7.5328593,6.359873,5.186886,5.7253356,6.261973,6.8004227,7.3370595,7.8755093,7.85738,7.83925,7.8229337,7.804804,7.7866745,6.7859187,5.7833505,4.780782,3.778214,2.7756457,3.0874753,3.3993049,3.7129474,4.024777,4.3366065,4.6593137,4.9820213,5.3047285,5.6274357,5.9501433,5.3554916,4.76084,4.164375,3.5697234,2.9750717,3.5751622,4.175253,4.7753434,5.375434,5.975525,6.48678,6.9998484,7.512917,8.024173,8.537241,8.435715,8.3323765,8.23085,8.127511,8.024173,8.000604,7.9752226,7.949841,7.9244595,7.900891,7.9208336,7.9407763,7.9607186,7.9806614,8.000604,7.6380115,7.2754188,6.9128265,6.550234,6.187641,6.6191263,7.0524244,7.4857225,7.9172077,8.350506,10.825199,13.299893,15.774588,18.24928,20.725788,18.048042,15.3702965,12.692551,10.014805,7.3370595,7.7141557,8.093065,8.470161,8.847258,9.224354,9.692098,10.1598425,10.627586,11.095331,11.563075,11.242181,10.9230995,10.602205,10.283124,9.96223,9.5597515,9.157274,8.754796,8.352319,7.949841,7.935337,7.9208336,7.9045167,7.890013,7.8755093,7.1448855,6.414262,5.6854506,4.954827,4.2242026,3.9921436,3.7600844,3.5280252,3.294153,3.0620937,3.0131438,2.962381,2.911618,2.8626678,2.811905,3.4953918,4.177066,4.860553,5.542227,6.2257137,6.249282,6.2746634,6.300045,6.3254266,6.350808,7.9298983,9.510801,11.089892,12.670795,14.249886,15.092914,15.934128,16.777155,17.620184,18.463211,17.863121,17.26303,16.66294,16.062849,15.462758,18.40701,21.353073,24.297325,27.24339,30.18764,28.570477,26.953314,25.33434,23.717176,22.100014,21.13008,20.160145,19.190208,18.220274,17.25034,16.38737,15.524399,14.663241,13.800271,12.937301,12.645414,12.351714,12.059827,11.7679405,11.47424,11.485118,11.494183,11.50506,11.514126,11.525003,11.062697,10.600392,10.138086,9.675781,9.211663,8.801933,8.392203,7.9824743,7.572745,7.1630154,7.7322855,8.303369,8.872639,9.441909,10.012992,10.391902,10.772624,11.153346,11.532255,11.912977,12.0145035,12.117842,12.219368,12.322706,12.4242325,12.5873995,12.750566,12.91192,13.075087,13.238253,13.394168,13.551895,13.709623,13.867351,14.025079,14.355038,14.684997,15.014956,15.344915,15.674874,15.4500675,15.22526,15.000452,14.775645,14.5508375,15.227073,15.905121,16.583168,17.259403,17.937452,17.087172,16.236893,15.386614,14.538147,13.687867,13.452183,13.21831,12.982625,12.74694,12.513068,11.922042,11.332829,10.741803,10.152591,9.563377,9.969481,10.377398,10.785315,11.193231,11.599335,12.645414,13.68968,14.73576,15.780026,16.824293,13.647983,10.469859,7.2917356,4.115425,0.93730164,0.7505665,0.5620184,0.37528324,0.18673515,0.0,2.469255,4.940323,7.409578,9.880646,12.349901,10.658407,8.9651,7.271793,5.580299,3.8869917,4.1081734,4.327542,4.5469103,4.7680917,4.98746,4.989273,4.992899,4.994712,4.9983377,5.0001507,5.3627434,5.7253356,6.0879283,6.450521,6.813113,7.7123427,8.611572,9.512614,10.411844,11.312886,11.3872175,11.463363,11.537694,11.612025,11.6881695,9.440096,7.192023,4.945762,2.6976883,0.44961473,1.4594349,2.469255,3.4808881,4.4907084,5.5005283,5.3500524,5.199577,5.049101,4.900438,4.749962,4.059223,3.3702974,2.6795588,1.9906329,1.2998942,1.9743162,2.6505513,3.3249733,3.9993954,4.6756306,5.5531044,6.430578,7.308052,8.185526,9.063,8.829127,8.597069,8.365009,8.13295,7.900891,7.902704,7.9045167,7.9081426,7.909956,7.911769,8.46291,9.012237,9.563377,10.112705,10.662033,10.879588,11.097144,11.314699,11.532255,11.74981,13.33434,14.920682,16.50521,18.08974,19.67427,19.920834,20.165583,20.410334,20.655083,20.899832,21.247921,21.594198,21.942286,22.290375,22.63665,21.035805,19.433146,17.830486,16.227829,14.625169,13.716875,12.810393,11.9021,10.995618,10.087324,10.348391,10.607644,10.866898,11.127964,11.3872175,10.674724,9.96223,9.249735,8.537241,7.8247466,8.384952,8.945157,9.5053625,10.065568,10.625773,10.903157,11.18054,11.457924,11.735307,12.012691,11.711739,11.4126,11.111648,10.812509,10.51337,11.5503845,12.5873995,13.6244135,14.663241,15.700256,15.522586,15.344915,15.167245,14.989574,14.811904,16.597672,18.381628,20.167397,21.953163,23.73712,29.199575,34.662033,40.12449,45.586945,51.0494,46.97386,42.900135,38.824593,34.749054,30.675327,25.82384,20.975977,16.124489,11.274815,6.4251394,6.9055743,7.3841968,7.8646317,8.345067,8.825501,8.9052725,8.985043,9.064813,9.144584,9.224354,10.085511,10.944855,11.804199,12.665357,13.524701,12.957244,12.389787,11.822329,11.254871,10.687414,10.636651,10.587702,10.536939,10.487988,10.437225,8.9324665,7.4277077,5.922949,4.41819,2.911618,2.4058013,1.8981718,1.3905423,0.88291276,0.37528324,1.9743162,3.5751622,5.1741953,6.775041,8.375887,9.189907,10.00574,10.81976,11.635593,12.449615,13.225562,13.999697,14.775645,15.54978,16.325727,15.014956,13.704185,12.395226,11.084454,9.775495,9.052122,8.330563,7.607191,6.885632,6.16226,6.11331,6.0625467,6.011784,5.962834,5.9120708,5.1578784,4.401873,3.6476808,2.8916752,2.137483,2.4456866,2.752077,3.0602808,3.3666716,3.6748753,4.1099863,4.5450974,4.9802084,5.4153194,5.8504305,6.472276,7.0941224,7.7177815,8.339628,8.963287,8.985043,9.006798,9.030367,9.052122,9.07569,8.9052725,8.734854,8.564435,8.39583,8.225411,8.580752,8.934279,9.28962,9.644961,10.000301,9.420154,8.840006,8.259857,7.6797094,7.0995617,6.8221784,6.544795,6.2674117,5.9900284,5.712645,5.7398396,5.767034,5.7942286,5.823236,5.8504305,7.2609153,8.669587,10.080072,11.490557,12.899229,12.119655,11.340081,10.560507,9.77912,8.999546,8.98323,8.9651,8.94697,8.930654,8.912524,8.705847,8.497355,8.290678,8.082188,7.8755093,8.238102,8.600695,8.963287,9.325879,9.686659,10.212419,10.738177,11.262123,11.787883,12.311829,12.377095,12.442362,12.507628,12.572895,12.638163,11.965553,11.292944,10.620335,9.947725,9.275117,8.644206,8.015107,7.3841968,6.755099,6.1241875,6.588306,7.0506115,7.512917,7.9752226,8.437528,9.623205,10.80707,11.992747,13.176612,14.362289,14.61973,14.877171,15.134612,15.392053,15.649493,16.80979,17.970085,19.13038,20.290678,21.44916,23.537693,25.624413,27.712946,29.799665,31.888199,31.077805,30.26741,29.457016,28.648436,27.838041,27.022207,26.208187,25.392353,24.578333,23.7625,24.85209,25.94168,27.033085,28.122675,29.212267,29.877623,30.54298,31.208338,31.871881,32.53724,31.574556,30.611874,29.64919,28.68832,27.725637,26.65055,25.575462,24.500376,23.42529,22.350203,24.56927,26.790148,29.009214,31.230093,33.44916,33.097446,32.74573,32.392204,32.04049,31.68696,30.08974,28.49252,26.8953,25.29808,23.70086,24.021753,24.344461,24.66717,24.989876,25.312584,25.069647,24.82671,24.585585,24.34265,24.099712,23.019186,21.940474,20.859947,19.77942,18.700708,19.502039,20.305182,21.108324,21.909653,22.712795,26.719442,30.727903,34.73455,38.74301,42.749657,39.89424,37.038826,34.185223,31.329807,28.47439,27.738327,27.000452,26.262575,25.5247,24.786825,3.1618068,3.7618973,4.361988,4.9620786,5.562169,6.16226,6.981719,7.802991,8.62245,9.441909,10.263181,9.197159,8.13295,7.066928,6.002719,4.936697,5.674573,6.412449,7.1503243,7.8882003,8.624263,8.192778,7.75948,7.327995,6.8946967,6.4632115,5.727149,4.992899,4.256836,3.5225863,2.7883365,3.2506418,3.7129474,4.175253,4.6375585,5.0998635,5.5023413,5.904819,6.3072968,6.7097745,7.112252,6.345369,5.576673,4.8097897,4.0429068,3.2742105,3.8126602,4.349297,4.8877473,5.424384,5.962834,6.736969,7.512917,8.287052,9.063,9.837135,9.365765,8.892582,8.419398,7.948028,7.474845,7.5872483,7.699652,7.8120556,7.9244595,8.036863,8.054993,8.073122,8.089439,8.107569,8.125698,7.949841,7.7757964,7.5999393,7.4258947,7.250037,7.7177815,8.185526,8.653271,9.119202,9.5869465,11.450671,13.312584,15.174497,17.038223,18.900135,16.57773,14.255324,11.9329195,9.610515,7.28811,7.5981264,7.9081426,8.21816,8.528176,8.838193,8.881703,8.927028,8.972352,9.017676,9.063,8.970539,8.8780775,8.785617,8.693155,8.600695,8.551744,8.504607,8.457471,8.410334,8.363196,8.152893,7.9425893,7.7322855,7.5219817,7.311678,6.604623,5.8975673,5.1905117,4.4816437,3.774588,3.5951047,3.4156215,3.2343252,3.054842,2.8753586,2.811905,2.7502642,2.6868105,2.6251698,2.561716,3.0167696,3.4718235,3.926877,4.3819304,4.836984,5.163317,5.487838,5.812358,6.1368785,6.4632115,7.7195945,8.977791,10.234174,11.49237,12.750566,14.095784,15.439189,16.784407,18.129625,19.474844,18.849373,18.225714,17.60024,16.97477,16.349297,19.743162,23.135216,26.52727,29.919321,33.313187,30.941832,28.57229,26.202747,23.833206,21.461851,20.582563,19.703278,18.822178,17.94289,17.06179,16.175253,15.2869005,14.400362,13.512011,12.625471,12.268318,11.909351,11.552197,11.195044,10.837891,10.926725,11.017374,11.108022,11.1968565,11.287505,10.912222,10.536939,10.161655,9.788185,9.412902,8.885329,8.357758,7.8301854,7.3026133,6.775041,7.2808576,7.7848616,8.290678,8.794682,9.300498,9.795437,10.290376,10.785315,11.280253,11.775192,12.248375,12.719746,13.192928,13.664299,14.137483,14.05046,13.961625,13.874602,13.7875805,13.700559,13.754947,13.809336,13.865538,13.919927,13.974316,14.29521,14.614291,14.935185,15.254267,15.575162,15.299591,15.025834,14.750263,14.474693,14.199123,15.172684,16.144432,17.117992,18.08974,19.063301,17.812357,16.563227,15.312282,14.06315,12.812206,12.884725,12.957244,13.029762,13.102281,13.174799,12.427858,11.680918,10.932164,10.185224,9.438283,9.704789,9.973107,10.239613,10.507931,10.774437,11.555823,12.335398,13.114971,13.894546,14.674119,11.86584,9.055748,6.245656,3.435564,0.62547207,0.50037766,0.37528324,0.25018883,0.12509441,0.0,2.079468,4.160749,6.240217,8.319685,10.399154,8.917963,7.4349594,5.9519563,4.4707656,2.9877625,3.491766,3.9975824,4.503399,5.0074024,5.5132194,5.660069,5.806919,5.955582,6.1024323,6.249282,6.338117,6.4251394,6.5121617,6.599184,6.688019,7.8882003,9.086569,10.28675,11.486931,12.687112,12.186734,11.6881695,11.187792,10.687414,10.1870365,8.221786,6.258347,4.2930956,2.327844,0.36259252,1.93987,3.5171473,5.0944247,6.6717024,8.2507925,8.024173,7.799365,7.574558,7.3497505,7.124943,6.089741,5.0545397,4.019338,2.9841363,1.9507477,2.675933,3.3993049,4.12449,4.8496747,5.57486,6.6100616,7.645263,8.680465,9.715667,10.750868,10.145339,9.539809,8.934279,8.330563,7.7250338,7.8229337,7.9208336,8.01692,8.1148205,8.212721,8.649645,9.088382,9.525306,9.96223,10.399154,10.857833,11.314699,11.773379,12.230246,12.687112,14.440247,16.191568,17.944704,19.697838,21.44916,21.441908,21.434656,21.427404,21.420153,21.4129,22.15259,22.892279,23.631968,24.371656,25.113157,22.99018,20.867199,18.74422,16.623055,14.500074,13.832905,13.165734,12.496751,11.829581,11.162411,11.539507,11.916603,12.295512,12.672608,13.049705,12.137785,11.225864,10.312131,9.400211,8.488291,8.589817,8.693155,8.794682,8.898021,8.999546,9.460039,9.920531,10.37921,10.839704,11.300196,11.274815,11.249433,11.225864,11.200482,11.175101,12.32452,13.475751,14.625169,15.774588,16.92582,17.264843,17.60568,17.944704,18.285542,18.624565,20.165583,21.704788,23.245806,24.785011,26.324217,31.801176,37.27451,42.749657,48.224804,53.69995,49.774887,45.849823,41.92476,37.999695,34.07463,28.41275,22.750868,17.087172,11.42529,5.7615952,6.3707504,6.978093,7.5854354,8.192778,8.80012,8.669587,8.540867,8.410334,8.2798,8.149267,9.639522,11.129777,12.620032,14.110288,15.600543,14.280706,12.96087,11.63922,10.319383,8.999546,9.438283,9.875207,10.312131,10.750868,11.187792,9.791811,8.397643,7.0016613,5.6074934,4.213325,3.4192474,2.6269827,1.8347181,1.0424535,0.25018883,1.7875811,3.3249733,4.8623657,6.399758,7.93715,9.035806,10.1326475,11.22949,12.328146,13.424988,13.762199,14.09941,14.436621,14.775645,15.112856,13.635292,12.157727,10.680162,9.202598,7.7250338,7.059676,6.394319,5.730775,5.0654173,4.40006,4.550536,4.699199,4.8496747,5.0001507,5.1506267,4.405499,3.6603715,2.9152439,2.1701162,1.4249886,1.6298534,1.8347181,2.039583,2.2444477,2.4493124,2.752077,3.054842,3.3576066,3.6603715,3.9631362,4.802538,5.6419396,6.4831543,7.322556,8.161958,8.602508,9.043057,9.481794,9.922344,10.362894,9.933222,9.501737,9.072064,8.642392,8.212721,8.270736,8.326937,8.384952,8.442966,8.499168,7.9679704,7.4349594,6.9019485,6.3707504,5.8377395,5.7779117,5.718084,5.658256,5.5966153,5.5367875,5.621997,5.7072062,5.7924156,5.8776245,5.962834,7.039734,8.116633,9.195346,10.272246,11.349146,11.22949,11.109835,10.990179,10.870523,10.750868,10.629399,10.509744,10.390089,10.270433,10.150778,9.719293,9.28962,8.859948,8.430276,8.000604,8.312433,8.624263,8.937905,9.249735,9.563377,10.199727,10.837891,11.47424,12.112403,12.750566,12.910107,13.069647,13.229188,13.390542,13.550082,12.835775,12.119655,11.405348,10.689227,9.97492,9.567003,9.1609,8.752983,8.345067,7.93715,8.312433,8.6877165,9.063,9.438283,9.811753,11.00287,12.192173,13.383289,14.572594,15.761897,15.992143,16.22239,16.452635,16.682882,16.913128,18.227526,19.541924,20.858135,22.172533,23.48693,25.49932,27.511707,29.52591,31.536484,33.550686,32.247166,30.945457,29.64194,28.34023,27.03671,26.315151,25.59178,24.87022,24.146849,23.42529,24.659918,25.894545,27.129171,28.365612,29.60024,30.109682,30.619125,31.13038,31.639824,32.149265,31.211964,30.274662,29.33736,28.400059,27.462757,26.275267,25.087776,23.900286,22.712795,21.525305,23.642845,25.760386,27.877926,29.995466,32.113007,31.940775,31.766731,31.5945,31.422268,31.250036,30.096992,28.94576,27.792717,26.639671,25.486628,25.827465,26.168303,26.507326,26.848164,27.187187,26.77927,26.373167,25.96525,25.557333,25.149418,24.516693,23.885782,23.253057,22.620335,21.98761,22.522434,23.057259,23.592083,24.126905,24.66173,28.392807,32.12207,35.85315,39.582413,43.311676,40.191566,37.07146,33.953163,30.833055,27.712946,26.674118,25.637104,24.60009,23.563074,22.524246,2.9877625,3.53709,4.0882306,4.6375585,5.186886,5.7380266,6.484967,7.231908,7.9806614,8.727602,9.474543,8.517298,7.560054,6.60281,5.6455655,4.688321,5.6256227,6.5629244,7.500226,8.437528,9.374829,8.528176,7.6797094,6.833056,5.9845896,5.137936,4.670192,4.2024474,3.7347028,3.2669585,2.7992141,3.4119956,4.024777,4.6375585,5.2503395,5.863121,6.345369,6.827617,7.309865,7.7921133,8.274362,7.3352466,6.394319,5.4552045,4.514277,3.5751622,4.0501585,4.5251546,5.0001507,5.475147,5.9501433,6.987158,8.024173,9.063,10.100015,11.137029,10.2958145,9.452786,8.609759,7.7667317,6.925517,7.175706,7.4258947,7.6742706,7.9244595,8.174648,8.189152,8.205468,8.219973,8.234476,8.2507925,8.26167,8.274362,8.287052,8.299743,8.312433,8.814624,9.316814,9.820818,10.323009,10.825199,12.07433,13.325275,14.574407,15.825351,17.074482,15.107417,13.140353,11.173288,9.2044115,7.2373466,7.4802837,7.723221,7.9643445,8.207282,8.450218,8.073122,7.6942134,7.317117,6.9400206,6.5629244,6.697084,6.833056,6.967215,7.1031876,7.2373466,7.5455503,7.851941,8.160145,8.4683485,8.774739,8.370448,7.9643445,7.560054,7.155763,6.7496595,6.0643597,5.3808727,4.695573,4.0102735,3.3249733,3.198066,3.0693457,2.9424384,2.8155308,2.6868105,2.612479,2.5381477,2.4620032,2.3876717,2.3133402,2.5399606,2.7683938,2.9950142,3.2216346,3.4500678,4.07554,4.699199,5.3246713,5.9501433,6.5756154,7.509291,8.444779,9.380268,10.315757,11.249433,13.096842,14.94425,16.79166,18.64088,20.48829,19.837437,19.188396,18.537542,17.886688,17.237648,21.077503,24.917358,28.757212,32.59707,36.43692,33.315,30.193079,27.069344,23.947422,20.8255,20.03505,19.244598,18.454145,17.665508,16.875055,15.963136,15.049402,14.137483,13.225562,12.311829,11.889409,11.466989,11.044568,10.622148,10.199727,10.370146,10.540565,10.70917,10.879588,11.050007,10.761745,10.475298,10.1870365,9.900589,9.612328,8.966913,8.323311,7.6778965,7.0324817,6.3870673,6.827617,7.268167,7.706904,8.147454,8.588004,9.197159,9.808127,10.417283,11.028252,11.637406,12.480434,13.321649,14.164677,15.007704,15.850732,15.511708,15.174497,14.837286,14.500074,14.162864,14.115726,14.066776,14.01964,13.972503,13.925365,14.235382,14.545399,14.855415,15.165432,15.475449,15.149116,14.824595,14.500074,14.175554,13.849221,15.118295,16.385555,17.652817,18.920078,20.187338,18.537542,16.887747,15.23795,13.588155,11.938358,12.317267,12.697989,13.0769,13.457622,13.838344,12.931862,12.027194,11.122525,10.217857,9.313189,9.440096,9.567003,9.695724,9.822631,9.949538,10.46442,10.979301,11.494183,12.010877,12.525759,10.081885,7.6398244,5.197764,2.7557032,0.31182957,0.25018883,0.18673515,0.12509441,0.06164073,0.0,1.6896812,3.3793623,5.0708566,6.7605376,8.450218,7.177519,5.904819,4.632119,3.3594196,2.08672,2.8771715,3.6676233,4.458075,5.2467136,6.037165,6.3308654,6.622752,6.9146395,7.208339,7.500226,7.311678,7.124943,6.9382076,6.7496595,6.5629244,8.062244,9.561564,11.062697,12.562017,14.06315,12.988064,11.912977,10.837891,9.762803,8.6877165,7.0052876,5.3228583,3.6404288,1.9579996,0.2755703,2.420305,4.5650396,6.7097745,8.854509,10.999244,10.700105,10.399154,10.100015,9.800876,9.499924,8.120259,6.740595,5.3591175,3.9794528,2.5997884,3.3757362,4.1498713,4.9258194,5.6999545,6.4759026,7.667019,8.859948,10.052877,11.245807,12.436923,11.459737,10.48255,9.5053625,8.528176,7.549176,7.743163,7.935337,8.127511,8.319685,8.511859,8.838193,9.162713,9.487233,9.811753,10.138086,10.834265,11.532255,12.230246,12.928236,13.6244135,15.544341,17.464268,19.384195,21.304123,23.225864,22.964798,22.705544,22.444477,22.185223,21.924156,23.057259,24.19036,25.321648,26.45475,27.587852,24.944551,22.303066,19.659767,17.01828,14.37498,13.947122,13.519262,13.093216,12.665357,12.237497,12.732436,13.227375,13.722314,14.217253,14.712192,13.599032,12.487686,11.374527,10.263181,9.1500225,8.794682,8.439341,8.0858135,7.7304726,7.3751316,8.01692,8.660522,9.302311,9.945912,10.587702,10.837891,11.088079,11.338268,11.586644,11.836833,13.100468,14.362289,15.625924,16.887747,18.149569,19.0071,19.864632,20.722162,21.579693,22.437225,23.73168,25.027948,26.322403,27.61686,28.913128,34.400967,39.88699,45.37483,50.862667,56.350502,52.5741,48.799515,45.024925,41.25034,37.47575,30.999847,24.525759,18.049856,11.575767,5.0998635,5.8359265,6.5701766,7.304426,8.040489,8.774739,8.435715,8.094878,7.755854,7.415017,7.07418,9.195346,11.314699,13.435865,15.555219,17.674572,15.602356,13.53014,11.457924,9.385707,7.311678,8.238102,9.162713,10.087324,11.011934,11.938358,10.652968,9.367578,8.082188,6.796797,5.5132194,4.4345064,3.3576066,2.280707,1.2019942,0.12509441,1.6008459,3.0747845,4.550536,6.0244746,7.500226,8.87989,10.259555,11.63922,13.020698,14.400362,14.300649,14.199123,14.09941,13.999697,13.899984,12.255627,10.609457,8.9651,7.320743,5.674573,5.06723,4.459888,3.8525455,3.245203,2.6378605,2.9877625,3.3376641,3.6875658,4.0374675,4.3873696,3.6531196,2.9170568,2.182807,1.4467441,0.7124943,0.81583315,0.91735905,1.020698,1.1222239,1.2255627,1.3941683,1.5645868,1.7350051,1.9054236,2.0758421,3.1327994,4.1897564,5.2467136,6.305484,7.362441,8.219973,9.077503,9.935035,10.792566,11.650098,10.959359,10.270433,9.579695,8.890768,8.200029,7.9607186,7.7195945,7.4802837,7.2391596,6.9998484,6.5157876,6.0299134,5.5458527,5.0599785,4.574105,4.7318325,4.88956,5.047288,5.2050157,5.3627434,5.504154,5.6473784,5.7906027,5.9320135,6.0752378,6.8203654,7.5654926,8.31062,9.055748,9.800876,10.339326,10.879588,11.419851,11.9601145,12.500377,12.277383,12.054388,11.833207,11.610212,11.3872175,10.734551,10.081885,9.429218,8.778365,8.125698,8.386765,8.649645,8.912524,9.175404,9.438283,10.1870365,10.937603,11.6881695,12.436923,13.1874895,13.443117,13.696932,13.95256,14.208188,14.462003,13.704185,12.948178,12.19036,11.432542,10.674724,10.489801,10.304879,10.119957,9.935035,9.750113,10.038374,10.324821,10.613083,10.899531,11.187792,12.382534,13.577277,14.772019,15.966762,17.163317,17.364555,17.567608,17.770658,17.971897,18.17495,19.645262,21.115576,22.585888,24.054388,25.5247,27.462757,29.400814,31.337059,33.275116,35.213173,33.416527,31.621693,29.82686,28.032028,26.237194,25.608097,24.977186,24.348087,23.717176,23.088078,24.467743,25.847408,27.227072,28.606737,29.988214,30.341742,30.697083,31.052423,31.407764,31.763105,30.849371,29.93745,29.025532,28.111797,27.199877,25.899984,24.60009,23.300196,22.000301,20.700407,22.71461,24.730623,26.744823,28.759026,30.77504,30.782291,30.789543,30.796795,30.80586,30.813112,30.104244,29.397188,28.690132,27.983078,27.27421,27.633175,27.99033,28.347483,28.704636,29.06179,28.490707,27.91781,27.344915,26.772018,26.199121,26.0142,25.829277,25.644356,25.459433,25.274511,25.54283,25.809336,26.077654,26.34416,26.612478,30.064358,33.51805,36.969933,40.421814,43.875507,40.48889,37.10409,33.71929,30.33449,26.949688,25.611723,24.27557,22.937603,21.599636,20.26167,2.811905,3.3122826,3.8126602,4.313038,4.8116026,5.3119802,5.9882154,6.6626377,7.3370595,8.013294,8.6877165,7.837437,6.987158,6.1368785,5.2865987,4.4381323,5.57486,6.7115874,7.850128,8.9868555,10.125396,8.861761,7.5999393,6.338117,5.0744824,3.8126602,3.6132345,3.4119956,3.2125697,3.0131438,2.811905,3.5751622,4.3366065,5.0998635,5.863121,6.624565,7.1883965,7.750415,8.312433,8.874452,9.438283,8.325124,7.211965,6.1006193,4.98746,3.874301,4.2876563,4.699199,5.1125546,5.52591,5.9374523,7.2373466,8.537241,9.837135,11.137029,12.436923,11.225864,10.012992,8.80012,7.5872483,6.3743763,6.7623506,7.1503243,7.5382986,7.9244595,8.312433,8.325124,8.337815,8.350506,8.363196,8.375887,8.575313,8.774739,8.974165,9.175404,9.374829,9.91328,10.449916,10.988366,11.525003,12.06164,12.699803,13.337966,13.974316,14.612478,15.250641,13.637105,12.025381,10.411844,8.80012,7.1883965,7.362441,7.5382986,7.7123427,7.8882003,8.062244,7.262728,6.4632115,5.661882,4.8623657,4.062849,4.4254417,4.788034,5.1506267,5.5132194,5.8758116,6.5375433,7.1992745,7.8628187,8.52455,9.188094,8.588004,7.987913,7.3878226,6.787732,6.187641,5.52591,4.8623657,4.2006345,3.53709,2.8753586,2.7992141,2.7248828,2.6505513,2.5744069,2.5000753,2.4130533,2.324218,2.2371957,2.1501737,2.0631514,2.0631514,2.0631514,2.0631514,2.0631514,2.0631514,2.9877625,3.9123733,4.836984,5.763408,6.688019,7.3008003,7.911769,8.52455,9.137331,9.750113,12.099712,14.449312,16.800724,19.150324,21.499924,20.8255,20.149265,19.474844,18.800423,18.124187,22.411844,26.6995,30.987156,35.274815,39.56247,35.688168,31.812054,27.937754,24.06164,20.187338,19.487535,18.787731,18.087927,17.388124,16.68832,15.749206,14.811904,13.874602,12.937301,11.999999,11.512312,11.024626,10.536939,10.049252,9.563377,9.811753,10.061942,10.312131,10.56232,10.812509,10.613083,10.411844,10.212419,10.012992,9.811753,9.050309,8.287052,7.5256076,6.7623506,6.000906,6.3743763,6.7496595,7.124943,7.500226,7.8755093,8.600695,9.325879,10.049252,10.774437,11.499621,12.712494,13.925365,15.138238,16.349297,17.562168,16.97477,16.38737,15.799969,15.212569,14.625169,14.474693,14.324218,14.175554,14.025079,13.874602,14.175554,14.474693,14.775645,15.074784,15.375735,15.000452,14.625169,14.249886,13.874602,13.499319,15.062093,16.624866,18.187641,19.750414,21.313189,19.262728,17.212267,15.161806,13.113158,11.062697,11.74981,12.436923,13.125849,13.812962,14.500074,13.437678,12.375282,11.312886,10.25049,9.188094,9.175404,9.162713,9.1500225,9.137331,9.12464,9.374829,9.625018,9.875207,10.125396,10.375585,8.299743,6.2257137,4.1498713,2.0758421,0.0,0.0,0.0,0.0,0.0,0.0,1.2998942,2.5997884,3.8996825,5.199577,6.4994707,5.4370747,4.3746786,3.3122826,2.2498865,1.1874905,2.2625773,3.3376641,4.4127507,5.487838,6.5629244,6.9998484,7.4367723,7.8755093,8.312433,8.749357,8.287052,7.8247466,7.362441,6.9001355,6.43783,8.238102,10.036561,11.836833,13.637105,15.437376,13.7875805,12.137785,10.487988,8.838193,7.1883965,5.7869763,4.3873696,2.9877625,1.5881553,0.18673515,2.9007401,5.612932,8.325124,11.037316,13.749508,13.374225,13.000754,12.625471,12.250188,11.874905,10.150778,8.424837,6.70071,4.974769,3.2506418,4.07554,4.900438,5.7253356,6.550234,7.3751316,8.725789,10.074633,11.42529,12.774135,14.124791,12.774135,11.42529,10.074633,8.725789,7.3751316,7.663393,7.949841,8.238102,8.52455,8.812811,9.024928,9.237044,9.449161,9.663091,9.875207,10.812509,11.74981,12.687112,13.6244135,14.561715,16.650248,18.736969,20.8255,22.912222,25.000753,24.487686,23.974617,23.463362,22.950293,22.437225,23.961926,25.486628,27.013142,28.537844,30.062546,26.898926,23.73712,20.575312,17.411694,14.249886,14.06315,13.874602,13.687867,13.499319,13.312584,13.925365,14.538147,15.149116,15.761897,16.374678,15.062093,13.749508,12.436923,11.124338,9.811753,8.999546,8.187339,7.3751316,6.5629244,5.750717,6.5756154,7.400513,8.225411,9.050309,9.875207,10.399154,10.924912,11.450671,11.974618,12.500377,13.874602,15.250641,16.624866,18.000906,19.375132,20.749357,22.125395,23.49962,24.87566,26.249886,27.299591,28.349297,29.400814,30.45052,31.500225,37.00075,42.49947,47.999996,53.500526,58.99924,55.37513,51.75102,48.12509,44.49917,40.875053,33.586945,26.300648,19.012539,11.724429,4.4381323,5.2992897,6.16226,7.02523,7.8882003,8.749357,8.200029,7.650702,7.0995617,6.550234,6.000906,8.749357,11.499621,14.249886,17.00015,19.750414,16.924006,14.09941,11.274815,8.450218,5.6256227,7.037921,8.450218,9.862516,11.274815,12.687112,11.512312,10.337513,9.162713,7.987913,6.813113,5.4497657,4.0882306,2.7248828,1.3633479,0.0,1.4122978,2.8245957,4.2368937,5.6491914,7.063302,8.725789,10.388275,12.050762,13.713249,15.375735,14.837286,14.300649,13.762199,13.225562,12.687112,10.874149,9.063,7.250037,5.4370747,3.6241121,3.0747845,2.525457,1.9743162,1.4249886,0.87566096,1.4249886,1.9743162,2.525457,3.0747845,3.6241121,2.9007401,2.175555,1.4503701,0.72518504,0.0,0.0,0.0,0.0,0.0,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,1.4630609,2.7375734,4.0120864,5.2884116,6.5629244,7.837437,9.11195,10.388275,11.662788,12.937301,11.9873085,11.037316,10.087324,9.137331,8.187339,7.650702,7.112252,6.5756154,6.037165,5.5005283,5.0617914,4.6248674,4.1879435,3.7492065,3.3122826,3.6875658,4.062849,4.4381323,4.8116026,5.186886,5.388125,5.5875506,5.7869763,5.9882154,6.187641,6.599184,7.0125394,7.4258947,7.837437,8.2507925,9.4509735,10.649343,11.849524,13.049705,14.249886,13.925365,13.600845,13.274512,12.949992,12.625471,11.74981,10.874149,10.000301,9.12464,8.2507925,8.46291,8.675026,8.887142,9.099259,9.313189,10.174346,11.037316,11.900287,12.763257,13.6244135,13.974316,14.324218,14.674119,15.025834,15.375735,14.574407,13.77489,12.975373,12.175857,11.374527,11.4126,11.450671,11.486931,11.525003,11.563075,11.762501,11.961927,12.163166,12.362592,12.562017,13.762199,14.96238,16.162561,17.362743,18.562923,18.736969,18.912827,19.08687,19.262728,19.436771,21.063,22.687414,24.311829,25.938055,27.56247,29.424383,31.288109,33.15002,35.011932,36.87566,34.5877,32.29974,30.011782,27.725637,25.437677,24.89923,24.36259,23.82414,23.287504,22.750868,24.27557,25.80027,27.324972,28.849674,30.374374,30.575613,30.77504,30.974466,31.175705,31.37513,30.486778,29.60024,28.71189,27.82535,26.936998,25.5247,24.112402,22.700104,21.287807,19.87551,21.788185,23.70086,25.611723,27.524399,29.437073,29.625622,29.812357,30.000904,30.18764,30.374374,30.113308,29.85043,29.58755,29.324669,29.06179,29.437073,29.812357,30.18764,30.562923,30.938206,30.20033,29.462456,28.724579,27.986704,27.25064,27.511707,27.774588,28.037466,28.300346,28.563225,28.563225,28.563225,28.563225,28.563225,28.563225,31.737722,34.91222,38.08672,41.263027,44.437527,40.788033,37.136726,33.487232,29.837738,26.188244,24.549326,22.912222,21.275116,19.63801,18.000906,2.663242,3.005892,3.346729,3.6893787,4.0320287,4.3746786,5.027345,5.6800117,6.3326783,6.985345,7.6380115,7.0306687,6.4233265,5.814171,5.2068286,4.599486,5.527723,6.454147,7.382384,8.31062,9.237044,8.033237,6.827617,5.621997,4.41819,3.2125697,3.1726844,3.1327994,3.092914,3.053029,3.0131438,3.8126602,4.612177,5.411693,6.2130227,7.0125394,7.407765,7.802991,8.198216,8.59163,8.9868555,8.31062,7.6325727,6.9545245,6.2782893,5.600241,5.57486,5.5494785,5.524097,5.5005283,5.475147,6.6155005,7.755854,8.894395,10.034748,11.175101,10.31757,9.460039,8.602508,7.744976,6.887445,7.2482243,7.607191,7.9679704,8.326937,8.6877165,8.620637,8.551744,8.484665,8.417585,8.350506,8.354132,8.3595705,8.365009,8.370448,8.375887,9.026741,9.679407,10.332074,10.98474,11.637406,12.132345,12.627284,13.122223,13.617162,14.112101,12.730623,11.347333,9.965856,8.582565,7.1992745,7.124943,7.0506115,6.9744673,6.9001355,6.825804,6.1822023,5.540414,4.896812,4.255023,3.6132345,3.8833659,4.1516843,4.421816,4.691947,4.9620786,5.612932,6.261973,6.9128265,7.5618668,8.212721,7.8102427,7.407765,7.0052876,6.60281,6.200332,5.4969025,4.795286,4.0918565,3.39024,2.6868105,2.5870976,2.4873846,2.3876717,2.2879589,2.1882458,2.2081885,2.228131,2.2480736,2.268016,2.2879589,2.2353828,2.182807,2.1302311,2.077655,2.0250793,2.7847104,3.5443418,4.305786,5.0654173,5.825049,6.599184,7.3751316,8.149267,8.925215,9.699349,11.856775,14.014201,16.173439,18.330864,20.48829,20.100317,19.712341,19.324368,18.938208,18.550234,23.220425,27.890615,32.560806,37.229187,41.89938,37.999695,34.100014,30.20033,26.300648,22.399153,21.664904,20.930653,20.19459,19.46034,18.724277,17.4407,16.15531,14.869919,13.584529,12.299138,11.965553,11.630155,11.294757,10.959359,10.625773,10.812509,10.999244,11.187792,11.374527,11.563075,11.563075,11.563075,11.563075,11.563075,11.563075,10.73999,9.916905,9.0956335,8.272549,7.4494634,7.5854354,7.7195945,7.855567,7.989726,8.125698,8.865387,9.605076,10.344765,11.084454,11.8241415,12.902855,13.979754,15.056654,16.135366,17.212267,16.691946,16.171627,15.653119,15.132799,14.612478,14.353225,14.092158,13.832905,13.571837,13.312584,13.742256,14.171928,14.603414,15.033086,15.462758,15.072971,14.683184,14.291584,13.901797,13.512011,14.935185,16.358362,17.779724,19.2029,20.624262,18.715212,16.80435,14.895301,12.984438,11.075388,11.570327,12.065266,12.5602045,13.055143,13.550082,12.872034,12.195799,11.517752,10.839704,10.161655,9.731983,9.302311,8.872639,8.442966,8.013294,8.074935,8.138389,8.200029,8.26167,8.325124,6.6698895,5.0146546,3.3594196,1.7041848,0.05076295,0.22480737,0.40066472,0.5747091,0.7505665,0.9246109,2.0577126,3.1908143,4.322103,5.4552045,6.588306,5.5494785,4.512464,3.4754493,2.4366217,1.3996071,2.6505513,3.8996825,5.1506267,6.399758,7.650702,7.855567,8.0604315,8.265296,8.470161,8.675026,8.210908,7.744976,7.2808576,6.814926,6.350808,7.699652,9.050309,10.399154,11.74981,13.100468,11.680918,10.259555,8.840006,7.420456,5.999093,4.8297324,3.6603715,2.4891977,1.3198367,0.15047589,2.962381,5.774286,8.588004,11.399909,14.211814,13.925365,13.637105,13.3506565,13.062395,12.774135,10.765372,8.754796,6.7442207,4.7354584,2.7248828,3.5534067,4.3801174,5.2068286,6.035352,6.8620634,8.406708,9.953164,11.497808,13.042453,14.587097,13.727753,12.868408,12.007251,11.147907,10.28675,9.882459,9.4781685,9.072064,8.667774,8.26167,8.830941,9.396585,9.965856,10.533313,11.10077,11.769753,12.440549,13.109532,13.780329,14.449312,15.814472,17.179634,18.544794,19.909956,21.275116,20.705845,20.134762,19.565493,18.99441,18.425138,19.739536,21.055748,22.370146,23.684544,25.000753,22.930351,20.859947,18.789545,16.719141,14.650551,14.68681,14.724882,14.762955,14.799213,14.837286,14.762955,14.68681,14.612478,14.538147,14.462003,13.220123,11.978244,10.734551,9.492672,8.2507925,7.746789,7.2445984,6.742408,6.240217,5.7380266,6.4269524,7.117691,7.806617,8.497355,9.188094,10.125396,11.062697,11.999999,12.937301,13.874602,15.854358,17.834112,19.815681,21.795437,23.77519,24.737875,25.700558,26.66324,27.625923,28.586794,29.536787,30.486778,31.436771,32.386765,33.336758,38.077652,42.81674,47.557636,52.29672,57.037617,53.475143,49.912674,46.3502,42.78773,39.225258,32.27255,25.319836,18.367125,11.4144125,4.461701,5.177821,5.8921285,6.6082487,7.322556,8.036863,7.804804,7.572745,7.3406854,7.1068134,6.874754,9.104698,11.334642,13.564586,15.79453,18.024473,15.838041,13.649796,11.46155,9.275117,7.0868707,8.247167,9.407463,10.567759,11.728055,12.888351,11.419851,9.953164,8.484665,7.017978,5.5494785,4.8641787,4.1806917,3.4953918,2.810092,2.124792,2.904366,3.6857529,4.465327,5.2449007,6.0244746,8.06587,10.1054535,12.145037,14.184619,16.224201,15.181748,14.139296,13.096842,12.054388,11.011934,9.400211,7.7866745,6.1749506,4.5632267,2.94969,2.5472124,2.1447346,1.742257,1.3397794,0.93730164,1.5101979,2.0830941,2.6541772,3.2270734,3.7999697,3.0403383,2.280707,1.5192627,0.75963134,0.0,0.0,0.0,0.0,0.0,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,1.2291887,2.3097143,3.39024,4.4707656,5.5494785,6.6644506,7.7794223,8.894395,10.009366,11.124338,10.435412,9.744674,9.055748,8.365009,7.6742706,7.322556,6.970841,6.6173134,6.265599,5.9120708,5.6818247,5.4533916,5.223145,4.992899,4.762653,4.933071,5.101677,5.272095,5.4425135,5.612932,5.9392653,6.2674117,6.5955577,6.921891,7.250037,8.013294,8.774739,9.537996,10.29944,11.062697,11.827768,12.592838,13.357908,14.122978,14.888049,14.9877615,15.087475,15.187187,15.2869005,15.386614,14.46019,13.531953,12.605529,11.677292,10.750868,10.752681,10.754494,10.75812,10.7599325,10.761745,11.354585,11.947423,12.540262,13.1331005,13.724127,13.874602,14.025079,14.175554,14.324218,14.474693,13.812962,13.149418,12.487686,11.8241415,11.162411,11.285692,11.407161,11.530442,11.651911,11.775192,12.077957,12.380721,12.681673,12.984438,13.287203,14.26439,15.241576,16.220575,17.197763,18.17495,18.76235,19.34975,19.93715,20.52455,21.11195,22.489801,23.867653,25.245504,26.621542,27.999393,29.09805,30.194891,31.291735,32.39039,33.487232,31.68152,29.877623,28.071913,26.268015,24.462305,24.03807,23.612024,23.187792,22.761745,22.337511,23.577578,24.817644,26.05771,27.297777,28.537844,28.316662,28.097294,27.877926,27.656744,27.437376,26.835472,26.231756,25.629852,25.027948,24.424232,23.38903,22.355642,21.32044,20.285238,19.250036,20.675026,22.100014,23.525002,24.949991,26.374979,26.949688,27.524399,28.099108,28.675629,29.250338,29.15244,29.054539,28.956638,28.860552,28.762651,29.06179,29.362741,29.66188,29.962833,30.26197,29.30654,28.352922,27.397491,26.442059,25.486628,25.96525,26.442059,26.920681,27.397491,27.8743,27.61686,27.359419,27.101978,26.844538,26.587097,28.70101,30.813112,32.925213,35.037315,37.149418,34.06738,30.985344,27.901495,24.819458,21.737421,20.502794,19.268166,18.031725,16.797098,15.56247,2.5127661,2.6976883,2.8826106,3.0675328,3.2524548,3.437377,4.068288,4.6973863,5.328297,5.957395,6.588306,6.2220874,5.857682,5.4932766,5.127058,4.762653,5.480586,6.1967063,6.9146395,7.6325727,8.350506,7.2029004,6.055295,4.9076896,3.7600844,2.612479,2.7321346,2.8517902,2.9732587,3.092914,3.2125697,4.0501585,4.8877473,5.7253356,6.5629244,7.400513,7.6271334,7.855567,8.082188,8.31062,8.537241,8.294304,8.05318,7.8102427,7.567306,7.324369,6.8620634,6.399758,5.9374523,5.475147,5.0128417,5.9918413,6.972654,7.951654,8.9324665,9.91328,9.409276,8.907085,8.404895,7.902704,7.400513,7.7322855,8.06587,8.397643,8.729415,9.063,8.914337,8.767487,8.620637,8.471974,8.325124,8.134763,7.944402,7.755854,7.5654926,7.3751316,8.1420145,8.910711,9.677594,10.444477,11.213174,11.564888,11.916603,12.270131,12.621845,12.975373,11.822329,10.669285,9.518054,8.365009,7.211965,6.887445,6.5629244,6.2365913,5.9120708,5.5875506,5.101677,4.6176157,4.1317415,3.6476808,3.1618068,3.339477,3.5171473,3.6948178,3.872488,4.0501585,4.688321,5.3246713,5.962834,6.599184,7.2373466,7.0324817,6.827617,6.622752,6.4178877,6.2130227,5.469708,4.7282066,3.9848917,3.24339,2.5000753,2.374981,2.2498865,2.124792,1.9996977,1.8746033,2.0033236,2.1302311,2.2571385,2.3858588,2.5127661,2.4076142,2.3024626,2.1973107,2.0921588,1.987007,2.5816586,3.1781235,3.7727752,4.367427,4.9620786,5.89938,6.836682,7.7757964,8.713099,9.6504,11.615651,13.57909,15.544341,17.509592,19.474844,19.375132,19.275417,19.175705,19.074179,18.974466,24.027193,29.07992,34.132645,39.18537,44.2381,40.313038,36.387974,32.46291,28.537844,24.61278,23.842272,23.071762,22.303066,21.532557,20.762047,19.13038,17.496902,15.865235,14.231756,12.60009,12.416981,12.235684,12.052575,11.869466,11.6881695,11.813264,11.938358,12.06164,12.186734,12.311829,12.513068,12.712494,12.91192,13.113158,13.312584,12.429671,11.546759,10.665659,9.782746,8.899834,8.794682,8.689529,8.584378,8.479226,8.375887,9.130079,9.884272,10.640278,11.39447,12.1504755,13.093216,14.034143,14.976884,15.919624,16.862366,16.409124,15.957697,15.504456,15.053028,14.599788,14.229943,13.860099,13.490254,13.12041,12.750566,13.310771,13.8691635,14.429369,14.989574,15.54978,15.14549,14.739386,14.335095,13.930804,13.524701,14.808278,16.090042,17.371807,18.655384,19.93715,18.167698,16.398247,14.626982,12.857531,11.088079,11.390844,11.691795,11.99456,12.297325,12.60009,12.308203,12.0145035,11.722616,11.430729,11.137029,10.290376,9.441909,8.595256,7.746789,6.9001355,6.775041,6.6499467,6.5248523,6.399758,6.2746634,5.040036,3.8054085,2.570781,1.3343405,0.099712946,0.44961473,0.7995165,1.1494182,1.49932,1.8492218,2.8155308,3.780027,4.744523,5.710832,6.6753283,5.661882,4.650249,3.636803,2.6251698,1.6117238,3.0367124,4.461701,5.8866897,7.311678,8.736667,8.709473,8.682278,8.655084,8.627889,8.600695,8.13295,7.665206,7.1974616,6.7297173,6.261973,7.1630154,8.062244,8.963287,9.862516,10.761745,9.572442,8.383139,7.192023,6.002719,4.8116026,3.872488,2.9333735,1.9924458,1.0533313,0.11240368,3.0258346,5.9374523,8.8508835,11.762501,14.674119,14.474693,14.275268,14.075842,13.874602,13.675177,11.379966,9.084756,6.789545,4.494334,2.1991236,3.0294604,3.8597972,4.690134,5.520471,6.350808,8.089439,9.829884,11.570327,13.310771,15.049402,14.679558,14.309713,13.939869,13.5700245,13.200181,12.103338,11.004683,9.907841,8.809185,7.7123427,8.63514,9.557939,10.480737,11.401722,12.32452,12.726997,13.129475,13.531953,13.93443,14.336908,14.98051,15.622298,16.2659,16.907688,17.549479,16.922194,16.294909,15.667623,15.040338,14.413053,15.517147,16.623055,17.727148,18.833055,19.93715,18.959963,17.982777,17.005589,16.026588,15.049402,15.312282,15.575162,15.838041,16.100922,16.361988,15.600543,14.837286,14.075842,13.312584,12.549327,11.378153,10.205167,9.03218,7.859193,6.688019,6.495845,6.301858,6.109684,5.91751,5.7253356,6.2801023,6.834869,7.3896356,7.944402,8.499168,9.849826,11.200482,12.549327,13.899984,15.250641,17.835926,20.419397,23.004683,25.589968,28.175251,28.724579,29.27572,29.825047,30.374374,30.925516,31.775795,32.62426,33.47454,34.32482,35.1751,39.154552,43.134007,47.115273,51.094723,55.074177,51.57516,48.07433,44.57531,41.074482,37.575462,30.956337,24.340836,17.721708,11.104396,4.4870825,5.0545397,5.621997,6.189454,6.7569118,7.324369,7.409578,7.494787,7.5799966,7.665206,7.750415,9.460039,11.169662,12.879286,14.590723,16.300346,14.750263,13.200181,11.650098,10.100015,8.549932,9.458226,10.364707,11.273002,12.179482,13.087777,11.327391,9.567003,7.806617,6.0480433,4.2876563,4.2804046,4.273153,4.265901,4.256836,4.249584,4.3982472,4.5450974,4.691947,4.84061,4.98746,7.405952,9.822631,12.23931,14.657803,17.074482,15.528025,13.979754,12.433297,10.885027,9.336758,7.9244595,6.5121617,5.0998635,3.6875658,2.275268,2.0196402,1.7658255,1.5101979,1.2545701,1.0007553,1.5954071,2.1900587,2.7847104,3.3793623,3.975827,3.1799364,2.3858588,1.5899682,0.79589057,0.0,0.0,0.0,0.0,0.0,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.99712944,1.8818551,2.7683938,3.6531196,4.537845,5.4932766,6.446895,7.402326,8.357758,9.313189,8.881703,8.452031,8.02236,7.592687,7.1630154,6.9944096,6.827617,6.6608243,6.492219,6.3254266,6.301858,6.2801023,6.258347,6.2347784,6.2130227,6.1767635,6.1423173,6.107871,6.071612,6.037165,6.492219,6.947273,7.402326,7.85738,8.312433,9.425592,10.536939,11.650098,12.763257,13.874602,14.204562,14.534521,14.86448,15.194439,15.524399,16.050158,16.574104,17.099863,17.625622,18.149569,17.170568,16.189756,15.210756,14.229943,13.24913,13.042453,12.835775,12.627284,12.420607,12.212116,12.534823,12.857531,13.180238,13.502945,13.825653,13.77489,13.724127,13.675177,13.6244135,13.575464,13.049705,12.525759,11.999999,11.47424,10.950294,11.156972,11.365462,11.57214,11.780631,11.9873085,12.393413,12.797703,13.201994,13.608097,14.012388,14.7683935,15.522586,16.276777,17.032784,17.786976,18.787731,19.786674,20.78743,21.788185,22.787127,23.918415,25.047892,26.177366,27.306843,28.438131,28.769903,29.101675,29.43526,29.767033,30.100618,28.777155,27.455505,26.132042,24.810392,23.48693,23.1751,22.863272,22.54963,22.237799,21.924156,22.879587,23.835018,24.790451,25.744068,26.6995,26.059525,25.419548,24.779573,24.139597,23.49962,23.182352,22.865084,22.547815,22.230547,21.913279,21.255173,20.597069,19.940775,19.282671,18.624565,19.561867,20.50098,21.438282,22.375584,23.312885,24.27557,25.238253,26.199121,27.161806,28.124489,28.19338,28.26046,28.32754,28.39462,28.4617,28.68832,28.913128,29.137934,29.362741,29.58755,28.414562,27.241575,26.070402,24.897415,23.724428,24.41698,25.109531,25.802084,26.494635,27.187187,26.672306,26.157425,25.642542,25.12766,24.61278,25.662485,26.71219,27.761896,28.811602,29.86312,27.346727,24.832148,22.31757,19.80299,17.286598,16.454449,15.622298,14.790149,13.957999,13.125849,2.3622901,2.3894846,2.4166791,2.4456866,2.472881,2.5000753,3.1074178,3.7147603,4.322103,4.9294453,5.5367875,5.4153194,5.292038,5.1705694,5.047288,4.9258194,5.431636,5.9392653,6.446895,6.9545245,7.462154,6.3725634,5.282973,4.1915693,3.101979,2.0123885,2.2933977,2.572594,2.8517902,3.1327994,3.4119956,4.2876563,5.163317,6.037165,6.9128265,7.7866745,7.8483152,7.9081426,7.9679704,8.027799,8.087626,8.2798,8.471974,8.664148,8.858135,9.050309,8.149267,7.250037,6.350808,5.4497657,4.550536,5.369995,6.189454,7.0107265,7.8301854,8.649645,8.502794,8.354132,8.207282,8.0604315,7.911769,8.21816,8.5227375,8.827314,9.131892,9.438283,9.20985,8.98323,8.754796,8.528176,8.299743,7.915395,7.5292335,7.1448855,6.7605376,6.3743763,7.2572894,8.140202,9.023115,9.904215,10.7871275,10.997431,11.207735,11.418038,11.628342,11.836833,10.915848,9.99305,9.070251,8.147454,7.224656,6.6499467,6.0752378,5.5005283,4.9258194,4.349297,4.022964,3.6948178,3.3666716,3.0403383,2.712192,2.7974012,2.8826106,2.9678197,3.053029,3.1382382,3.7618973,4.3873696,5.0128417,5.638314,6.261973,6.2547207,6.247469,6.240217,6.2329655,6.2257137,5.4425135,4.6593137,3.877927,3.094727,2.3133402,2.1628644,2.0123885,1.8619126,1.7132497,1.5627737,1.7966459,2.032331,2.268016,2.5018883,2.7375734,2.5798457,2.422118,2.2643902,2.1066625,1.9507477,2.38042,2.810092,3.2397642,3.6694362,4.099108,5.199577,6.300045,7.400513,8.499168,9.599637,11.372714,13.145792,14.917056,16.690134,18.463211,18.649946,18.836681,19.025229,19.211964,19.400513,24.835773,30.269224,35.704487,41.139748,46.57501,42.624565,38.67593,34.725487,30.77504,26.824594,26.019638,25.214684,24.409729,23.604773,22.799818,20.820063,18.840307,16.860552,14.880796,12.899229,12.870221,12.839401,12.810393,12.779573,12.750566,12.812206,12.87566,12.937301,13.000754,13.062395,13.46306,13.861912,14.262577,14.663241,15.062093,14.119352,13.178425,12.235684,11.292944,10.3502035,10.00574,9.659465,9.3150015,8.970539,8.624263,9.394773,10.165281,10.93579,11.704487,12.474996,13.281764,14.090345,14.897114,15.705695,16.512463,16.128115,15.741954,15.357606,14.973258,14.587097,14.106662,13.628039,13.147605,12.66717,12.186734,12.877473,13.568212,14.257137,14.947877,15.636803,15.218008,14.7974,14.376793,13.957999,13.537392,14.679558,15.821725,16.965704,18.10787,19.250036,17.620184,15.99033,14.3604765,12.730623,11.10077,11.209548,11.320138,11.430729,11.539507,11.650098,11.7425585,11.83502,11.927481,12.019942,12.112403,10.846955,9.583321,8.317872,7.0524244,5.7869763,5.475147,5.163317,4.8496747,4.537845,4.2242026,3.4101827,2.5943494,1.7803292,0.9644961,0.15047589,0.6744221,1.2001812,1.7241274,2.2498865,2.7756457,3.5733492,4.36924,5.1669436,5.964647,6.7623506,5.774286,4.788034,3.7999697,2.811905,1.8256533,3.4246864,5.0255322,6.624565,8.225411,9.824444,9.56519,9.304124,9.04487,8.785617,8.52455,8.054993,7.5854354,7.115878,6.644508,6.1749506,6.624565,7.07418,7.5256076,7.9752226,8.424837,7.46578,6.5049095,5.5458527,4.5849824,3.6241121,2.9152439,2.2045624,1.4956942,0.7850128,0.07433146,3.0874753,6.1006193,9.11195,12.125093,15.138238,15.025834,14.911617,14.799213,14.68681,14.574407,11.99456,9.414715,6.834869,4.255023,1.6751775,2.5073273,3.339477,4.171627,5.0055895,5.8377395,7.7721705,9.706602,11.642846,13.577277,15.511708,15.633177,15.752831,15.872487,15.992143,16.1118,14.322405,12.5330105,10.741803,8.952409,7.1630154,8.439341,9.71748,10.995618,12.271944,13.550082,13.684241,13.820213,13.954373,14.090345,14.224504,14.144734,14.064963,13.985193,13.905423,13.825653,13.140353,12.455053,11.769753,11.084454,10.399154,11.294757,12.19036,13.084151,13.979754,14.875358,14.989574,15.105604,15.219821,15.335851,15.4500675,15.937754,16.425442,16.913128,17.400814,17.886688,16.438131,14.9877615,13.537392,12.087022,10.636651,9.53437,8.432089,7.3298078,6.2275267,5.125245,5.243088,5.3591175,5.47696,5.5948024,5.712645,6.1332526,6.552047,6.972654,7.3932614,7.8120556,9.574255,11.338268,13.100468,14.862667,16.624866,19.815681,23.004683,26.195496,29.384497,32.575314,32.713097,32.850883,32.986855,33.124638,33.262424,34.012993,34.761745,35.51231,36.26288,37.01163,40.233265,43.453087,46.67291,49.89273,53.112553,49.675175,46.237797,42.80042,39.363045,35.925667,29.64194,23.360023,17.078108,10.794379,4.512464,4.933071,5.351866,5.772473,6.19308,6.6118746,7.0143523,7.41683,7.819308,8.221786,8.624263,9.815379,11.004683,12.195799,13.385102,14.574407,13.662486,12.750566,11.836833,10.924912,10.012992,10.667472,11.321951,11.978244,12.632723,13.287203,11.234929,9.182655,7.130382,5.0781083,3.0258346,3.6948178,4.365614,5.034597,5.7053933,6.3743763,5.8903155,5.4044414,4.9203806,4.4345064,3.9504454,6.7460337,9.539809,12.335398,15.129172,17.92476,15.872487,13.820213,11.7679405,9.715667,7.663393,6.450521,5.237649,4.024777,2.811905,1.6008459,1.4920682,1.3851035,1.2781386,1.1693609,1.062396,1.6806163,2.2970235,2.9152439,3.531651,4.1498713,3.3195345,2.4891977,1.6606737,0.83033687,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.7650702,1.455809,2.1447346,2.8354735,3.5243993,4.3202896,5.1143675,5.910258,6.7043357,7.500226,7.3298078,7.159389,6.9907837,6.8203654,6.6499467,6.6680765,6.684393,6.7025228,6.720652,6.736969,6.921891,7.1068134,7.2917356,7.476658,7.663393,7.422269,7.1829576,6.9418335,6.7025228,6.4632115,7.0451727,7.6271334,8.210908,8.792869,9.374829,10.837891,12.299138,13.762199,15.22526,16.68832,16.583168,16.478018,16.372866,16.267714,16.162561,17.112555,18.062546,19.012539,19.96253,20.912523,19.879135,18.847559,17.81417,16.782595,15.749206,15.332225,14.915243,14.498261,14.079468,13.662486,13.715062,13.767638,13.820213,13.872789,13.925365,13.675177,13.424988,13.174799,12.92461,12.674421,12.28826,11.900287,11.512312,11.124338,10.738177,11.030065,11.321951,11.615651,11.907538,12.199425,12.707055,13.2146845,13.722314,14.229943,14.737573,15.270584,15.801782,16.334793,16.867804,17.400814,18.813112,20.22541,21.637709,23.050007,24.462305,25.345217,26.22813,27.10923,27.992142,28.875055,28.441757,28.010271,27.576973,27.145489,26.71219,25.87279,25.033388,24.192173,23.352772,22.513369,22.31213,22.112705,21.913279,21.71204,21.512613,22.18341,22.852394,23.52319,24.192173,24.862968,23.802385,22.741802,21.683033,20.62245,19.561867,19.529232,19.4966,19.465778,19.433146,19.400513,19.119503,18.840307,18.559298,18.280102,17.999092,18.45052,18.900135,19.34975,19.799364,20.250792,21.599636,22.950293,24.299137,25.649796,27.000452,27.232512,27.464571,27.696629,27.930502,28.162561,28.313036,28.4617,28.612175,28.762651,28.913128,27.522585,26.132042,24.743313,23.352772,21.962229,22.870523,23.777004,24.685299,25.59178,26.500074,25.727753,24.95543,24.183107,23.410786,22.63665,22.625772,22.613083,22.600391,22.5877,22.57501,20.627888,18.678953,16.731833,14.78471,12.837588,12.407916,11.978244,11.546759,11.117086,10.687414,2.2118144,2.0830941,1.9525607,1.8220274,1.693307,1.5627737,2.1483607,2.7321346,3.3177216,3.9033084,4.4870825,4.606738,4.7282066,4.847862,4.9675174,5.087173,5.384499,5.6818247,5.979151,6.2782893,6.5756154,5.542227,4.510651,3.4772623,2.4456866,1.4122978,1.8528478,2.2915847,2.7321346,3.1726844,3.6132345,4.5251546,5.4370747,6.350808,7.262728,8.174648,8.067683,7.9607186,7.851941,7.744976,7.6380115,8.265296,8.892582,9.519867,10.147152,10.774437,9.438283,8.100317,6.7623506,5.424384,4.0882306,4.748149,5.408067,6.0679855,6.7279043,7.3878226,7.5945,7.802991,8.009668,8.21816,8.424837,8.70222,8.979604,9.256987,9.53437,9.811753,9.5053625,9.197159,8.890768,8.582565,8.274362,7.6942134,7.115878,6.53573,5.955582,5.375434,6.3725634,7.369693,8.366822,9.365765,10.362894,10.429974,10.497053,10.564133,10.633025,10.700105,10.007553,9.3150015,8.62245,7.9298983,7.2373466,6.412449,5.5875506,4.762653,3.9377546,3.1128569,2.9424384,2.7720199,2.6016014,2.4329958,2.2625773,2.2553256,2.2480736,2.2408218,2.231757,2.2245052,2.8372865,3.4500678,4.062849,4.6756306,5.2865987,5.47696,5.667321,5.857682,6.0480433,6.2384043,5.4153194,4.592234,3.7691493,2.9478772,2.124792,1.9507477,1.7748904,1.6008459,1.4249886,1.2491312,1.5917811,1.9344311,2.277081,2.619731,2.962381,2.752077,2.5417736,2.333283,2.1229792,1.9126755,2.1773682,2.4420607,2.7067533,2.9732587,3.2379513,4.499773,5.7615952,7.02523,8.287052,9.550687,11.129777,12.710681,14.289771,15.870674,17.449764,17.92476,18.399757,18.874754,19.34975,19.824745,25.642542,31.46034,37.278137,43.095932,48.91192,44.937904,40.96208,36.988064,33.012238,29.038221,28.197006,27.357605,26.518204,25.676989,24.837587,22.509743,20.1819,17.854055,15.528025,13.200181,13.321649,13.44493,13.568212,13.68968,13.812962,13.812962,13.812962,13.812962,13.812962,13.812962,14.413053,15.013144,15.613234,16.213324,16.811602,15.810846,14.808278,13.80571,12.803142,11.800573,11.214987,10.629399,10.045626,9.460039,8.874452,9.659465,10.444477,11.22949,12.0145035,12.799516,13.472125,14.144734,14.817343,15.489952,16.162561,15.845293,15.528025,15.210756,14.891675,14.574407,13.985193,13.394168,12.804955,12.215742,11.624716,12.444175,13.265448,14.084907,14.904366,15.725637,15.290526,14.855415,14.420304,13.985193,13.550082,14.55265,15.555219,16.557787,17.560356,18.562923,17.072668,15.582414,14.092158,12.601903,11.111648,11.030065,10.946668,10.865085,10.781689,10.700105,11.176914,11.655537,12.132345,12.609155,13.087777,11.405348,9.7229185,8.040489,6.35806,4.6756306,4.175253,3.6748753,3.1744974,2.6741197,2.175555,1.7803292,1.3851035,0.9898776,0.5946517,0.19942589,0.89922947,1.6008459,2.3006494,3.000453,3.7002566,4.329355,4.9602656,5.5893636,6.2202744,6.849373,5.8866897,4.9258194,3.9631362,3.000453,2.03777,3.8126602,5.5875506,7.362441,9.137331,10.912222,10.420909,9.927783,9.434657,8.943344,8.450218,7.9770355,7.5056653,7.0324817,6.5592985,6.0879283,6.0879283,6.0879283,6.0879283,6.0879283,6.0879283,5.3573046,4.6266804,3.8978696,3.1672456,2.4366217,1.9579996,1.4775645,0.99712944,0.5166943,0.038072214,3.149116,6.261973,9.374829,12.487686,15.600543,15.575162,15.54978,15.524399,15.50083,15.475449,12.609155,9.744674,6.880193,4.0157123,1.1494182,1.9851941,2.819157,3.6549325,4.4907084,5.3246713,7.454902,9.585134,11.715364,13.845595,15.975826,16.584982,17.194138,17.805105,18.41426,19.025229,16.541471,14.059525,11.5775795,9.0956335,6.6118746,8.245354,9.87702,11.510499,13.142166,14.775645,14.643299,14.50914,14.376793,14.244447,14.112101,13.310771,12.507628,11.704487,10.903157,10.100015,9.3567,8.615198,7.8718834,7.130382,6.3870673,7.072367,7.757667,8.442966,9.128266,9.811753,11.019187,12.22662,13.435865,14.643299,15.850732,16.563227,17.27572,17.988214,18.700708,19.413204,17.27572,15.138238,13.000754,10.863272,8.725789,7.6924005,6.6608243,5.6274357,4.59586,3.5624714,3.9903307,4.41819,4.844236,5.272095,5.6999545,5.9845896,6.2692246,6.5556726,6.8403077,7.124943,9.300498,11.47424,13.649796,15.825351,17.999092,21.795437,25.589968,29.384497,33.18084,36.975372,36.699802,36.424232,36.150475,35.874905,35.599335,36.250187,36.899227,37.55008,38.199123,38.849976,41.310165,43.770355,46.230545,48.690735,51.149113,47.77519,44.399452,41.02553,37.649796,34.27587,28.32754,22.381023,16.432693,10.484363,4.537845,4.8097897,5.081734,5.3554916,5.6274357,5.89938,6.6209393,7.3406854,8.0604315,8.780178,9.499924,10.17072,10.839704,11.510499,12.179482,12.850279,12.574709,12.299138,12.025381,11.74981,11.47424,11.876718,12.279196,12.681673,13.084151,13.486629,11.142468,8.798307,6.452334,4.1081734,1.7621996,3.1092308,4.458075,5.805106,7.1521373,8.499168,7.382384,6.265599,5.147001,4.0302157,2.911618,6.0843024,9.256987,12.429671,15.602356,18.77504,16.21695,13.660673,11.102583,8.544493,5.9882154,4.974769,3.9631362,2.94969,1.938057,0.9246109,0.9644961,1.0043813,1.0442665,1.0841516,1.1258497,1.7658255,2.4058013,3.045777,3.6857529,4.325729,3.4591327,2.5943494,1.7295663,0.86478317,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.533011,1.0279498,1.5228885,2.0178273,2.5127661,3.147303,3.7818398,4.41819,5.0527267,5.6872635,5.7779117,5.866747,5.957395,6.0480433,6.1368785,6.33993,6.542982,6.7442207,6.947273,7.1503243,7.5419245,7.935337,8.326937,8.72035,9.11195,8.667774,8.221786,7.7776093,7.3316207,6.887445,7.5981264,8.306994,9.017676,9.728357,10.437225,12.250188,14.06315,15.8743,17.687263,19.500225,18.959963,18.4197,17.879436,17.339174,16.800724,18.17495,19.549175,20.925215,22.29944,23.675478,22.589514,21.505362,20.419397,19.335245,18.24928,17.621996,16.99471,16.367426,15.740141,15.112856,14.895301,14.677745,14.46019,14.242634,14.025079,13.575464,13.125849,12.674421,12.224807,11.775192,11.525003,11.274815,11.024626,10.774437,10.524248,10.903157,11.280253,11.65735,12.034446,12.413355,13.022511,13.631665,14.242634,14.851789,15.462758,15.772775,16.08279,16.392807,16.702824,17.01284,18.838493,20.662334,22.487988,24.311829,26.137482,26.772018,27.40837,28.042906,28.677443,29.31198,28.115423,26.917055,25.7205,24.522131,23.325577,22.96661,22.609457,22.252302,21.89515,21.537996,21.44916,21.362139,21.275116,21.188093,21.099258,21.48542,21.869768,22.254116,22.640276,23.024624,21.545248,20.06587,18.584679,17.105303,15.624111,15.877926,16.129929,16.38193,16.635744,16.887747,16.985647,17.081734,17.179634,17.277533,17.375433,17.33736,17.29929,17.26303,17.224958,17.186886,18.925516,20.662334,22.400965,24.137783,25.874601,26.27164,26.670492,27.067532,27.464571,27.861609,27.937754,28.012085,28.08823,28.162561,28.236893,26.630608,25.022509,23.414412,21.808126,20.20003,21.322252,22.444477,23.5667,24.690737,25.812962,24.7832,23.751623,22.72186,21.692097,20.662334,19.587248,18.512161,17.437075,16.361988,15.2869005,13.907236,12.527572,11.147907,9.768243,8.386765,8.3595705,8.3323765,8.3051815,8.2779875,8.2507925,2.0631514,1.7748904,1.4866294,1.2001812,0.9119202,0.62547207,1.1874905,1.7495089,2.3133402,2.8753586,3.437377,3.7999697,4.162562,4.5251546,4.8877473,5.2503395,5.337362,5.424384,5.5132194,5.600241,5.6872635,4.7118897,3.738329,2.762955,1.7875811,0.8122072,1.4122978,2.0123885,2.612479,3.2125697,3.8126602,4.762653,5.712645,6.6626377,7.61263,8.562622,8.287052,8.013294,7.7377243,7.462154,7.1883965,8.2507925,9.313189,10.375585,11.437981,12.500377,10.725487,8.950596,7.175706,5.4008155,3.6241121,4.12449,4.6248674,5.125245,5.6256227,6.1241875,6.688019,7.250037,7.8120556,8.375887,8.937905,9.188094,9.438283,9.686659,9.936848,10.1870365,9.800876,9.412902,9.024928,8.636953,8.2507925,7.474845,6.70071,5.924762,5.1506267,4.3746786,5.487838,6.599184,7.7123427,8.825501,9.936848,9.862516,9.788185,9.712041,9.637709,9.563377,9.099259,8.636953,8.174648,7.7123427,7.250037,6.1749506,5.0998635,4.024777,2.94969,1.8746033,1.8619126,1.8492218,1.8383441,1.8256533,1.8129625,1.7132497,1.6117238,1.5120108,1.4122978,1.3125849,1.9126755,2.5127661,3.1128569,3.7129474,4.313038,4.699199,5.087173,5.475147,5.863121,6.249282,5.388125,4.5251546,3.6621845,2.7992141,1.938057,1.7368182,1.5373923,1.3379664,1.1367276,0.93730164,1.3869164,1.8383441,2.2879589,2.7375734,3.1871881,2.9243085,2.663242,2.4003625,2.137483,1.8746033,1.9743162,2.0758421,2.175555,2.275268,2.374981,3.7999697,5.224958,6.6499467,8.074935,9.499924,10.88684,12.27557,13.662486,15.049402,16.438131,17.199575,17.962833,18.724277,19.487535,20.250792,26.44931,32.649643,38.849976,45.05031,51.25064,47.24943,43.250034,39.25064,35.24943,31.250036,30.374374,29.500526,28.624866,27.749205,26.875357,24.199425,21.525305,18.849373,16.175253,13.499319,13.77489,14.05046,14.324218,14.599788,14.875358,14.811904,14.750263,14.68681,14.625169,14.561715,15.363045,16.162561,16.962078,17.763407,18.562923,17.500528,16.438131,15.375735,14.313339,13.24913,12.4242325,11.599335,10.774437,9.949538,9.12464,9.924157,10.725487,11.525003,12.32452,13.125849,13.662486,14.199123,14.737573,15.27421,15.812659,15.56247,15.312282,15.062093,14.811904,14.561715,13.861912,13.162108,12.462305,11.762501,11.062697,12.012691,12.962683,13.912675,14.862667,15.812659,15.363045,14.911617,14.462003,14.012388,13.562773,14.425743,15.2869005,16.14987,17.01284,17.87581,16.525154,15.174497,13.825653,12.474996,11.124338,10.850581,10.57501,10.29944,10.025683,9.750113,10.613083,11.47424,12.337211,13.200181,14.06315,11.961927,9.862516,7.763106,5.661882,3.5624714,2.8753586,2.1882458,1.49932,0.8122072,0.12509441,0.15047589,0.17585737,0.19942589,0.22480737,0.25018883,1.1258497,1.9996977,2.8753586,3.7492065,4.6248674,5.087173,5.5494785,6.011784,6.4759026,6.9382076,6.000906,5.0617914,4.12449,3.1871881,2.2498865,4.2006345,6.149569,8.100317,10.049252,11.999999,11.274815,10.549629,9.824444,9.099259,8.375887,7.900891,7.4258947,6.9490857,6.474089,6.000906,5.5494785,5.0998635,4.650249,4.2006345,3.7492065,3.2506418,2.7502642,2.2498865,1.7495089,1.2491312,1.0007553,0.7505665,0.50037766,0.25018883,0.0,3.2125697,6.4251394,9.637709,12.850279,16.062849,16.124489,16.187943,16.249584,16.313038,16.374678,13.225562,10.074633,6.925517,3.774588,0.62547207,1.4630609,2.3006494,3.1382382,3.975827,4.8116026,7.137634,9.461852,11.787883,14.112101,16.438131,17.536787,18.637255,19.737724,20.838192,21.936848,18.76235,15.5878525,12.411542,9.237044,6.0625467,8.049554,10.036561,12.025381,14.012388,15.999394,15.600543,15.199879,14.799213,14.400362,13.999697,12.474996,10.950294,9.425592,7.899078,6.3743763,5.57486,4.7753434,3.975827,3.1744974,2.374981,2.8499773,3.3249733,3.7999697,4.274966,4.749962,7.0506115,9.349448,11.650098,13.9507475,16.249584,17.186886,18.124187,19.063301,20.000603,20.937904,18.111496,15.2869005,12.462305,9.637709,6.813113,5.8504305,4.8877473,3.925064,2.962381,1.9996977,2.7375734,3.4754493,4.213325,4.949388,5.6872635,5.8377395,5.9882154,6.1368785,6.2873545,6.43783,9.024928,11.612025,14.200936,16.788034,19.375132,23.77519,28.175251,32.575314,36.975372,41.37543,40.68832,39.999393,39.31228,38.625168,37.938053,38.48738,39.03671,39.587852,40.13718,40.68832,42.387066,44.087624,45.78818,47.486927,49.18749,45.875206,42.562923,39.25064,35.93836,32.62426,27.01133,21.40021,15.787278,10.174346,4.5632267,4.688321,4.8116026,4.936697,5.0617914,5.186886,6.2257137,7.262728,8.299743,9.336758,10.375585,10.524248,10.674724,10.825199,10.975676,11.124338,11.486931,11.849524,12.212116,12.574709,12.937301,13.087777,13.238253,13.386916,13.537392,13.687867,11.050007,8.412147,5.774286,3.1382382,0.50037766,2.525457,4.550536,6.5756154,8.600695,10.625773,8.874452,7.124943,5.375434,3.6241121,1.8746033,5.424384,8.974165,12.525759,16.075539,19.62532,16.561413,13.499319,10.437225,7.3751316,4.313038,3.5008307,2.6868105,1.8746033,1.062396,0.25018883,0.43692398,0.62547207,0.8122072,1.0007553,1.1874905,1.8492218,2.5127661,3.1744974,3.8380418,4.499773,3.6005437,2.6995013,1.8002719,0.89922947,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.2991388,0.6000906,0.89922947,1.2001812,1.49932,1.9743162,2.4493124,2.9243085,3.3993049,3.874301,4.2242026,4.574105,4.9258194,5.275721,5.6256227,6.011784,6.399758,6.787732,7.175706,7.5618668,8.161958,8.762048,9.362139,9.96223,10.56232,9.91328,9.262425,8.613385,7.9625316,7.311678,8.149267,8.9868555,9.824444,10.662033,11.499621,13.662486,15.825351,17.988214,20.149265,22.31213,21.336756,20.363195,19.387821,18.412449,17.437075,19.237347,21.037619,22.837889,24.63816,26.43662,25.299892,24.163166,23.024624,21.887897,20.749357,19.911768,19.074179,18.236591,17.400814,16.563227,16.075539,15.5878525,15.100165,14.612478,14.124791,13.475751,12.824898,12.175857,11.525003,10.874149,10.761745,10.649343,10.536939,10.424535,10.312131,10.774437,11.236742,11.700861,12.163166,12.625471,13.337966,14.05046,14.762955,15.475449,16.187943,16.274965,16.361988,16.450823,16.537846,16.624866,18.862062,21.099258,23.338266,25.575462,27.812658,28.200632,28.586794,28.974768,29.362741,29.750715,27.787277,25.825651,23.862213,21.900587,19.93715,20.062244,20.187338,20.312433,20.437527,20.562622,20.588003,20.613384,20.636953,20.662334,20.687716,20.78743,20.887142,20.986855,21.08838,21.188093,19.288109,17.388124,15.488139,13.588155,11.6881695,12.224807,12.763257,13.299893,13.838344,14.37498,14.849977,15.324973,15.799969,16.274965,16.749962,16.224201,15.700256,15.174497,14.650551,14.124791,16.249584,18.374376,20.499168,22.625772,24.750565,25.312584,25.874601,26.43662,27.000452,27.56247,27.56247,27.56247,27.56247,27.56247,27.56247,25.736816,23.912977,22.087322,20.263483,18.43783,19.775795,21.11195,22.449915,23.787882,25.125849,23.836832,22.54963,21.262424,19.975222,18.688019,16.550535,14.413053,12.27557,10.138086,8.000604,7.1865835,6.3743763,5.562169,4.749962,3.9377546,4.313038,4.688321,5.0617914,5.4370747,5.812358,2.8372865,2.4801328,2.1229792,1.7658255,1.4068589,1.0497054,1.4648738,1.8800422,2.2952106,2.7103791,3.1255474,3.4101827,3.6948178,3.9794528,4.265901,4.550536,4.7771564,5.0055895,5.23221,5.4606433,5.6872635,4.7155156,3.7419548,2.770207,1.7966459,0.824898,1.7295663,2.6342347,3.540716,4.445384,5.3500524,5.9519563,6.5556726,7.157576,7.75948,8.363196,8.10213,7.842876,7.5818095,7.322556,7.063302,7.7848616,8.508233,9.229793,9.953164,10.674724,9.2606125,7.844689,6.430578,5.0146546,3.6005437,4.0302157,4.459888,4.88956,5.319232,5.750717,6.147756,6.544795,6.9418335,7.3406854,7.7377243,7.987913,8.238102,8.488291,8.736667,8.9868555,8.945157,8.901647,8.859948,8.81825,8.774739,7.844689,6.9146395,5.9845896,5.0545397,4.12449,5.2503395,6.3743763,7.500226,8.624263,9.750113,9.585134,9.420154,9.255174,9.090195,8.925215,8.363196,7.799365,7.2373466,6.6753283,6.11331,5.315606,4.517903,3.720199,2.9224956,2.124792,2.079468,2.034144,1.9906329,1.9453088,1.8999848,1.7767034,1.6552348,1.5319533,1.4104849,1.2872034,2.0250793,2.762955,3.5008307,4.2368937,4.974769,5.0001507,5.0255322,5.049101,5.0744824,5.0998635,4.3946214,3.6893787,2.9841363,2.280707,1.5754645,1.4231756,1.2708868,1.1167849,0.9644961,0.8122072,1.1747998,1.5373923,1.8999848,2.2625773,2.6251698,2.467442,2.3097143,2.1519866,1.9942589,1.8383441,2.1102884,2.382233,2.6541772,2.9279346,3.199879,4.5269675,5.8540564,7.1829576,8.510046,9.837135,11.325577,12.812206,14.300649,15.787278,17.27572,18.577427,19.879135,21.182655,22.484362,23.787882,28.202446,32.61701,37.033386,41.447952,45.862514,42.998035,40.13174,37.267258,34.40278,31.538298,30.260159,28.98202,27.705694,26.427555,25.149418,22.859646,20.569874,18.280102,15.99033,13.700559,14.188245,14.674119,15.161806,15.649493,16.13718,15.879739,15.622298,15.364858,15.107417,14.849977,15.40293,15.955884,16.507025,17.059978,17.612932,16.777155,15.9431925,15.107417,14.271642,13.437678,12.581961,11.728055,10.872336,10.016619,9.162713,9.6504,10.138086,10.625773,11.111648,11.599335,12.291886,12.984438,13.67699,14.369541,15.062093,14.953316,14.842725,14.732134,14.623356,14.512766,14.157425,13.802084,13.446743,13.093216,12.737875,13.21831,13.696932,14.177367,14.657803,15.138238,14.73576,14.333282,13.930804,13.528327,13.125849,13.820213,14.514579,15.210756,15.905121,16.599485,15.760084,14.920682,14.079468,13.240066,12.400664,12.474996,12.549327,12.625471,12.699803,12.774135,12.74694,12.719746,12.692551,12.665357,12.638163,10.689227,8.7421055,6.794984,4.847862,2.9007401,2.5055144,2.1102884,1.7150626,1.3198367,0.9246109,0.9554313,0.98443866,1.015259,1.0442665,1.0750868,1.6171626,2.1592383,2.7031271,3.245203,3.787279,4.401873,5.0182805,5.632875,6.247469,6.8620634,6.1405044,5.4171324,4.695573,3.972201,3.2506418,4.7390842,6.2293396,7.7195945,9.20985,10.700105,10.1054535,9.510801,8.914337,8.319685,7.7250338,7.2482243,6.7696023,6.2927933,5.814171,5.337362,5.2158933,5.092612,4.9693303,4.847862,4.7245803,4.137181,3.5497808,2.962381,2.374981,1.7875811,1.4467441,1.1077201,0.7668832,0.42785916,0.0870222,2.9678197,5.846804,8.727602,11.608399,14.487384,14.389484,14.293397,14.195497,14.097597,13.999697,11.379966,8.760235,6.1405044,3.5207734,0.89922947,1.5754645,2.2498865,2.9243085,3.6005437,4.274966,6.70071,9.12464,11.5503845,13.974316,16.400059,17.368181,18.33449,19.302612,20.270735,21.237043,18.577427,15.917811,13.258195,10.596766,7.93715,9.420154,10.903157,12.384347,13.867351,15.350354,14.657803,13.965251,13.272699,12.580148,11.887595,10.654781,9.421967,8.189152,6.9581504,5.7253356,5.1741953,4.6248674,4.07554,3.5243993,2.9750717,3.6658103,4.3547363,5.045475,5.7344007,6.4251394,8.100317,9.775495,11.450671,13.125849,14.799213,15.569723,16.34023,17.11074,17.879436,18.649946,16.22239,13.794832,11.367275,8.939718,6.5121617,6.104245,5.6981416,5.290225,4.882308,4.4743915,5.0744824,5.674573,6.2746634,6.874754,7.474845,7.705091,7.935337,8.165584,8.39583,8.624263,11.245807,13.865538,16.48527,19.105,21.724731,25.085964,28.445383,31.804802,35.164223,38.525455,39.069344,39.615044,40.160748,40.704636,41.25034,41.89938,42.550232,43.199272,43.850124,44.49917,44.859947,45.220726,45.579693,45.94047,46.29944,43.074177,39.85073,36.62547,33.40021,30.17495,25.095028,20.015106,14.935185,9.855265,4.7753434,5.8794374,6.985345,8.089439,9.195346,10.29944,10.304879,10.310318,10.315757,10.319383,10.324821,10.410031,10.49524,10.58045,10.665659,10.750868,11.091705,11.434355,11.777005,12.119655,12.462305,12.493125,12.522133,12.552953,12.581961,12.612781,10.8415165,9.072064,7.3026133,5.5331616,3.7618973,5.2104545,6.6571984,8.105756,9.5525,10.999244,9.211663,7.4258947,5.638314,3.8507326,2.0631514,4.93851,7.8120556,10.687414,13.562773,16.438131,14.097597,11.757062,9.416528,7.077806,4.7372713,3.8851788,3.0330863,2.179181,1.3270886,0.4749962,0.56927025,0.6653573,0.75963134,0.8557183,0.9499924,1.4848163,2.0196402,2.5544643,3.0892882,3.6241121,2.9007401,2.175555,1.4503701,0.72518504,0.0,0.0,0.0,0.0,0.0,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.3825351,0.6526665,0.922798,1.1929294,1.4630609,1.8292793,2.1973107,2.565342,2.9333735,3.299592,3.540716,3.780027,4.019338,4.2604623,4.499773,5.029158,5.560356,6.089741,6.6191263,7.1503243,7.6180687,8.0858135,8.551744,9.019489,9.487233,8.963287,8.437528,7.911769,7.3878226,6.8620634,7.460341,8.056806,8.655084,9.253361,9.849826,11.784257,13.720501,15.654932,17.589363,19.525606,18.546608,17.56942,16.592234,15.6150465,14.63786,16.142618,17.647377,19.152136,20.656897,22.161655,21.262424,20.363195,19.462152,18.562923,17.661882,16.936697,16.213324,15.488139,14.762955,14.037769,13.749508,13.46306,13.174799,12.888351,12.60009,12.222994,11.845898,11.466989,11.089892,10.712796,10.667472,10.622148,10.576823,10.533313,10.487988,10.939416,11.392657,11.845898,12.297325,12.750566,13.464873,14.17918,14.895301,15.609608,16.325727,16.757214,17.190512,17.621996,18.055294,18.48678,20.11482,21.74286,23.370901,24.997128,26.625168,26.617916,26.610664,26.6016,26.594349,26.587097,24.917358,23.24762,21.57788,19.908142,18.236591,18.595556,18.952711,19.309864,19.667019,20.024172,20.044115,20.06587,20.085812,20.105755,20.125698,20.085812,20.044115,20.004229,19.964344,19.92446,18.454145,16.985647,15.515334,14.045021,12.574709,12.839401,13.1059065,13.370599,13.635292,13.899984,14.030518,14.159238,14.289771,14.420304,14.5508375,14.190058,13.829279,13.470312,13.109532,12.750566,14.200936,15.649493,17.099863,18.550234,20.000603,20.464722,20.930653,21.394772,21.860703,22.324821,22.859646,23.394468,23.929293,24.464117,25.000753,23.807825,22.614895,21.421967,20.23085,19.03792,20.713097,22.388275,24.063452,25.736816,27.411995,25.093216,22.772623,20.45203,18.133251,15.812659,14.112101,12.411542,10.712796,9.012237,7.311678,6.622752,5.9320135,5.243088,4.552349,3.8616104,4.177066,4.4925213,4.8079767,5.121619,5.4370747,3.6132345,3.1853752,2.7575161,2.3296568,1.9017978,1.4757515,1.742257,2.0105755,2.277081,2.5453994,2.811905,3.0203958,3.2270734,3.435564,3.6422417,3.8507326,4.216951,4.5849824,4.953014,5.319232,5.6872635,4.7173285,3.7473936,2.7774587,1.8075237,0.8375887,2.0468347,3.2578938,4.4671397,5.678199,6.887445,7.1430726,7.3968873,7.652515,7.9081426,8.161958,7.9172077,7.6724577,7.4277077,7.1829576,6.9382076,7.320743,7.703278,8.0858135,8.4683485,8.8508835,7.795739,6.740595,5.6854506,4.6303062,3.5751622,3.9341288,4.2949085,4.655688,5.0146546,5.375434,5.6074934,5.8395524,6.071612,6.305484,6.5375433,6.787732,7.037921,7.28811,7.5382986,7.7866745,8.089439,8.392203,8.694968,8.997733,9.300498,8.214534,7.130382,6.0444174,4.9602656,3.874301,5.0128417,6.149569,7.28811,8.424837,9.563377,9.30775,9.052122,8.798307,8.54268,8.287052,7.6253204,6.9617763,6.300045,5.638314,4.974769,4.454449,3.9341288,3.4156215,2.8953013,2.374981,2.2970235,2.220879,2.1429217,2.0649643,1.987007,1.84197,1.696933,1.551896,1.4068589,1.261822,2.137483,3.0131438,3.8869917,4.762653,5.638314,5.2992897,4.9620786,4.6248674,4.2876563,3.9504454,3.4029307,2.855416,2.3079014,1.7603867,1.2128719,1.1077201,1.0025684,0.8974165,0.79226464,0.6871128,0.96268314,1.2382535,1.5120108,1.7875811,2.0631514,2.0105755,1.9579996,1.9054236,1.8528478,1.8002719,2.2444477,2.6904364,3.1346123,3.5806012,4.024777,5.2557783,6.484967,7.7141557,8.945157,10.174346,11.762501,13.3506565,14.936998,16.525154,18.11331,19.955278,21.797249,23.63922,25.483002,27.324972,29.955582,32.584377,35.214985,37.845592,40.47439,38.744823,37.01526,35.28569,33.55431,31.824745,30.144129,28.465326,26.78471,25.104094,23.42529,21.519865,19.614443,17.71083,15.805408,13.899984,14.599788,15.299591,15.999394,16.699198,17.400814,16.947575,16.494333,16.042906,15.589665,15.138238,15.442815,15.747393,16.051971,16.358362,16.66294,16.055597,15.448255,14.839099,14.231756,13.6244135,12.739688,11.854962,10.970237,10.085511,9.200785,9.374829,9.550687,9.724731,9.900589,10.074633,10.9230995,11.769753,12.618219,13.464873,14.313339,14.342347,14.373167,14.402175,14.432995,14.462003,14.452938,14.4420595,14.432995,14.422117,14.413053,14.422117,14.432995,14.4420595,14.452938,14.462003,14.106662,13.753134,13.397794,13.042453,12.687112,13.2146845,13.742256,14.269829,14.7974,15.324973,14.995013,14.665054,14.335095,14.005136,13.675177,14.09941,14.525456,14.94969,15.375735,15.799969,14.882609,13.965251,13.047892,12.130532,11.213174,9.418341,7.6216946,5.826862,4.0320287,2.2371957,2.13567,2.032331,1.9308052,1.8274662,1.7241274,1.7603867,1.794833,1.8292793,1.8655385,1.8999848,2.1102884,2.3205922,2.5308957,2.7393866,2.94969,3.7183862,4.4852695,5.2521524,6.0208488,6.787732,6.2801023,5.772473,5.2648435,4.7572136,4.249584,5.279347,6.3091097,7.3406854,8.370448,9.400211,8.934279,8.470161,8.00423,7.5401115,7.07418,6.5955577,6.115123,5.634688,5.1542525,4.6756306,4.880495,5.08536,5.290225,5.4950895,5.6999545,5.0255322,4.349297,3.6748753,3.000453,2.324218,1.8945459,1.4648738,1.0352017,0.6055295,0.17585737,2.72307,5.2702823,7.817495,10.364707,12.91192,12.654479,12.397038,12.139598,11.882156,11.624716,9.53437,7.4458375,5.3554916,3.2651455,1.1747998,1.6878681,2.1991236,2.712192,3.2252605,3.738329,6.261973,8.78743,11.312886,13.838344,16.361988,17.197763,18.031725,18.867502,19.703278,20.537241,18.392506,16.24777,14.103036,11.958302,9.811753,10.790753,11.7679405,12.745127,13.722314,14.699501,13.715062,12.730623,11.744371,10.7599325,9.775495,8.834567,7.895452,6.9545245,6.01541,5.0744824,4.7753434,4.4743915,4.175253,3.874301,3.5751622,4.4798307,5.384499,6.2891674,7.1956487,8.100317,9.1500225,10.199727,11.249433,12.299138,13.3506565,13.95256,14.554463,15.15818,15.760084,16.361988,14.33147,12.302764,10.272246,8.241728,6.2130227,6.359873,6.506723,6.6553855,6.8022356,6.9508986,7.413204,7.8755093,8.337815,8.80012,9.262425,9.572442,9.882459,10.192475,10.502492,10.812509,13.464873,16.117237,18.769602,21.421967,24.07433,26.394922,28.715515,31.034294,33.354885,35.675476,37.452183,39.230698,41.0074,42.785915,44.562622,45.313187,46.06194,46.812508,47.563072,48.31183,47.33283,46.352013,45.373016,44.3922,43.4132,40.274963,37.136726,34.0003,30.862062,27.725637,23.176914,18.630003,14.083094,9.53437,4.98746,7.072367,9.157274,11.242181,13.327088,15.411995,14.385859,13.357908,12.329959,11.302009,10.275872,10.2958145,10.315757,10.3357,10.355642,10.375585,10.698292,11.019187,11.341894,11.664601,11.9873085,11.896661,11.807825,11.717177,11.628342,11.537694,10.634838,9.731983,8.829127,7.9280853,7.02523,7.895452,8.765674,9.635896,10.504305,11.374527,9.550687,7.7250338,5.89938,4.07554,2.2498865,4.4508233,6.6499467,8.8508835,11.050007,13.24913,11.631968,10.014805,8.397643,6.78048,5.163317,4.269527,3.3775494,2.4855716,1.5917811,0.69980353,0.7016165,0.70524246,0.7070554,0.7106813,0.7124943,1.1204109,1.5283275,1.9344311,2.3423476,2.7502642,2.1991236,1.649796,1.1004683,0.5493277,0.0,0.0,0.0,0.0,0.0,0.0,0.045324065,0.09064813,0.13415924,0.1794833,0.22480737,0.46411842,0.70524246,0.9445535,1.1856775,1.4249886,1.6842422,1.9453088,2.2045624,2.465629,2.7248828,2.855416,2.9841363,3.1146698,3.245203,3.3757362,4.0483456,4.7191415,5.391751,6.0643597,6.736969,7.072367,7.407765,7.743163,8.076748,8.412147,8.013294,7.61263,7.211965,6.813113,6.412449,6.7696023,7.1267557,7.4857225,7.842876,8.200029,9.907841,11.615651,13.321649,15.02946,16.73727,15.758271,14.777458,13.796645,12.817645,11.836833,13.047892,14.257137,15.468197,16.677443,17.886688,17.224958,16.563227,15.899682,15.23795,14.574407,13.961625,13.3506565,12.737875,12.125093,11.512312,11.42529,11.338268,11.249433,11.162411,11.075388,10.970237,10.865085,10.7599325,10.654781,10.549629,10.573197,10.594954,10.616709,10.640278,10.662033,11.104396,11.546759,11.989121,12.433297,12.87566,13.591781,14.309713,15.027647,15.74558,16.4617,17.239462,18.017221,18.794983,19.572744,20.350506,21.367577,22.38465,23.401722,24.420607,25.437677,25.0352,24.632723,24.230246,23.827766,23.42529,22.047438,20.669586,19.291735,17.915697,16.537846,17.127058,17.718082,18.307297,18.898321,19.487535,19.502039,19.518354,19.53286,19.547363,19.561867,19.382383,19.2029,19.021603,18.84212,18.662638,17.621996,16.583168,15.542528,14.501887,13.46306,13.455809,13.446743,13.439491,13.43224,13.424988,13.209246,12.995316,12.779573,12.565643,12.349901,12.154101,11.9601145,11.764315,11.570327,11.374527,12.1504755,12.92461,13.700559,14.474693,15.250641,15.616859,15.984891,16.352922,16.719141,17.087172,18.15682,19.228281,20.29793,21.367577,22.437225,21.87702,21.316814,20.756609,20.198215,19.63801,21.650398,23.662788,25.675177,27.687565,29.699953,26.347786,22.993805,19.641636,16.289469,12.937301,11.675479,10.411844,9.1500225,7.8882003,6.624565,6.057108,5.4896507,4.9221935,4.3547363,3.787279,4.0429068,4.2967215,4.552349,4.8079767,5.0617914,4.3873696,3.8906176,3.392053,2.8953013,2.3967366,1.8999848,2.0196402,2.1392958,2.2607644,2.38042,2.5000753,2.6306088,2.759329,2.8898623,3.0203958,3.149116,3.6567454,4.164375,4.6720047,5.179634,5.6872635,4.7191415,3.7528327,2.7847104,1.8165885,0.85027945,2.3641033,3.87974,5.3953767,6.9092,8.424837,8.3323765,8.239915,8.147454,8.054993,7.9625316,7.7322855,7.502039,7.271793,7.0433598,6.813113,6.8548117,6.8983226,6.9400206,6.981719,7.02523,6.3308654,5.634688,4.940323,4.2441454,3.5497808,3.8398547,4.1299286,4.420003,4.710077,5.0001507,5.06723,5.1343102,5.2032027,5.2702823,5.337362,5.5875506,5.8377395,6.0879283,6.338117,6.588306,7.2355337,7.8827615,8.529989,9.177217,9.824444,8.584378,7.344311,6.104245,4.8641787,3.6241121,4.7753434,5.924762,7.07418,8.225411,9.374829,9.030367,8.685904,8.339628,7.995165,7.650702,6.887445,6.1241875,5.3627434,4.599486,3.8380418,3.5951047,3.3521678,3.1092308,2.8681068,2.6251698,2.514579,2.4058013,2.2952106,2.18462,2.0758421,1.9072367,1.7404441,1.5718386,1.405046,1.2382535,2.2498865,3.2633326,4.274966,5.2884116,6.300045,5.600241,4.900438,4.2006345,3.5008307,2.7992141,2.4094272,2.0196402,1.6298534,1.2400664,0.85027945,0.79226464,0.73424983,0.678048,0.6200332,0.5620184,0.7505665,0.93730164,1.1258497,1.3125849,1.49932,1.551896,1.6044719,1.6570477,1.7096237,1.7621996,2.38042,2.9968271,3.6150475,4.233268,4.8496747,5.9827766,7.114065,8.247167,9.380268,10.51337,12.199425,13.887294,15.575162,17.26303,18.950897,21.33313,23.715364,26.097597,28.47983,30.862062,31.706903,32.551743,33.398396,34.243237,35.088078,34.49161,33.89696,33.30231,32.707657,32.113007,30.029913,27.946817,25.865538,23.782444,21.699348,20.180086,18.660824,17.139748,15.620485,14.09941,15.013144,15.925063,16.836983,17.750717,18.662638,18.01541,17.368181,16.719141,16.071913,15.4246855,15.4827,15.540715,15.596917,15.654932,15.712947,15.332225,14.953316,14.572594,14.191871,13.812962,12.897416,11.98187,11.068136,10.152591,9.237044,9.099259,8.963287,8.825501,8.6877165,8.549932,9.5525,10.555068,11.557636,12.5602045,13.562773,13.7331915,13.901797,14.072216,14.242634,14.413053,14.746637,15.082036,15.417434,15.752831,16.08823,15.627737,15.167245,14.706753,14.248073,13.7875805,13.479377,13.172986,12.864782,12.558392,12.250188,12.609155,12.969934,13.330714,13.68968,14.05046,14.229943,14.409427,14.590723,14.770206,14.94969,15.725637,16.499773,17.27572,18.049856,18.825804,17.01828,15.210756,13.403233,11.595709,9.788185,8.145641,6.5030966,4.860553,3.2180085,1.5754645,1.7658255,1.9543737,2.1447346,2.335096,2.525457,2.565342,2.6052272,2.6451125,2.6849976,2.7248828,2.6016014,2.4801328,2.3568513,2.2353828,2.1121013,3.0330863,3.9522583,4.8732433,5.7924156,6.7134004,6.4197006,6.1278133,5.8341136,5.542227,5.2503395,5.81961,6.390693,6.9599633,7.5292335,8.100317,7.764919,7.4295206,7.0941224,6.7605376,6.4251394,5.942891,5.4606433,4.976582,4.494334,4.0120864,4.5450974,5.0781083,5.6093063,6.1423173,6.6753283,5.9120708,5.1506267,4.3873696,3.6241121,2.8626678,2.3423476,1.8220274,1.3017071,0.78319985,0.26287958,2.47832,4.691947,6.9073873,9.122828,11.338268,10.919474,10.502492,10.085511,9.666717,9.249735,7.690587,6.1296263,4.5704784,3.009518,1.4503701,1.8002719,2.1501737,2.5000753,2.8499773,3.199879,5.825049,8.450218,11.075388,13.700559,16.325727,17.027344,17.730774,18.43239,19.13582,19.837437,18.207582,16.57773,14.947877,13.318023,11.6881695,12.15954,12.632723,13.1059065,13.577277,14.05046,12.772322,11.494183,10.217857,8.939718,7.663393,7.0143523,6.3671246,5.719897,5.0726695,4.4254417,4.3746786,4.325729,4.274966,4.2242026,4.175253,5.295664,6.414262,7.5346723,8.655084,9.775495,10.199727,10.625773,11.050007,11.47424,11.900287,12.335398,12.770509,13.20562,13.640731,14.075842,12.442362,10.810696,9.177217,7.5455503,5.9120708,6.6155005,7.317117,8.020547,8.722163,9.425592,9.750113,10.074633,10.399154,10.725487,11.050007,11.439794,11.829581,12.219368,12.609155,13.000754,15.685752,18.37075,21.055748,23.740746,26.425743,27.705694,28.985645,30.265598,31.54555,32.8255,35.83502,38.844536,41.855865,44.865383,47.874905,48.72518,49.575462,50.425743,51.274208,52.12449,49.80571,47.485115,45.164524,42.845745,40.525154,37.473938,34.424534,31.37513,28.325727,25.274511,21.260612,17.2449,13.229188,9.215289,5.199577,8.265296,11.329204,14.394923,17.460642,20.52455,18.465023,16.405499,14.34416,12.284635,10.225109,10.179785,10.13446,10.089137,10.045626,10.000301,10.303066,10.605831,10.906783,11.209548,11.512312,11.302009,11.091705,10.883214,10.672911,10.462607,10.428161,10.391902,10.357455,10.323009,10.28675,10.58045,10.872336,11.164224,11.457924,11.74981,9.8878975,8.024173,6.16226,4.3003473,2.4366217,3.9631362,5.487838,7.0125394,8.537241,10.061942,9.168152,8.272549,7.3769445,6.4831543,5.5875506,4.655688,3.7220123,2.7901495,1.8582866,0.9246109,0.83577573,0.7451276,0.6544795,0.5656443,0.4749962,0.7541924,1.0352017,1.3143979,1.5954071,1.8746033,1.49932,1.1258497,0.7505665,0.37528324,0.0,0.0,0.0,0.0,0.0,0.0,0.06707962,0.13415924,0.2030518,0.27013144,0.33721104,0.5475147,0.75781834,0.968122,1.1766127,1.3869164,1.5392052,1.693307,1.845596,1.9978848,2.1501737,2.1701162,2.1900587,2.2100015,2.229944,2.2498865,3.0657198,3.87974,4.695573,5.5095935,6.3254266,6.526665,6.7297173,6.932769,7.135821,7.3370595,7.063302,6.787732,6.5121617,6.2365913,5.962834,6.0806766,6.1967063,6.3145485,6.432391,6.550234,8.029612,9.510801,10.990179,12.469557,13.9507475,12.968122,11.985496,11.00287,10.020245,9.037619,9.953164,10.866898,11.782444,12.697989,13.611723,13.1874895,12.763257,12.337211,11.912977,11.486931,10.988366,10.487988,9.987611,9.487233,8.9868555,9.099259,9.211663,9.325879,9.438283,9.550687,9.71748,9.884272,10.052877,10.21967,10.388275,10.477111,10.567759,10.658407,10.747242,10.837891,11.269376,11.702674,12.134158,12.567456,13.000754,13.720501,14.440247,15.159993,15.879739,16.599485,17.721708,18.845747,19.96797,21.090193,22.212418,22.620335,23.028252,23.434355,23.842272,24.250187,23.452484,22.654781,21.857077,21.059374,20.26167,19.177519,18.093367,17.007402,15.92325,14.837286,15.660371,16.481644,17.304728,18.127813,18.950897,18.959963,18.97084,18.979906,18.990784,18.999847,18.680767,18.359873,18.04079,17.719896,17.400814,16.789846,16.18069,15.569723,14.960567,14.349599,14.070402,13.789393,13.510198,13.229188,12.949992,12.389787,11.829581,11.269376,10.70917,10.150778,10.119957,10.089137,10.060129,10.029309,10.000301,10.100015,10.199727,10.29944,10.399154,10.500679,10.770811,11.039129,11.30926,11.579392,11.849524,13.455809,15.06028,16.664753,18.269224,19.87551,19.948027,20.020546,20.093063,20.165583,20.238102,22.5877,24.9373,27.2869,29.6365,31.987911,27.602356,23.216799,18.833055,14.447499,10.061942,9.237044,8.412147,7.5872483,6.7623506,5.9374523,5.4932766,5.047288,4.603112,4.157123,3.7129474,3.9069343,4.102734,4.2967215,4.4925213,4.688321,5.163317,4.59586,4.028403,3.4591327,2.8916752,2.324218,2.2970235,2.269829,2.2426348,2.2154403,2.1882458,2.2408218,2.2933977,2.3441606,2.3967366,2.4493124,3.0983531,3.7455807,4.3928084,5.040036,5.6872635,4.7227674,3.7582715,2.7919624,1.8274662,0.8629702,2.6831846,4.501586,6.3218007,8.1420145,9.96223,9.52168,9.082943,8.642392,8.201842,7.763106,7.5473633,7.3316207,7.117691,6.9019485,6.688019,6.390693,6.093367,5.7942286,5.4969025,5.199577,4.8641787,4.5305934,4.195195,3.8597972,3.5243993,3.7455807,3.9649491,4.1843176,4.405499,4.6248674,4.5269675,4.4308805,4.3329806,4.2350807,4.137181,4.3873696,4.6375585,4.8877473,5.137936,5.388125,6.379815,7.3733187,8.365009,9.3567,10.3502035,8.954222,7.560054,6.164073,4.7699046,3.3757362,4.537845,5.6999545,6.8620634,8.024173,9.188094,8.752983,8.317872,7.8827615,7.4476504,7.0125394,6.149569,5.2884116,4.4254417,3.5624714,2.6995013,2.7357605,2.770207,2.8046532,2.8390994,2.8753586,2.7321346,2.5907235,2.4474995,2.3042755,2.1628644,1.9725033,1.7821422,1.5917811,1.403233,1.2128719,2.3622901,3.5117085,4.6629395,5.812358,6.9617763,5.89938,4.836984,3.774588,2.712192,1.649796,1.4177368,1.1856775,0.95180535,0.7197462,0.48768693,0.47680917,0.46774435,0.45686656,0.44780177,0.43692398,0.53663695,0.63816285,0.73787576,0.8375887,0.93730164,1.0950294,1.2527572,1.4104849,1.5682126,1.7241274,2.514579,3.3050308,4.0954823,4.8841214,5.674573,6.7097745,7.744976,8.780178,9.815379,10.850581,12.638163,14.425743,16.213324,18.000906,19.786674,22.70917,25.631664,28.555973,31.476656,34.39915,33.460037,32.520924,31.579996,30.64088,29.699953,30.240215,30.78048,31.320742,31.859192,32.399456,29.915695,27.430124,24.944551,22.460793,19.975222,18.840307,17.705393,16.570478,15.435563,14.300649,15.4246855,16.550535,17.674572,18.800423,19.92446,19.083244,18.240217,17.397188,16.554161,15.712947,15.522586,15.332225,15.141864,14.953316,14.762955,14.610665,14.458377,14.304275,14.151986,13.999697,13.055143,12.11059,11.164224,10.21967,9.275117,8.825501,8.375887,7.9244595,7.474845,7.02523,8.1819,9.340384,10.497053,11.655537,12.812206,13.122223,13.43224,13.742256,14.052273,14.362289,15.0421505,15.722012,16.401873,17.081734,17.761595,16.833357,15.903308,14.973258,14.043208,13.113158,12.852092,12.592838,12.331772,12.072517,11.813264,12.005438,12.197612,12.389787,12.581961,12.774135,13.464873,14.155612,14.844538,15.535276,16.224201,17.350052,18.474089,19.59994,20.725788,21.849825,19.152136,16.454449,13.75676,11.059072,8.363196,6.872941,5.382686,3.8924308,2.4021754,0.9119202,1.3941683,1.8782293,2.3604772,2.8427253,3.3249733,3.3702974,3.4156215,3.4591327,3.5044568,3.5497808,3.094727,2.6396735,2.18462,1.7295663,1.2745126,2.3477864,3.4192474,4.4925213,5.565795,6.637256,6.5592985,6.4831543,6.4051967,6.3272395,6.249282,6.359873,6.4704633,6.5792413,6.6898317,6.8004227,6.5955577,6.390693,6.185828,5.979151,5.774286,5.290225,4.804351,4.3202896,3.834416,3.350355,4.209699,5.0708566,5.9302006,6.789545,7.650702,6.8004227,5.9501433,5.0998635,4.249584,3.3993049,2.7901495,2.179181,1.5700256,0.96087015,0.34990177,2.231757,4.115425,5.99728,7.8791356,9.762803,9.184468,8.607946,8.029612,7.453089,6.874754,5.844991,4.8152285,3.785466,2.7557032,1.7241274,1.9126755,2.0994108,2.2879589,2.474694,2.663242,5.388125,8.113008,10.837891,13.562773,16.287657,16.856926,17.428009,17.99728,18.568363,19.137632,18.022661,16.907688,15.792717,14.677745,13.562773,13.53014,13.497506,13.464873,13.43224,13.399607,11.829581,10.259555,8.689529,7.119504,5.5494785,5.1941376,4.84061,4.4852695,4.1299286,3.774588,3.975827,4.175253,4.3746786,4.574105,4.7753434,6.109684,7.4458375,8.780178,10.114518,11.450671,11.249433,11.050007,10.850581,10.649343,10.449916,10.718235,10.98474,11.253058,11.519565,11.787883,10.553255,9.316814,8.082188,6.8475595,5.612932,6.869315,8.127511,9.385707,10.642091,11.900287,12.087022,12.27557,12.462305,12.650853,12.837588,13.307145,13.776703,14.248073,14.71763,15.187187,17.904818,20.62245,23.34008,26.05771,28.775343,29.014652,29.255777,29.495089,29.7344,29.975523,34.217857,38.46019,42.702522,46.944855,51.187187,52.137177,53.08717,54.037163,54.987156,55.93715,52.276775,48.618217,44.957848,41.297474,37.637104,34.67472,31.712341,28.74996,25.78758,22.8252,19.342497,15.859797,12.377095,8.894395,5.411693,9.458226,13.502945,17.547665,21.592384,25.637104,22.54419,19.453089,16.360174,13.267261,10.174346,10.065568,9.954978,9.844387,9.735609,9.625018,9.907841,10.190662,10.471672,10.754494,11.037316,10.707357,10.377398,10.047439,9.71748,9.38752,10.21967,11.05182,11.885782,12.717933,13.550082,13.265448,12.980812,12.694364,12.409729,12.125093,10.225109,8.325124,6.4251394,4.5251546,2.6251698,3.4754493,4.325729,5.1741953,6.0244746,6.874754,6.7025228,6.530291,6.35806,6.185828,6.011784,5.040036,4.068288,3.094727,2.1229792,1.1494182,0.968122,0.7850128,0.60190356,0.42060733,0.2374981,0.38978696,0.5420758,0.69436467,0.8466535,1.0007553,0.7995165,0.6000906,0.40066472,0.19942589,0.0,0.0,0.0,0.0,0.0,0.0,0.09064813,0.1794833,0.27013144,0.36077955,0.44961473,0.630911,0.8103943,0.9898776,1.1693609,1.3506571,1.3941683,1.4394923,1.4848163,1.5301404,1.5754645,1.4848163,1.3941683,1.305333,1.214685,1.1258497,2.0830941,3.0403383,3.9975824,4.954827,5.9120708,5.9827766,6.051669,6.1223745,6.19308,6.261973,6.11331,5.962834,5.812358,5.661882,5.5132194,5.389938,5.2666564,5.145188,5.0219064,4.900438,6.153195,7.404139,8.656897,9.909654,11.162411,10.177972,9.19172,8.207282,7.2228427,6.2384043,6.8584375,7.476658,8.096691,8.716724,9.336758,9.1500225,8.963287,8.774739,8.588004,8.399456,8.013294,7.6253204,7.2373466,6.849373,6.4632115,6.775041,7.0868707,7.400513,7.7123427,8.024173,8.464723,8.9052725,9.345822,9.784559,10.225109,10.382836,10.540565,10.698292,10.854207,11.011934,11.434355,11.856775,12.279196,12.701616,13.125849,13.847408,14.57078,15.292339,16.01571,16.73727,18.20577,19.672457,21.139143,22.607643,24.07433,23.87309,23.67004,23.466988,23.265749,23.062696,21.869768,20.676838,19.485722,18.292793,17.099863,16.307598,15.515334,14.723069,13.930804,13.136727,14.191871,15.247015,16.30216,17.357304,18.412449,18.417887,18.423326,18.426952,18.43239,18.43783,17.977337,17.516844,17.058165,16.597672,16.13718,15.957697,15.7782135,15.596917,15.417434,15.23795,14.684997,14.132043,13.57909,13.027949,12.474996,11.570327,10.665659,9.759177,8.854509,7.949841,8.0858135,8.219973,8.354132,8.490104,8.624263,8.049554,7.474845,6.9001355,6.3254266,5.750717,5.922949,6.09518,6.2674117,6.439643,6.6118746,8.752983,10.89228,13.033388,15.172684,17.31198,18.017221,18.722466,19.427708,20.13295,20.838192,23.525002,26.213627,28.900436,31.587248,34.27587,28.856926,23.439793,18.022661,12.605529,7.1883965,6.8004227,6.412449,6.0244746,5.638314,5.2503395,4.9276323,4.604925,4.2822175,3.9595103,3.636803,3.7727752,3.9069343,4.0429068,4.177066,4.313038,5.9374523,5.2992897,4.6629395,4.024777,3.386614,2.7502642,2.5744069,2.4003625,2.2245052,2.0504606,1.8746033,1.8492218,1.8256533,1.8002719,1.7748904,1.7495089,2.5381477,3.3249733,4.1117992,4.900438,5.6872635,4.7245803,3.7618973,2.7992141,1.8383441,0.87566096,3.000453,5.125245,7.250037,9.374829,11.499621,10.712796,9.924157,9.137331,8.350506,7.5618668,7.362441,7.1630154,6.9617763,6.7623506,6.5629244,5.924762,5.2884116,4.650249,4.0120864,3.3757362,3.3993049,3.4246864,3.4500678,3.4754493,3.5008307,3.6494937,3.7999697,3.9504454,4.099108,4.249584,3.9867048,3.7256382,3.4627585,3.199879,2.9369993,3.1871881,3.437377,3.6875658,3.9377546,4.1879435,5.524097,6.8620634,8.200029,9.537996,10.874149,9.325879,7.7757964,6.2257137,4.6756306,3.1255474,4.3003473,5.475147,6.6499467,7.8247466,8.999546,8.4756,7.949841,7.424082,6.9001355,6.3743763,5.411693,4.4508233,3.48814,2.525457,1.5627737,1.8746033,2.1882458,2.5000753,2.811905,3.1255474,2.94969,2.7756457,2.5997884,2.4257438,2.2498865,2.03777,1.8256533,1.6117238,1.3996071,1.1874905,2.474694,3.7618973,5.050914,6.338117,7.6253204,6.200332,4.7753434,3.350355,1.9253663,0.50037766,0.42423326,0.34990177,0.2755703,0.19942589,0.12509441,0.16316663,0.19942589,0.2374981,0.2755703,0.31182957,0.3245203,0.33721104,0.34990177,0.36259252,0.37528324,0.63816285,0.89922947,1.162109,1.4249886,1.6878681,2.6505513,3.6132345,4.5759177,5.5367875,6.4994707,7.4367723,8.374074,9.313189,10.25049,11.187792,13.075087,14.96238,16.849674,18.736969,20.624262,24.08702,27.54978,31.012537,34.475296,37.938053,35.213173,32.48829,29.761593,27.03671,24.311829,25.987005,27.662184,29.33736,31.012537,32.687714,29.799665,26.91343,24.025381,21.137331,18.24928,17.500528,16.749962,15.999394,15.250641,14.500074,15.838041,17.174194,18.512161,19.850128,21.188093,20.149265,19.112251,18.075237,17.038223,15.999394,15.56247,15.125546,14.68681,14.249886,13.812962,13.887294,13.961625,14.037769,14.112101,14.188245,13.212872,12.237497,11.262123,10.28675,9.313189,8.549932,7.7866745,7.02523,6.261973,5.5005283,6.813113,8.125698,9.438283,10.750868,12.06164,12.513068,12.962683,13.412297,13.861912,14.313339,15.337664,16.361988,17.388124,18.412449,19.436771,18.037165,16.637558,15.23795,13.838344,12.436923,12.224807,12.012691,11.800573,11.586644,11.374527,11.399909,11.42529,11.450671,11.47424,11.499621,12.699803,13.899984,15.100165,16.300346,17.500528,18.974466,20.450218,21.924156,23.399908,24.87566,21.287807,17.699953,14.112101,10.524248,6.9382076,5.600241,4.262275,2.9243085,1.5881553,0.25018883,1.0243238,1.8002719,2.5744069,3.350355,4.12449,4.175253,4.2242026,4.274966,4.325729,4.3746786,3.587853,2.7992141,2.0123885,1.2255627,0.43692398,1.6624867,2.8880494,4.1117992,5.337362,6.5629244,6.70071,6.836682,6.9744673,7.112252,7.250037,6.9001355,6.550234,6.200332,5.8504305,5.5005283,5.424384,5.3500524,5.275721,5.199577,5.125245,4.6375585,4.1498713,3.6621845,3.1744974,2.6868105,3.874301,5.0617914,6.249282,7.4367723,8.624263,7.686961,6.7496595,5.812358,4.8750563,3.9377546,3.2379513,2.5381477,1.8383441,1.1367276,0.43692398,1.987007,3.53709,5.087173,6.637256,8.187339,7.4494634,6.7134004,5.975525,5.237649,4.499773,3.9993954,3.5008307,3.000453,2.5000753,1.9996977,2.0250793,2.0504606,2.0758421,2.0994108,2.124792,4.949388,7.7757964,10.600392,13.424988,16.249584,16.68832,17.125244,17.562168,18.000906,18.43783,17.837738,17.237648,16.637558,16.037468,15.437376,14.90074,14.362289,13.825653,13.287203,12.750566,10.88684,9.024928,7.1630154,5.2992897,3.437377,3.3757362,3.3122826,3.2506418,3.1871881,3.1255474,3.5751622,4.024777,4.4743915,4.9258194,5.375434,6.925517,8.4756,10.025683,11.575767,13.125849,12.299138,11.47424,10.649343,9.824444,8.999546,9.099259,9.200785,9.300498,9.400211,9.499924,8.662335,7.8247466,6.987158,6.149569,5.3119802,7.124943,8.937905,10.750868,12.562017,14.37498,14.425743,14.474693,14.525456,14.574407,14.625169,15.174497,15.725637,16.274965,16.824293,17.375433,20.125698,22.87415,25.624413,28.374678,31.12494,30.325424,29.52591,28.724579,27.925062,27.125546,32.600693,38.074028,43.550987,49.024323,54.49947,55.549175,56.600693,57.6504,58.700104,59.74981,54.749657,49.749508,44.749355,39.749203,34.750866,31.875507,29.000149,26.12479,23.249432,20.375887,17.424383,14.474693,11.525003,8.575313,5.6256227,10.651155,15.674874,20.700407,25.725939,30.749659,26.625168,22.500679,18.374376,14.249886,10.125396,9.949538,9.775495,9.599637,9.425592,9.249735,9.512614,9.775495,10.038374,10.29944,10.56232,10.112705,9.663091,9.211663,8.762048,8.312433,10.012992,11.711739,13.412297,15.112856,16.811602,15.950445,15.087475,14.224504,13.363347,12.500377,10.56232,8.624263,6.688019,4.749962,2.811905,2.9877625,3.1618068,3.3376641,3.5117085,3.6875658,4.2368937,4.788034,5.337362,5.8866897,6.43783,5.424384,4.4127507,3.3993049,2.3876717,1.3742256,1.1004683,0.824898,0.5493277,0.2755703,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.11240368,0.22480737,0.33721104,0.44961473,0.5620184,0.7124943,0.8629702,1.0116332,1.162109,1.3125849,1.2491312,1.1874905,1.1258497,1.062396,1.0007553,0.7995165,0.6000906,0.40066472,0.19942589,0.0,1.1004683,2.1991236,3.299592,4.40006,5.5005283,5.4370747,5.375434,5.3119802,5.2503395,5.186886,5.163317,5.137936,5.1125546,5.087173,5.0617914,4.699199,4.3366065,3.975827,3.6132345,3.2506418,4.274966,5.2992897,6.3254266,7.3497505,8.375887,7.3878226,6.399758,5.411693,4.4254417,3.437377,3.7618973,4.0882306,4.4127507,4.7372713,5.0617914,5.1125546,5.163317,5.2122674,5.2630305,5.3119802,5.038223,4.762653,4.4870825,4.213325,3.9377546,4.4508233,4.9620786,5.475147,5.9882154,6.4994707,7.211965,7.9244595,8.636953,9.349448,10.061942,10.28675,10.51337,10.738177,10.962985,11.187792,11.599335,12.012691,12.4242325,12.837588,13.24913,13.974316,14.699501,15.4246855,16.14987,16.875055,18.688019,20.499168,22.31213,24.125093,25.938055,25.125849,24.311829,23.49962,22.687414,21.875206,20.287052,18.700708,17.112555,15.524399,13.938056,13.437678,12.937301,12.436923,11.938358,11.437981,12.725184,14.012388,15.299591,16.586794,17.87581,17.87581,17.87581,17.87581,17.87581,17.87581,17.27572,16.67563,16.075539,15.475449,14.875358,15.125546,15.375735,15.624111,15.8743,16.124489,15.299591,14.474693,13.649796,12.824898,11.999999,10.749055,9.499924,8.2507925,6.9998484,5.750717,6.049856,6.350808,6.6499467,6.9490857,7.250037,5.999093,4.749962,3.5008307,2.2498865,1.0007553,1.0750868,1.1494182,1.2255627,1.2998942,1.3742256,4.0501585,6.7260914,9.400211,12.07433,14.750263,16.08823,17.424383,18.76235,20.100317,21.438282,24.462305,27.488138,30.51216,33.537994,36.562016,30.111496,23.660975,17.212267,10.763558,4.313038,4.361988,4.4127507,4.461701,4.512464,4.5632267,4.361988,4.162562,3.9631362,3.7618973,3.5624714,3.636803,3.7129474,3.787279,3.8616104,3.9377546,5.2992897,4.7372713,4.175253,3.6132345,3.049403,2.4873846,2.3006494,2.1121013,1.9253663,1.7368182,1.550083,1.5319533,1.5156367,1.4975071,1.4793775,1.4630609,2.2245052,2.9877625,3.7492065,4.512464,5.275721,4.512464,3.7492065,2.9877625,2.2245052,1.4630609,3.4174345,5.371808,7.327995,9.282369,11.236742,10.502492,9.768243,9.03218,8.29793,7.5618668,7.4875355,7.413204,7.3370595,7.262728,7.1883965,6.5629244,5.9374523,5.3119802,4.688321,4.062849,3.9051213,3.7473936,3.589666,3.4319382,3.2742105,3.680314,4.0846047,4.4907084,4.894999,5.2992897,4.9076896,4.514277,4.122677,3.729264,3.3376641,3.4591327,3.5824142,3.7056956,3.827164,3.9504454,5.1741953,6.399758,7.6253204,8.8508835,10.074633,8.714911,7.3551893,5.995467,4.6357455,3.2742105,4.3946214,5.5150323,6.635443,7.755854,8.874452,8.317872,7.75948,7.2029004,6.644508,6.0879283,5.121619,4.157123,3.1926272,2.228131,1.261822,1.6008459,1.938057,2.275268,2.612479,2.94969,2.855416,2.759329,2.665055,2.570781,2.474694,2.7357605,2.9950142,3.254268,3.5153344,3.774588,4.2405195,4.704638,5.1705694,5.634688,6.1006193,4.9602656,3.8199122,2.6795588,1.5392052,0.40066472,0.34264994,0.28463513,0.22662032,0.17041849,0.11240368,0.14684997,0.18310922,0.21755551,0.2520018,0.28826106,0.2955129,0.30276474,0.3100166,0.31726846,0.3245203,0.71430725,1.1040943,1.4956942,1.8854811,2.275268,3.1074178,3.9395678,4.7717175,5.6056805,6.43783,7.554615,8.673213,9.789998,10.906783,12.025381,13.555521,15.085662,16.615803,18.144129,19.67427,22.814322,25.954372,29.094423,32.234474,35.374527,32.82006,30.265598,27.70932,25.154856,22.600391,24.290073,25.979753,27.669436,29.359116,31.05061,28.499771,25.950747,23.399908,20.84907,18.300045,17.772472,17.2449,16.717327,16.189756,15.662184,16.494333,17.328297,18.160446,18.992596,19.824745,19.054237,18.285542,17.515032,16.744522,15.975826,15.662184,15.350354,15.036712,14.724882,14.413053,14.282519,14.151986,14.023266,13.892733,13.762199,12.984438,12.206677,11.430729,10.652968,9.875207,9.316814,8.760235,8.201842,7.645263,7.0868707,8.227224,9.367578,10.507931,11.648285,12.786825,13.192928,13.597219,14.003323,14.407614,14.811904,15.702069,16.592234,17.482399,18.372562,19.262728,17.99184,16.722767,15.45188,14.182806,12.91192,12.9427395,12.971747,13.002567,13.033388,13.062395,12.922797,12.783199,12.6417885,12.50219,12.362592,13.290829,14.217253,15.14549,16.071913,17.00015,18.216648,19.43496,20.653269,21.869768,23.088078,19.579996,16.071913,12.565643,9.057561,5.5494785,4.4798307,3.4101827,2.3405347,1.2708868,0.19942589,1.2346275,2.269829,3.3050308,4.3402324,5.375434,5.484212,5.5948024,5.7053933,5.814171,5.924762,5.045475,4.164375,3.2850883,2.4058013,1.5247015,2.4366217,3.350355,4.262275,5.1741953,6.0879283,6.48678,6.887445,7.28811,7.686961,8.087626,7.610817,7.132195,6.6553855,6.1767635,5.6999545,5.5531044,5.4044414,5.2575917,5.1107416,4.9620786,4.4508233,3.9377546,3.4246864,2.911618,2.4003625,3.4283123,4.454449,5.482399,6.510349,7.5382986,6.6608243,5.7833505,4.9040637,4.02659,3.149116,2.960568,2.770207,2.5798457,2.3894846,2.1991236,3.3050308,4.409125,5.5150323,6.6191263,7.7250338,7.1902094,6.6553855,6.1205616,5.5857377,5.049101,5.4497657,5.8504305,6.249282,6.6499467,7.0506115,6.0317264,5.0146546,3.9975824,2.9805105,1.9616255,4.6720047,7.382384,10.092763,12.803142,15.511708,15.6150465,15.718386,15.819912,15.92325,16.024776,15.934128,15.845293,15.754644,15.66581,15.575162,15.335851,15.094727,14.855415,14.614291,14.37498,12.74694,11.120712,9.492672,7.8646317,6.2384043,6.3344913,6.432391,6.530291,6.628191,6.7242785,7.1648283,7.605378,8.045928,8.484665,8.925215,9.7773075,10.629399,11.483305,12.335398,13.1874895,12.574709,11.961927,11.349146,10.738177,10.125396,10.484363,10.845142,11.205922,11.564888,11.925668,11.379966,10.834265,10.290376,9.744674,9.200785,10.667472,12.134158,13.602658,15.0693445,16.537846,16.83517,17.132496,17.429823,17.727148,18.024473,18.809486,19.5945,20.379513,21.164526,21.949537,24.143223,26.335094,28.526966,30.720652,32.91252,32.859947,32.80737,32.754795,32.70222,32.649643,36.884724,41.119804,45.354885,49.589966,53.825047,53.87037,53.915695,53.959206,54.004528,54.049854,49.41411,44.780174,40.144432,35.510498,30.874752,28.532406,26.190058,23.84771,21.505362,19.163015,16.432693,13.702372,10.97205,8.241728,5.5132194,9.644961,13.776703,17.910257,22.042,26.175554,23.057259,19.940775,16.82248,13.704185,10.587702,10.555068,10.522435,10.489801,10.457169,10.424535,10.397341,10.370146,10.342952,10.315757,10.28675,10.491614,10.698292,10.903157,11.108022,11.312886,12.308203,13.301706,14.297023,15.292339,16.287657,15.477262,14.666867,13.858286,13.047892,12.237497,10.337513,8.437528,6.5375433,4.6375585,2.7375734,3.3757362,4.0120864,4.650249,5.2884116,5.924762,6.2275267,6.530291,6.833056,7.135821,7.4367723,6.2257137,5.0128417,3.7999697,2.5870976,1.3742256,1.1022812,0.83033687,0.55839247,0.28463513,0.012690738,0.032633327,0.052575916,0.072518505,0.092461094,0.11240368,0.09064813,0.06707962,0.045324065,0.02175555,0.0,0.0,0.0,0.0,0.0,0.0,0.09064813,0.1794833,0.27013144,0.36077955,0.44961473,0.56927025,0.69073874,0.8103943,0.9300498,1.0497054,1.0007553,0.9499924,0.89922947,0.85027945,0.7995165,0.6399758,0.48043507,0.3208944,0.15954071,0.0,0.88291276,1.7658255,2.6469254,3.529838,4.4127507,4.3982472,4.3819304,4.367427,4.3529234,4.3366065,4.3003473,4.262275,4.2242026,4.1879435,4.1498713,3.8416677,3.5352771,3.2270734,2.9206827,2.612479,3.4301252,4.2477713,5.0654173,5.883064,6.70071,5.9845896,5.2702823,4.554162,3.8398547,3.1255474,3.3122826,3.5008307,3.6875658,3.874301,4.062849,4.102734,4.1426196,4.1825047,4.2223897,4.262275,4.0392804,3.8180993,3.5951047,3.3721104,3.149116,3.6096084,4.070101,4.5305934,4.989273,5.4497657,6.149569,6.849373,7.549176,8.2507925,8.950596,9.117389,9.284182,9.452786,9.619579,9.788185,10.094576,10.40278,10.70917,11.017374,11.325577,12.005438,12.685299,13.36516,14.045021,14.724882,16.22239,17.719896,19.217403,20.71491,22.212418,21.626831,21.043056,20.45747,19.871883,19.288109,17.805105,16.322102,14.839099,13.357908,11.874905,11.499621,11.124338,10.750868,10.375585,10.000301,11.195044,12.389787,13.584529,14.779271,15.975826,15.979452,15.984891,15.99033,15.995769,15.999394,15.363045,14.724882,14.0867195,13.45037,12.812206,12.91192,13.011633,13.113158,13.212872,13.312584,12.701616,12.092461,11.483305,10.872336,10.263181,9.162713,8.062244,6.9617763,5.863121,4.762653,4.98746,5.2122674,5.4370747,5.661882,5.8866897,4.876869,3.8670492,2.857229,1.8474089,0.8375887,0.89560354,0.95180535,1.0098201,1.067835,1.1258497,3.2633326,5.4008155,7.5382986,9.673968,11.813264,13.064208,14.316965,15.569723,16.82248,18.075237,20.410334,22.745428,25.080524,27.41562,29.750715,24.552952,19.355188,14.157425,8.9596615,3.7618973,3.9431937,4.122677,4.3021603,4.4816437,4.6629395,4.4725785,4.2822175,4.0918565,3.9033084,3.7129474,3.7147603,3.7183862,3.720199,3.7220123,3.7256382,4.6629395,4.175253,3.6875658,3.199879,2.712192,2.2245052,2.0250793,1.8256533,1.6244144,1.4249886,1.2255627,1.214685,1.2056202,1.1947423,1.1856775,1.1747998,1.9126755,2.6505513,3.386614,4.12449,4.8623657,4.3003473,3.738329,3.1744974,2.612479,2.0504606,3.834416,5.620184,7.405952,9.189907,10.975676,10.292189,9.610515,8.927028,8.245354,7.5618668,7.61263,7.663393,7.7123427,7.763106,7.8120556,7.1992745,6.588306,5.975525,5.3627434,4.749962,4.409125,4.070101,3.729264,3.39024,3.049403,3.7093215,4.36924,5.029158,5.6908894,6.350808,5.826862,5.3047285,4.782595,4.2604623,3.738329,3.73289,3.727451,3.7220123,3.7183862,3.7129474,4.8242936,5.9374523,7.0506115,8.161958,9.275117,8.105756,6.9345818,5.765221,4.59586,3.4246864,4.4907084,5.5549173,6.6191263,7.6851482,8.749357,8.160145,7.569119,6.979906,6.390693,5.7996674,4.8333583,3.8652363,2.8971143,1.9308052,0.96268314,1.3252757,1.6878681,2.0504606,2.4130533,2.7756457,2.759329,2.7448254,2.7303216,2.715818,2.6995013,3.4319382,4.164375,4.896812,5.6292486,6.3616858,6.004532,5.6473784,5.290225,4.933071,4.574105,3.720199,2.864481,2.0105755,1.1548572,0.2991388,0.25925365,0.21936847,0.1794833,0.13959812,0.099712946,0.13234627,0.16497959,0.19761293,0.23024625,0.26287958,0.26469254,0.26831847,0.27013144,0.27194437,0.2755703,0.79226464,1.310772,1.8274662,2.3441606,2.8626678,3.5642843,4.267714,4.9693303,5.67276,6.3743763,7.6724577,8.970539,10.266808,11.564888,12.862969,14.034143,15.20713,16.380117,17.553104,18.724277,21.541622,24.360779,27.178122,29.995466,32.81281,30.42695,28.042906,25.657047,23.273,20.887142,22.59314,24.297325,26.003323,27.707508,29.411692,27.199877,24.988064,22.774435,20.562622,18.350807,18.044416,17.73984,17.43526,17.130684,16.824293,17.15244,17.480585,17.80692,18.135065,18.463211,17.959208,17.457016,16.954826,16.452635,15.950445,15.761897,15.575162,15.386614,15.199879,15.013144,14.677745,14.342347,14.006948,13.673364,13.337966,12.757817,12.17767,11.597522,11.017374,10.437225,10.085511,9.731983,9.380268,9.026741,8.675026,9.643148,10.609457,11.5775795,12.545701,13.512011,13.872789,14.231756,14.592536,14.953316,15.312282,16.068287,16.82248,17.576672,18.332678,19.08687,17.94833,16.807976,15.667623,14.527269,13.386916,13.660673,13.932617,14.204562,14.478319,14.750263,14.445685,14.139296,13.834718,13.53014,13.225562,13.880041,14.534521,15.190813,15.845293,16.499773,17.460642,18.4197,19.38057,20.339626,21.300497,17.872185,14.445685,11.017374,7.5890613,4.162562,3.3594196,2.5580902,1.7549478,0.95180535,0.15047589,1.4449311,2.7393866,4.0356545,5.33011,6.624565,6.794984,6.965402,7.135821,7.304426,7.474845,6.5030966,5.529536,4.557788,3.584227,2.612479,3.2125697,3.8126602,4.4127507,5.0128417,5.612932,6.2746634,6.9382076,7.5999393,8.26167,8.925215,8.319685,7.7141557,7.1104393,6.5049095,5.89938,5.6800117,5.4606433,5.239462,5.0200934,4.800725,4.262275,3.7256382,3.1871881,2.6505513,2.1121013,2.9805105,3.8471067,4.7155156,5.582112,6.450521,5.632875,4.8152285,3.9975824,3.1799364,2.3622901,2.6831846,3.002266,3.3231604,3.6422417,3.9631362,4.6230545,5.282973,5.942891,6.60281,7.262728,6.929143,6.5973706,6.265599,5.9320135,5.600241,6.9001355,8.200029,9.499924,10.799818,12.099712,10.040187,7.9806614,5.919323,3.8597972,1.8002719,4.3946214,6.9907837,9.585134,12.179482,14.775645,14.541773,14.309713,14.077655,13.845595,13.611723,14.0323305,14.452938,14.871732,15.292339,15.712947,15.769149,15.827164,15.885179,15.9431925,15.999394,14.607039,13.2146845,11.822329,10.429974,9.037619,9.295059,9.5525,9.80994,10.067381,10.324821,10.754494,11.184166,11.615651,12.045323,12.474996,12.63091,12.785012,12.939114,13.095029,13.24913,12.850279,12.449615,12.050762,11.650098,11.249433,11.869466,12.489499,13.109532,13.729566,14.349599,14.097597,13.845595,13.591781,13.339779,13.087777,14.210001,15.332225,16.454449,17.576672,18.700708,19.244598,19.7903,20.334188,20.87989,21.425592,22.444477,23.465176,24.485872,25.504757,26.525455,28.160748,29.794228,31.42952,33.06481,34.700104,35.39447,36.090645,36.78501,37.479374,38.175552,41.170567,44.16558,47.160595,50.15561,53.150623,52.189754,51.230698,50.269825,49.31077,48.3499,44.08037,39.810844,35.539505,31.26998,27.000452,25.189302,23.379965,21.57063,19.75948,17.950142,15.439189,12.930049,10.419096,7.909956,5.4008155,8.640579,11.880343,15.120108,18.359873,21.599636,19.489347,17.380873,15.270584,13.1602955,11.050007,11.160598,11.269376,11.379966,11.490557,11.599335,11.282066,10.964798,10.64753,10.330261,10.012992,10.872336,11.731681,12.592838,13.452183,14.313339,14.603414,14.891675,15.181748,15.471823,15.761897,15.004078,14.248073,13.490254,12.732436,11.974618,10.112705,8.2507925,6.3870673,4.5251546,2.663242,3.7618973,4.8623657,5.962834,7.063302,8.161958,8.21816,8.272549,8.326937,8.383139,8.437528,7.02523,5.612932,4.2006345,2.7883365,1.3742256,1.1040943,0.83577573,0.5656443,0.2955129,0.025381476,0.03988518,0.054388877,0.07070554,0.08520924,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0,0.0,0.0,0.0,0.0,0.06707962,0.13415924,0.2030518,0.27013144,0.33721104,0.42785916,0.5166943,0.6073425,0.6979906,0.7868258,0.7505665,0.7124943,0.6744221,0.63816285,0.6000906,0.48043507,0.36077955,0.23931105,0.11965553,0.0,0.6653573,1.3307146,1.9942589,2.659616,3.3249733,3.3576066,3.39024,3.4228733,3.4555066,3.48814,3.437377,3.386614,3.3376641,3.2869012,3.2379513,2.9841363,2.7321346,2.4801328,2.228131,1.9743162,2.5852847,3.1944401,3.8054085,4.4145637,5.0255322,4.5831695,4.1408067,3.6966307,3.254268,2.811905,2.8626678,2.911618,2.962381,3.0131438,3.0620937,3.092914,3.1219215,3.152742,3.1817493,3.2125697,3.0421512,2.8717327,2.7031271,2.5327086,2.3622901,2.770207,3.1781235,3.584227,3.9921436,4.40006,5.087173,5.774286,6.4632115,7.1503243,7.837437,7.948028,8.056806,8.167397,8.2779875,8.386765,8.589817,8.792869,8.994107,9.197159,9.400211,10.034748,10.669285,11.3056345,11.940171,12.574709,13.75676,14.940624,16.122677,17.304728,18.48678,18.129625,17.772472,17.41532,17.058165,16.699198,15.32316,13.945308,12.567456,11.189605,9.811753,9.561564,9.313189,9.063,8.812811,8.562622,9.664904,10.767185,11.869466,12.971747,14.075842,14.084907,14.095784,14.104849,14.115726,14.124791,13.45037,12.774135,12.099712,11.42529,10.750868,10.700105,10.649343,10.600392,10.549629,10.500679,10.1054535,9.710228,9.3150015,8.919776,8.52455,7.574558,6.624565,5.674573,4.7245803,3.774588,3.925064,4.07554,4.2242026,4.3746786,4.5251546,3.7546456,2.9841363,2.2154403,1.4449311,0.6744221,0.71430725,0.7541924,0.79589057,0.83577573,0.87566096,2.474694,4.07554,5.674573,7.2754188,8.874452,10.042,11.209548,12.377095,13.544643,14.712192,16.358362,18.002718,19.647076,21.293245,22.937603,18.992596,15.047589,11.102583,7.157576,3.2125697,3.5225863,3.832603,4.1426196,4.4526362,4.762653,4.5831695,4.401873,4.2223897,4.0429068,3.8616104,3.7927177,3.7220123,3.6531196,3.5824142,3.5117085,4.024777,3.6132345,3.199879,2.7883365,2.374981,1.9616255,1.7495089,1.5373923,1.3252757,1.1131591,0.89922947,0.8974165,0.89560354,0.8919776,0.8901646,0.8883517,1.6008459,2.3133402,3.0258346,3.738329,4.4508233,4.0882306,3.7256382,3.3630457,3.000453,2.6378605,4.25321,5.866747,7.4820967,9.097446,10.712796,10.081885,9.452786,8.821876,8.192778,7.5618668,7.7377243,7.911769,8.087626,8.26167,8.437528,7.837437,7.2373466,6.637256,6.037165,5.4370747,4.914942,4.3928084,3.870675,3.346729,2.8245957,3.7401419,4.655688,5.569421,6.484967,7.400513,6.7478466,6.09518,5.4425135,4.7898474,4.137181,4.004834,3.872488,3.7401419,3.6077955,3.4754493,4.4743915,5.475147,6.4759026,7.474845,8.4756,7.494787,6.5157876,5.5349746,4.554162,3.5751622,4.5849824,5.5948024,6.604623,7.614443,8.624263,8.002417,7.380571,6.7569118,6.1350656,5.5132194,4.5432844,3.5733492,2.6016014,1.6316663,0.66173136,1.0497054,1.4376793,1.8256533,2.2118144,2.5997884,2.665055,2.7303216,2.7955883,2.8608549,2.9243085,4.1299286,5.335549,6.539356,7.744976,8.950596,7.7703576,6.590119,5.40988,4.229642,3.049403,2.4801328,1.9108626,1.3397794,0.7705091,0.19942589,0.17767033,0.15410182,0.13234627,0.11059072,0.0870222,0.11784257,0.14684997,0.17767033,0.20667773,0.2374981,0.23568514,0.23205921,0.23024625,0.22662032,0.22480737,0.87022203,1.5156367,2.1592383,2.8046532,3.4500678,4.022964,4.59586,5.1669436,5.7398396,6.3127356,7.7903004,9.267865,10.745429,12.222994,13.700559,14.514579,15.330412,16.144432,16.960264,17.774284,20.270735,22.765371,25.260008,27.754644,30.24928,28.035654,25.820213,23.604773,21.389332,19.175705,20.894394,22.614895,24.335396,26.055899,27.774588,25.899984,24.025381,22.150776,20.27436,18.399757,18.318174,18.234777,18.153194,18.069798,17.988214,17.810545,17.632874,17.455204,17.277533,17.099863,16.864178,16.630306,16.39462,16.160748,15.925063,15.861609,15.799969,15.738328,15.674874,15.613234,15.072971,14.532708,13.992445,13.452183,12.91192,12.529385,12.14685,11.764315,11.381779,10.999244,10.852394,10.705544,10.556881,10.410031,10.263181,11.057259,11.853149,12.647227,13.443117,14.237195,14.55265,14.868106,15.181748,15.497204,15.812659,16.432693,17.052727,17.67276,18.292793,18.912827,17.903006,16.893185,15.883366,14.871732,13.861912,14.376793,14.891675,15.408369,15.92325,16.438131,15.966762,15.497204,15.027647,14.558089,14.0867195,14.4692545,14.851789,15.234324,15.616859,15.999394,16.702824,17.40444,18.10787,18.809486,19.512917,16.164375,12.817645,9.469104,6.1223745,2.7756457,2.2408218,1.7041848,1.1693609,0.6345369,0.099712946,1.6552348,3.2107568,4.764466,6.319988,7.8755093,8.105756,8.334189,8.564435,8.794682,9.024928,7.9607186,6.8946967,5.8304877,4.764466,3.7002566,3.9867048,4.274966,4.5632267,4.8496747,5.137936,6.0625467,6.987158,7.911769,8.838193,9.762803,9.030367,8.29793,7.5654926,6.833056,6.1006193,5.806919,5.5150323,5.223145,4.9294453,4.6375585,4.07554,3.5117085,2.94969,2.3876717,1.8256533,2.5327086,3.2397642,3.9468195,4.655688,5.3627434,4.604925,3.8471067,3.0892882,2.333283,1.5754645,2.4058013,3.2343252,4.064662,4.894999,5.7253356,5.9392653,6.155008,6.3707504,6.58468,6.8004227,6.6698895,6.539356,6.4106355,6.2801023,6.149569,8.350506,10.549629,12.750566,14.94969,17.150625,14.046834,10.944855,7.842876,4.7390842,1.6371052,4.117238,6.5973706,9.077503,11.557636,14.037769,13.470312,12.902855,12.335398,11.7679405,11.200482,12.130532,13.060582,13.990632,14.920682,15.850732,16.20426,16.5596,16.914942,17.27028,17.625622,16.467138,15.310469,14.151986,12.995316,11.836833,12.255627,12.672608,13.08959,13.508384,13.925365,14.34416,14.764768,15.185374,15.604169,16.024776,15.4827,14.940624,14.396736,13.85466,13.312584,13.125849,12.937301,12.750566,12.562017,12.375282,13.254569,14.13567,15.014956,15.894243,16.775343,16.815228,16.855114,16.894999,16.934883,16.97477,17.75253,18.53029,19.308052,20.085812,20.861761,21.655838,22.448103,23.240368,24.032633,24.824896,26.079466,27.33585,28.59042,29.84499,31.09956,32.178272,33.255173,34.332073,35.410786,36.487686,37.9308,39.37211,40.815228,42.258347,43.69965,45.454597,47.209545,48.964493,50.71944,52.47439,50.509136,48.5457,46.58045,44.615196,42.649944,38.744823,34.839703,30.93458,27.029459,23.124338,21.848013,20.569874,19.291735,18.01541,16.73727,14.447499,12.157727,9.867955,7.5781837,5.2865987,7.6343856,9.982172,12.329959,14.677745,17.025532,15.92325,14.819156,13.716875,12.6145935,11.512312,11.764315,12.018129,12.270131,12.522133,12.774135,12.166792,11.559449,10.952107,10.344765,9.737422,11.253058,12.766883,14.282519,15.798156,17.31198,16.89681,16.481644,16.068287,15.653119,15.23795,14.532708,13.827466,13.122223,12.416981,11.711739,9.8878975,8.062244,6.2365913,4.4127507,2.5870976,4.1498713,5.712645,7.2754188,8.838193,10.399154,10.20698,10.014805,9.822631,9.630457,9.438283,7.8247466,6.2130227,4.599486,2.9877625,1.3742256,1.1077201,0.83940166,0.5728962,0.3045777,0.038072214,0.047137026,0.058014803,0.06707962,0.07795739,0.0870222,0.07070554,0.052575916,0.034446288,0.018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.045324065,0.09064813,0.13415924,0.1794833,0.22480737,0.28463513,0.3444629,0.40429065,0.46411842,0.52575916,0.50037766,0.4749962,0.44961473,0.42423326,0.40066472,0.3208944,0.23931105,0.15954071,0.07977036,0.0,0.44780177,0.89560354,1.3434052,1.789394,2.2371957,2.3169663,2.3967366,2.47832,2.5580902,2.6378605,2.5744069,2.5127661,2.4493124,2.3876717,2.324218,2.126605,1.9308052,1.7331922,1.5355793,1.3379664,1.7404441,2.1429217,2.5453994,2.9478772,3.350355,3.1799364,3.009518,2.8390994,2.6704938,2.5000753,2.4130533,2.324218,2.2371957,2.1501737,2.0631514,2.0830941,2.1030366,2.1229792,2.1429217,2.1628644,2.0450218,1.9271792,1.8093367,1.693307,1.5754645,1.9308052,2.2843328,2.6396735,2.9950142,3.350355,4.024777,4.699199,5.375434,6.049856,6.7242785,6.776854,6.82943,6.882006,6.9345818,6.987158,7.0850577,7.1829576,7.2808576,7.3769445,7.474845,8.06587,8.655084,9.244296,9.835322,10.424535,11.292944,12.15954,13.027949,13.894546,14.762955,14.632421,14.501887,14.373167,14.242634,14.112101,12.839401,11.566701,10.2958145,9.023115,7.750415,7.6253204,7.500226,7.3751316,7.250037,7.124943,8.134763,9.144584,10.154404,11.164224,12.175857,12.19036,12.2048645,12.219368,12.235684,12.250188,11.537694,10.825199,10.112705,9.400211,8.6877165,8.488291,8.287052,8.087626,7.8882003,7.686961,7.507478,7.327995,7.1466985,6.967215,6.787732,5.9882154,5.186886,4.3873696,3.587853,2.7883365,2.8626678,2.9369993,3.0131438,3.0874753,3.1618068,2.6324217,2.1030366,1.5718386,1.0424535,0.51306844,0.53482395,0.55839247,0.58014804,0.60190356,0.62547207,1.6878681,2.7502642,3.8126602,4.8750563,5.9374523,7.019791,8.10213,9.184468,10.266808,11.349146,12.304577,13.260008,14.21544,15.169058,16.124489,13.43224,10.73999,8.047741,5.3554916,2.663242,3.101979,3.5425289,3.9830787,4.421816,4.8623657,4.691947,4.5233417,4.3529234,4.1825047,4.0120864,3.870675,3.727451,3.584227,3.442816,3.299592,3.386614,3.049403,2.712192,2.374981,2.03777,1.7005589,1.4757515,1.2491312,1.0243238,0.7995165,0.5747091,0.58014804,0.5855869,0.58921283,0.5946517,0.6000906,1.2872034,1.9743162,2.663242,3.350355,4.0374675,3.874301,3.7129474,3.5497808,3.386614,3.2252605,4.670192,6.115123,7.560054,9.004985,10.449916,9.873394,9.295059,8.716724,8.140202,7.5618668,7.8628187,8.161958,8.46291,8.762048,9.063,8.4756,7.8882003,7.3008003,6.7115874,6.1241875,5.4207582,4.7155156,4.0102735,3.3050308,2.5997884,3.7691493,4.940323,6.109684,7.2808576,8.450218,7.667019,6.885632,6.1024323,5.319232,4.537845,4.2767787,4.017525,3.7582715,3.4972048,3.2379513,4.12449,5.0128417,5.89938,6.787732,7.6742706,6.885632,6.09518,5.3047285,4.514277,3.7256382,4.6792564,5.634688,6.590119,7.5455503,8.499168,7.844689,7.1902094,6.53573,5.8794374,5.224958,4.25321,3.2796493,2.3079014,1.3343405,0.36259252,0.774135,1.1874905,1.6008459,2.0123885,2.4257438,2.570781,2.715818,2.8608549,3.005892,3.149116,4.8279195,6.5049095,8.1819,9.860703,11.537694,9.53437,7.5328593,5.529536,3.5280252,1.5247015,1.2400664,0.9554313,0.67079616,0.38434806,0.099712946,0.09427405,0.09064813,0.08520924,0.07977036,0.07433146,0.10333887,0.13053331,0.15772775,0.18492219,0.21211663,0.20486477,0.19761293,0.19036107,0.18310922,0.17585737,0.9481794,1.7205015,2.4928236,3.2651455,4.0374675,4.4798307,4.9221935,5.3645563,5.806919,6.249282,7.9081426,9.56519,11.222239,12.879286,14.538147,14.995013,15.45188,15.91056,16.367426,16.824293,18.998035,21.169964,23.341894,25.515635,27.687565,25.642542,23.59752,21.5525,19.507477,17.462456,19.19746,20.932467,22.66747,24.402477,26.137482,24.60009,23.062696,21.525305,19.987913,18.45052,18.590118,18.729717,18.869314,19.010725,19.150324,18.466837,17.785164,17.101677,16.420002,15.738328,15.769149,15.801782,15.834415,15.867048,15.899682,15.963136,16.024776,16.08823,16.14987,16.213324,15.468197,14.723069,13.9779415,13.232814,12.487686,12.302764,12.117842,11.9329195,11.747997,11.563075,11.619277,11.677292,11.735307,11.793322,11.849524,12.473183,13.095029,13.716875,14.340534,14.96238,15.2325115,15.502643,15.772775,16.042906,16.313038,16.797098,17.282972,17.767033,18.252907,18.736969,17.857681,16.978395,16.097294,15.218008,14.336908,15.094727,15.852545,16.610363,17.368181,18.124187,17.48965,16.855114,16.220575,15.584227,14.94969,15.06028,15.170871,15.279649,15.39024,15.50083,15.945006,16.389181,16.83517,17.279346,17.725336,14.458377,11.189605,7.9226465,4.655688,1.3869164,1.1204109,0.8520924,0.5855869,0.31726846,0.05076295,1.8655385,3.680314,5.4950895,7.309865,9.12464,9.414715,9.704789,9.994863,10.284937,10.57501,9.418341,8.259857,7.1031876,5.9447045,4.788034,4.762653,4.7372713,4.7118897,4.688321,4.6629395,5.8504305,7.037921,8.225411,9.412902,10.600392,9.739235,8.87989,8.020547,7.159389,6.300045,5.9356394,5.569421,5.2050157,4.84061,4.4743915,3.8869917,3.299592,2.712192,2.124792,1.5373923,2.084907,2.6324217,3.1799364,3.727451,4.274966,3.576975,2.8807976,2.182807,1.4848163,0.7868258,2.126605,3.4681973,4.8079767,6.147756,7.4875355,7.2572894,7.027043,6.796797,6.5683637,6.338117,6.4106355,6.4831543,6.5556726,6.628191,6.70071,9.800876,12.899229,15.999394,19.099562,22.199726,18.055294,13.910862,9.764616,5.620184,1.4757515,3.8398547,6.205771,8.569874,10.93579,13.299893,12.397038,11.494183,10.593141,9.690285,8.78743,10.226922,11.668227,13.107719,14.547212,15.986704,16.63937,17.292038,17.944704,10258.0,19.250036,18.327238,17.40444,16.481644,15.5606575,14.63786,15.214382,15.792717,16.36924,16.947575,17.524096,17.935638,18.345367,18.755098,19.164827,19.574556,18.33449,17.094423,15.854358,14.614291,13.374225,13.399607,13.424988,13.45037,13.475751,13.499319,14.639673,15.780026,16.92038,18.060734,19.199274,19.53286,19.864632,20.198215,20.529987,20.861761,21.29506,21.728357,22.159842,22.59314,23.024624,24.065266,25.104094,26.144733,27.185373,28.224201,29.714457,31.204712,32.694965,34.185223,35.675476,36.195797,36.714306,37.234627,37.754948,38.275265,40.465324,42.655384,44.845444,47.0355,49.22556,49.74044,50.25532,50.770203,51.285084,51.79997,48.830334,45.860703,42.889256,39.919624,36.94999,33.409275,29.87037,26.329655,22.790752,19.250036,18.50491,17.75978,17.014654,16.269526,15.524399,13.453996,11.385405,9.3150015,7.2445984,5.1741953,6.630004,8.0858135,9.539809,10.995618,12.449615,12.35534,12.259253,12.164979,12.070704,11.974618,12.3698435,12.76507,13.1602955,13.555521,13.9507475,13.05333,12.155914,11.256684,10.359268,9.461852,11.631968,13.802084,15.9722,18.142317,20.312433,19.192022,18.073423,16.953012,15.8326025,14.712192,14.059525,13.406858,12.754191,12.103338,11.450671,9.663091,7.8755093,6.0879283,4.3003473,2.5127661,4.537845,6.5629244,8.588004,10.613083,12.638163,12.197612,11.757062,11.318325,10.877775,10.437225,8.624263,6.813113,5.0001507,3.1871881,1.3742256,1.1095331,0.8448406,0.58014804,0.3154555,0.05076295,0.054388877,0.059827764,0.065266654,0.07070554,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.14322405,0.17223145,0.2030518,0.23205921,0.26287958,0.25018883,0.2374981,0.22480737,0.21211663,0.19942589,0.15954071,0.11965553,0.07977036,0.03988518,0.0,0.23024625,0.4604925,0.69073874,0.91917205,1.1494182,1.2781386,1.405046,1.5319533,1.6606737,1.7875811,1.7132497,1.6371052,1.5627737,1.4866294,1.4122978,1.2708868,1.1276628,0.98443866,0.8430276,0.69980353,0.89560354,1.0895905,1.2853905,1.4793775,1.6751775,1.7767034,1.8800422,1.983381,2.084907,2.1882458,1.9616255,1.7368182,1.5120108,1.2872034,1.062396,1.0732739,1.0823387,1.0932164,1.1022812,1.1131591,1.0478923,0.9826257,0.91735905,0.8520924,0.7868258,1.0895905,1.3923552,1.69512,1.9978848,2.3006494,2.962381,3.6241121,4.2876563,4.949388,5.612932,5.6074934,5.6020546,5.5966153,5.5929894,5.5875506,5.580299,5.573047,5.565795,5.5567303,5.5494785,6.09518,6.640882,7.1847706,7.7304726,8.274362,8.827314,9.380268,9.933222,10.484363,11.037316,11.135216,11.233116,11.329204,11.427103,11.525003,10.357455,9.189907,8.02236,6.8548117,5.6872635,5.6872635,5.6872635,5.6872635,5.6872635,5.6872635,6.604623,7.5219817,8.439341,9.3567,10.275872,10.2958145,10.315757,10.3357,10.355642,10.375585,9.625018,8.874452,8.125698,7.3751316,6.624565,6.2746634,5.924762,5.57486,5.224958,4.8750563,4.9095025,4.945762,4.9802084,5.0146546,5.049101,4.40006,3.7492065,3.100166,2.4493124,1.8002719,1.8002719,1.8002719,1.8002719,1.8002719,1.8002719,1.5101979,1.2201238,0.9300498,0.6399758,0.34990177,0.35534066,0.36077955,0.36440548,0.36984438,0.37528324,0.89922947,1.4249886,1.9507477,2.474694,3.000453,3.9975824,4.994712,5.9918413,6.9907837,7.987913,8.252605,8.517298,8.781991,9.046683,9.313189,7.8718834,6.432391,4.992899,3.5534067,2.1121013,2.6831846,3.2524548,3.8217251,4.3928084,4.9620786,4.802538,4.6429973,4.4816437,4.322103,4.162562,3.9468195,3.73289,3.5171473,3.303218,3.0874753,2.7502642,2.4873846,2.2245052,1.9616255,1.7005589,1.4376793,1.2001812,0.96268314,0.72518504,0.48768693,0.25018883,0.26287958,0.2755703,0.28826106,0.2991388,0.31182957,0.97537386,1.6371052,2.3006494,2.962381,3.6241121,3.6621845,3.7002566,3.738329,3.774588,3.8126602,5.087173,6.3616858,7.6380115,8.912524,10.1870365,9.663091,9.137331,8.613385,8.087626,7.5618668,7.987913,8.412147,8.838193,9.262425,9.686659,9.11195,8.537241,7.9625316,7.3878226,6.813113,5.924762,5.038223,4.1498713,3.2633326,2.374981,3.7999697,5.224958,6.6499467,8.074935,9.499924,8.588004,7.6742706,6.7623506,5.8504305,4.936697,4.550536,4.162562,3.774588,3.386614,3.000453,3.774588,4.550536,5.3246713,6.1006193,6.874754,6.2746634,5.674573,5.0744824,4.4743915,3.874301,4.7753434,5.674573,6.5756154,7.474845,8.375887,7.686961,6.9998484,6.3127356,5.6256227,4.936697,3.9631362,2.9877625,2.0123885,1.0370146,0.06164073,0.50037766,0.93730164,1.3742256,1.8129625,2.2498865,2.474694,2.6995013,2.9243085,3.149116,3.3757362,5.524097,7.6742706,9.824444,11.974618,14.124791,11.300196,8.4756,5.6491914,2.8245957,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.0870222,0.11240368,0.13778515,0.16316663,0.18673515,0.17585737,0.16316663,0.15047589,0.13778515,0.12509441,1.0243238,1.9253663,2.8245957,3.7256382,4.6248674,4.936697,5.2503395,5.562169,5.8758116,6.187641,8.024173,9.862516,11.700861,13.537392,15.375735,15.475449,15.575162,15.674874,15.774588,15.8743,17.725336,19.574556,21.425592,23.274813,25.125849,23.249432,21.374828,19.500225,17.625622,15.749206,17.500528,19.250036,20.999546,22.750868,24.500376,23.300196,22.100014,20.899832,19.699652,18.49947,18.862062,19.224655,19.587248,19.94984,20.312433,19.124943,17.937452,16.749962,15.56247,14.37498,14.674119,14.975071,15.27421,15.575162,15.8743,16.062849,16.249584,16.438131,16.624866,16.811602,15.861609,14.91343,13.961625,13.011633,12.06164,12.07433,12.087022,12.099712,12.112403,12.125093,12.387974,12.650853,12.91192,13.174799,13.437678,13.887294,14.336908,14.788336,15.23795,15.687565,15.912373,16.13718,16.361988,16.586794,16.811602,17.163317,17.513218,17.863121,18.213022,18.562923,17.812357,17.06179,16.313038,15.56247,14.811904,15.812659,16.811602,17.812357,18.813112,19.812056,19.012539,18.213022,17.411694,16.612177,15.812659,15.649493,15.488139,15.324973,15.161806,15.000452,15.187187,15.375735,15.56247,15.749206,15.937754,12.750566,9.563377,6.3743763,3.1871881,0.0,0.0,0.0,0.0,0.0,0.0,2.0758421,4.1498713,6.2257137,8.299743,10.375585,10.725487,11.075388,11.42529,11.775192,12.125093,10.874149,9.625018,8.374074,7.124943,5.8758116,5.5367875,5.199577,4.8623657,4.5251546,4.1879435,5.638314,7.0868707,8.537241,9.987611,11.437981,10.449916,9.461852,8.4756,7.4875355,6.4994707,6.0625467,5.6256227,5.186886,4.749962,4.313038,3.7002566,3.0874753,2.474694,1.8619126,1.2491312,1.6371052,2.0250793,2.4130533,2.7992141,3.1871881,2.5508385,1.9126755,1.2745126,0.63816285,0.0,1.8492218,3.7002566,5.5494785,7.400513,9.249735,8.575313,7.900891,7.224656,6.550234,5.8758116,6.149569,6.4251394,6.70071,6.9744673,7.250037,11.249433,15.250641,19.250036,23.249432,27.25064,22.061941,16.875055,11.6881695,6.4994707,1.3125849,3.5624714,5.812358,8.062244,10.312131,12.562017,11.325577,10.087324,8.849071,7.61263,6.3743763,8.325124,10.274059,12.224807,14.175554,16.124489,17.074482,18.024473,18.974466,19.92446,20.87445,20.187338,19.500225,18.813112,18.124187,17.437075,18.17495,18.912827,19.650702,20.386765,21.12464,21.525305,21.924156,22.324821,22.725487,23.124338,21.188093,19.250036,17.31198,15.375735,13.437678,13.675177,13.912675,14.150173,14.387671,14.625169,16.024776,17.424383,18.825804,20.22541,21.625017,22.25049,22.87415,23.49962,24.125093,24.750565,24.837587,24.92461,25.011631,25.100468,25.187489,26.474693,27.761896,29.050913,30.338116,31.625319,33.349445,35.075386,36.799515,38.525455,40.24958,40.21332,40.17525,40.13718,40.099106,40.062847,42.999847,45.936848,48.87566,51.812656,54.749657,54.02447,53.299286,52.5741,51.85073,51.125546,47.14972,43.175705,39.19988,35.22405,31.250036,28.075539,24.89923,21.724731,18.550234,15.375735,15.161806,14.94969,14.737573,14.525456,14.313339,12.462305,10.613083,8.762048,6.9128265,5.0617914,5.6256227,6.187641,6.7496595,7.311678,7.8755093,8.78743,9.699349,10.613083,11.525003,12.436923,12.975373,13.512011,14.05046,14.587097,15.125546,13.938056,12.750566,11.563075,10.375585,9.188094,12.012691,14.837286,17.661882,20.48829,23.312885,21.487232,19.663393,17.837738,16.012085,14.188245,13.588155,12.988064,12.387974,11.787883,11.187792,9.438283,7.686961,5.9374523,4.1879435,2.4366217,4.9258194,7.413204,9.900589,12.387974,14.875358,14.188245,13.499319,12.812206,12.125093,11.437981,9.425592,7.413204,5.4008155,3.386614,1.3742256,1.1131591,0.85027945,0.5873999,0.3245203,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.2374981,0.41335547,0.5873999,0.76325727,0.93730164,0.85027945,0.76325727,0.6744221,0.5873999,0.50037766,0.41335547,0.3245203,0.2374981,0.15047589,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.37528324,0.7505665,1.1258497,1.49932,1.8746033,1.5120108,1.1494182,0.7868258,0.42423326,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.25018883,0.50037766,0.7505665,1.0007553,1.2491312,1.8999848,2.5508385,3.199879,3.8507326,4.499773,4.4381323,4.3746786,4.313038,4.249584,4.1879435,4.07554,3.9631362,3.8507326,3.738329,3.6241121,4.12449,4.6248674,5.125245,5.6256227,6.1241875,6.3616858,6.599184,6.836682,7.07418,7.311678,7.6380115,7.9625316,8.287052,8.613385,8.937905,7.8755093,6.813113,5.750717,4.688321,3.6241121,3.7492065,3.874301,3.9993954,4.12449,4.249584,5.0744824,5.89938,6.7242785,7.549176,8.375887,8.399456,8.424837,8.450218,8.4756,8.499168,7.7123427,6.925517,6.1368785,5.3500524,4.5632267,4.062849,3.5624714,3.0620937,2.561716,2.0631514,2.3133402,2.561716,2.811905,3.0620937,3.3122826,2.811905,2.3133402,1.8129625,1.3125849,0.8122072,0.73787576,0.66173136,0.5873999,0.51306844,0.43692398,0.387974,0.33721104,0.28826106,0.2374981,0.18673515,0.17585737,0.16316663,0.15047589,0.13778515,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.97537386,1.887294,2.7992141,3.7129474,4.6248674,4.2006345,3.774588,3.350355,2.9243085,2.5000753,2.3133402,2.124792,1.938057,1.7495089,1.5627737,2.2625773,2.962381,3.6621845,4.361988,5.0617914,4.9131284,4.762653,4.612177,4.461701,4.313038,4.024777,3.738329,3.4500678,3.1618068,2.8753586,3.1255474,2.8826106,2.6396735,2.3967366,2.1556125,1.9126755,1.69512,1.4775645,1.260009,1.0424535,0.824898,0.8122072,0.7995165,0.7868258,0.774135,0.76325727,1.4249886,2.08672,2.7502642,3.4119956,4.07554,4.0120864,3.9504454,3.8869917,3.825351,3.7618973,4.9167547,6.071612,7.228282,8.383139,9.537996,9.03218,8.528176,8.02236,7.518356,7.0125394,7.4694057,7.9280853,8.384952,8.841819,9.300498,8.705847,8.109382,7.51473,6.9200783,6.3254266,5.638314,4.949388,4.262275,3.5751622,2.8880494,4.1444325,5.4026284,6.6608243,7.9172077,9.175404,8.357758,7.5401115,6.722465,5.904819,5.087173,4.74271,4.3982472,4.0519714,3.7075086,3.3630457,4.115425,4.8678045,5.620184,6.3725634,7.124943,6.6481338,6.169512,5.6927023,5.2158933,4.7372713,5.4932766,6.247469,7.0016613,7.757667,8.511859,7.7322855,6.9527116,6.1731377,5.391751,4.612177,3.7129474,2.811905,1.9126755,1.0116332,0.11240368,0.50037766,0.8883517,1.2745126,1.6624867,2.0504606,2.6451125,3.2397642,3.834416,4.4308805,5.0255322,6.5774283,8.129324,9.683033,11.234929,12.786825,10.232361,7.6778965,5.121619,2.5671551,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.07070554,0.09064813,0.11059072,0.13053331,0.15047589,0.24293698,0.33539808,0.42785916,0.52032024,0.61278135,1.2527572,1.892733,2.5327086,3.1726844,3.8126602,4.1444325,4.478018,4.8097897,5.143375,5.475147,6.9527116,8.430276,9.907841,11.385405,12.862969,13.182051,13.502945,13.822026,14.142921,14.462003,15.977639,17.493277,19.0071,20.522736,22.038374,20.736666,19.436771,18.136877,16.836983,15.537089,16.90225,18.26741,19.632572,20.997732,22.362894,21.327692,20.29249,19.257288,18.222088,17.186886,17.420757,17.652817,17.884876,18.116936,18.350807,17.3428,16.334793,15.326786,14.320591,13.312584,13.684241,14.057712,14.429369,14.802839,15.174497,15.437376,15.700256,15.963136,16.224201,16.487082,15.89243,15.297778,14.703127,14.106662,13.512011,13.452183,13.392355,13.332527,13.272699,13.212872,13.299893,13.386916,13.475751,13.562773,13.649796,14.13023,14.610665,15.089288,15.569723,16.050158,16.21695,16.385555,16.55235,16.719141,16.887747,17.50778,18.127813,18.747847,19.36788,19.987913,19.137632,18.287354,17.437075,16.586794,15.738328,16.478018,17.217705,17.957394,18.697083,19.436771,18.568363,17.698141,16.827919,15.957697,15.087475,15.408369,15.72745,16.048346,16.367426,16.68832,16.48527,16.282217,16.079165,15.877926,15.674874,12.627284,9.579695,6.532104,3.484514,0.43692398,0.44961473,0.46230546,0.4749962,0.48768693,0.50037766,2.324218,4.1498713,5.975525,7.799365,9.625018,9.869768,10.114518,10.359268,10.605831,10.850581,9.960417,9.070251,8.180087,7.2899227,6.399758,6.004532,5.6093063,5.2158933,4.8206677,4.4254417,5.542227,6.6608243,7.7776093,8.894395,10.012992,9.460039,8.907085,8.354132,7.802991,7.250037,6.775041,6.300045,5.825049,5.3500524,4.8750563,4.168001,3.4591327,2.752077,2.0450218,1.3379664,1.7368182,2.137483,2.5381477,2.9369993,3.3376641,2.6723068,2.0069497,1.3415923,0.678048,0.012690738,2.1991236,4.3873696,6.5756154,8.762048,10.950294,10.37921,9.80994,9.24067,8.669587,8.100317,7.8791356,7.6597667,7.440398,7.219217,6.9998484,10.0510645,13.100468,16.14987,19.199274,22.25049,18.25472,14.260764,10.264994,6.2692246,2.275268,4.0392804,5.805106,7.570932,9.334945,11.10077,10.172533,9.244296,8.317872,7.3896356,6.4632115,8.118446,9.771869,11.427103,13.082338,14.737573,15.622298,16.507025,17.39175,18.278288,19.163015,19.083244,19.001661,18.92189,18.84212,18.76235,19.222843,19.683334,20.142014,20.602507,21.063,21.070251,21.077503,21.084755,21.092007,21.099258,19.259102,17.420757,15.580601,13.740443,11.900287,12.766883,13.635292,14.501887,15.3702965,16.236893,17.125244,18.011784,18.900135,19.786674,20.675026,21.652212,22.629398,23.608398,24.585585,25.562773,25.577276,25.59178,25.608097,25.6226,25.637104,27.009516,28.38193,29.754341,31.126755,32.49917,33.98217,35.465176,36.948177,38.429367,39.912373,40.285843,40.657497,41.029156,41.402626,41.774284,43.81568,45.855263,47.894844,49.93443,51.975822,50.784706,49.595406,48.40429,47.214985,46.02568,42.361683,38.6995,35.037315,31.37513,27.712946,25.069647,22.42816,19.78486,17.141562,14.500074,14.297023,14.095784,13.892733,13.68968,13.486629,11.894848,10.303066,8.709473,7.117691,5.524097,6.09518,6.6644506,7.2355337,7.804804,8.375887,8.917963,9.460039,10.002114,10.54419,11.088079,11.539507,11.992747,12.444175,12.897416,13.3506565,12.572895,11.795135,11.017374,10.239613,9.461852,11.399909,13.337966,15.27421,17.212267,19.150324,18.20577,17.259403,16.31485,15.3702965,14.425743,13.36516,12.304577,11.245807,10.185224,9.12464,7.7340984,6.345369,4.954827,3.5642843,2.175555,4.555975,6.9345818,9.3150015,11.695421,14.075842,13.397794,12.719746,12.0416975,11.365462,10.687414,8.901647,7.117691,5.331923,3.5479677,1.7621996,1.4195497,1.0768998,0.73424983,0.39159992,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.34264994,0.6726091,1.0025684,1.3325275,1.6624867,1.9181144,2.1719291,2.427557,2.6831846,2.9369993,2.4402475,1.9416829,1.4449311,0.9481794,0.44961473,0.47318324,0.4949388,0.5166943,0.5402629,0.5620184,1.0225109,1.4830034,1.9416829,2.4021754,2.8626678,2.5907235,2.3169663,2.0450218,1.7730774,1.49932,1.214685,0.9300498,0.64541465,0.36077955,0.07433146,0.072518505,0.07070554,0.06707962,0.065266654,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.2030518,0.40429065,0.6073425,0.8103943,1.0116332,1.5355793,2.0577126,2.5798457,3.101979,3.6241121,3.5733492,3.5207734,3.4681973,3.4156215,3.3630457,3.2705846,3.1781235,3.0856624,2.9932013,2.9007401,3.299592,3.7002566,4.099108,4.499773,4.900438,5.090799,5.279347,5.469708,5.660069,5.8504305,6.109684,6.3707504,6.630004,6.889258,7.1503243,6.3072968,5.464269,4.6230545,3.780027,2.9369993,3.0294604,3.1219215,3.2143826,3.3068438,3.3993049,4.059223,4.7191415,5.3808727,6.0407915,6.70071,6.720652,6.740595,6.7605376,6.78048,6.8004227,6.1749506,5.5494785,4.9258194,4.3003473,3.6748753,3.2832751,2.8898623,2.4982624,2.1048496,1.7132497,1.9126755,2.1121013,2.3133402,2.5127661,2.712192,2.3097143,1.9072367,1.504759,1.1022812,0.69980353,0.6399758,0.58014804,0.52032024,0.4604925,0.40066472,0.36077955,0.3208944,0.27919623,0.23931105,0.19942589,0.19036107,0.1794833,0.17041849,0.15954071,0.15047589,0.13415924,0.11965553,0.10515183,0.09064813,0.07433146,0.8031424,1.5301404,2.2571385,2.9841363,3.7129474,3.3757362,3.0367124,2.6995013,2.3622901,2.0250793,1.8746033,1.7241274,1.5754645,1.4249886,1.2745126,1.8347181,2.3949237,2.955129,3.5153344,4.07554,3.972201,3.870675,3.7673361,3.6658103,3.5624714,3.3848011,3.207131,3.0294604,2.8517902,2.6741197,3.5008307,3.2778363,3.054842,2.8318477,2.610666,2.3876717,2.1900587,1.9924458,1.794833,1.5972201,1.3996071,1.3633479,1.3252757,1.2872034,1.2491312,1.2128719,1.8746033,2.5381477,3.199879,3.8616104,4.5251546,4.361988,4.2006345,4.0374675,3.874301,3.7129474,4.748149,5.7833505,6.816739,7.851941,8.887142,8.403082,7.9172077,7.4331465,6.947273,6.4632115,6.9527116,7.4422116,7.931711,8.423024,8.912524,8.29793,7.6833353,7.066928,6.452334,5.8377395,5.3500524,4.8623657,4.3746786,3.8869917,3.3993049,4.4907084,5.580299,6.6698895,7.75948,8.8508835,8.127511,7.404139,6.68258,5.959208,5.237649,4.934884,4.632119,4.329355,4.028403,3.7256382,4.454449,5.185073,5.915697,6.644508,7.3751316,7.019791,6.6644506,6.3091097,5.955582,5.600241,6.209397,6.8203654,7.4295206,8.040489,8.649645,7.7776093,6.9055743,6.0317264,5.1596913,4.2876563,3.4627585,2.6378605,1.8129625,0.9880646,0.16316663,0.50037766,0.8375887,1.1747998,1.5120108,1.8492218,2.8155308,3.780027,4.744523,5.710832,6.6753283,7.6307597,8.584378,9.539809,10.49524,11.450671,9.164526,6.880193,4.594047,2.3097143,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.052575916,0.06707962,0.08339628,0.09789998,0.11240368,0.3100166,0.5076295,0.70524246,0.90285534,1.1004683,1.4793775,1.8600996,2.2408218,2.619731,3.000453,3.3521678,3.7056956,4.0574102,4.409125,4.762653,5.8794374,6.9980354,8.1148205,9.231606,10.3502035,10.890467,11.430729,11.969179,12.509441,13.049705,14.229943,15.410182,16.59042,17.770658,18.949085,18.225714,17.500528,16.775343,16.050158,15.324973,16.305786,17.284784,18.265598,19.244598,20.22541,19.355188,18.484966,17.614744,16.744522,15.8743,15.977639,16.079165,16.182505,16.285843,16.38737,15.5606575,14.732134,13.905423,13.0769,12.250188,12.694364,13.140353,13.584529,14.030518,14.474693,14.811904,15.149116,15.488139,15.825351,16.162561,15.92325,15.682126,15.442815,15.201692,14.96238,14.830034,14.697688,14.565341,14.432995,14.300649,14.211814,14.124791,14.037769,13.9507475,13.861912,14.373167,14.882609,15.392053,15.903308,16.41275,16.52334,16.632118,16.74271,16.8533,16.962078,17.852243,18.742407,19.632572,20.522736,21.4129,20.462908,19.512917,18.562923,17.612932,16.66294,17.143373,17.621996,18.102432,18.582867,19.063301,18.122374,17.18326,16.242332,15.303217,14.362289,15.165432,15.966762,16.769903,17.573046,18.374376,17.78335,17.190512,16.597672,16.004833,15.411995,12.5058155,9.597824,6.6898317,3.7818398,0.87566096,0.89922947,0.9246109,0.9499924,0.97537386,1.0007553,2.5744069,4.1498713,5.7253356,7.3008003,8.874452,9.015862,9.155461,9.295059,9.434657,9.574255,9.04487,8.515485,7.9842873,7.454902,6.925517,6.472276,6.0208488,5.567608,5.1143675,4.6629395,5.4479527,6.2329655,7.017978,7.802991,8.588004,8.470161,8.352319,8.234476,8.116633,8.000604,7.4875355,6.9744673,6.4632115,5.9501433,5.4370747,4.6357455,3.832603,3.0294604,2.228131,1.4249886,1.8383441,2.2498865,2.663242,3.0747845,3.48814,2.7955883,2.1030366,1.4104849,0.7179332,0.025381476,2.5508385,5.0744824,7.5999393,10.125396,12.650853,12.184921,11.720803,11.254871,10.790753,10.324821,9.610515,8.894395,8.180087,7.46578,6.7496595,8.8508835,10.950294,13.049705,15.149116,17.25034,14.447499,11.644659,8.841819,6.0407915,3.2379513,4.517903,5.7978544,7.077806,8.357758,9.637709,9.019489,8.403082,7.7848616,7.166641,6.550234,7.909956,9.269678,10.629399,11.989121,13.3506565,14.170115,14.989574,15.810846,16.630306,17.449764,17.977337,18.50491,19.03248,19.560053,20.087626,20.270735,20.45203,20.63514,20.818249,20.999546,20.615198,20.23085,19.844688,19.46034,19.074179,17.331923,15.589665,13.847408,12.105151,10.362894,11.860401,13.357908,14.855415,16.352922,17.85043,18.225714,18.599184,18.974466,19.34975,19.725033,21.055748,22.38465,23.715364,25.044266,26.374979,26.316965,26.260763,26.202747,26.144733,26.08672,27.54434,29.001963,30.459585,31.917206,33.37483,34.614895,35.85496,37.095028,38.335094,39.57516,40.35836,41.139748,41.922947,42.704334,43.487534,44.6297,45.771866,46.915844,48.058014,49.20018,47.544945,45.88971,44.234474,42.57924,40.925816,37.575462,34.22511,30.874752,27.524399,24.175856,22.065567,19.955278,17.84499,15.734702,13.6244135,13.43224,13.240066,13.047892,12.855718,12.661731,11.327391,9.99305,8.656897,7.322556,5.9882154,6.5647373,7.1430726,7.7195945,8.29793,8.874452,9.046683,9.220728,9.39296,9.56519,9.737422,10.1054535,10.471672,10.839704,11.207735,11.575767,11.207735,10.839704,10.471672,10.1054535,9.737422,10.7871275,11.836833,12.888351,13.938056,14.9877615,14.922495,14.857228,14.791962,14.726695,14.663241,13.142166,11.622903,10.101828,8.582565,7.063302,6.0317264,5.0019636,3.972201,2.9424384,1.9126755,4.1843176,6.4577727,8.729415,11.00287,13.274512,12.607342,11.940171,11.273002,10.605831,9.936848,8.379513,6.8221784,5.2648435,3.7075086,2.1501737,1.7277533,1.305333,0.88291276,0.4604925,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.099712946,0.19942589,0.2991388,0.40066472,0.50037766,0.40066472,0.2991388,0.19942589,0.099712946,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.6726091,1.3198367,1.9670644,2.6142921,3.2633326,3.5969179,3.9323158,4.267714,4.603112,4.936697,4.0302157,3.1219215,2.2154403,1.3071461,0.40066472,0.533011,0.6653573,0.79770356,0.9300498,1.062396,1.9942589,2.9279346,3.8597972,4.7916603,5.7253356,4.804351,3.8851788,2.9641938,2.0450218,1.1258497,0.91735905,0.7106813,0.50219065,0.2955129,0.0870222,0.08339628,0.07795739,0.072518505,0.06707962,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.15591478,0.3100166,0.46411842,0.6200332,0.774135,1.1693609,1.5645868,1.9598125,2.3550384,2.7502642,2.7067533,2.665055,2.6233568,2.5798457,2.5381477,2.465629,2.3931105,2.3205922,2.2480736,2.175555,2.474694,2.7756457,3.0747845,3.3757362,3.6748753,3.8180993,3.9595103,4.102734,4.2441454,4.3873696,4.5831695,4.7771564,4.972956,5.1669436,5.3627434,4.7390842,4.117238,3.4953918,2.8717327,2.2498865,2.3097143,2.3695421,2.42937,2.4891977,2.5508385,3.045777,3.540716,4.0356545,4.5305934,5.0255322,5.040036,5.0545397,5.0708566,5.08536,5.0998635,4.6375585,4.175253,3.7129474,3.2506418,2.7883365,2.5018883,2.2172532,1.9326181,1.647983,1.3633479,1.5120108,1.6624867,1.8129625,1.9616255,2.1121013,1.8075237,1.502946,1.1983683,0.8919776,0.5873999,0.5420758,0.49675176,0.45324063,0.40791658,0.36259252,0.33177215,0.30276474,0.27194437,0.24293698,0.21211663,0.20486477,0.19761293,0.19036107,0.18310922,0.17585737,0.15772775,0.13959812,0.12328146,0.10515183,0.0870222,0.630911,1.1729867,1.7150626,2.2571385,2.7992141,2.5508385,2.3006494,2.0504606,1.8002719,1.550083,1.4376793,1.3252757,1.2128719,1.1004683,0.9880646,1.4068589,1.8274662,2.2480736,2.666868,3.0874753,3.0330863,2.9768846,2.9224956,2.8681068,2.811905,2.7448254,2.6777458,2.610666,2.5417736,2.474694,3.874301,3.673062,3.4700103,3.2669585,3.0657198,2.8626678,2.6849976,2.5073273,2.3296568,2.1519866,1.9743162,1.9126755,1.8492218,1.7875811,1.7241274,1.6624867,2.324218,2.9877625,3.6494937,4.313038,4.974769,4.7118897,4.4508233,4.1879435,3.925064,3.6621845,4.5777307,5.4932766,6.4070096,7.322556,8.238102,7.7721705,7.308052,6.8421206,6.378002,5.9120708,6.434204,6.9581504,7.4802837,8.002417,8.52455,7.890013,7.2554765,6.6191263,5.9845896,5.3500524,5.0617914,4.7753434,4.4870825,4.2006345,3.9123733,4.835171,5.7579694,6.680767,7.6017523,8.52455,7.897265,7.26998,6.642695,6.01541,5.388125,5.127058,4.8678045,4.606738,4.347484,4.0882306,4.795286,5.5023413,6.209397,6.9182653,7.6253204,7.3932614,7.159389,6.92733,6.695271,6.4632115,6.92733,7.3932614,7.85738,8.323311,8.78743,7.8229337,6.8566246,5.8921285,4.9276323,3.9631362,3.2125697,2.4620032,1.7132497,0.96268314,0.21211663,0.50037766,0.7868258,1.0750868,1.3633479,1.649796,2.9841363,4.3202896,5.65463,6.9907837,8.325124,8.682278,9.039432,9.398398,9.755551,10.112705,8.096691,6.0824895,4.068288,2.0522738,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.034446288,0.045324065,0.054388877,0.065266654,0.07433146,0.3770962,0.67986095,0.9826257,1.2853905,1.5881553,1.7078108,1.8274662,1.9471219,2.0667772,2.1882458,2.5599031,2.9333735,3.3050308,3.6766882,4.0501585,4.8079767,5.565795,6.3218007,7.079619,7.837437,8.597069,9.3567,10.118144,10.877775,11.637406,12.482247,13.327088,14.171928,15.016769,15.861609,15.712947,15.56247,15.411995,15.263332,15.112856,15.707508,16.30216,16.89681,17.493277,18.087927,17.382685,16.677443,15.9722,15.266958,14.561715,14.534521,14.507326,14.480132,14.452938,14.425743,13.776703,13.129475,12.482247,11.83502,11.187792,11.704487,12.222994,12.739688,13.258195,13.77489,14.188245,14.599788,15.013144,15.4246855,15.838041,15.952258,16.068287,16.182505,16.29672,16.41275,16.207886,16.003021,15.798156,15.593291,15.386614,15.125546,14.862667,14.599788,14.336908,14.075842,14.614291,15.154554,15.694818,16.23508,16.775343,16.827919,16.880495,16.933071,16.985647,17.038223,18.196705,19.357002,20.517298,21.677593,22.837889,21.788185,20.736666,19.68696,18.637255,17.58755,17.80692,18.0281,18.247469,18.466837,18.688019,17.678198,16.668379,15.656745,14.646925,13.637105,14.922495,16.207886,17.493277,18.776854,20.062244,19.079618,18.096992,17.114367,16.13174,15.149116,12.382534,9.615953,6.8475595,4.079166,1.3125849,1.3506571,1.3869164,1.4249886,1.4630609,1.49932,2.8245957,4.1498713,5.475147,6.8004227,8.125698,8.160145,8.194591,8.23085,8.265296,8.299743,8.129324,7.9607186,7.7903004,7.6198816,7.4494634,6.9400206,6.430578,5.919323,5.40988,4.900438,5.351866,5.805106,6.258347,6.7097745,7.1630154,7.4802837,7.797552,8.1148205,8.432089,8.749357,8.200029,7.650702,7.0995617,6.550234,6.000906,5.101677,4.2042603,3.3068438,2.4094272,1.5120108,1.938057,2.3622901,2.7883365,3.2125697,3.636803,2.9170568,2.1973107,1.4775645,0.75781834,0.038072214,2.9007401,5.7615952,8.624263,11.486931,14.349599,13.990632,13.629852,13.270886,12.910107,12.549327,11.340081,10.130835,8.919776,7.71053,6.4994707,7.650702,8.80012,9.949538,11.10077,12.250188,10.640278,9.030367,7.420456,5.810545,4.2006345,4.994712,5.7906027,6.58468,7.380571,8.174648,7.8682575,7.560054,7.25185,6.94546,6.637256,7.703278,8.767487,9.8316965,10.897718,11.961927,12.717933,13.472125,14.22813,14.982323,15.738328,16.873243,18.008158,19.143072,20.277987,21.4129,21.316814,21.22254,21.128265,21.032179,20.937904,20.160145,19.382383,18.604622,17.82686,17.0491,15.404743,13.760386,12.114216,10.469859,8.825501,10.952107,13.080525,15.20713,17.335548,19.462152,19.324368,19.188396,19.050611,18.912827,18.77504,20.45747,22.139898,23.822329,25.504757,27.187187,27.056654,26.927933,26.7974,26.666866,26.538147,28.080976,29.621996,31.164827,32.707657,34.25049,35.24762,36.244747,37.24188,38.240818,39.23795,40.430878,41.621994,42.814926,44.007854,45.200783,45.445534,45.690285,45.93503,46.179783,46.424534,44.30518,42.185825,40.06466,37.94531,35.824142,32.78743,29.750715,26.71219,23.675478,20.636953,19.059675,17.482399,15.905121,14.327844,12.750566,12.567456,12.384347,12.203052,12.019942,11.836833,10.7599325,9.683033,8.604321,7.5274205,6.450521,7.0342946,7.6198816,8.205468,8.789243,9.374829,9.177217,8.979604,8.781991,8.584378,8.386765,8.669587,8.952409,9.235231,9.518054,9.800876,9.842574,9.884272,9.927783,9.969481,10.012992,10.174346,10.337513,10.500679,10.662033,10.825199,11.63922,12.455053,13.270886,14.084907,14.90074,12.919171,10.939416,8.9596615,6.979906,5.0001507,4.329355,3.6603715,2.9895754,2.3205922,1.649796,3.8144734,5.979151,8.145641,10.310318,12.474996,11.81689,11.160598,10.502492,9.844387,9.188094,7.85738,6.526665,5.197764,3.8670492,2.5381477,2.034144,1.5319533,1.0297627,0.5275721,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.15047589,0.2991388,0.44961473,0.6000906,0.7505665,0.6000906,0.44961473,0.2991388,0.15047589,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,1.0025684,1.9670644,2.9333735,3.8978696,4.8623657,5.277534,5.6927023,6.107871,6.5230393,6.9382076,5.620184,4.3021603,2.9841363,1.6679256,0.34990177,0.59283876,0.83577573,1.0768998,1.3198367,1.5627737,2.9678197,4.3728657,5.7779117,7.1829576,8.588004,7.019791,5.4533916,3.8851788,2.3169663,0.7505665,0.6200332,0.4894999,0.36077955,0.23024625,0.099712946,0.092461094,0.08520924,0.07795739,0.07070554,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.10696479,0.21574254,0.32270733,0.42967212,0.53663695,0.80495536,1.0732739,1.3397794,1.6080978,1.8746033,1.84197,1.8093367,1.7767034,1.745883,1.7132497,1.6606737,1.6080978,1.5555218,1.502946,1.4503701,1.649796,1.8492218,2.0504606,2.2498865,2.4493124,2.5453994,2.6396735,2.7357605,2.8300345,2.9243085,3.054842,3.1853752,3.3140955,3.444629,3.5751622,3.1726844,2.770207,2.3677292,1.9652514,1.5627737,1.5899682,1.6171626,1.6443571,1.6733645,1.7005589,2.030518,2.3604772,2.6904364,3.0203958,3.350355,3.3594196,3.3702974,3.3793623,3.39024,3.3993049,3.100166,2.7992141,2.5000753,2.1991236,1.8999848,1.7223145,1.5446441,1.3669738,1.1893034,1.0116332,1.1131591,1.2128719,1.3125849,1.4122978,1.5120108,1.305333,1.0968424,0.8901646,0.68167394,0.4749962,0.44417584,0.41516843,0.38434806,0.35534066,0.3245203,0.3045777,0.28463513,0.26469254,0.24474995,0.22480737,0.21936847,0.21574254,0.21030366,0.20486477,0.19942589,0.1794833,0.15954071,0.13959812,0.11965553,0.099712946,0.45686656,0.81583315,1.1729867,1.5301404,1.887294,1.7241274,1.5627737,1.3996071,1.2382535,1.0750868,1.0007553,0.9246109,0.85027945,0.774135,0.69980353,0.9808127,1.260009,1.5392052,1.8202144,2.0994108,2.0921588,2.084907,2.077655,2.0704033,2.0631514,2.1048496,2.1483607,2.1900587,2.231757,2.275268,4.249584,4.068288,3.8851788,3.7020695,3.5207734,3.3376641,3.1799364,3.0222087,2.864481,2.7067533,2.5508385,2.4620032,2.374981,2.2879589,2.1991236,2.1121013,2.7756457,3.437377,4.100921,4.762653,5.424384,5.0617914,4.699199,4.3366065,3.975827,3.6132345,4.407312,5.2032027,5.99728,6.793171,7.5872483,7.1430726,6.697084,6.2529078,5.806919,5.3627434,5.91751,6.472276,7.027043,7.5818095,8.138389,7.4820967,6.827617,6.1731377,5.516845,4.8623657,4.7753434,4.688321,4.599486,4.512464,4.4254417,5.179634,5.9356394,6.6898317,7.4458375,8.200029,7.667019,7.135821,6.60281,6.069799,5.5367875,5.319232,5.101677,4.8841214,4.668379,4.4508233,5.1343102,5.81961,6.5049095,7.1902094,7.8755093,7.764919,7.654328,7.5455503,7.4349594,7.324369,7.645263,7.9643445,8.285239,8.604321,8.925215,7.8682575,6.8094873,5.75253,4.695573,3.636803,2.962381,2.2879589,1.6117238,0.93730164,0.26287958,0.50037766,0.73787576,0.97537386,1.2128719,1.4503701,3.1545548,4.860553,6.5647373,8.270736,9.97492,9.735609,9.494485,9.255174,9.015862,8.774739,7.0306687,5.2847857,3.540716,1.794833,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.018129626,0.02175555,0.027194439,0.032633327,0.038072214,0.44417584,0.8520924,1.260009,1.6679256,2.0758421,1.9344311,1.794833,1.6552348,1.5156367,1.3742256,1.7676386,2.1592383,2.5526514,2.9442513,3.3376641,3.7347028,4.1317415,4.5305934,4.9276323,5.3246713,6.305484,7.2844834,8.265296,9.244296,10.225109,10.734551,11.245807,11.755249,12.264692,12.774135,13.200181,13.6244135,14.05046,14.474693,14.90074,15.10923,15.319533,15.529838,15.740141,15.950445,15.410182,14.869919,14.329657,13.789393,13.24913,13.093216,12.935488,12.7777605,12.620032,12.462305,11.99456,11.526816,11.060884,10.593141,10.125396,10.714609,11.3056345,11.894848,12.485873,13.075087,13.562773,14.05046,14.538147,15.025834,15.511708,15.983078,16.452635,16.922194,17.39175,17.863121,17.585737,17.308353,17.029158,16.751774,16.474392,16.037468,15.600543,15.161806,14.724882,14.287958,14.857228,15.428311,15.9975815,16.566853,17.137936,17.132496,17.127058,17.121618,17.117992,17.112555,18.542982,19.971596,21.402023,22.83245,24.262878,23.111647,21.962229,20.81281,19.66158,18.512161,18.472277,18.43239,18.392506,18.352621,18.312735,17.23221,16.151684,15.072971,13.992445,12.91192,14.679558,16.447197,18.214834,19.982473,21.750113,20.377699,19.005287,17.632874,16.260462,14.888049,12.259253,9.63227,7.0052876,4.3783045,1.7495089,1.8002719,1.8492218,1.8999848,1.9507477,1.9996977,3.0747845,4.1498713,5.224958,6.300045,7.3751316,7.304426,7.2355337,7.1648283,7.0941224,7.02523,7.215591,7.404139,7.5945,7.7848616,7.9752226,7.407765,6.8403077,6.2728505,5.7053933,5.137936,5.2575917,5.377247,5.4969025,5.618371,5.7380266,6.490406,7.2427855,7.995165,8.747544,9.499924,8.912524,8.325124,7.7377243,7.1503243,6.5629244,5.569421,4.5777307,3.584227,2.5925364,1.6008459,2.03777,2.474694,2.911618,3.350355,3.787279,3.0403383,2.2933977,1.5446441,0.79770356,0.05076295,3.2506418,6.450521,9.6504,12.850279,16.050158,15.79453,15.540715,15.285088,15.02946,14.775645,13.069647,11.365462,9.659465,7.95528,6.249282,6.450521,6.6499467,6.849373,7.0506115,7.250037,6.833056,6.414262,5.99728,5.580299,5.163317,5.473334,5.7833505,6.093367,6.4033837,6.7134004,6.7152133,6.717026,6.720652,6.722465,6.7242785,7.494787,8.265296,9.035806,9.804502,10.57501,11.26575,11.954676,12.645414,13.33434,14.025079,15.767336,17.509592,19.25185,20.99592,22.738176,22.364706,21.99305,21.61958,21.247921,20.87445,19.70509,18.53573,17.364555,16.195194,15.025834,13.477564,11.929294,10.382836,8.834567,7.28811,10.045626,12.803142,15.5606575,18.318174,21.07569,20.424837,19.775795,19.124943,18.474089,17.825048,19.861006,21.89515,23.929293,25.96525,27.999393,27.798155,27.595104,27.392052,27.190813,26.98776,28.6158,30.24203,31.87007,33.498108,35.124336,35.88034,36.634537,37.39054,38.144733,38.900738,40.5034,42.104244,43.7069,45.309563,46.91222,46.259552,45.606888,44.95422,44.303368,43.6507,41.065414,38.48013,35.894848,33.309563,30.724277,27.999393,25.274511,22.54963,19.824745,17.099863,16.055597,15.009518,13.965251,12.919171,11.874905,11.702674,11.530442,11.358211,11.184166,11.011934,10.192475,9.373016,8.551744,7.7322855,6.9128265,7.5056653,8.096691,8.689529,9.282369,9.875207,9.30775,8.740293,8.172835,7.605378,7.037921,7.2355337,7.4331465,7.6307597,7.8283725,8.024173,8.477413,8.930654,9.382081,9.835322,10.28675,9.561564,8.838193,8.113008,7.3878226,6.6626377,8.357758,10.052877,11.747997,13.443117,15.138238,12.697989,10.257742,7.817495,5.377247,2.9369993,2.6269827,2.3169663,2.0069497,1.696933,1.3869164,3.444629,5.5023413,7.560054,9.617766,11.675479,11.028252,10.37921,9.731983,9.084756,8.437528,7.3352466,6.2329655,5.130684,4.02659,2.9243085,2.3423476,1.7603867,1.1766127,0.5946517,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.19942589,0.40066472,0.6000906,0.7995165,1.0007553,0.7995165,0.6000906,0.40066472,0.19942589,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,1.3325275,2.6142921,3.8978696,5.179634,6.4632115,6.9581504,7.453089,7.948028,8.442966,8.937905,7.210152,5.482399,3.7546456,2.0268922,0.2991388,0.6526665,1.0043813,1.357909,1.7096237,2.0631514,3.9395678,5.8177967,7.6942134,9.572442,11.450671,9.235231,7.019791,4.804351,2.5907235,0.37528324,0.32270733,0.27013144,0.21755551,0.16497959,0.11240368,0.10333887,0.092461094,0.08339628,0.072518505,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.059827764,0.11965553,0.1794833,0.23931105,0.2991388,0.4405499,0.58014804,0.7197462,0.85934424,1.0007553,0.97718686,0.9554313,0.9318628,0.9101072,0.8883517,0.8557183,0.823085,0.7904517,0.75781834,0.72518504,0.824898,0.9246109,1.0243238,1.1258497,1.2255627,1.2726997,1.3198367,1.3669738,1.4141108,1.4630609,1.5283275,1.5917811,1.6570477,1.7223145,1.7875811,1.6044719,1.4231756,1.2400664,1.0569572,0.87566096,0.87022203,0.86478317,0.85934424,0.8557183,0.85027945,1.015259,1.1802386,1.3452182,1.5101979,1.6751775,1.6806163,1.6842422,1.6896812,1.69512,1.7005589,1.5627737,1.4249886,1.2872034,1.1494182,1.0116332,0.94274056,0.872035,0.8031424,0.7324369,0.66173136,0.7124943,0.76325727,0.8122072,0.8629702,0.9119202,0.8031424,0.69255173,0.581961,0.47318324,0.36259252,0.3480888,0.33177215,0.31726846,0.30276474,0.28826106,0.27738327,0.26831847,0.2574407,0.24837588,0.2374981,0.23568514,0.23205921,0.23024625,0.22662032,0.22480737,0.2030518,0.1794833,0.15772775,0.13415924,0.11240368,0.28463513,0.45686656,0.630911,0.8031424,0.97537386,0.89922947,0.824898,0.7505665,0.6744221,0.6000906,0.5620184,0.52575916,0.48768693,0.44961473,0.41335547,0.5529536,0.69255173,0.8321498,0.97174793,1.1131591,1.1530442,1.1929294,1.2328146,1.2726997,1.3125849,1.4648738,1.6171626,1.7694515,1.9217403,2.0758421,4.6248674,4.461701,4.3003473,4.137181,3.975827,3.8126602,3.6748753,3.53709,3.3993049,3.2633326,3.1255474,3.0131438,2.9007401,2.7883365,2.6741197,2.561716,3.2252605,3.8869917,4.550536,5.2122674,5.8758116,5.411693,4.949388,4.4870825,4.024777,3.5624714,4.2368937,4.9131284,5.5875506,6.261973,6.9382076,6.5121617,6.0879283,5.661882,5.237649,4.8116026,5.4008155,5.9882154,6.5756154,7.1630154,7.750415,7.07418,6.399758,5.7253356,5.049101,4.3746786,4.4870825,4.599486,4.7118897,4.8242936,4.936697,5.524097,6.11331,6.70071,7.28811,7.8755093,7.4367723,6.9998484,6.5629244,6.1241875,5.6872635,5.5132194,5.337362,5.163317,4.98746,4.8116026,5.475147,6.1368785,6.8004227,7.462154,8.125698,8.138389,8.149267,8.161958,8.174648,8.187339,8.363196,8.537241,8.713099,8.887142,9.063,7.911769,6.7623506,5.612932,4.461701,3.3122826,2.712192,2.1121013,1.5120108,0.9119202,0.31182957,0.50037766,0.6871128,0.87566096,1.062396,1.2491312,3.3249733,5.4008155,7.474845,9.550687,11.624716,10.7871275,9.949538,9.11195,8.274362,7.4367723,5.962834,4.4870825,3.0131438,1.5373923,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.51306844,1.0243238,1.5373923,2.0504606,2.561716,2.1628644,1.7621996,1.3633479,0.96268314,0.5620184,0.97537386,1.3869164,1.8002719,2.2118144,2.6251698,2.663242,2.6995013,2.7375734,2.7756457,2.811905,4.0120864,5.2122674,6.412449,7.61263,8.812811,8.9868555,9.162713,9.336758,9.512614,9.686659,10.687414,11.6881695,12.687112,13.687867,14.68681,14.512766,14.336908,14.162864,13.987006,13.812962,13.437678,13.062395,12.687112,12.311829,11.938358,11.650098,11.361836,11.075388,10.7871275,10.500679,10.212419,9.924157,9.637709,9.349448,9.063,9.724731,10.388275,11.050007,11.711739,12.375282,12.937301,13.499319,14.06315,14.625169,15.187187,16.012085,16.836983,17.661882,18.48678,19.311678,18.961775,18.611874,18.261972,17.912071,17.562168,16.949387,16.338419,15.725637,15.112856,14.500074,15.100165,15.700256,16.300346,16.900436,17.500528,17.437075,17.375433,17.31198,17.25034,17.186886,18.887444,20.588003,22.286749,23.987309,25.687866,24.436922,23.187792,21.936848,20.687716,19.436771,19.137632,18.836681,18.537542,18.236591,17.937452,16.788034,15.636803,14.487384,13.337966,12.186734,14.436621,16.68832,18.938208,21.188093,23.43798,21.675781,19.911768,18.149569,16.38737,14.625169,12.137785,9.6504,7.1630154,4.6756306,2.1882458,2.2498865,2.3133402,2.374981,2.4366217,2.5000753,3.3249733,4.1498713,4.974769,5.7996674,6.624565,6.450521,6.2746634,6.1006193,5.924762,5.750717,6.300045,6.849373,7.400513,7.949841,8.499168,7.8755093,7.250037,6.624565,5.999093,5.375434,5.163317,4.949388,4.7372713,4.5251546,4.313038,5.5005283,6.688019,7.8755093,9.063,10.25049,9.625018,8.999546,8.375887,7.750415,7.124943,6.037165,4.949388,3.8616104,2.7756457,1.6878681,2.137483,2.5870976,3.0367124,3.48814,3.9377546,3.1618068,2.3876717,1.6117238,0.8375887,0.06164073,3.6005437,7.137634,10.674724,14.211814,17.750717,17.60024,17.449764,17.29929,17.150625,17.00015,14.799213,12.60009,10.399154,8.200029,6.000906,5.2503395,4.499773,3.7492065,3.000453,2.2498865,3.0258346,3.7999697,4.5759177,5.3500524,6.1241875,5.9501433,5.774286,5.600241,5.424384,5.2503395,5.562169,5.8758116,6.187641,6.4994707,6.813113,7.28811,7.763106,8.238102,8.713099,9.188094,9.811753,10.437225,11.062697,11.6881695,12.311829,14.663241,17.01284,19.36244,21.71204,24.06164,23.4126,22.761745,22.112705,21.461851,20.81281,19.250036,17.687263,16.124489,14.561715,13.000754,11.5503845,10.100015,8.649645,7.1992745,5.750717,9.137331,12.525759,15.912373,19.3008,22.687414,21.525305,20.363195,19.199274,18.037165,16.875055,19.262728,21.650398,24.03807,26.425743,28.811602,28.537844,28.262274,27.986704,27.712946,27.437376,29.150625,30.862062,32.575314,34.286747,35.999996,36.513065,37.024323,37.53739,38.050457,38.561714,40.575916,42.588303,44.600693,46.61308,48.62547,47.075386,45.525303,43.97522,42.425137,40.875053,37.825653,34.774437,31.725033,28.675629,25.624413,23.213173,20.80012,18.387066,15.975826,13.562773,13.049705,12.536636,12.025381,11.512312,10.999244,10.837891,10.674724,10.51337,10.3502035,10.1870365,9.625018,9.063,8.499168,7.93715,7.3751316,7.9752226,8.575313,9.175404,9.775495,10.375585,9.438283,8.499168,7.5618668,6.624565,5.6872635,5.7996674,5.9120708,6.0244746,6.1368785,6.249282,7.112252,7.9752226,8.838193,9.699349,10.56232,8.950596,7.3370595,5.7253356,4.1117992,2.5000753,5.0744824,7.650702,10.225109,12.799516,15.375735,12.474996,9.574255,6.6753283,3.774588,0.87566096,0.9246109,0.97537386,1.0243238,1.0750868,1.1258497,3.0747845,5.0255322,6.9744673,8.925215,10.874149,10.2378,9.599637,8.963287,8.325124,7.686961,6.813113,5.9374523,5.0617914,4.1879435,3.3122826,2.6505513,1.987007,1.3252757,0.66173136,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.25018883,0.50037766,0.7505665,1.0007553,1.2491312,1.0007553,0.7505665,0.50037766,0.25018883,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,1.6624867,3.2633326,4.8623657,6.4632115,8.062244,8.636953,9.211663,9.788185,10.362894,10.937603,8.80012,6.6626377,4.5251546,2.3876717,0.25018883,0.7124943,1.1747998,1.6371052,2.0994108,2.561716,4.9131284,7.262728,9.612328,11.961927,14.313339,11.450671,8.588004,5.7253356,2.8626678,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.16316663,0.19942589,0.2374981,0.2755703,0.31182957,0.31182957,0.31182957,0.31182957,0.31182957,0.31182957,0.2991388,0.28826106,0.2755703,0.26287958,0.25018883,0.25018883,0.25018883,0.25018883,0.25018883,0.25018883,0.25018883,0.25018883,0.25018883,0.25018883,0.25018883,0.25018883,0.25018883,0.25018883,0.25018883,0.25018883,0.22480737,0.19942589,0.17585737,0.15047589,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.21211663,0.2991388,0.387974,0.4749962,0.5620184,0.824898,1.0877775,1.3506571,1.6117238,1.8746033,4.4127507,4.2876563,4.162562,4.0374675,3.9123733,3.787279,3.63499,3.482701,3.3304121,3.1781235,3.0258346,2.9369993,2.8499773,2.762955,2.6741197,2.5870976,3.1128569,3.636803,4.162562,4.688321,5.2122674,4.835171,4.458075,4.079166,3.7020695,3.3249733,4.0320287,4.7390842,5.4479527,6.155008,6.8620634,6.6082487,6.352621,6.096993,5.8431783,5.5875506,6.3272395,7.066928,7.8084297,8.548119,9.287807,8.375887,7.462154,6.550234,5.638314,4.7245803,4.9657044,5.2050157,5.4443264,5.6854506,5.924762,6.2220874,6.5194135,6.816739,7.115878,7.413204,7.0052876,6.5973706,6.189454,5.7833505,5.375434,5.335549,5.295664,5.2557783,5.2158933,5.1741953,5.6945157,6.2148356,6.735156,7.2554765,7.7757964,8.221786,8.669587,9.117389,9.56519,10.012992,9.7773075,9.541622,9.30775,9.072064,8.838193,7.650702,6.4632115,5.275721,4.0882306,2.9007401,2.373168,1.845596,1.3180238,0.7904517,0.26287958,0.4169814,0.5728962,0.726998,0.88291276,1.0370146,3.6295512,6.2220874,8.814624,11.407161,13.999697,12.496751,10.995618,9.492672,7.989726,6.48678,5.199577,3.9123733,2.6251698,1.3379664,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.41516843,0.83033687,1.2455053,1.6606737,2.0758421,2.124792,2.175555,2.2245052,2.275268,2.324218,2.1646774,2.0051367,1.845596,1.6842422,1.5247015,1.9471219,2.3695421,2.7919624,3.2143826,3.636803,3.6549325,3.673062,3.6893787,3.7075086,3.7256382,4.59586,5.464269,6.3344913,7.2047133,8.074935,8.39039,8.705847,9.019489,9.334945,9.6504,10.46442,11.280253,12.094274,12.910107,13.724127,13.435865,13.145792,12.855718,12.565643,12.27557,12.114216,11.954676,11.795135,11.635593,11.47424,11.447045,11.419851,11.392657,11.365462,11.338268,10.93579,10.533313,10.130835,9.728357,9.325879,9.857078,10.390089,10.9230995,11.454298,11.9873085,12.621845,13.258195,13.892733,14.527269,15.161806,15.792717,16.421816,17.052727,17.681824,18.312735,17.951956,17.592989,17.23221,16.873243,16.512463,16.305786,16.097294,15.890617,15.682126,15.475449,15.872487,16.269526,16.668379,17.065416,17.462456,17.513218,17.562168,17.612932,17.661882,17.712645,19.235533,20.756609,22.279497,23.802385,25.325274,24.652666,23.980057,23.307447,22.634838,21.962229,21.857077,21.751925,21.646772,21.541622,21.438282,20.074934,18.7134,17.350052,15.986704,14.625169,16.563227,18.49947,20.437527,22.375584,24.311829,22.451729,20.593443,18.733343,16.873243,15.013144,13.270886,11.526816,9.784559,8.042302,6.300045,6.495845,6.6898317,6.885632,7.079619,7.2754188,7.0904965,6.9055743,6.720652,6.53573,6.350808,6.089741,5.8304877,5.569421,5.3101673,5.049101,5.5367875,6.0244746,6.5121617,6.9998484,7.4875355,7.208339,6.92733,6.6481338,6.3671246,6.0879283,5.67276,5.2575917,4.842423,4.4272547,4.0120864,5.06723,6.1223745,7.177519,8.232663,9.287807,8.709473,8.13295,7.554615,6.978093,6.399758,5.5005283,4.599486,3.7002566,2.7992141,1.8999848,2.1501737,2.4003625,2.6505513,2.9007401,3.149116,3.2016919,3.254268,3.3068438,3.3594196,3.4119956,5.826862,8.241728,10.658407,13.073273,15.488139,15.442815,15.397491,15.352167,15.306843,15.263332,13.464873,11.668227,9.869768,8.073122,6.2746634,5.40988,4.5450974,3.680314,2.8155308,1.9507477,2.5526514,3.1545548,3.7582715,4.360175,4.9620786,4.8623657,4.762653,4.6629395,4.5632267,4.461701,4.9131284,5.3627434,5.812358,6.261973,6.7134004,7.2482243,7.783048,8.317872,8.852696,9.38752,9.824444,10.263181,10.700105,11.137029,11.575767,13.555521,15.535276,17.515032,19.494787,21.474543,20.852695,20.23085,19.607191,18.985344,18.361685,17.515032,16.668379,15.819912,14.973258,14.124791,13.245504,12.364405,11.485118,10.605831,9.724731,12.549327,15.375735,18.20033,21.024927,23.849524,22.725487,21.599636,20.4756,19.34975,18.225714,20.345066,22.464418,24.585585,26.704939,28.824291,28.300346,27.774588,27.25064,26.724882,26.199121,28.41275,30.624563,32.838192,35.050007,37.26182,37.076897,36.891975,36.707054,36.522133,36.337208,37.510197,38.68318,39.854355,41.027344,42.20033,40.73002,39.259705,37.78939,36.31908,34.85058,32.363194,29.87581,27.386612,24.89923,22.411844,20.397642,18.38344,16.367426,14.353225,12.337211,12.103338,11.867653,11.631968,11.398096,11.162411,10.932164,10.701918,10.471672,10.243238,10.012992,9.557939,9.102885,8.647832,8.192778,7.7377243,8.225411,8.713099,9.200785,9.686659,10.174346,9.066626,7.9607186,6.8529987,5.7452784,4.6375585,4.860553,5.081734,5.3047285,5.527723,5.750717,6.5157876,7.2808576,8.044115,8.809185,9.574255,8.70222,7.8301854,6.9581504,6.0843024,5.2122674,6.885632,8.557183,10.230548,11.9021,13.575464,11.4416065,9.309563,7.177519,5.045475,2.911618,2.6469254,2.382233,2.1175404,1.8528478,1.5881553,3.3195345,5.0527267,6.7859187,8.517298,10.25049,9.440096,8.629702,7.819308,7.0107265,6.200332,5.4950895,4.7898474,4.0846047,3.3793623,2.6741197,2.1392958,1.6044719,1.0696479,0.53482395,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.21574254,0.42967212,0.64541465,0.85934424,1.0750868,0.90285534,0.7306239,0.55839247,0.38434806,0.21211663,0.7904517,1.3669738,1.9453088,2.521831,3.100166,2.4873846,1.8746033,1.261822,0.6508536,0.038072214,0.07795739,0.11784257,0.15772775,0.19761293,0.2374981,1.7857682,3.3322253,4.880495,6.4269524,7.9752226,8.165584,8.354132,8.544493,8.734854,8.925215,7.315304,5.7053933,4.0954823,2.4855716,0.87566096,1.1457924,1.4141108,1.6842422,1.9543737,2.2245052,4.070101,5.915697,7.75948,9.605076,11.450671,9.159087,6.869315,4.5795436,2.2897718,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.11421664,0.13053331,0.14503701,0.15954071,0.17585737,0.14503701,0.11421664,0.08520924,0.054388877,0.025381476,0.032633327,0.03988518,0.047137026,0.054388877,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.04169814,0.072518505,0.10333887,0.13234627,0.16316663,0.13234627,0.10333887,0.072518505,0.04169814,0.012690738,0.014503701,0.018129626,0.01994259,0.02175555,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.13415924,0.17041849,0.20486477,0.23931105,0.2755703,0.27738327,0.27919623,0.28282216,0.28463513,0.28826106,0.27738327,0.26831847,0.2574407,0.24837588,0.2374981,0.2374981,0.2374981,0.2374981,0.2374981,0.2374981,0.23568514,0.23205921,0.23024625,0.22662032,0.22480737,0.23024625,0.23568514,0.23931105,0.24474995,0.25018883,0.23024625,0.21030366,0.19036107,0.17041849,0.15047589,0.13959812,0.13053331,0.11965553,0.11059072,0.099712946,0.10696479,0.11421664,0.12328146,0.13053331,0.13778515,0.13234627,0.12690738,0.12328146,0.11784257,0.11240368,0.11240368,0.11240368,0.11240368,0.11240368,0.11240368,0.18310922,0.2520018,0.32270733,0.39159992,0.46230546,0.6726091,0.88291276,1.0932164,1.3017071,1.5120108,4.2006345,4.1117992,4.024777,3.9377546,3.8507326,3.7618973,3.5951047,3.4283123,3.2597067,3.092914,2.9243085,2.8626678,2.7992141,2.7375734,2.6741197,2.612479,3.000453,3.386614,3.774588,4.162562,4.550536,4.256836,3.9649491,3.673062,3.3793623,3.0874753,3.827164,4.5668526,5.3083544,6.0480433,6.787732,6.7025228,6.6173134,6.532104,6.446895,6.3616858,7.2554765,8.147454,9.039432,9.933222,10.825199,9.675781,8.52455,7.3751316,6.2257137,5.0744824,5.4425135,5.810545,6.1767635,6.544795,6.9128265,6.9200783,6.92733,6.9345818,6.9418335,6.9508986,6.5719895,6.1948934,5.8177967,5.4407005,5.0617914,5.1578784,5.2521524,5.3482394,5.4425135,5.5367875,5.915697,6.2927933,6.6698895,7.0469856,7.4258947,8.306994,9.189907,10.07282,10.955733,11.836833,11.193231,10.547816,9.902402,9.256987,8.613385,7.3878226,6.16226,4.936697,3.7129474,2.4873846,2.032331,1.5772774,1.1222239,0.6671702,0.21211663,0.33539808,0.45686656,0.58014804,0.7016165,0.824898,3.9341288,7.0451727,10.154404,13.265448,16.374678,14.208188,12.039885,9.871581,7.705091,5.5367875,4.4381323,3.3376641,2.2371957,1.1367276,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.83033687,1.6606737,2.4891977,3.3195345,4.1498713,3.738329,3.3249733,2.911618,2.5000753,2.08672,2.1683033,2.2480736,2.327844,2.4076142,2.4873846,2.9206827,3.3521678,3.785466,4.216951,4.650249,4.646623,4.64481,4.6429973,4.6393714,4.6375585,5.177821,5.718084,6.258347,6.796797,7.3370595,7.7921133,8.247167,8.70222,9.157274,9.612328,10.243238,10.872336,11.503247,12.132345,12.763257,12.357153,11.952863,11.546759,11.142468,10.738177,10.792566,10.846955,10.903157,10.957546,11.011934,11.245807,11.477866,11.709926,11.941984,12.175857,11.65735,11.1406555,10.622148,10.1054535,9.5869465,9.989424,10.391902,10.794379,11.1968565,11.599335,12.308203,13.015259,13.722314,14.429369,15.138238,15.573349,16.006647,16.441757,16.87687,17.31198,16.942135,16.57229,16.202446,15.8326025,15.462758,15.660371,15.857984,16.055597,16.25321,16.450823,16.64481,16.840609,17.034595,17.230396,17.424383,17.58755,17.750717,17.912071,18.075237,18.238403,19.581808,20.927027,22.272245,23.617464,24.962683,24.868408,24.77232,24.678047,24.581959,24.487686,24.578333,24.66717,24.757816,24.846653,24.9373,23.361835,21.788185,20.212719,18.637255,17.06179,18.688019,20.312433,21.936848,23.563074,25.187489,23.22949,21.273302,19.315304,17.357304,15.399304,14.402175,13.4050455,12.407916,11.410787,10.411844,10.73999,11.068136,11.39447,11.722616,12.050762,10.854207,9.659465,8.464723,7.26998,6.0752378,5.730775,5.384499,5.040036,4.695573,4.349297,4.7753434,5.199577,5.6256227,6.049856,6.474089,6.539356,6.604623,6.6698895,6.735156,6.8004227,6.1822023,5.565795,4.947575,4.329355,3.7129474,4.6357455,5.5567303,6.4795284,7.402326,8.325124,7.795739,7.264541,6.735156,6.205771,5.674573,4.9620786,4.249584,3.53709,2.8245957,2.1121013,2.1628644,2.2118144,2.2625773,2.3133402,2.3622901,3.24339,4.122677,5.0019636,5.883064,6.7623506,8.054993,9.347635,10.640278,11.9329195,13.225562,13.28539,13.345218,13.4050455,13.464873,13.524701,12.130532,10.734551,9.340384,7.944402,6.550234,5.569421,4.590421,3.6096084,2.6306088,1.649796,2.079468,2.5091403,2.9406252,3.3702974,3.7999697,3.774588,3.7492065,3.7256382,3.7002566,3.6748753,4.262275,4.8496747,5.4370747,6.0244746,6.6118746,7.208339,7.802991,8.397643,8.992294,9.5869465,9.837135,10.087324,10.337513,10.587702,10.837891,12.447801,14.057712,15.667623,17.277533,18.887444,18.292793,17.698141,17.101677,16.507025,15.912373,15.780026,15.64768,15.515334,15.382988,15.250641,14.940624,14.630608,14.320591,14.010575,13.700559,15.963136,18.225714,20.48829,22.750868,25.011631,23.925667,22.837889,21.750113,20.662334,19.574556,21.427404,23.280252,25.1331,26.984135,28.836983,28.062847,27.2869,26.512764,25.736816,24.962683,27.674873,30.387066,33.09926,35.813263,38.525455,37.642544,36.75963,35.876717,34.995617,34.112705,34.444477,34.77806,35.109833,35.441605,35.775192,34.384647,32.994106,31.605377,30.214834,28.824291,26.90074,24.975372,23.050007,21.12464,19.199274,17.582111,15.964949,14.347786,12.730623,11.111648,11.155159,11.1968565,11.240368,11.282066,11.325577,11.028252,10.729113,10.431787,10.13446,9.837135,9.490859,9.142771,8.794682,8.446592,8.100317,8.4756,8.8508835,9.224354,9.599637,9.97492,8.696781,7.420456,6.1423173,4.8641787,3.587853,3.919625,4.25321,4.5849824,4.9167547,5.2503395,5.91751,6.58468,7.25185,7.9208336,8.588004,8.455658,8.323311,8.189152,8.056806,7.9244595,8.694968,9.465478,10.234174,11.004683,11.775192,10.410031,9.04487,7.6797094,6.3145485,4.949388,4.36924,3.7909048,3.2107568,2.6306088,2.0504606,3.5642843,5.0799212,6.5955577,8.109382,9.625018,8.642392,7.6597667,6.677141,5.6945157,4.7118897,4.177066,3.6422417,3.1074178,2.572594,2.03777,1.6298534,1.2219368,0.81583315,0.40791658,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1794833,0.36077955,0.5402629,0.7197462,0.89922947,0.80495536,0.7106813,0.61459434,0.52032024,0.42423326,1.5809034,2.7357605,3.8906176,5.045475,6.200332,4.974769,3.7492065,2.525457,1.2998942,0.07433146,0.14322405,0.21030366,0.27738327,0.3444629,0.41335547,1.9072367,3.4029307,4.896812,6.392506,7.8882003,7.6924005,7.4966,7.3026133,7.1068134,6.9128265,5.8304877,4.748149,3.6658103,2.5816586,1.49932,1.5772774,1.6552348,1.7331922,1.8093367,1.887294,3.2270734,4.5668526,5.906632,7.2482243,8.588004,6.869315,5.1524396,3.435564,1.7168756,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.11784257,0.15954071,0.2030518,0.24474995,0.28826106,0.23931105,0.19217403,0.14503701,0.09789998,0.05076295,0.052575916,0.054388877,0.058014803,0.059827764,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.047137026,0.07070554,0.092461094,0.11421664,0.13778515,0.11421664,0.092461094,0.07070554,0.047137026,0.025381476,0.030820364,0.034446288,0.03988518,0.045324065,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.10696479,0.13959812,0.17223145,0.20486477,0.2374981,0.24293698,0.24837588,0.2520018,0.2574407,0.26287958,0.25562772,0.24837588,0.23931105,0.23205921,0.22480737,0.22480737,0.22480737,0.22480737,0.22480737,0.22480737,0.21936847,0.21574254,0.21030366,0.20486477,0.19942589,0.21030366,0.21936847,0.23024625,0.23931105,0.25018883,0.23568514,0.21936847,0.20486477,0.19036107,0.17585737,0.16679256,0.15954071,0.15228885,0.14503701,0.13778515,0.13959812,0.14322405,0.14503701,0.14684997,0.15047589,0.13959812,0.13053331,0.11965553,0.11059072,0.099712946,0.099712946,0.099712946,0.099712946,0.099712946,0.099712946,0.15228885,0.20486477,0.2574407,0.3100166,0.36259252,0.52032024,0.678048,0.83577573,0.9916905,1.1494182,3.9867048,3.9377546,3.8869917,3.8380418,3.787279,3.738329,3.5552197,3.3721104,3.1908143,3.007705,2.8245957,2.7883365,2.7502642,2.712192,2.6741197,2.6378605,2.8880494,3.1382382,3.386614,3.636803,3.8869917,3.680314,3.4718235,3.2651455,3.056655,2.8499773,3.6222992,4.3946214,5.1669436,5.9392653,6.7134004,6.796797,6.882006,6.967215,7.0524244,7.137634,8.1819,9.22798,10.272246,11.318325,12.362592,10.975676,9.5869465,8.200029,6.813113,5.424384,5.919323,6.414262,6.9092,7.404139,7.900891,7.6180687,7.3352466,7.0524244,6.7696023,6.48678,6.1405044,5.7924156,5.4443264,5.0980506,4.749962,4.9802084,5.2104545,5.4407005,5.669134,5.89938,6.1350656,6.3707504,6.604623,6.8403077,7.07418,8.392203,9.710228,11.028252,12.344462,13.662486,12.607342,11.552197,10.497053,9.441909,8.386765,7.124943,5.863121,4.599486,3.3376641,2.0758421,1.693307,1.310772,0.92823684,0.54570174,0.16316663,0.2520018,0.34264994,0.43329805,0.52213323,0.61278135,4.2405195,7.8682575,11.4959955,15.121921,18.749659,15.917811,13.085964,10.252303,7.420456,4.5867953,3.6748753,2.762955,1.8492218,0.93730164,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,1.2455053,2.4891977,3.7347028,4.9802084,6.2257137,5.3500524,4.4743915,3.6005437,2.7248828,1.8492218,2.1701162,2.4891977,2.810092,3.1291735,3.4500678,3.8924308,4.3347936,4.7771564,5.219519,5.661882,5.6401267,5.618371,5.5948024,5.573047,5.5494785,5.7597823,5.9700856,6.1803894,6.390693,6.599184,7.1956487,7.7903004,8.384952,8.979604,9.574255,10.020245,10.46442,10.910409,11.354585,11.800573,11.280253,10.7599325,10.239613,9.719293,9.200785,9.469104,9.739235,10.009366,10.279498,10.549629,11.042755,11.535881,12.027194,12.52032,13.011633,12.380721,11.747997,11.115273,10.48255,9.849826,10.12177,10.395528,10.667472,10.939416,11.213174,11.992747,12.772322,13.551895,14.333282,15.112856,15.352167,15.593291,15.8326025,16.071913,16.313038,15.932315,15.553406,15.172684,14.791962,14.413053,15.014956,15.616859,16.220575,16.82248,17.424383,17.417131,17.40988,17.402628,17.395376,17.388124,17.661882,17.937452,18.213022,18.48678,18.76235,19.929897,21.097446,22.264994,23.43254,24.60009,25.082336,25.564585,26.046833,26.530895,27.013142,27.297777,27.582413,27.867048,28.151684,28.438131,26.65055,24.862968,23.075388,21.287807,19.500225,20.81281,22.125395,23.43798,24.750565,26.06315,24.00725,21.953163,19.897264,17.843178,15.787278,15.535276,15.283275,15.02946,14.777458,14.525456,14.984136,15.444629,15.905121,16.365614,16.824293,14.61973,12.415168,10.210606,8.00423,5.7996674,5.369995,4.940323,4.510651,4.079166,3.6494937,4.0120864,4.3746786,4.7372713,5.0998635,5.462456,5.8721857,6.281915,6.6916447,7.1031876,7.512917,6.6916447,5.8721857,5.0527267,4.233268,3.4119956,4.2024474,4.992899,5.7833505,6.5719895,7.362441,6.880193,6.397945,5.915697,5.431636,4.949388,4.4254417,3.8996825,3.3757362,2.8499773,2.324218,2.175555,2.0250793,1.8746033,1.7241274,1.5754645,3.2832751,4.989273,6.697084,8.404895,10.112705,10.283124,10.451729,10.622148,10.792566,10.962985,11.127964,11.292944,11.457924,11.622903,11.787883,10.794379,9.802689,8.809185,7.817495,6.825804,5.730775,4.6357455,3.540716,2.4456866,1.3506571,1.6080978,1.8655385,2.1229792,2.38042,2.6378605,2.6868105,2.7375734,2.7883365,2.8372865,2.8880494,3.6132345,4.3366065,5.0617914,5.7869763,6.5121617,7.166641,7.8229337,8.477413,9.131892,9.788185,9.849826,9.91328,9.97492,10.038374,10.100015,11.340081,12.580148,13.820213,15.06028,16.300346,15.732889,15.165432,14.597975,14.030518,13.46306,14.045021,14.626982,15.210756,15.792717,16.374678,16.635744,16.894999,17.154251,17.41532,17.674572,19.375132,21.07569,22.774435,24.474995,26.175554,25.124035,24.07433,23.024624,21.97492,20.925215,22.509743,24.094273,25.680614,27.265144,28.849674,27.82535,26.799213,25.774889,24.750565,23.724428,26.936998,30.149569,33.362137,36.574707,39.787277,38.208187,36.62728,35.04819,33.46729,31.888199,31.38057,30.87294,30.36531,29.857681,29.350052,28.03928,26.73032,25.419548,24.11059,22.799818,21.438282,20.074934,18.711586,17.350052,15.986704,14.766581,13.548269,12.328146,11.108022,9.8878975,10.20698,10.527874,10.846955,11.16785,11.486931,11.122525,10.75812,10.391902,10.027496,9.663091,9.421967,9.182655,8.943344,8.70222,8.46291,8.725789,8.9868555,9.249735,9.512614,9.775495,8.326937,6.880193,5.431636,3.9848917,2.5381477,2.9805105,3.4228733,3.8652363,4.307599,4.749962,5.319232,5.8903155,6.4595857,7.0306687,7.5999393,8.207282,8.814624,9.421967,10.029309,10.636651,10.504305,10.371959,10.239613,10.107266,9.97492,9.376642,8.780178,8.1819,7.5854354,6.987158,6.091554,5.197764,4.3021603,3.4083695,2.5127661,3.8108473,5.1071157,6.4051967,7.703278,8.999546,7.844689,6.6898317,5.5349746,4.3801174,3.2252605,2.8608549,2.4946365,2.1302311,1.7658255,1.3996071,1.1204109,0.83940166,0.56020546,0.27919623,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14503701,0.29007402,0.43511102,0.58014804,0.72518504,0.7070554,0.69073874,0.6726091,0.6544795,0.63816285,2.3695421,4.102734,5.8359265,7.567306,9.300498,7.462154,5.6256227,3.787279,1.9507477,0.11240368,0.20667773,0.30276474,0.39703882,0.49312583,0.5873999,2.030518,3.4718235,4.914942,6.35806,7.799365,7.219217,6.640882,6.060734,5.480586,4.900438,4.345671,3.7909048,3.2343252,2.6795588,2.124792,2.0105755,1.8945459,1.7803292,1.6642996,1.550083,2.3858588,3.2198215,4.0555973,4.88956,5.7253356,4.5795436,3.435564,2.2897718,1.1457924,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.11965553,0.19036107,0.25925365,0.32995918,0.40066472,0.33539808,0.27013144,0.20486477,0.13959812,0.07433146,0.072518505,0.07070554,0.06707962,0.065266654,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.052575916,0.06707962,0.08339628,0.09789998,0.11240368,0.09789998,0.08339628,0.06707962,0.052575916,0.038072214,0.045324065,0.052575916,0.059827764,0.06707962,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.07977036,0.11059072,0.13959812,0.17041849,0.19942589,0.20667773,0.21574254,0.2229944,0.23024625,0.2374981,0.23205921,0.22662032,0.2229944,0.21755551,0.21211663,0.21211663,0.21211663,0.21211663,0.21211663,0.21211663,0.20486477,0.19761293,0.19036107,0.18310922,0.17585737,0.19036107,0.20486477,0.21936847,0.23568514,0.25018883,0.23931105,0.23024625,0.21936847,0.21030366,0.19942589,0.19579996,0.19036107,0.18492219,0.1794833,0.17585737,0.17223145,0.17041849,0.16679256,0.16497959,0.16316663,0.14684997,0.13234627,0.11784257,0.10333887,0.0870222,0.0870222,0.0870222,0.0870222,0.0870222,0.0870222,0.12328146,0.15772775,0.19217403,0.22662032,0.26287958,0.3680314,0.47318324,0.57833505,0.68167394,0.7868258,3.774588,3.7618973,3.7492065,3.738329,3.7256382,3.7129474,3.5153344,3.3177216,3.1201086,2.9224956,2.7248828,2.712192,2.6995013,2.6868105,2.6741197,2.663242,2.7756457,2.8880494,3.000453,3.1128569,3.2252605,3.101979,2.9805105,2.857229,2.7357605,2.612479,3.4174345,4.2223897,5.027345,5.8323007,6.637256,6.892884,7.1466985,7.402326,7.6579537,7.911769,9.110137,10.306692,11.50506,12.701616,13.899984,12.27557,10.649343,9.024928,7.400513,5.774286,6.397945,7.019791,7.6416373,8.265296,8.887142,8.314246,7.743163,7.170267,6.5973706,6.0244746,5.7072062,5.389938,5.0726695,4.7554007,4.4381323,4.802538,5.1669436,5.5331616,5.8975673,6.261973,6.354434,6.446895,6.539356,6.6318173,6.7242785,8.477413,10.230548,11.98187,13.735004,15.488139,14.023266,12.558392,11.091705,9.626831,8.161958,6.8620634,5.562169,4.262275,2.962381,1.6624867,1.35247,1.0424535,0.7324369,0.4224203,0.11240368,0.17041849,0.22662032,0.28463513,0.34264994,0.40066472,4.5450974,8.689529,12.835775,16.980207,21.12464,17.627436,14.13023,10.633025,7.135821,3.636803,2.911618,2.1882458,1.4630609,0.73787576,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,1.6606737,3.3195345,4.9802084,6.640882,8.299743,6.9617763,5.6256227,4.2876563,2.94969,1.6117238,2.1719291,2.7321346,3.29234,3.8525455,4.4127507,4.8641787,5.317419,5.77066,6.2220874,6.6753283,6.6318173,6.590119,6.546608,6.5049095,6.4632115,6.341743,6.2220874,6.1024323,5.9827766,5.863121,6.5973706,7.3316207,8.067683,8.801933,9.537996,9.79725,10.058316,10.31757,10.576823,10.837891,10.203354,9.567003,8.9324665,8.29793,7.663393,8.147454,8.6333275,9.117389,9.603263,10.087324,10.839704,11.592083,12.344462,13.096842,13.849221,13.102281,12.35534,11.606586,10.859646,10.112705,10.254116,10.397341,10.540565,10.681975,10.825199,11.677292,12.529385,13.383289,14.235382,15.087475,15.132799,15.1781225,15.221634,15.266958,15.312282,14.922495,14.532708,14.142921,13.753134,13.363347,14.369541,15.377548,16.385555,17.39175,18.399757,18.189453,17.97915,17.770658,17.560356,17.350052,17.738026,18.124187,18.512161,18.900135,19.288109,20.277987,21.267864,22.257742,23.24762,24.237497,25.29808,26.35685,27.417433,28.478016,29.536787,30.017221,30.497656,30.978092,31.456715,31.93715,29.93745,27.937754,25.938055,23.938358,21.936848,22.937603,23.938358,24.9373,25.938055,26.936998,24.785011,22.633024,20.479225,18.327238,16.175253,16.668379,17.15969,17.652817,18.144129,18.637255,19.230095,19.822933,20.415771,21.006798,21.599636,18.385254,15.170871,11.954676,8.740293,5.524097,5.009216,4.494334,3.9794528,3.4645715,2.94969,3.2506418,3.5497808,3.8507326,4.1498713,4.4508233,5.2050157,5.959208,6.7152133,7.4694057,8.225411,7.2029004,6.1803894,5.1578784,4.135368,3.1128569,3.7691493,4.4272547,5.08536,5.7416525,6.399758,5.964647,5.529536,5.0944247,4.6593137,4.2242026,3.8869917,3.5497808,3.2125697,2.8753586,2.5381477,2.1882458,1.8383441,1.4866294,1.1367276,0.7868258,3.3231604,5.857682,8.392203,10.926725,13.46306,12.509441,11.557636,10.605831,9.652213,8.700407,8.970539,9.24067,9.510801,9.77912,10.049252,9.460039,8.870826,8.2798,7.690587,7.0995617,5.8903155,4.6792564,3.4700103,2.2607644,1.0497054,1.1349145,1.2201238,1.305333,1.3905423,1.4757515,1.6008459,1.7241274,1.8492218,1.9743162,2.0994108,2.962381,3.825351,4.688321,5.5494785,6.412449,7.1267557,7.842876,8.557183,9.273304,9.987611,9.862516,9.737422,9.612328,9.487233,9.362139,10.232361,11.102583,11.972805,12.843027,13.713249,13.172986,12.632723,12.092461,11.552197,11.011934,12.310016,13.608097,14.904366,16.202446,17.500528,18.330864,19.15939,19.989725,20.820063,21.650398,22.787127,23.925667,25.062395,26.199121,27.337664,26.324217,25.312584,24.299137,23.287504,22.275871,23.592083,24.910107,26.22813,27.54434,28.862364,27.587852,26.31334,25.037014,23.7625,22.487988,26.200935,29.91207,33.625015,37.337963,41.0491,38.77202,36.494938,34.217857,31.940775,29.66188,28.31485,26.96782,25.620787,24.271942,22.924911,21.695723,20.464722,19.235533,18.004532,16.775343,15.975826,15.174497,14.37498,13.575464,12.774135,11.952863,11.129777,10.306692,9.48542,8.662335,9.2606125,9.857078,10.455356,11.05182,11.650098,11.2168,10.785315,10.352016,9.920531,9.487233,9.354887,9.222541,9.090195,8.957849,8.825501,8.974165,9.12464,9.275117,9.425592,9.574255,7.957093,6.33993,4.7227674,3.105605,1.4866294,2.039583,2.5925364,3.1454902,3.6966307,4.249584,4.7227674,5.1941376,5.667321,6.1405044,6.6118746,7.9607186,9.30775,10.654781,12.001812,13.3506565,12.3154545,11.280253,10.245051,9.20985,8.174648,8.345067,8.515485,8.685904,8.854509,9.024928,7.8156815,6.604623,5.3953767,4.1843176,2.9750717,4.0555973,5.1343102,6.2148356,7.2953615,8.375887,7.0469856,5.719897,4.3928084,3.0657198,1.7368182,1.5428312,1.3470312,1.1530442,0.9572442,0.76325727,0.6091554,0.45686656,0.3045777,0.15228885,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.11059072,0.21936847,0.32995918,0.4405499,0.5493277,0.6091554,0.67079616,0.7306239,0.7904517,0.85027945,3.159994,5.469708,7.7794223,10.089137,12.400664,9.949538,7.500226,5.049101,2.5997884,0.15047589,0.27194437,0.39522585,0.5166943,0.6399758,0.76325727,2.1519866,3.5425289,4.933071,6.3218007,7.7123427,6.7478466,5.7833505,4.8170414,3.8525455,2.8880494,2.8608549,2.8318477,2.8046532,2.7774587,2.7502642,2.4420607,2.13567,1.8274662,1.5192627,1.2128719,1.5428312,1.8727903,2.2027495,2.5327086,2.8626678,2.2897718,1.7168756,1.1457924,0.5728962,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.12328146,0.21936847,0.31726846,0.41516843,0.51306844,0.42967212,0.3480888,0.26469254,0.18310922,0.099712946,0.092461094,0.08520924,0.07795739,0.07070554,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.058014803,0.065266654,0.072518505,0.07977036,0.0870222,0.07977036,0.072518505,0.065266654,0.058014803,0.05076295,0.059827764,0.07070554,0.07977036,0.09064813,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.052575916,0.07977036,0.10696479,0.13415924,0.16316663,0.17223145,0.18310922,0.19217403,0.2030518,0.21211663,0.21030366,0.20667773,0.20486477,0.2030518,0.19942589,0.19942589,0.19942589,0.19942589,0.19942589,0.19942589,0.19036107,0.1794833,0.17041849,0.15954071,0.15047589,0.17041849,0.19036107,0.21030366,0.23024625,0.25018883,0.24474995,0.23931105,0.23568514,0.23024625,0.22480737,0.2229944,0.21936847,0.21755551,0.21574254,0.21211663,0.20486477,0.19761293,0.19036107,0.18310922,0.17585737,0.15410182,0.13415924,0.11421664,0.09427405,0.07433146,0.07433146,0.07433146,0.07433146,0.07433146,0.07433146,0.092461094,0.11059072,0.12690738,0.14503701,0.16316663,0.21574254,0.26831847,0.3208944,0.37165734,0.42423326,3.5624714,3.587853,3.6132345,3.636803,3.6621845,3.6875658,3.4754493,3.2633326,3.049403,2.8372865,2.6251698,2.6378605,2.6505513,2.663242,2.6741197,2.6868105,2.663242,2.6378605,2.612479,2.5870976,2.561716,2.525457,2.4873846,2.4493124,2.4130533,2.374981,3.2125697,4.0501585,4.8877473,5.7253356,6.5629244,6.987158,7.413204,7.837437,8.26167,8.6877165,10.038374,11.3872175,12.737875,14.0867195,15.437376,13.575464,11.711739,9.849826,7.987913,6.1241875,6.874754,7.6253204,8.375887,9.12464,9.875207,9.012237,8.149267,7.28811,6.4251394,5.562169,5.275721,4.98746,4.699199,4.4127507,4.12449,4.6248674,5.125245,5.6256227,6.1241875,6.624565,6.5756154,6.5248523,6.4759026,6.4251394,6.3743763,8.562622,10.749055,12.937301,15.125546,17.31198,15.437376,13.562773,11.6881695,9.811753,7.93715,6.599184,5.2630305,3.925064,2.5870976,1.2491312,1.0116332,0.774135,0.53663695,0.2991388,0.06164073,0.0870222,0.11240368,0.13778515,0.16316663,0.18673515,4.8496747,9.512614,14.175554,18.836681,23.49962,19.337059,15.174497,11.011934,6.849373,2.6868105,2.1501737,1.6117238,1.0750868,0.53663695,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.0758421,4.1498713,6.2257137,8.299743,10.375585,8.575313,6.775041,4.974769,3.1744974,1.3742256,2.175555,2.9750717,3.774588,4.5759177,5.375434,5.8377395,6.300045,6.7623506,7.224656,7.686961,7.6253204,7.5618668,7.500226,7.4367723,7.3751316,6.925517,6.4759026,6.0244746,5.57486,5.125245,5.999093,6.874754,7.750415,8.624263,9.499924,9.574255,9.6504,9.724731,9.800876,9.875207,9.12464,8.375887,7.6253204,6.874754,6.1241875,6.825804,7.5256076,8.225411,8.925215,9.625018,10.636651,11.650098,12.661731,13.675177,14.68681,13.825653,12.962683,12.099712,11.236742,10.375585,10.388275,10.399154,10.411844,10.424535,10.437225,11.361836,12.28826,13.212872,14.137483,15.062093,14.911617,14.762955,14.612478,14.462003,14.313339,13.912675,13.512011,13.113158,12.712494,12.311829,13.724127,15.138238,16.550535,17.962833,19.375132,18.961775,18.550234,18.136877,17.725336,17.31198,17.812357,18.312735,18.813112,19.311678,19.812056,20.624262,21.438282,22.25049,23.062696,23.874905,25.512009,27.149115,28.788033,30.425138,32.062244,32.736664,33.4129,34.087322,34.761745,35.43798,33.224354,31.012537,28.800724,26.587097,24.375282,25.062395,25.749508,26.43662,27.125546,27.812658,25.562773,23.312885,21.063,18.813112,16.563227,17.799667,19.03792,20.27436,21.512613,22.750868,23.47424,24.199425,24.92461,25.649796,26.374979,22.150776,17.92476,13.700559,9.474543,5.2503395,4.650249,4.0501585,3.4500678,2.8499773,2.2498865,2.4873846,2.7248828,2.962381,3.199879,3.437377,4.537845,5.638314,6.736969,7.837437,8.937905,7.7123427,6.48678,5.2630305,4.0374675,2.811905,3.3376641,3.8616104,4.3873696,4.9131284,5.4370747,5.049101,4.6629395,4.274966,3.8869917,3.5008307,3.350355,3.199879,3.049403,2.9007401,2.7502642,2.1991236,1.649796,1.1004683,0.5493277,0.0,3.3630457,6.7242785,10.087324,13.45037,16.811602,14.737573,12.661731,10.587702,8.511859,6.43783,6.813113,7.1865835,7.5618668,7.93715,8.312433,8.125698,7.93715,7.750415,7.5618668,7.3751316,6.049856,4.7245803,3.3993049,2.0758421,0.7505665,0.66173136,0.5747091,0.48768693,0.40066472,0.31182957,0.51306844,0.7124943,0.9119202,1.1131591,1.3125849,2.3133402,3.3122826,4.313038,5.3119802,6.3127356,7.0868707,7.8628187,8.636953,9.412902,10.1870365,9.875207,9.563377,9.249735,8.937905,8.624263,9.12464,9.625018,10.125396,10.625773,11.124338,10.613083,10.100015,9.5869465,9.07569,8.562622,10.57501,12.5873995,14.599788,16.612177,18.624565,20.025984,21.425592,22.8252,24.224806,25.624413,26.200935,26.775644,27.350353,27.925062,28.499771,27.524399,26.550837,25.575462,24.60009,23.624716,24.674421,25.724127,26.775644,27.82535,28.875055,27.350353,25.825651,24.299137,22.774435,21.249735,25.46306,29.674572,33.887897,38.099407,42.312733,39.33766,36.36259,33.38752,30.412447,27.437376,25.24913,23.062696,20.87445,18.688019,16.499773,15.350354,14.200936,13.049705,11.900287,10.750868,10.51337,10.275872,10.038374,9.800876,9.563377,9.137331,8.713099,8.287052,7.8628187,7.4367723,8.312433,9.188094,10.061942,10.937603,11.813264,11.312886,10.812509,10.312131,9.811753,9.313189,9.287807,9.262425,9.237044,9.211663,9.188094,9.224354,9.262425,9.300498,9.336758,9.374829,7.5872483,5.7996674,4.0120864,2.2245052,0.43692398,1.1004683,1.7621996,2.4257438,3.0874753,3.7492065,4.12449,4.499773,4.8750563,5.2503395,5.6256227,7.7123427,9.799063,11.887595,13.974316,16.062849,14.124791,12.186734,10.25049,8.312433,6.3743763,7.311678,8.2507925,9.188094,10.125396,11.062697,9.537996,8.013294,6.48678,4.9620786,3.437377,4.3003473,5.163317,6.0244746,6.887445,7.750415,6.249282,4.749962,3.2506418,1.7495089,0.25018883,0.22480737,0.19942589,0.17585737,0.15047589,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07433146,0.15047589,0.22480737,0.2991388,0.37528324,0.51306844,0.6508536,0.7868258,0.9246109,1.062396,3.9504454,6.836682,9.724731,12.612781,15.50083,12.436923,9.374829,6.3127356,3.2506418,0.18673515,0.33721104,0.48768693,0.63816285,0.7868258,0.93730164,2.275268,3.6132345,4.949388,6.2873545,7.6253204,6.2746634,4.9258194,3.5751622,2.2245052,0.87566096,1.3742256,1.8746033,2.374981,2.8753586,3.3757362,2.8753586,2.374981,1.8746033,1.3742256,0.87566096,0.69980353,0.52575916,0.34990177,0.17585737,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.12509441,0.25018883,0.37528324,0.50037766,0.62547207,0.52575916,0.42423326,0.3245203,0.22480737,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.13778515,0.15047589,0.16316663,0.17585737,0.18673515,0.18673515,0.18673515,0.18673515,0.18673515,0.18673515,0.18673515,0.18673515,0.18673515,0.18673515,0.18673515,0.17585737,0.16316663,0.15047589,0.13778515,0.12509441,0.15047589,0.17585737,0.19942589,0.22480737,0.25018883,0.25018883,0.25018883,0.25018883,0.25018883,0.25018883,0.25018883,0.25018883,0.25018883,0.25018883,0.25018883,0.2374981,0.22480737,0.21211663,0.19942589,0.18673515,0.16316663,0.13778515,0.11240368,0.0870222,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,3.6748753,3.6476808,3.6204863,3.5932918,3.5642843,3.53709,3.3648586,3.1926272,3.0203958,2.8481643,2.6741197,2.8626678,3.049403,3.2379513,3.4246864,3.6132345,3.489953,3.3666716,3.245203,3.1219215,3.000453,3.005892,3.009518,3.0149567,3.0203958,3.0258346,3.6676233,4.309412,4.953014,5.5948024,6.2384043,6.6499467,7.063302,7.474845,7.8882003,8.299743,9.712041,11.124338,12.538449,13.9507475,15.363045,13.789393,12.217555,10.645717,9.072064,7.500226,7.8791356,8.259857,8.640579,9.019489,9.400211,8.812811,8.225411,7.6380115,7.0506115,6.4632115,6.202145,5.942891,5.6818247,5.422571,5.163317,5.3953767,5.6274357,5.859495,6.093367,6.3254266,6.2293396,6.1350656,6.0407915,5.9447045,5.8504305,8.232663,10.614896,12.9971285,15.379361,17.763407,15.640429,13.517449,11.39447,9.273304,7.1503243,5.9283876,4.704638,3.482701,2.2607644,1.0370146,0.8430276,0.64722764,0.45324063,0.2574407,0.06164073,0.08520924,0.10696479,0.13053331,0.15228885,0.17585737,4.7300196,9.284182,13.840157,18.394318,22.950293,18.990784,15.02946,11.069949,7.1104393,3.149116,2.561716,1.9743162,1.3869164,0.7995165,0.21211663,0.17041849,0.12690738,0.08520924,0.04169814,0.0,0.13053331,0.25925365,0.38978696,0.52032024,0.6508536,2.2915847,3.9341288,5.576673,7.219217,8.861761,7.663393,6.4632115,5.2630305,4.062849,2.8626678,3.5443418,4.227829,4.9095025,5.5929894,6.2746634,6.530291,6.784106,7.039734,7.2953615,7.549176,7.4258947,7.3008003,7.175706,7.0506115,6.925517,6.755099,6.58468,6.414262,6.245656,6.0752378,6.7623506,7.4494634,8.138389,8.825501,9.512614,9.822631,10.1326475,10.442664,10.752681,11.062697,10.230548,9.398398,8.564435,7.7322855,6.9001355,7.304426,7.71053,8.1148205,8.519112,8.925215,9.893337,10.859646,11.827768,12.79589,13.762199,13.037014,12.311829,11.586644,10.863272,10.138086,10.303066,10.468046,10.633025,10.798005,10.962985,11.9021,12.843027,13.782142,14.723069,15.662184,15.277836,14.891675,14.507326,14.122978,13.736817,13.439491,13.142166,12.84484,12.547514,12.250188,13.539205,14.830034,16.120863,17.40988,18.700708,18.526665,18.354433,18.182201,18.00997,17.837738,18.285542,18.733343,19.17933,19.627132,20.074934,20.564434,21.055748,21.545248,22.034748,22.524246,24.235683,25.945307,27.654932,29.364555,31.074179,31.920832,32.765675,33.61051,34.455353,35.300194,33.16815,31.034294,28.90225,26.770205,24.63816,24.66173,24.68711,24.712494,24.737875,24.763256,23.32195,21.882458,20.442966,19.001661,17.562168,18.651758,19.743162,20.832752,21.922344,23.011934,25.379663,27.747393,30.115122,32.48285,34.85058,29.371807,23.894846,18.417887,12.939114,7.462154,6.5248523,5.5875506,4.650249,3.7129474,2.7756457,2.909805,3.045777,3.1799364,3.3159087,3.4500678,4.5432844,5.634688,6.7279043,7.819308,8.912524,8.013294,7.112252,6.2130227,5.3119802,4.4127507,4.668379,4.9221935,5.177821,5.431636,5.6872635,5.185073,4.6828823,4.1806917,3.6766882,3.1744974,3.149116,3.1255474,3.100166,3.0747845,3.049403,3.4119956,3.774588,4.137181,4.499773,4.8623657,7.066928,9.273304,11.477866,13.682428,15.8869915,13.7875805,11.6881695,9.5869465,7.4875355,5.388125,5.6401267,5.8921285,6.14413,6.397945,6.6499467,6.755099,6.8602505,6.965402,7.0705543,7.175706,5.903006,4.6303062,3.3576066,2.084907,0.8122072,0.8466535,0.88291276,0.91735905,0.95180535,0.9880646,1.0750868,1.162109,1.2491312,1.3379664,1.4249886,2.520018,3.6150475,4.710077,5.805106,6.9001355,7.4277077,7.95528,8.482852,9.010424,9.537996,9.24067,8.943344,8.644206,8.34688,8.049554,8.615198,9.180842,9.744674,10.310318,10.874149,11.452485,12.03082,12.607342,13.185677,13.762199,15.435563,17.107115,18.78048,20.45203,22.125395,22.765371,23.405348,24.045322,24.685299,25.325274,25.807522,26.28977,26.772018,27.254267,27.738327,27.290525,26.842724,26.394922,25.94712,25.49932,25.785767,26.070402,26.355038,26.639671,26.924307,25.80027,24.674421,23.550385,22.424534,21.300497,24.52757,27.754644,30.981718,34.210606,37.437675,34.854206,32.27255,29.689075,27.107416,24.525759,22.500679,20.4756,18.45052,16.425442,14.400362,13.392355,12.384347,11.378153,10.370146,9.362139,9.175404,8.9868555,8.80012,8.613385,8.424837,8.087626,7.750415,7.413204,7.07418,6.736969,7.4277077,8.116633,8.807372,9.498111,10.1870365,9.73017,9.273304,8.814624,8.357758,7.900891,8.227224,8.55537,8.881703,9.20985,9.537996,9.510801,9.481794,9.4546,9.427405,9.400211,7.6851482,5.9700856,4.255023,2.5399606,0.824898,1.5283275,2.229944,2.9333735,3.63499,4.3366065,4.507025,4.6774435,4.847862,5.0182805,5.186886,6.827617,8.4683485,10.107266,11.747997,13.386916,11.813264,10.2378,8.662335,7.0868707,5.5132194,6.3725634,7.231908,8.093065,8.952409,9.811753,8.694968,7.5781837,6.4595857,5.3428006,4.2242026,4.695573,5.1651306,5.634688,6.104245,6.5756154,5.3047285,4.0356545,2.764768,1.4956942,0.22480737,0.20486477,0.18492219,0.16497959,0.14503701,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.059827764,0.11965553,0.1794833,0.23931105,0.2991388,0.40972954,0.52032024,0.629098,0.73968875,0.85027945,3.6458678,6.439643,9.235231,12.03082,14.824595,11.99456,9.164526,6.3344913,3.5044568,0.6744221,1.0605831,1.4449311,1.8292793,2.2154403,2.5997884,3.7546456,4.9095025,6.0643597,7.219217,8.375887,6.978093,5.580299,4.1825047,2.7847104,1.3869164,1.6534219,1.9181144,2.182807,2.4474995,2.712192,2.3097143,1.9072367,1.504759,1.1022812,0.69980353,0.56020546,0.42060733,0.27919623,0.13959812,0.0,0.12690738,0.25562772,0.3825351,0.5094425,0.63816285,0.5094425,0.3825351,0.25562772,0.12690738,0.0,0.17041849,0.34083697,0.5094425,0.67986095,0.85027945,0.7016165,0.55476654,0.40791658,0.25925365,0.11240368,0.10696479,0.10333887,0.09789998,0.092461094,0.0870222,0.09064813,0.092461094,0.09427405,0.09789998,0.099712946,0.09064813,0.07977036,0.07070554,0.059827764,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.059827764,0.058014803,0.054388877,0.052575916,0.05076295,0.052575916,0.054388877,0.058014803,0.059827764,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.10333887,0.07977036,0.058014803,0.034446288,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.12509441,0.13778515,0.15047589,0.16316663,0.17585737,0.17767033,0.1794833,0.18310922,0.18492219,0.18673515,0.18492219,0.18310922,0.1794833,0.17767033,0.17585737,0.16316663,0.15047589,0.13778515,0.12509441,0.11240368,0.13415924,0.15772775,0.1794833,0.2030518,0.22480737,0.22662032,0.23024625,0.23205921,0.23568514,0.2374981,0.23568514,0.23205921,0.23024625,0.22662032,0.22480737,0.2229944,0.21936847,0.21755551,0.21574254,0.21211663,0.18310922,0.15228885,0.12328146,0.092461094,0.06164073,0.059827764,0.058014803,0.054388877,0.052575916,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,3.787279,3.7075086,3.6277382,3.5479677,3.4681973,3.386614,3.254268,3.1219215,2.9895754,2.857229,2.7248828,3.0874753,3.4500678,3.8126602,4.175253,4.537845,4.3166637,4.0972953,3.877927,3.6567454,3.437377,3.484514,3.531651,3.5806012,3.6277382,3.6748753,4.122677,4.5704784,5.0182805,5.464269,5.9120708,6.3127356,6.7115874,7.112252,7.512917,7.911769,9.38752,10.863272,12.337211,13.812962,15.2869005,14.005136,12.7233715,11.439794,10.15803,8.874452,8.885329,8.894395,8.9052725,8.914337,8.925215,8.613385,8.299743,7.987913,7.6742706,7.362441,7.130382,6.8983226,6.6644506,6.432391,6.200332,6.165886,6.1296263,6.09518,6.060734,6.0244746,5.8848767,5.7452784,5.6056805,5.464269,5.3246713,7.902704,10.480737,13.056956,15.63499,18.213022,15.841667,13.472125,11.102583,8.733041,6.3616858,5.2557783,4.1480584,3.0403383,1.9326181,0.824898,0.6726091,0.52032024,0.3680314,0.21574254,0.06164073,0.08339628,0.10333887,0.12328146,0.14322405,0.16316663,4.610364,9.057561,13.504758,17.951956,22.399153,18.642694,14.884423,11.127964,7.369693,3.6132345,2.9750717,2.3369088,1.7005589,1.062396,0.42423326,0.34083697,0.25562772,0.17041849,0.08520924,0.0,0.25925365,0.52032024,0.7795739,1.0406405,1.2998942,2.5091403,3.720199,4.9294453,6.1405044,7.3497505,6.7496595,6.149569,5.5494785,4.949388,4.349297,4.914942,5.480586,6.0444174,6.6100616,7.175706,7.2228427,7.26998,7.317117,7.364254,7.413204,7.224656,7.037921,6.849373,6.6626377,6.4759026,6.58468,6.695271,6.8058615,6.9146395,7.02523,7.5256076,8.024173,8.52455,9.024928,9.525306,10.069194,10.614896,11.160598,11.704487,12.250188,11.334642,10.420909,9.5053625,8.589817,7.6742706,7.7848616,7.895452,8.00423,8.1148205,8.225411,9.14821,10.069194,10.991992,11.91479,12.837588,12.250188,11.662788,11.075388,10.487988,9.900589,10.217857,10.535126,10.852394,11.169662,11.486931,12.442362,13.397794,14.353225,15.306843,16.262274,15.6422415,15.022208,14.402175,13.782142,13.162108,12.968122,12.772322,12.578335,12.382534,12.186734,13.354282,14.521831,15.689378,16.856926,18.024473,18.093367,18.160446,18.227526,18.294605,18.361685,18.75691,19.152136,19.547363,19.942589,20.337814,20.504606,20.673212,20.840004,21.006798,21.175404,22.957544,24.739687,26.52183,28.305784,30.087927,31.103186,32.11663,33.13189,34.147152,35.16241,33.110134,31.057861,29.005589,26.953314,24.89923,24.262878,23.624716,22.988365,22.350203,21.71204,21.082941,20.45203,19.822933,19.192022,18.562923,19.505665,20.446592,21.389332,22.332073,23.274813,27.285088,31.29536,35.305634,39.315907,43.324368,36.59465,29.864933,23.135216,16.405499,9.675781,8.399456,7.124943,5.8504305,4.574105,3.299592,3.3322253,3.3648586,3.397492,3.4301252,3.4627585,4.5469103,5.632875,6.717026,7.802991,8.887142,8.312433,7.7377243,7.1630154,6.588306,6.011784,5.99728,5.9827766,5.9682727,5.9519563,5.9374523,5.319232,4.702825,4.0846047,3.4681973,2.8499773,2.94969,3.049403,3.149116,3.2506418,3.350355,4.6248674,5.89938,7.175706,8.450218,9.724731,10.772624,11.820516,12.868408,13.914488,14.96238,12.837588,10.712796,8.588004,6.4632115,4.3366065,4.4671397,4.597673,4.7282066,4.856927,4.98746,5.384499,5.7833505,6.1803894,6.5774283,6.9744673,5.754343,4.5342193,3.3140955,2.0957847,0.87566096,1.0333886,1.1893034,1.3470312,1.504759,1.6624867,1.6371052,1.6117238,1.5881553,1.5627737,1.5373923,2.7266958,3.917812,5.1071157,6.298232,7.4875355,7.7667317,8.047741,8.326937,8.607946,8.887142,8.604321,8.323311,8.040489,7.757667,7.474845,8.105756,8.734854,9.365765,9.994863,10.625773,12.291886,13.959812,15.627737,17.295664,18.961775,20.294304,21.626831,22.959358,24.291885,25.624413,25.504757,25.385101,25.265446,25.14579,25.024323,25.415922,25.80571,26.195496,26.585283,26.97507,27.05484,27.134611,27.214382,27.294151,27.375734,26.8953,26.414865,25.93443,25.455807,24.975372,24.250187,23.525002,22.799818,22.074633,21.349447,23.592083,25.834717,28.07735,30.319986,32.562622,30.372562,28.182503,25.992445,23.802385,21.612328,19.750414,17.886688,16.024776,14.162864,12.299138,11.434355,10.5695715,9.704789,8.840006,7.9752226,7.837437,7.699652,7.5618668,7.4258947,7.28811,7.037921,6.787732,6.5375433,6.2873545,6.037165,6.542982,7.0469856,7.552802,8.056806,8.562622,8.147454,7.7322855,7.317117,6.9019485,6.48678,7.166641,7.8483152,8.528176,9.208037,9.8878975,9.795437,9.702975,9.610515,9.518054,9.425592,7.783048,6.1405044,4.49796,2.855416,1.2128719,1.9543737,2.6976883,3.43919,4.1825047,4.9258194,4.88956,4.855114,4.8206677,4.784408,4.749962,5.942891,7.135821,8.326937,9.519867,10.712796,9.499924,8.287052,7.07418,5.863121,4.650249,5.431636,6.2148356,6.9980354,7.7794223,8.562622,7.851941,7.1430726,6.432391,5.7217097,5.0128417,5.090799,5.1669436,5.2449007,5.3228583,5.4008155,4.360175,3.3195345,2.280707,1.2400664,0.19942589,0.18492219,0.17041849,0.15410182,0.13959812,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.045324065,0.09064813,0.13415924,0.1794833,0.22480737,0.30820364,0.38978696,0.47318324,0.55476654,0.63816285,3.339477,6.0426044,8.745731,11.447045,14.150173,11.552197,8.954222,6.35806,3.7600844,1.162109,1.7821422,2.4021754,3.0222087,3.6422417,4.262275,5.235836,6.207584,7.179332,8.152893,9.12464,7.6797094,6.2347784,4.7898474,3.3449159,1.8999848,1.9308052,1.9598125,1.9906329,2.0196402,2.0504606,1.745883,1.4394923,1.1349145,0.83033687,0.52575916,0.42060733,0.3154555,0.21030366,0.10515183,0.0,0.25562772,0.5094425,0.7650702,1.020698,1.2745126,1.020698,0.7650702,0.5094425,0.25562772,0.0,0.21574254,0.42967212,0.64541465,0.85934424,1.0750868,0.8792868,0.6852999,0.4894999,0.2955129,0.099712946,0.10333887,0.10515183,0.10696479,0.11059072,0.11240368,0.10515183,0.09789998,0.09064813,0.08339628,0.07433146,0.06707962,0.059827764,0.052575916,0.045324065,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.058014803,0.052575916,0.047137026,0.04169814,0.038072214,0.04169814,0.047137026,0.052575916,0.058014803,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.10515183,0.08520924,0.065266654,0.045324065,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.11240368,0.12509441,0.13778515,0.15047589,0.16316663,0.16679256,0.17223145,0.17767033,0.18310922,0.18673515,0.18310922,0.17767033,0.17223145,0.16679256,0.16316663,0.15047589,0.13778515,0.12509441,0.11240368,0.099712946,0.11965553,0.13959812,0.15954071,0.1794833,0.19942589,0.20486477,0.21030366,0.21574254,0.21936847,0.22480737,0.21936847,0.21574254,0.21030366,0.20486477,0.19942589,0.20667773,0.21574254,0.2229944,0.23024625,0.2374981,0.2030518,0.16679256,0.13234627,0.09789998,0.06164073,0.058014803,0.052575916,0.047137026,0.04169814,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,3.8996825,3.7673361,3.63499,3.5026438,3.3702974,3.2379513,3.1454902,3.053029,2.960568,2.8681068,2.7756457,3.3122826,3.8507326,4.3873696,4.9258194,5.462456,5.145188,4.8279195,4.510651,4.1933823,3.874301,3.9649491,4.0555973,4.1444325,4.2350807,4.325729,4.5777307,4.8297324,5.081734,5.335549,5.5875506,5.975525,6.3616858,6.7496595,7.137634,7.5256076,9.063,10.600392,12.137785,13.675177,15.212569,14.220879,13.227375,12.235684,11.242181,10.25049,9.88971,9.530745,9.169965,8.809185,8.450218,8.412147,8.375887,8.337815,8.299743,8.26167,8.056806,7.851941,7.647076,7.4422116,7.2373466,6.9345818,6.6318173,6.3308654,6.0281005,5.7253356,5.540414,5.3554916,5.1705694,4.985647,4.800725,7.572745,10.344765,13.116784,15.890617,18.662638,16.04472,13.426801,10.810696,8.192778,5.57486,4.5831695,3.589666,2.5979755,1.6044719,0.61278135,0.50219065,0.39159992,0.28282216,0.17223145,0.06164073,0.07977036,0.09789998,0.11421664,0.13234627,0.15047589,4.4907084,8.829127,13.16936,17.509592,21.849825,18.294605,14.739386,11.184166,7.6307597,4.07554,3.386614,2.6995013,2.0123885,1.3252757,0.63816285,0.5094425,0.3825351,0.25562772,0.12690738,0.0,0.38978696,0.7795739,1.1693609,1.5591478,1.9507477,2.7266958,3.5044568,4.2822175,5.0599785,5.8377395,5.8377395,5.8377395,5.8377395,5.8377395,5.8377395,6.285541,6.733343,7.179332,7.6271334,8.074935,7.915395,7.755854,7.5945,7.4349594,7.2754188,7.02523,6.775041,6.5248523,6.2746634,6.0244746,6.414262,6.8058615,7.1956487,7.5854354,7.9752226,8.287052,8.600695,8.912524,9.224354,9.537996,10.31757,11.097144,11.876718,12.658105,13.437678,12.440549,11.443419,10.444477,9.447348,8.450218,8.265296,8.080374,7.895452,7.71053,7.5256076,8.403082,9.280556,10.15803,11.035503,11.912977,11.463363,11.011934,10.56232,10.112705,9.663091,10.1326475,10.602205,11.071762,11.543133,12.012691,12.982625,13.95256,14.922495,15.89243,16.862366,16.006647,15.152741,14.297023,13.443117,12.5873995,12.494938,12.402477,12.310016,12.217555,12.125093,13.16936,14.21544,15.2597065,16.305786,17.350052,17.658255,17.964645,18.27285,18.57924,18.887444,19.230095,19.572744,19.915394,20.258043,20.600695,20.444778,20.290678,20.134762,19.980661,19.824745,21.679407,23.534067,25.390541,27.245201,29.099863,30.28554,31.469404,32.655083,33.84076,35.024624,33.05212,31.079618,29.107115,27.134611,25.162107,23.862213,22.562319,21.262424,19.96253,18.662638,18.84212,19.021603,19.2029,19.382383,19.561867,20.357758,21.151834,21.947725,22.741802,23.537693,29.19051,34.841515,40.49433,46.14715,51.79997,43.817493,35.83502,27.852545,19.87007,11.887595,10.275872,8.662335,7.0506115,5.4370747,3.825351,3.7546456,3.6857529,3.6150475,3.5443418,3.4754493,4.552349,5.6292486,6.7079616,7.7848616,8.861761,8.613385,8.363196,8.113008,7.8628187,7.61263,7.327995,7.0433598,6.7569118,6.472276,6.187641,5.4552045,4.7227674,3.9903307,3.2578938,2.525457,2.7502642,2.9750717,3.199879,3.4246864,3.6494937,5.8377395,8.024173,10.212419,12.400664,14.587097,14.478319,14.367728,14.257137,14.14836,14.037769,11.887595,9.737422,7.5872483,5.4370747,3.2869012,3.294153,3.303218,3.3104696,3.3177216,3.3249733,4.0157123,4.704638,5.3953767,6.0843024,6.775041,5.6074934,4.439945,3.2723975,2.1048496,0.93730164,1.2183108,1.4975071,1.7767034,2.0577126,2.3369088,2.1991236,2.0631514,1.9253663,1.7875811,1.649796,2.9351864,4.220577,5.504154,6.789545,8.074935,8.107569,8.140202,8.172835,8.205468,8.238102,7.9697833,7.703278,7.4349594,7.166641,6.9001355,7.5945,8.290678,8.985043,9.679407,10.375585,13.1331005,15.890617,18.648132,21.40565,24.163166,25.154856,26.146545,27.140049,28.13174,29.125244,28.244144,27.364857,26.48557,25.604471,24.725183,25.022509,25.319836,25.61716,25.914488,26.211813,26.819155,27.42831,28.035654,28.642996,29.250338,28.004833,26.759327,25.515635,24.27013,23.024624,22.700104,22.375584,22.049252,21.724731,21.40021,22.658407,23.91479,25.172985,26.429369,27.687565,25.889105,24.09246,22.295815,20.497355,18.700708,17.00015,15.299591,13.600845,11.900287,10.199727,9.4781685,8.754796,8.033237,7.309865,6.588306,6.4994707,6.412449,6.3254266,6.2384043,6.149569,5.9882154,5.825049,5.661882,5.5005283,5.337362,5.658256,5.977338,6.298232,6.6173134,6.9382076,6.5647373,6.19308,5.81961,5.4479527,5.0744824,6.107871,7.1394467,8.172835,9.2044115,10.2378,10.080072,9.922344,9.764616,9.606889,9.449161,7.8791356,6.3109226,4.7390842,3.1708715,1.6008459,2.382233,3.1654327,3.9468195,4.7300196,5.5132194,5.272095,5.032784,4.7916603,4.552349,4.313038,5.0581656,5.803293,6.548421,7.2917356,8.036863,7.1865835,6.338117,5.487838,4.6375585,3.787279,4.4925213,5.197764,5.903006,6.6082487,7.311678,7.0107265,6.7079616,6.4051967,6.1024323,5.7996674,5.484212,5.1705694,4.855114,4.539658,4.2242026,3.4156215,2.6052272,1.794833,0.98443866,0.17585737,0.16497959,0.15410182,0.14503701,0.13415924,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.20486477,0.25925365,0.3154555,0.36984438,0.42423326,3.0348995,5.6455655,8.254418,10.865085,13.475751,11.109835,8.745731,6.379815,4.0157123,1.649796,2.5055144,3.3594196,4.215138,5.0708566,5.924762,6.7152133,7.5056653,8.294304,9.084756,9.875207,8.383139,6.889258,5.3971896,3.9051213,2.4130533,2.2081885,2.0033236,1.7966459,1.5917811,1.3869164,1.1802386,0.97174793,0.7650702,0.55839247,0.34990177,0.27919623,0.21030366,0.13959812,0.07070554,0.0,0.3825351,0.7650702,1.1476053,1.5301404,1.9126755,1.5301404,1.1476053,0.7650702,0.3825351,0.0,0.25925365,0.52032024,0.7795739,1.0406405,1.2998942,1.0569572,0.81583315,0.5728962,0.32995918,0.0870222,0.09789998,0.10696479,0.11784257,0.12690738,0.13778515,0.11965553,0.10333887,0.08520924,0.06707962,0.05076295,0.045324065,0.03988518,0.034446288,0.030820364,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.054388877,0.047137026,0.03988518,0.032633327,0.025381476,0.032633327,0.03988518,0.047137026,0.054388877,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.10696479,0.09064813,0.072518505,0.054388877,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.018129626,0.034446288,0.052575916,0.07070554,0.0870222,0.099712946,0.11240368,0.12509441,0.13778515,0.15047589,0.15772775,0.16497959,0.17223145,0.1794833,0.18673515,0.1794833,0.17223145,0.16497959,0.15772775,0.15047589,0.13778515,0.12509441,0.11240368,0.099712946,0.0870222,0.10515183,0.12328146,0.13959812,0.15772775,0.17585737,0.18310922,0.19036107,0.19761293,0.20486477,0.21211663,0.20486477,0.19761293,0.19036107,0.18310922,0.17585737,0.19217403,0.21030366,0.22662032,0.24474995,0.26287958,0.2229944,0.18310922,0.14322405,0.10333887,0.06164073,0.054388877,0.047137026,0.03988518,0.032633327,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,4.0120864,3.827164,3.6422417,3.4573197,3.2723975,3.0874753,3.0348995,2.9823234,2.9297476,2.8771715,2.8245957,3.53709,4.249584,4.9620786,5.674573,6.3870673,5.9718986,5.5567303,5.143375,4.7282066,4.313038,4.445384,4.5777307,4.710077,4.842423,4.974769,5.032784,5.090799,5.147001,5.2050157,5.2630305,5.638314,6.011784,6.3870673,6.7623506,7.137634,8.736667,10.337513,11.938358,13.537392,15.138238,14.434808,13.7331915,13.029762,12.328146,11.624716,10.8959055,10.165281,9.434657,8.705847,7.9752226,8.212721,8.450218,8.6877165,8.925215,9.162713,8.985043,8.807372,8.629702,8.452031,8.274362,7.705091,7.135821,6.5647373,5.995467,5.424384,5.1941376,4.9657044,4.7354584,4.505212,4.274966,7.2427855,10.210606,13.178425,16.144432,19.112251,16.24777,13.383289,10.516996,7.652515,4.788034,3.9105604,3.0330863,2.1556125,1.2781386,0.40066472,0.33177215,0.26469254,0.19761293,0.13053331,0.06164073,0.07795739,0.092461094,0.10696479,0.12328146,0.13778515,4.36924,8.602508,12.835775,17.06723,21.300497,17.94833,14.594349,11.242181,7.890013,4.537845,3.7999697,3.0620937,2.324218,1.5881553,0.85027945,0.67986095,0.5094425,0.34083697,0.17041849,0.0,0.52032024,1.0406405,1.5591478,2.079468,2.5997884,2.9442513,3.290527,3.63499,3.9794528,4.325729,4.9258194,5.524097,6.1241875,6.7242785,7.324369,7.654328,7.9842873,8.314246,8.644206,8.974165,8.607946,8.239915,7.8718834,7.5056653,7.137634,6.825804,6.5121617,6.200332,5.8866897,5.57486,6.245656,6.9146395,7.5854354,8.254418,8.925215,9.050309,9.175404,9.300498,9.425592,9.550687,10.564133,11.579392,12.594651,13.60991,14.625169,13.544643,12.465931,11.385405,10.304879,9.224354,8.745731,8.265296,7.7848616,7.304426,6.825804,7.6579537,8.490104,9.322253,10.154404,10.988366,10.674724,10.362894,10.049252,9.737422,9.425592,10.047439,10.669285,11.292944,11.91479,12.536636,13.522888,14.507326,15.491765,16.478018,17.462456,16.372866,15.283275,14.191871,13.102281,12.012691,12.021755,12.032633,12.0416975,12.052575,12.06164,12.984438,13.907236,14.830034,15.752831,16.67563,17.223145,17.770658,18.318174,18.865688,19.413204,19.703278,19.993351,20.281612,20.571686,20.861761,20.38495,19.908142,19.42952,18.952711,18.475903,20.40308,22.33026,24.257439,26.184618,28.111797,29.467894,30.822176,32.178272,33.532555,34.88684,32.99592,31.103186,29.210453,27.31772,25.424988,23.463362,21.499924,19.538298,17.57486,15.613234,16.603111,17.592989,18.582867,19.572744,20.562622,21.209848,21.857077,22.504305,23.153345,23.800573,31.094122,38.389484,45.684845,52.980206,60.275566,51.040337,41.805103,32.569874,23.33464,14.09941,12.1504755,10.199727,8.2507925,6.300045,4.349297,4.177066,4.004834,3.832603,3.6603715,3.48814,4.557788,5.6274357,6.697084,7.7667317,8.838193,8.912524,8.9868555,9.063,9.137331,9.211663,8.656897,8.10213,7.5473633,6.9925966,6.43783,5.5893636,4.74271,3.8942437,3.04759,2.1991236,2.5508385,2.9007401,3.2506418,3.6005437,3.9504454,7.0506115,10.150778,13.250943,16.349297,19.449463,18.182201,16.914942,15.64768,14.380419,13.113158,10.937603,8.762048,6.588306,4.4127507,2.2371957,2.1229792,2.0069497,1.892733,1.7767034,1.6624867,2.6451125,3.6277382,4.610364,5.5929894,6.5756154,5.4606433,4.345671,3.2306993,2.1157274,1.0007553,1.403233,1.8057107,2.2081885,2.610666,3.0131438,2.762955,2.5127661,2.2625773,2.0123885,1.7621996,3.141864,4.5233417,5.903006,7.2826705,8.662335,8.446592,8.232663,8.01692,7.802991,7.5872483,7.3352466,7.083245,6.82943,6.5774283,6.3254266,7.0850577,7.844689,8.604321,9.365765,10.125396,13.972503,17.819609,21.666716,25.515635,29.362741,30.015408,30.668076,31.320742,31.971596,32.62426,30.985344,29.344612,27.705694,26.064962,24.424232,24.630909,24.835773,25.04064,25.245504,25.450369,26.585283,27.720198,28.855112,29.990026,31.12494,29.114367,27.105604,25.095028,23.084452,21.07569,21.15002,21.224354,21.300497,21.374828,21.44916,21.722918,21.994862,22.266806,22.540564,22.812508,21.407463,20.002417,10258.0,17.192324,15.787278,14.249886,12.712494,11.175101,9.637709,8.100317,7.520169,6.9400206,6.359873,5.7797246,5.199577,5.163317,5.125245,5.087173,5.049101,5.0128417,4.936697,4.8623657,4.788034,4.7118897,4.6375585,4.7717175,4.9076896,5.041849,5.177821,5.3119802,4.9820213,4.652062,4.322103,3.9921436,3.6621845,5.047288,6.432391,7.817495,9.202598,10.587702,10.364707,10.141713,9.920531,9.697536,9.474543,7.9770355,6.4795284,4.9820213,3.484514,1.987007,2.810092,3.633177,4.454449,5.277534,6.1006193,5.65463,5.2104545,4.764466,4.3202896,3.874301,4.171627,4.4707656,4.7680917,5.0654173,5.3627434,4.8750563,4.3873696,3.8996825,3.4119956,2.9243085,3.5534067,4.1806917,4.8079767,5.4352617,6.0625467,6.167699,6.2728505,6.378002,6.4831543,6.588306,5.8794374,5.1723824,4.465327,3.7582715,3.049403,2.469255,1.8909199,1.310772,0.7306239,0.15047589,0.14503701,0.13959812,0.13415924,0.13053331,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.10333887,0.13053331,0.15772775,0.18492219,0.21211663,2.7303216,5.2467136,7.764919,10.283124,12.799516,10.667472,8.535428,6.401571,4.269527,2.137483,3.2270734,4.3166637,5.408067,6.497658,7.5872483,8.194591,8.801933,9.409276,10.016619,10.625773,9.084756,7.5455503,6.004532,4.465327,2.9243085,2.4855716,2.0450218,1.6044719,1.1657349,0.72518504,0.61459434,0.5058166,0.39522585,0.28463513,0.17585737,0.13959812,0.10515183,0.07070554,0.034446288,0.0,0.5094425,1.020698,1.5301404,2.039583,2.5508385,2.039583,1.5301404,1.020698,0.5094425,0.0,0.3045777,0.6091554,0.9155461,1.2201238,1.5247015,1.2346275,0.9445535,0.6544795,0.36440548,0.07433146,0.092461094,0.11059072,0.12690738,0.14503701,0.16316663,0.13415924,0.10696479,0.07977036,0.052575916,0.025381476,0.02175555,0.01994259,0.018129626,0.014503701,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.052575916,0.04169814,0.032633327,0.02175555,0.012690738,0.02175555,0.032633327,0.04169814,0.052575916,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.11059072,0.09427405,0.07977036,0.065266654,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.13778515,0.14684997,0.15772775,0.16679256,0.17767033,0.18673515,0.17767033,0.16679256,0.15772775,0.14684997,0.13778515,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.09064813,0.10515183,0.11965553,0.13415924,0.15047589,0.15954071,0.17041849,0.1794833,0.19036107,0.19942589,0.19036107,0.1794833,0.17041849,0.15954071,0.15047589,0.17767033,0.20486477,0.23205921,0.25925365,0.28826106,0.24293698,0.19761293,0.15228885,0.10696479,0.06164073,0.052575916,0.04169814,0.032633327,0.02175555,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,4.12449,3.8869917,3.6494937,3.4119956,3.1744974,2.9369993,2.9243085,2.911618,2.9007401,2.8880494,2.8753586,3.7618973,4.650249,5.5367875,6.4251394,7.311678,6.8004227,6.2873545,5.774286,5.2630305,4.749962,4.9258194,5.0998635,5.275721,5.4497657,5.6256227,5.487838,5.3500524,5.2122674,5.0744824,4.936697,5.2992897,5.661882,6.0244746,6.3870673,6.7496595,8.412147,10.074633,11.73712,13.399607,15.062093,14.650551,14.237195,13.825653,13.412297,13.000754,11.900287,10.799818,9.699349,8.600695,7.500226,8.013294,8.52455,9.037619,9.550687,10.061942,9.91328,9.762803,9.612328,9.461852,9.313189,8.4756,7.6380115,6.8004227,5.962834,5.125245,4.8496747,4.574105,4.3003473,4.024777,3.7492065,6.9128265,10.074633,13.238253,16.400059,19.561867,16.450823,13.337966,10.225109,7.112252,3.9993954,3.2379513,2.474694,1.7132497,0.9499924,0.18673515,0.16316663,0.13778515,0.11240368,0.0870222,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,4.249584,8.374074,12.500377,16.624866,20.749357,17.60024,14.449312,11.300196,8.149267,5.0001507,4.213325,3.4246864,2.6378605,1.8492218,1.062396,0.85027945,0.63816285,0.42423326,0.21211663,0.0,0.6508536,1.2998942,1.9507477,2.5997884,3.2506418,3.1618068,3.0747845,2.9877625,2.9007401,2.811905,4.0120864,5.2122674,6.412449,7.61263,8.812811,9.024928,9.237044,9.449161,9.663091,9.875207,9.300498,8.725789,8.149267,7.574558,6.9998484,6.624565,6.249282,5.8758116,5.5005283,5.125245,6.0752378,7.02523,7.9752226,8.925215,9.875207,9.811753,9.750113,9.686659,9.625018,9.563377,10.812509,12.06164,13.312584,14.561715,15.812659,14.650551,13.488441,12.32452,11.162411,10.000301,9.224354,8.450218,7.6742706,6.9001355,6.1241875,6.9128265,7.699652,8.488291,9.275117,10.061942,9.8878975,9.712041,9.537996,9.362139,9.188094,9.96223,10.738177,11.512312,12.28826,13.062395,14.06315,15.062093,16.062849,17.06179,18.062546,16.73727,15.411995,14.0867195,12.763257,11.437981,11.5503845,11.662788,11.775192,11.887595,11.999999,12.799516,13.600845,14.400362,15.199879,15.999394,16.788034,17.57486,18.361685,19.150324,19.93715,20.174648,20.412146,20.649643,20.887142,21.12464,20.325123,19.525606,18.724277,17.92476,17.125244,19.124943,21.12464,23.124338,25.125849,27.125546,28.650248,30.17495,31.69965,33.224354,34.750866,32.937904,31.12494,29.31198,27.50083,25.687866,23.062696,20.437527,17.812357,15.187187,12.562017,14.362289,16.162561,17.962833,19.763105,21.563377,22.061941,22.562319,23.062696,23.563074,24.06164,32.999546,41.93745,50.875355,59.813263,68.74935,58.26318,47.77519,37.2872,26.799213,16.313038,14.025079,11.73712,9.449161,7.1630154,4.8750563,4.599486,4.325729,4.0501585,3.774588,3.5008307,4.5632267,5.6256227,6.688019,7.750415,8.812811,9.211663,9.612328,10.012992,10.411844,10.812509,9.987611,9.162713,8.337815,7.512917,6.688019,5.7253356,4.762653,3.7999697,2.8372865,1.8746033,2.3495996,2.8245957,3.299592,3.774588,4.249584,8.26167,12.27557,16.287657,20.299742,24.311829,21.887897,19.462152,17.038223,14.612478,12.186734,9.987611,7.7866745,5.5875506,3.386614,1.1874905,0.9499924,0.7124943,0.4749962,0.2374981,0.0,1.2745126,2.5508385,3.825351,5.0998635,6.3743763,5.3119802,4.249584,3.1871881,2.124792,1.062396,1.5881553,2.1121013,2.6378605,3.1618068,3.6875658,3.3249733,2.962381,2.5997884,2.2371957,1.8746033,3.350355,4.8242936,6.300045,7.7757964,9.249735,8.78743,8.325124,7.8628187,7.400513,6.9382076,6.70071,6.4632115,6.2257137,5.9882154,5.750717,6.5756154,7.400513,8.225411,9.050309,9.875207,14.811904,19.750414,24.68711,29.625622,34.562317,34.87415,35.18779,35.49962,35.813263,36.12509,33.72473,31.324368,28.925817,26.525455,24.125093,24.237497,24.349901,24.462305,24.574707,24.68711,26.349598,28.012085,29.674572,31.337059,32.999546,30.225712,27.450066,24.674421,21.900587,19.124943,19.59994,20.074934,20.54993,21.024927,21.499924,20.78743,20.074934,19.36244,18.649946,17.937452,16.92582,15.912373,14.90074,13.887294,12.87566,11.499621,10.125396,8.749357,7.3751316,6.000906,5.562169,5.125245,4.688321,4.249584,3.8126602,3.825351,3.8380418,3.8507326,3.8616104,3.874301,3.8869917,3.8996825,3.9123733,3.925064,3.9377546,3.8869917,3.8380418,3.787279,3.738329,3.6875658,3.3993049,3.1128569,2.8245957,2.5381477,2.2498865,3.9867048,5.7253356,7.462154,9.200785,10.937603,10.649343,10.362894,10.074633,9.788185,9.499924,8.074935,6.6499467,5.224958,3.7999697,2.374981,3.2379513,4.099108,4.9620786,5.825049,6.688019,6.037165,5.388125,4.7372713,4.0882306,3.437377,3.2869012,3.1382382,2.9877625,2.8372865,2.6868105,2.561716,2.4366217,2.3133402,2.1882458,2.0631514,2.612479,3.1618068,3.7129474,4.262275,4.8116026,5.3246713,5.8377395,6.350808,6.8620634,7.3751316,6.2746634,5.1741953,4.07554,2.9750717,1.8746033,1.5247015,1.1747998,0.824898,0.4749962,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.4257438,4.8496747,7.2754188,9.699349,12.125093,10.225109,8.325124,6.4251394,4.5251546,2.6251698,3.9504454,5.275721,6.599184,7.9244595,9.249735,9.675781,10.100015,10.524248,10.950294,11.374527,9.788185,8.200029,6.6118746,5.0255322,3.437377,2.762955,2.08672,1.4122978,0.73787576,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.63816285,1.2745126,1.9126755,2.5508385,3.1871881,2.5508385,1.9126755,1.2745126,0.63816285,0.0,0.34990177,0.69980353,1.0497054,1.3996071,1.7495089,1.4122978,1.0750868,0.73787576,0.40066472,0.06164073,0.0870222,0.11240368,0.13778515,0.16316663,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.13778515,0.15047589,0.16316663,0.17585737,0.18673515,0.17585737,0.16316663,0.15047589,0.13778515,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.13778515,0.15047589,0.16316663,0.17585737,0.18673515,0.17585737,0.16316663,0.15047589,0.13778515,0.12509441,0.16316663,0.19942589,0.2374981,0.2755703,0.31182957,0.26287958,0.21211663,0.16316663,0.11240368,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,3.8616104,3.673062,3.482701,3.29234,3.101979,2.911618,3.005892,3.0983531,3.1908143,3.2832751,3.3757362,4.0320287,4.690134,5.3482394,6.004532,6.6626377,6.4269524,6.19308,5.957395,5.7217097,5.487838,5.6274357,5.767034,5.906632,6.0480433,6.187641,6.0480433,5.906632,5.767034,5.6274357,5.487838,5.7017674,5.91751,6.1332526,6.347182,6.5629244,7.8755093,9.188094,10.500679,11.813264,13.125849,12.754191,12.384347,12.0145035,11.644659,11.274815,10.573197,9.869768,9.168152,8.464723,7.763106,8.189152,8.617011,9.04487,9.47273,9.900589,9.770056,9.639522,9.510801,9.380268,9.249735,8.384952,7.520169,6.6553855,5.7906027,4.9258194,4.947575,4.9693303,4.992899,5.0146546,5.038223,7.4966,9.956791,12.416981,14.877171,17.33736,14.50914,11.682731,8.854509,6.0281005,3.199879,2.5907235,1.9797552,1.3705997,0.75963134,0.15047589,0.13053331,0.11059072,0.09064813,0.07070554,0.05076295,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,3.8054085,7.4966,11.189605,14.882609,18.575615,15.720199,12.864782,10.009366,7.155763,4.3003473,3.6096084,2.9206827,2.229944,1.5392052,0.85027945,0.67986095,0.5094425,0.34083697,0.17041849,0.0,0.55839247,1.114972,1.6733645,2.229944,2.7883365,2.7103791,2.6324217,2.5544643,2.47832,2.4003625,3.5026438,4.604925,5.7072062,6.8094873,7.911769,8.13295,8.352319,8.571687,8.792869,9.012237,8.716724,8.423024,8.127511,7.8319983,7.5382986,7.271793,7.0071006,6.742408,6.4777155,6.2130227,6.9073873,7.6017523,8.29793,8.992294,9.686659,9.579695,9.47273,9.365765,9.256987,9.1500225,10.179785,11.209548,12.23931,13.270886,14.300649,13.417736,12.534823,11.651911,10.770811,9.8878975,9.460039,9.03218,8.604321,8.178274,7.750415,8.23085,8.709473,9.189907,9.670342,10.150778,10.027496,9.904215,9.782746,9.659465,9.537996,10.130835,10.721861,11.314699,11.907538,12.500377,13.524701,14.5508375,15.575162,16.599485,17.625622,16.557787,15.489952,14.422117,13.354282,12.28826,12.295512,12.302764,12.310016,12.317267,12.32452,12.975373,13.6244135,14.275268,14.924308,15.575162,16.327541,17.07992,17.8323,18.584679,19.337059,19.755854,20.172834,20.589815,21.006798,21.425592,20.992294,20.560808,20.12751,19.694212,19.262728,20.945156,22.627586,24.310015,25.992445,27.674873,28.94576,30.214834,31.485722,32.754795,34.02568,32.419395,30.814924,29.210453,27.604168,25.999697,25.185677,24.369843,23.555822,22.73999,21.924156,23.011934,24.099712,25.187489,26.275267,27.363045,27.937754,28.512463,29.087172,29.66188,30.238403,37.37966,44.522736,51.665806,58.807068,65.95014,57.012234,48.07614,39.136425,30.20033,21.262424,18.417887,15.573349,12.726997,9.882459,7.037921,6.432391,5.826862,5.223145,4.6176157,4.0120864,4.936697,5.863121,6.787732,7.7123427,8.636953,8.870826,9.102885,9.334945,9.567003,9.800876,9.055748,8.31062,7.5654926,6.8203654,6.0752378,5.411693,4.749962,4.0882306,3.4246864,2.762955,2.8898623,3.0167696,3.1454902,3.2723975,3.3993049,6.8946967,10.390089,13.885481,17.380873,20.87445,18.677141,16.47983,14.282519,12.085209,9.8878975,8.397643,6.9073873,5.4171324,3.926877,2.4366217,2.1574254,1.8782293,1.5972201,1.3180238,1.0370146,1.9453088,2.8517902,3.7600844,4.668379,5.57486,5.3391747,5.105303,4.8696175,4.6357455,4.40006,4.461701,4.5251546,4.5867953,4.650249,4.7118897,4.2876563,3.8616104,3.437377,3.0131438,2.5870976,3.8525455,5.1179934,6.3834414,7.647076,8.912524,8.3595705,7.806617,7.2554765,6.7025228,6.149569,6.0244746,5.89938,5.774286,5.6491914,5.524097,6.5592985,7.5945,8.629702,9.664904,10.700105,14.884423,19.070553,23.254871,27.439188,31.625319,31.85194,32.08037,32.30699,32.535427,32.762047,30.688017,28.612175,26.538147,24.462305,22.388275,22.582262,22.778063,22.97205,23.167849,23.361835,24.89923,26.43662,27.975826,29.513218,31.05061,28.284029,25.51926,22.754494,19.989725,17.224958,17.687263,18.149569,18.611874,19.074179,19.538298,18.840307,18.142317,17.444326,16.748148,16.050158,15.062093,14.075842,13.087777,12.099712,11.111648,9.851639,8.59163,7.3316207,6.071612,4.8116026,4.478018,4.1426196,3.8072214,3.4718235,3.1382382,3.2053177,3.2723975,3.339477,3.4083695,3.4754493,3.4319382,3.39024,3.346729,3.3050308,3.2633326,3.2125697,3.1618068,3.1128569,3.0620937,3.0131438,2.7792716,2.5472124,2.3151531,2.0830941,1.8492218,3.5080826,5.1651306,6.8221784,8.479226,10.138086,9.719293,9.302311,8.885329,8.4683485,8.049554,7.0306687,6.009971,4.989273,3.9703882,2.94969,3.5171473,4.0846047,4.652062,5.219519,5.7869763,5.23221,4.6774435,4.122677,3.5679104,3.0131438,3.0348995,3.056655,3.0802233,3.101979,3.1255474,2.8517902,2.5798457,2.3079014,2.034144,1.7621996,2.1882458,2.612479,3.0367124,3.4627585,3.8869917,4.3891826,4.893186,5.3953767,5.8975673,6.399758,5.462456,4.5251546,3.587853,2.6505513,1.7132497,1.3923552,1.0732739,0.7523795,0.43329805,0.11240368,0.11059072,0.10696479,0.10515183,0.10333887,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,2.1048496,4.022964,5.9392653,7.85738,9.775495,8.352319,6.929143,5.5077806,4.0846047,2.663242,4.0574102,5.4515786,6.8475595,8.241728,9.637709,10.435412,11.233116,12.03082,12.826711,13.6244135,11.631968,9.639522,7.647076,5.65463,3.6621845,3.2325122,2.8028402,2.373168,1.9416829,1.5120108,1.209246,0.90829426,0.6055295,0.30276474,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.6091554,1.1457924,1.6806163,2.2154403,2.7502642,2.1991236,1.649796,1.1004683,0.5493277,0.0,0.47318324,0.9445535,1.4177368,1.889107,2.3622901,1.9072367,1.452183,0.99712944,0.5420758,0.0870222,0.11059072,0.13234627,0.15410182,0.17767033,0.19942589,0.15954071,0.11965553,0.07977036,0.03988518,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.059827764,0.07070554,0.07977036,0.09064813,0.099712946,0.09064813,0.07977036,0.07070554,0.059827764,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.059827764,0.07070554,0.07977036,0.09064813,0.099712946,0.11240368,0.12509441,0.13778515,0.15047589,0.16316663,0.15410182,0.14684997,0.13959812,0.13234627,0.12509441,0.11421664,0.10515183,0.09427405,0.08520924,0.07433146,0.08339628,0.09064813,0.09789998,0.10515183,0.11240368,0.12328146,0.13234627,0.14322405,0.15228885,0.16316663,0.15410182,0.14684997,0.13959812,0.13234627,0.12509441,0.16679256,0.21030366,0.2520018,0.2955129,0.33721104,0.29732585,0.2574407,0.21755551,0.17767033,0.13778515,0.11784257,0.09789998,0.07795739,0.058014803,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,3.6005437,3.4573197,3.3159087,3.1726844,3.0294604,2.8880494,3.0856624,3.2832751,3.4808881,3.6766882,3.874301,4.3021603,4.7300196,5.1578784,5.5857377,6.011784,6.055295,6.096993,6.1405044,6.1822023,6.2257137,6.3308654,6.434204,6.539356,6.644508,6.7496595,6.6082487,6.4650245,6.3218007,6.1803894,6.037165,6.104245,6.1731377,6.240217,6.3072968,6.3743763,7.3370595,8.299743,9.262425,10.225109,11.187792,10.859646,10.533313,10.205167,9.87702,9.550687,9.244296,8.939718,8.63514,8.330563,8.024173,8.366822,8.709473,9.052122,9.394773,9.737422,9.626831,9.518054,9.407463,9.296872,9.188094,8.294304,7.402326,6.510349,5.618371,4.7245803,5.045475,5.3645563,5.6854506,6.004532,6.3254266,8.082188,9.840761,11.597522,13.354282,15.112856,12.569269,10.027496,7.4857225,4.942136,2.4003625,1.9416829,1.4848163,1.0279498,0.56927025,0.11240368,0.09789998,0.08339628,0.06707962,0.052575916,0.038072214,0.05076295,0.06164073,0.07433146,0.0870222,0.099712946,3.3594196,6.6191263,9.880646,13.140353,16.400059,13.840157,11.280253,8.72035,6.1604466,3.6005437,3.007705,2.4148662,1.8220274,1.2291887,0.63816285,0.5094425,0.3825351,0.25562772,0.12690738,0.0,0.46411842,0.9300498,1.3941683,1.8600996,2.324218,2.2571385,2.1900587,2.1229792,2.0558996,1.987007,2.9932013,3.9975824,5.0019636,6.008158,7.0125394,7.2391596,7.4675927,7.6942134,7.9226465,8.149267,8.134763,8.120259,8.105756,8.089439,8.074935,7.9208336,7.764919,7.610817,7.454902,7.3008003,7.7395372,8.180087,8.620637,9.059374,9.499924,9.347635,9.195346,9.043057,8.890768,8.736667,9.547061,10.357455,11.16785,11.978244,12.786825,12.184921,11.583018,10.979301,10.377398,9.775495,9.695724,9.6141405,9.53437,9.4546,9.374829,9.547061,9.719293,9.893337,10.065568,10.2378,10.167094,10.098202,10.027496,9.956791,9.8878975,10.297627,10.707357,11.117086,11.526816,11.938358,12.988064,14.037769,15.087475,16.13718,17.186886,16.378304,15.567909,14.757515,13.947122,13.136727,13.04064,12.9427395,12.84484,12.74694,12.650853,13.149418,13.649796,14.150173,14.650551,15.149116,15.867048,16.584982,17.302916,18.020847,18.736969,19.335245,19.931711,20.529987,21.128265,21.724731,21.659464,21.594198,21.530745,21.465477,21.40021,22.765371,24.130531,25.495693,26.860853,28.224201,29.23946,30.254719,31.26998,32.285236,33.300495,31.902702,30.504908,29.107115,27.70932,26.31334,27.306843,28.302158,29.297476,30.292791,31.288109,31.663391,32.03686,32.412144,32.78743,33.162712,33.811752,34.462605,35.11346,35.7625,36.413353,41.75978,47.10802,52.454445,57.802685,63.149113,55.763103,48.375282,40.987457,33.599636,26.211813,22.810696,19.407764,16.004833,12.601903,9.200785,8.265296,7.3298078,6.394319,5.4606433,4.5251546,5.3119802,6.1006193,6.887445,7.6742706,8.46291,8.528176,8.59163,8.656897,8.722163,8.78743,8.122072,7.456715,6.793171,6.1278133,5.462456,5.0998635,4.7372713,4.3746786,4.0120864,3.6494937,3.4301252,3.2107568,2.9895754,2.770207,2.5508385,5.527723,8.504607,11.483305,14.46019,17.437075,15.468197,13.497506,11.526816,9.557939,7.5872483,6.8076744,6.0281005,5.2467136,4.4671397,3.6875658,3.3648586,3.0421512,2.7194438,2.3967366,2.0758421,2.6142921,3.1545548,3.6948178,4.2350807,4.7753434,5.368182,5.959208,6.552047,7.1448855,7.7377243,7.3370595,6.9382076,6.5375433,6.1368785,5.7380266,5.2503395,4.762653,4.274966,3.787279,3.299592,4.3547363,5.40988,6.4650245,7.520169,8.575313,7.931711,7.2899227,6.6481338,6.004532,5.3627434,5.3500524,5.337362,5.3246713,5.3119802,5.2992897,6.544795,7.7903004,9.035806,10.279498,11.525003,14.956942,18.390692,21.82263,25.254568,28.68832,28.829731,28.972956,29.114367,29.25759,29.400814,27.649492,25.899984,24.150475,22.399153,20.649643,20.927027,21.20441,21.481794,21.759176,22.038374,23.45067,24.862968,26.275267,27.687565,29.099863,26.34416,23.59027,20.834566,18.080675,15.324973,15.774588,16.224201,16.67563,17.125244,17.57486,16.893185,16.209698,15.528025,14.844538,14.162864,13.200181,12.237497,11.274815,10.312131,9.349448,8.205468,7.059676,5.915697,4.7699046,3.6241121,3.392053,3.159994,2.9279346,2.6958754,2.4620032,2.5852847,2.7067533,2.8300345,2.953316,3.0747845,2.9768846,2.8807976,2.7828975,2.6849976,2.5870976,2.5381477,2.4873846,2.4366217,2.3876717,2.3369088,2.1592383,1.983381,1.8057107,1.6280404,1.4503701,3.0276475,4.604925,6.1822023,7.75948,9.336758,8.789243,8.241728,7.6942134,7.1466985,6.599184,5.9845896,5.369995,4.7554007,4.1408067,3.5243993,3.7981565,4.070101,4.3420453,4.615803,4.8877473,4.4272547,3.966762,3.5080826,3.04759,2.5870976,2.7828975,2.9768846,3.1726844,3.3666716,3.5624714,3.141864,2.72307,2.3024626,1.8818551,1.4630609,1.7621996,2.0631514,2.3622901,2.663242,2.962381,3.4555066,3.9468195,4.439945,4.933071,5.424384,4.650249,3.874301,3.100166,2.324218,1.550083,1.260009,0.969935,0.67986095,0.38978696,0.099712946,0.09427405,0.09064813,0.08520924,0.07977036,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07433146,0.15047589,0.22480737,0.2991388,0.37528324,1.7857682,3.1944401,4.604925,6.01541,7.424082,6.4795284,5.5349746,4.590421,3.6458678,2.6995013,4.164375,5.6292486,7.0959353,8.560809,10.025683,11.195044,12.364405,13.535579,14.70494,15.8743,13.477564,11.080828,8.682278,6.285541,3.8869917,3.7020695,3.5171473,3.3322253,3.147303,2.962381,2.3695421,1.7767034,1.1856775,0.59283876,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.581961,1.015259,1.4467441,1.8800422,2.3133402,1.8492218,1.3869164,0.9246109,0.46230546,0.0,0.5946517,1.1893034,1.7857682,2.38042,2.9750717,2.4021754,1.8292793,1.258196,0.6852999,0.11240368,0.13234627,0.15228885,0.17223145,0.19217403,0.21211663,0.17041849,0.12690738,0.08520924,0.04169814,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.045324065,0.052575916,0.059827764,0.06707962,0.07433146,0.06707962,0.059827764,0.052575916,0.045324065,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.045324065,0.052575916,0.059827764,0.06707962,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.13778515,0.13415924,0.13234627,0.13053331,0.12690738,0.12509441,0.11784257,0.11059072,0.10333887,0.09427405,0.0870222,0.09064813,0.092461094,0.09427405,0.09789998,0.099712946,0.10696479,0.11421664,0.12328146,0.13053331,0.13778515,0.13415924,0.13234627,0.13053331,0.12690738,0.12509441,0.17223145,0.21936847,0.26831847,0.3154555,0.36259252,0.33177215,0.30276474,0.27194437,0.24293698,0.21211663,0.18492219,0.15772775,0.13053331,0.10333887,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,3.3376641,3.24339,3.147303,3.053029,2.956942,2.8626678,3.1654327,3.4681973,3.7691493,4.071914,4.3746786,4.572292,4.7699046,4.9675174,5.1651306,5.3627434,5.6818247,6.002719,6.3218007,6.642695,6.9617763,7.0324817,7.1031876,7.17208,7.2427855,7.311678,7.166641,7.021604,6.87838,6.733343,6.588306,6.506723,6.4269524,6.347182,6.2674117,6.187641,6.8004227,7.413204,8.024173,8.636953,9.249735,8.9651,8.680465,8.39583,8.109382,7.8247466,7.9172077,8.009668,8.10213,8.194591,8.287052,8.544493,8.801933,9.059374,9.316814,9.574255,9.48542,9.394773,9.304124,9.215289,9.12464,8.205468,7.2844834,6.3653116,5.4443264,4.5251546,5.143375,5.7597823,6.378002,6.9944096,7.61263,8.667774,9.7229185,10.778063,11.833207,12.888351,10.629399,8.372261,6.115123,3.8579843,1.6008459,1.2944553,0.9898776,0.6852999,0.38072214,0.07433146,0.065266654,0.054388877,0.045324065,0.034446288,0.025381476,0.038072214,0.05076295,0.06164073,0.07433146,0.0870222,2.9152439,5.7416525,8.569874,11.398096,14.224504,11.9601145,9.695724,7.4295206,5.1651306,2.9007401,2.4058013,1.9108626,1.4141108,0.91917205,0.42423326,0.34083697,0.25562772,0.17041849,0.08520924,0.0,0.37165734,0.7451276,1.1167849,1.4902552,1.8619126,1.8057107,1.7476959,1.6896812,1.6316663,1.5754645,2.4819458,3.39024,4.2967215,5.2050157,6.11331,6.347182,6.582867,6.816739,7.0524244,7.28811,7.552802,7.817495,8.082188,8.34688,8.613385,8.568061,8.5227375,8.477413,8.432089,8.386765,8.571687,8.756609,8.943344,9.128266,9.313189,9.115576,8.917963,8.72035,8.5227375,8.325124,8.914337,9.5053625,10.094576,10.685601,11.274815,10.952107,10.629399,10.306692,9.985798,9.663091,9.929596,10.197914,10.46442,10.7327385,10.999244,10.865085,10.729113,10.594954,10.460794,10.324821,10.306692,10.290376,10.272246,10.254116,10.2378,10.46442,10.692853,10.919474,11.147907,11.374527,12.449615,13.524701,14.599788,15.674874,16.749962,16.197008,15.645867,15.092914,14.53996,13.987006,13.785768,13.582716,13.379663,13.176612,12.975373,13.325275,13.675177,14.025079,14.37498,14.724882,15.408369,16.090042,16.771717,17.455204,18.136877,18.914639,19.6924,20.470161,21.247921,22.025682,22.326633,22.629398,22.932163,23.234928,23.537693,24.585585,25.631664,26.679558,27.72745,28.775343,29.534973,30.294605,31.054235,31.81568,32.575314,31.384195,30.194891,29.005589,27.814472,26.625168,29.429821,32.234474,35.04094,37.845592,40.650246,40.313038,39.975826,39.636803,39.29959,38.96238,39.687565,40.41275,41.137936,41.863117,42.588303,46.139896,49.69149,53.2449,56.798306,60.3499,54.512157,48.67442,42.83668,37.00075,31.163013,27.20169,23.24218,19.282671,15.32316,11.361836,10.098202,8.832754,7.567306,6.301858,5.038223,5.6872635,6.338117,6.987158,7.6380115,8.287052,8.185526,8.082188,7.9806614,7.877322,7.7757964,7.1902094,6.604623,6.0208488,5.4352617,4.8496747,4.788034,4.7245803,4.6629395,4.599486,4.537845,3.9703882,3.4029307,2.8354735,2.268016,1.7005589,4.160749,6.6191263,9.079316,11.539507,13.999697,12.25744,10.515183,8.772926,7.0306687,5.2884116,5.217706,5.147001,5.0781083,5.0074024,4.936697,4.572292,4.207886,3.8416677,3.4772623,3.1128569,3.2850883,3.4573197,3.6295512,3.8017826,3.975827,5.3953767,6.814926,8.234476,9.655839,11.075388,10.212419,9.349448,8.488291,7.6253204,6.7623506,6.2130227,5.661882,5.1125546,4.5632267,4.0120864,4.856927,5.7017674,6.548421,7.3932614,8.238102,7.5056653,6.773228,6.0407915,5.3083544,4.574105,4.6756306,4.7753434,4.8750563,4.974769,5.0744824,6.530291,7.9842873,9.440096,10.8959055,12.349901,15.02946,17.709019,20.39039,23.069948,25.749508,25.807522,25.865538,25.92174,25.979753,26.03777,24.61278,23.187792,21.762802,20.337814,18.912827,19.271791,19.632572,19.993351,20.352318,20.713097,22.000301,23.287504,24.574707,25.861912,27.149115,24.40429,21.659464,18.914639,16.169813,13.424988,13.861912,14.300649,14.737573,15.174497,15.613234,14.94425,14.277081,13.60991,12.9427395,12.27557,11.338268,10.399154,9.461852,8.52455,7.5872483,6.5574856,5.527723,4.49796,3.4681973,2.4366217,2.3079014,2.1773682,2.0468347,1.9181144,1.7875811,1.9652514,2.1429217,2.3205922,2.4982624,2.6741197,2.521831,2.3695421,2.2172532,2.0649643,1.9126755,1.8619126,1.8129625,1.7621996,1.7132497,1.6624867,1.5392052,1.4177368,1.2944553,1.1729867,1.0497054,2.5472124,4.0447197,5.542227,7.039734,8.537241,7.859193,7.1829576,6.5049095,5.826862,5.1506267,4.940323,4.7300196,4.519716,4.309412,4.099108,4.077353,4.0555973,4.0320287,4.0102735,3.9867048,3.6222992,3.2578938,2.8916752,2.5272698,2.1628644,2.5308957,2.8971143,3.2651455,3.633177,3.9993954,3.4319382,2.864481,2.2970235,1.7295663,1.162109,1.3379664,1.5120108,1.6878681,1.8619126,2.03777,2.520018,3.002266,3.484514,3.966762,4.4508233,3.8380418,3.2252605,2.612479,1.9996977,1.3869164,1.1276628,0.8684091,0.6073425,0.3480888,0.0870222,0.07977036,0.072518505,0.065266654,0.058014803,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.11240368,0.22480737,0.33721104,0.44961473,0.5620184,1.4648738,2.3677292,3.2705846,4.171627,5.0744824,4.606738,4.1408067,3.673062,3.2053177,2.7375734,4.273153,5.806919,7.3424983,8.8780775,10.411844,11.954676,13.497506,15.040338,16.583168,18.124187,15.32316,12.52032,9.71748,6.9146395,4.1117992,4.171627,4.233268,4.2930956,4.3529234,4.4127507,3.529838,2.6469254,1.7658255,0.88291276,0.0,0.045324065,0.09064813,0.13415924,0.1794833,0.22480737,0.55476654,0.88472575,1.214685,1.5446441,1.8746033,1.49932,1.1258497,0.7505665,0.37528324,0.0,0.7179332,1.4358664,2.1519866,2.8699198,3.587853,2.8971143,2.2081885,1.5174497,0.82671094,0.13778515,0.15410182,0.17223145,0.19036107,0.20667773,0.22480737,0.1794833,0.13415924,0.09064813,0.045324065,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.030820364,0.034446288,0.03988518,0.045324065,0.05076295,0.045324065,0.03988518,0.034446288,0.030820364,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.030820364,0.034446288,0.03988518,0.045324065,0.05076295,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.11421664,0.11784257,0.11965553,0.12328146,0.12509441,0.11965553,0.11421664,0.11059072,0.10515183,0.099712946,0.09789998,0.09427405,0.092461094,0.09064813,0.0870222,0.092461094,0.09789998,0.10333887,0.10696479,0.11240368,0.11421664,0.11784257,0.11965553,0.12328146,0.12509441,0.17767033,0.23024625,0.28282216,0.33539808,0.387974,0.3680314,0.3480888,0.32814622,0.30820364,0.28826106,0.2520018,0.21755551,0.18310922,0.14684997,0.11240368,0.09064813,0.06707962,0.045324065,0.02175555,0.0,0.0,0.0,0.0,0.0,0.0,3.0747845,3.0276475,2.9805105,2.9333735,2.8844235,2.8372865,3.245203,3.6531196,4.059223,4.4671397,4.8750563,4.842423,4.8097897,4.7771564,4.744523,4.7118897,5.3101673,5.906632,6.5049095,7.1031876,7.699652,7.7340984,7.7703576,7.804804,7.83925,7.8755093,7.7268467,7.5799966,7.4331465,7.2844834,7.137634,6.9092,6.68258,6.454147,6.2275267,6.000906,6.261973,6.5248523,6.787732,7.0506115,7.311678,7.0705543,6.827617,6.58468,6.341743,6.1006193,6.590119,7.079619,7.569119,8.0604315,8.549932,8.722163,8.894395,9.066626,9.24067,9.412902,9.342196,9.273304,9.202598,9.131892,9.063,8.1148205,7.166641,6.2202744,5.272095,4.325729,5.239462,6.155008,7.0705543,7.9842873,8.899834,9.253361,9.605076,9.956791,10.310318,10.662033,8.689529,6.717026,4.744523,2.7720199,0.7995165,0.64722764,0.4949388,0.34264994,0.19036107,0.038072214,0.032633327,0.027194439,0.02175555,0.018129626,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.07433146,2.469255,4.8641787,7.2609153,9.655839,12.050762,10.080072,8.109382,6.1405044,4.169814,2.1991236,1.8020848,1.405046,1.0080072,0.6091554,0.21211663,0.17041849,0.12690738,0.08520924,0.04169814,0.0,0.27919623,0.56020546,0.83940166,1.1204109,1.3996071,1.35247,1.305333,1.258196,1.209246,1.162109,1.9725033,2.7828975,3.5932918,4.401873,5.2122674,5.4552045,5.6981416,5.9392653,6.1822023,6.4251394,6.970841,7.51473,8.0604315,8.604321,9.1500225,9.215289,9.280556,9.345822,9.409276,9.474543,9.40565,9.334945,9.264238,9.195346,9.12464,8.881703,8.640579,8.397643,8.154706,7.911769,8.281613,8.653271,9.023115,9.39296,9.762803,9.719293,9.677594,9.635896,9.592385,9.550687,10.165281,10.779876,11.39447,12.010877,12.625471,12.183108,11.740746,11.298383,10.854207,10.411844,10.448103,10.48255,10.516996,10.553255,10.587702,10.633025,10.6783495,10.721861,10.767185,10.812509,11.912977,13.011633,14.112101,15.212569,16.313038,16.017525,15.722012,15.428311,15.132799,14.837286,14.530895,14.222692,13.914488,13.608097,13.299893,13.499319,13.700559,13.899984,14.09941,14.300649,14.947877,15.595104,16.242332,16.889559,17.536787,18.495844,19.453089,20.410334,21.367577,22.324821,22.995617,23.6646,24.335396,25.00438,25.675177,26.4058,27.134611,27.865234,28.59586,29.324669,29.830486,30.33449,30.840307,31.34431,31.850126,30.8675,29.884874,28.90225,27.919624,26.936998,31.552801,36.16679,40.782593,45.398396,50.012386,48.96268,47.912975,46.86327,45.811752,44.762047,45.56156,46.362892,47.162407,47.961926,48.763256,50.520016,52.276775,54.03535,55.79211,57.550686,53.263027,48.975372,44.687714,40.40006,36.1124,31.5945,27.07841,22.560507,18.042604,13.524701,11.929294,10.3357,8.740293,7.1448855,5.5494785,6.0625467,6.5756154,7.0868707,7.5999393,8.113008,7.842876,7.572745,7.3026133,7.0324817,6.7623506,6.258347,5.75253,5.2467136,4.74271,4.2368937,4.4743915,4.7118897,4.949388,5.186886,5.424384,4.510651,3.5951047,2.6795588,1.7658255,0.85027945,2.7919624,4.7354584,6.677141,8.620637,10.56232,9.046683,7.5328593,6.017223,4.501586,2.9877625,3.6277382,4.267714,4.9076896,5.5476656,6.187641,5.7797246,5.371808,4.9657044,4.557788,4.1498713,3.9558845,3.7600844,3.5642843,3.3702974,3.1744974,5.422571,7.6706448,9.916905,12.164979,14.413053,13.087777,11.762501,10.437225,9.11195,7.7866745,7.175706,6.5629244,5.9501433,5.337362,4.7245803,5.3609304,5.995467,6.630004,7.264541,7.900891,7.077806,6.2547207,5.431636,4.610364,3.787279,3.9993954,4.213325,4.4254417,4.6375585,4.8496747,6.5157876,8.180087,9.844387,11.510499,13.174799,15.101978,17.029158,18.958149,20.885328,22.812508,22.785315,22.75812,22.729113,22.701918,22.674723,21.574255,20.4756,19.375132,18.274662,17.174194,17.61837,18.060734,18.503096,18.94546,19.387821,20.54993,21.71204,22.87415,24.03807,25.20018,22.464418,19.730473,16.99471,14.260764,11.525003,11.949236,12.375282,12.799516,13.225562,13.649796,12.9971285,12.344462,11.691795,11.039129,10.388275,9.474543,8.562622,7.650702,6.736969,5.825049,4.9095025,3.9957695,3.0802233,2.1646774,1.2491312,1.2219368,1.1947423,1.167548,1.1403534,1.1131591,1.3452182,1.5772774,1.8093367,2.0432088,2.275268,2.0667772,1.8600996,1.651609,1.4449311,1.2382535,1.1874905,1.1367276,1.0877775,1.0370146,0.9880646,0.91917205,0.8520924,0.7850128,0.7179332,0.6508536,2.0667772,3.484514,4.902251,6.319988,7.7377243,6.929143,6.1223745,5.315606,4.507025,3.7002566,3.8942437,4.0900435,4.2858434,4.4798307,4.6756306,4.358362,4.0392804,3.7220123,3.4047437,3.0874753,2.817344,2.5472124,2.277081,2.0069497,1.7368182,2.277081,2.817344,3.3576066,3.8978696,4.4381323,3.7220123,3.007705,2.2915847,1.5772774,0.8629702,0.9119202,0.96268314,1.0116332,1.062396,1.1131591,1.5845293,2.0577126,2.5308957,3.002266,3.4754493,3.0258346,2.5744069,2.124792,1.6751775,1.2255627,0.99531645,0.7650702,0.53482395,0.3045777,0.07433146,0.065266654,0.054388877,0.045324065,0.034446288,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.15047589,0.2991388,0.44961473,0.6000906,0.7505665,1.1457924,1.5392052,1.9344311,2.3296568,2.7248828,2.7357605,2.7448254,2.7557032,2.764768,2.7756457,4.3801174,5.9845896,7.590874,9.195346,10.799818,12.714307,14.630608,16.545097,18.459585,20.375887,17.166943,13.959812,10.752681,7.5455503,4.3366065,4.6429973,4.947575,5.2521524,5.5567303,5.863121,4.690134,3.5171473,2.3441606,1.1729867,0.0,0.059827764,0.11965553,0.1794833,0.23931105,0.2991388,0.5275721,0.7541924,0.9826257,1.209246,1.4376793,1.1494182,0.8629702,0.5747091,0.28826106,0.0,0.83940166,1.6806163,2.520018,3.3594196,4.2006345,3.392053,2.5852847,1.7767034,0.969935,0.16316663,0.17767033,0.19217403,0.20667773,0.2229944,0.2374981,0.19036107,0.14322405,0.09427405,0.047137026,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.014503701,0.018129626,0.01994259,0.02175555,0.025381476,0.02175555,0.01994259,0.018129626,0.014503701,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.014503701,0.018129626,0.01994259,0.02175555,0.025381476,0.038072214,0.05076295,0.06164073,0.07433146,0.0870222,0.09427405,0.10333887,0.11059072,0.11784257,0.12509441,0.12328146,0.11965553,0.11784257,0.11421664,0.11240368,0.10515183,0.09789998,0.09064813,0.08339628,0.07433146,0.07795739,0.07977036,0.08339628,0.08520924,0.0870222,0.09427405,0.10333887,0.11059072,0.11784257,0.12509441,0.18310922,0.23931105,0.29732585,0.35534066,0.41335547,0.40247768,0.39159992,0.3825351,0.37165734,0.36259252,0.3208944,0.27738327,0.23568514,0.19217403,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.0,0.0,0.0,0.0,0.0,2.811905,2.811905,2.811905,2.811905,2.811905,2.811905,3.3249733,3.8380418,4.349297,4.8623657,5.375434,5.1125546,4.8496747,4.5867953,4.325729,4.062849,4.936697,5.812358,6.688019,7.5618668,8.437528,8.437528,8.437528,8.437528,8.437528,8.437528,8.287052,8.138389,7.987913,7.837437,7.686961,7.311678,6.9382076,6.5629244,6.187641,5.812358,5.7253356,5.638314,5.5494785,5.462456,5.375434,5.1741953,4.974769,4.7753434,4.574105,4.3746786,5.2630305,6.149569,7.037921,7.9244595,8.812811,8.899834,8.9868555,9.07569,9.162713,9.249735,9.200785,9.1500225,9.099259,9.050309,8.999546,8.024173,7.0506115,6.0752378,5.0998635,4.12449,5.337362,6.550234,7.763106,8.974165,10.1870365,9.837135,9.487233,9.137331,8.78743,8.437528,6.7496595,5.0617914,3.3757362,1.6878681,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,2.0250793,3.9867048,5.9501433,7.911769,9.875207,8.200029,6.5248523,4.8496747,3.1744974,1.49932,1.2001812,0.89922947,0.6000906,0.2991388,0.0,0.0,0.0,0.0,0.0,0.0,0.18673515,0.37528324,0.5620184,0.7505665,0.93730164,0.89922947,0.8629702,0.824898,0.7868258,0.7505665,1.4630609,2.175555,2.8880494,3.6005437,4.313038,4.5632267,4.8116026,5.0617914,5.3119802,5.562169,6.3870673,7.211965,8.036863,8.861761,9.686659,9.862516,10.038374,10.212419,10.388275,10.56232,10.2378,9.91328,9.5869465,9.262425,8.937905,8.649645,8.363196,8.074935,7.7866745,7.500226,7.650702,7.799365,7.949841,8.100317,8.2507925,8.488291,8.725789,8.963287,9.200785,9.438283,10.399154,11.361836,12.32452,13.287203,14.249886,13.499319,12.750566,11.999999,11.249433,10.500679,10.587702,10.674724,10.761745,10.850581,10.937603,10.799818,10.662033,10.524248,10.388275,10.25049,11.374527,12.500377,13.6244135,14.750263,15.8743,15.838041,15.799969,15.761897,15.725637,15.687565,15.27421,14.862667,14.449312,14.037769,13.6244135,13.675177,13.724127,13.77489,13.825653,13.874602,14.487384,15.100165,15.712947,16.325727,16.936697,18.075237,19.211964,20.350506,21.487232,22.625772,23.662788,24.699802,25.736816,26.775644,27.812658,28.224201,28.637556,29.050913,29.462456,29.87581,30.124186,30.374374,30.624563,30.874752,31.12494,30.350807,29.574858,28.800724,28.024776,27.25064,33.67578,40.099106,46.52606,52.949387,59.374523,57.612324,55.850124,54.087925,52.325726,50.561714,51.437374,52.313034,53.186882,54.062546,54.938206,54.90013,54.86206,54.8258,54.787727,54.749657,52.012085,49.27451,46.536938,43.799362,41.06179,35.98731,30.912825,25.83653,20.762047,15.687565,13.762199,11.836833,9.91328,7.987913,6.0625467,6.43783,6.813113,7.1883965,7.5618668,7.93715,7.500226,7.063302,6.624565,6.187641,5.750717,5.3246713,4.900438,4.4743915,4.0501585,3.6241121,4.162562,4.699199,5.237649,5.774286,6.3127356,5.050914,3.787279,2.525457,1.261822,0.0,1.4249886,2.8499773,4.274966,5.6999545,7.124943,5.8377395,4.550536,3.2633326,1.9743162,0.6871128,2.03777,3.386614,4.7372713,6.0879283,7.4367723,6.987158,6.5375433,6.0879283,5.638314,5.186886,4.6248674,4.062849,3.5008307,2.9369993,2.374981,5.4497657,8.52455,11.599335,14.675932,17.750717,15.963136,14.175554,12.387974,10.600392,8.812811,8.136576,7.462154,6.787732,6.11331,5.4370747,5.863121,6.2873545,6.7134004,7.137634,7.5618668,6.6499467,5.7380266,4.8242936,3.9123733,3.000453,3.3249733,3.6494937,3.975827,4.3003473,4.6248674,6.4994707,8.374074,10.25049,12.125093,13.999697,15.174497,16.349297,17.52591,18.700708,19.87551,19.763105,19.650702,19.538298,19.425894,19.311678,18.537542,17.763407,16.98746,16.213324,15.437376,15.963136,16.487082,17.01284,17.536787,18.062546,19.099562,20.136576,21.175404,22.212418,23.249432,20.52455,17.799667,15.074784,12.349901,9.625018,10.038374,10.449916,10.863272,11.274815,11.6881695,11.050007,10.411844,9.775495,9.137331,8.499168,7.61263,6.7242785,5.8377395,4.949388,4.062849,3.2633326,2.4620032,1.6624867,0.8629702,0.06164073,0.13778515,0.21211663,0.28826106,0.36259252,0.43692398,0.72518504,1.0116332,1.2998942,1.5881553,1.8746033,1.6117238,1.3506571,1.0877775,0.824898,0.5620184,0.51306844,0.46230546,0.41335547,0.36259252,0.31182957,0.2991388,0.28826106,0.2755703,0.26287958,0.25018883,1.5881553,2.9243085,4.262275,5.600241,6.9382076,5.999093,5.0617914,4.12449,3.1871881,2.2498865,2.8499773,3.4500678,4.0501585,4.650249,5.2503395,4.6375585,4.024777,3.4119956,2.7992141,2.1882458,2.0123885,1.8383441,1.6624867,1.4866294,1.3125849,2.0250793,2.7375734,3.4500678,4.162562,4.8750563,4.0120864,3.150929,2.2879589,1.4249886,0.5620184,0.48768693,0.41335547,0.33721104,0.26287958,0.18673515,0.6508536,1.1131591,1.5754645,2.03777,2.5000753,2.2118144,1.9253663,1.6371052,1.3506571,1.062396,0.8629702,0.66173136,0.46230546,0.26287958,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.18673515,0.37528324,0.5620184,0.7505665,0.93730164,0.824898,0.7124943,0.6000906,0.48768693,0.37528324,0.8629702,1.3506571,1.8383441,2.324218,2.811905,4.4870825,6.16226,7.837437,9.512614,11.187792,13.475751,15.761897,18.049856,20.337814,22.625772,19.012539,15.399304,11.787883,8.174648,4.5632267,5.1125546,5.661882,6.2130227,6.7623506,7.311678,5.8504305,4.3873696,2.9243085,1.4630609,0.0,0.07433146,0.15047589,0.22480737,0.2991388,0.37528324,0.50037766,0.62547207,0.7505665,0.87566096,1.0007553,0.7995165,0.6000906,0.40066472,0.19942589,0.0,0.96268314,1.9253663,2.8880494,3.8507326,4.8116026,3.8869917,2.962381,2.03777,1.1131591,0.18673515,0.19942589,0.21211663,0.22480737,0.2374981,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.18673515,0.25018883,0.31182957,0.37528324,0.43692398,0.43692398,0.43692398,0.43692398,0.43692398,0.43692398,0.387974,0.33721104,0.28826106,0.2374981,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.0,0.0,0.0,0.0,0.0,3.5117085,3.4718235,3.4319382,3.392053,3.3521678,3.3122826,3.8108473,4.307599,4.804351,5.3029156,5.7996674,5.614745,5.429823,5.2449007,5.0599785,4.8750563,5.678199,6.4795284,7.2826705,8.0858135,8.887142,8.760235,8.6333275,8.504607,8.3777,8.2507925,8.187339,8.125698,8.062244,8.000604,7.93715,7.5872483,7.2373466,6.887445,6.5375433,6.187641,6.051669,5.91751,5.7833505,5.6473784,5.5132194,5.368182,5.223145,5.0781083,4.933071,4.788034,5.67276,6.5574856,7.4422116,8.326937,9.211663,9.137331,9.063,8.9868555,8.912524,8.838193,8.829127,8.821876,8.814624,8.807372,8.80012,7.9770355,7.155763,6.3326783,5.5095935,4.688321,6.816739,8.94697,11.077202,13.207433,15.337664,13.620788,11.9021,10.185224,8.4683485,6.7496595,5.4008155,4.0501585,2.6995013,1.3506571,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,1.789394,3.4681973,5.145188,6.8221784,8.499168,7.0469856,5.5948024,4.1426196,2.6904364,1.2382535,0.9898776,0.7433147,0.4949388,0.24837588,0.0,0.0,0.0,0.0,0.0,0.0,0.16497959,0.32995918,0.4949388,0.65991837,0.824898,0.78319985,0.73968875,0.6979906,0.6544795,0.61278135,1.2328146,1.8528478,2.472881,3.092914,3.7129474,4.0302157,4.347484,4.664753,4.9820213,5.2992897,6.1223745,6.94546,7.7667317,8.589817,9.412902,9.445535,9.4781685,9.510801,9.541622,9.574255,9.296872,9.019489,8.7421055,8.464723,8.187339,8.2798,8.372261,8.464723,8.557183,8.649645,8.762048,8.874452,8.9868555,9.099259,9.211663,9.334945,9.458226,9.579695,9.702975,9.824444,10.54419,11.26575,11.985496,12.705242,13.424988,12.757817,12.090648,11.421664,10.754494,10.087324,10.275872,10.462607,10.649343,10.837891,11.024626,10.830639,10.634838,10.440851,10.245051,10.049252,10.952107,11.854962,12.757817,13.660673,14.561715,14.86448,15.167245,15.47001,15.772775,16.075539,15.825351,15.575162,15.324973,15.074784,14.824595,14.5508375,14.275268,13.999697,13.724127,13.45037,14.057712,14.665054,15.272397,15.879739,16.487082,17.638313,18.787731,19.93715,21.08838,22.237799,23.195044,24.152288,25.109531,26.066776,27.025833,27.799969,28.574102,29.350052,30.124186,30.900135,31.123129,31.34431,31.567305,31.790298,32.013294,30.929142,29.846804,28.764463,27.682125,26.599787,31.706903,36.81402,41.922947,47.030064,52.137177,51.279648,50.422115,49.564583,48.707054,47.84952,48.799515,49.749508,50.699497,51.64949,52.599483,52.604923,52.610363,52.6158,52.619427,52.624866,50.550835,48.474995,46.39915,44.325123,42.24928,37.299892,32.350506,27.399303,22.449915,17.500528,15.732889,13.965251,12.197612,10.429974,8.662335,8.511859,8.363196,8.212721,8.062244,7.911769,7.382384,6.8529987,6.3218007,5.7924156,5.2630305,4.7898474,4.3166637,3.8452935,3.3721104,2.9007401,3.397492,3.8942437,4.3928084,4.88956,5.388125,4.503399,3.6168604,2.7321346,1.8474089,0.96268314,1.9326181,2.902553,3.872488,4.842423,5.812358,4.8242936,3.8380418,2.8499773,1.8619126,0.87566096,1.889107,2.904366,3.919625,4.934884,5.9501433,5.9120708,5.8758116,5.8377395,5.7996674,5.763408,5.1343102,4.507025,3.87974,3.2524548,2.6251698,5.277534,7.9298983,10.582263,13.234627,15.8869915,14.646925,13.406858,12.166792,10.926725,9.686659,8.974165,8.26167,7.549176,6.836682,6.1241875,6.147756,6.169512,6.19308,6.2148356,6.2365913,5.529536,4.8224807,4.115425,3.4083695,2.6995013,3.1708715,3.6404288,4.1099863,4.5795436,5.049101,6.78048,8.510046,10.239613,11.969179,13.700559,14.599788,15.50083,16.400059,17.29929,18.20033,18.347181,18.495844,18.642694,18.789545,18.938208,18.087927,17.237648,16.38737,15.537089,14.68681,15.0693445,15.45188,15.834415,16.21695,16.599485,17.384499,18.169512,18.954523,19.739536,20.52455,18.189453,15.854358,13.519262,11.184166,8.8508835,9.131892,9.414715,9.697536,9.980359,10.263181,9.659465,9.057561,8.455658,7.851941,7.250037,6.4831543,5.714458,4.947575,4.1806917,3.4119956,2.7466383,2.0830941,1.4177368,0.7523795,0.0870222,0.13959812,0.19217403,0.24474995,0.29732585,0.34990177,0.7106813,1.0696479,1.4304274,1.789394,2.1501737,1.84197,1.5355793,1.2273756,0.91917205,0.61278135,0.5529536,0.49312583,0.43329805,0.37165734,0.31182957,0.29732585,0.28282216,0.26831847,0.2520018,0.2374981,1.3180238,2.3967366,3.4772623,4.557788,5.638314,4.8750563,4.1117992,3.350355,2.5870976,1.8256533,2.4021754,2.9805105,3.5570326,4.135368,4.7118897,4.157123,3.6023567,3.04759,2.4928236,1.938057,1.7603867,1.5827163,1.405046,1.2273756,1.0497054,1.6606737,2.269829,2.8807976,3.489953,4.099108,3.3793623,2.659616,1.93987,1.2201238,0.50037766,0.42967212,0.36077955,0.29007402,0.21936847,0.15047589,0.5946517,1.0406405,1.4848163,1.9308052,2.374981,2.126605,1.8800422,1.6316663,1.3851035,1.1367276,0.91917205,0.7016165,0.48587397,0.26831847,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.15047589,0.2991388,0.44961473,0.6000906,0.7505665,0.65991837,0.56927025,0.48043507,0.38978696,0.2991388,1.0478923,1.794833,2.5417736,3.290527,4.0374675,7.5654926,11.091705,14.61973,18.147755,21.675781,21.003172,20.330563,19.657953,18.985344,18.312735,16.175253,14.037769,11.900287,9.762803,7.6253204,7.567306,7.509291,7.453089,7.3950744,7.3370595,5.9900284,4.6429973,3.294153,1.9471219,0.6000906,0.6653573,0.7306239,0.79589057,0.85934424,0.9246109,0.90466833,0.88472575,0.86478317,0.8448406,0.824898,0.66173136,0.50037766,0.33721104,0.17585737,0.012690738,0.92823684,1.84197,2.7575161,3.673062,4.5867953,3.7056956,2.8227828,1.93987,1.0569572,0.17585737,0.18673515,0.19942589,0.21211663,0.22480737,0.2374981,0.19036107,0.14322405,0.09427405,0.047137026,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.072518505,0.08339628,0.092461094,0.10333887,0.11240368,0.11784257,0.12328146,0.12690738,0.13234627,0.13778515,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.07433146,0.07433146,0.07433146,0.07433146,0.07433146,0.08520924,0.09427405,0.10515183,0.11421664,0.12509441,0.1794833,0.23568514,0.29007402,0.3444629,0.40066472,0.40066472,0.40066472,0.40066472,0.40066472,0.40066472,0.36077955,0.3208944,0.27919623,0.23931105,0.19942589,0.16497959,0.13053331,0.09427405,0.059827764,0.025381476,0.02175555,0.01994259,0.018129626,0.014503701,0.012690738,4.213325,4.1317415,4.0519714,3.972201,3.8924308,3.8126602,4.2949085,4.7771564,5.2594047,5.7416525,6.2257137,6.1169357,6.009971,5.903006,5.7942286,5.6872635,6.4178877,7.1466985,7.877322,8.607946,9.336758,9.082943,8.827314,8.571687,8.317872,8.062244,8.087626,8.113008,8.138389,8.161958,8.187339,7.8628187,7.5382986,7.211965,6.887445,6.5629244,6.379815,6.1967063,6.01541,5.8323007,5.6491914,5.560356,5.469708,5.3808727,5.290225,5.199577,6.0824895,6.965402,7.8483152,8.729415,9.612328,9.374829,9.137331,8.899834,8.662335,8.424837,8.459284,8.495543,8.529989,8.564435,8.600695,7.9298983,7.2609153,6.590119,5.919323,5.2503395,8.29793,11.34552,14.39311,17.4407,20.48829,17.402628,14.316965,11.233116,8.147454,5.0617914,4.0501585,3.0367124,2.0250793,1.0116332,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.032633327,0.065266654,0.09789998,0.13053331,0.16316663,1.5555218,2.9478772,4.3402324,5.732588,7.124943,5.8957543,4.664753,3.435564,2.2045624,0.97537386,0.7795739,0.5855869,0.38978696,0.19579996,0.0,0.0,0.0,0.0,0.0,0.0,0.14322405,0.28463513,0.42785916,0.56927025,0.7124943,0.6653573,0.61822027,0.56927025,0.52213323,0.4749962,1.0025684,1.5301404,2.0577126,2.5852847,3.1128569,3.4972048,3.8833659,4.267714,4.652062,5.038223,5.857682,6.677141,7.498413,8.317872,9.137331,9.026741,8.917963,8.807372,8.696781,8.588004,8.357758,8.127511,7.897265,7.667019,7.4367723,7.909956,8.383139,8.854509,9.327692,9.800876,9.875207,9.949538,10.025683,10.100015,10.174346,10.183411,10.190662,10.197914,10.205167,10.212419,10.689227,11.16785,11.644659,12.123281,12.60009,12.0145035,11.430729,10.845142,10.259555,9.675781,9.96223,10.25049,10.536939,10.825199,11.111648,10.859646,10.607644,10.355642,10.101828,9.849826,10.529687,11.209548,11.889409,12.569269,13.24913,13.892733,14.534521,15.1781225,15.819912,16.4617,16.374678,16.287657,16.200634,16.1118,16.024776,15.4246855,14.824595,14.224504,13.6244135,13.024323,13.628039,14.229943,14.831847,15.435563,16.037468,17.199575,18.361685,19.525606,20.687716,21.849825,22.727299,23.604773,24.482246,25.35972,26.237194,27.375734,28.512463,29.64919,30.787731,31.924458,32.12026,32.314243,32.510044,32.705845,32.899834,31.509289,30.12056,28.730019,27.339476,25.950747,29.739838,33.530743,37.319836,41.11074,44.89983,44.946968,44.994106,45.043056,45.09019,45.13733,46.16165,47.18779,48.212112,49.23825,50.262573,50.30971,50.35685,50.4058,50.452934,50.500072,49.087776,47.675476,46.26318,44.85088,43.43677,38.612476,33.788185,28.962078,24.137783,19.311678,17.701767,16.091856,14.481945,12.872034,11.262123,10.587702,9.91328,9.237044,8.562622,7.8882003,7.264541,6.642695,6.0208488,5.3971896,4.7753434,4.255023,3.7347028,3.2143826,2.6958754,2.175555,2.6324217,3.0892882,3.5479677,4.004834,4.461701,3.9558845,3.4482548,2.9406252,2.4329958,1.9253663,2.4402475,2.955129,3.4700103,3.9848917,4.499773,3.8126602,3.1255474,2.4366217,1.7495089,1.062396,1.742257,2.422118,3.101979,3.7818398,4.461701,4.836984,5.2122674,5.5875506,5.962834,6.338117,5.6455655,4.953014,4.2604623,3.5679104,2.8753586,5.105303,7.3352466,9.56519,11.795135,14.025079,13.332527,12.639976,11.947423,11.254871,10.56232,9.811753,9.063,8.312433,7.5618668,6.813113,6.432391,6.051669,5.67276,5.292038,4.9131284,4.409125,3.9069343,3.4047437,2.902553,2.4003625,3.0149567,3.6295512,4.2441454,4.860553,5.475147,7.059676,8.644206,10.230548,11.815077,13.399607,14.025079,14.650551,15.27421,15.899682,16.525154,16.933071,17.339174,17.747091,18.155006,18.562923,17.638313,16.71189,15.787278,14.862667,13.938056,14.177367,14.416678,14.657803,14.897114,15.138238,15.6694355,16.202446,16.735458,17.266655,17.799667,15.854358,13.910862,11.965553,10.020245,8.074935,8.227224,8.379513,8.531802,8.684091,8.838193,8.270736,7.703278,7.135821,6.5683637,5.999093,5.351866,4.704638,4.0574102,3.4101827,2.762955,2.231757,1.7023718,1.1729867,0.6417888,0.11240368,0.14322405,0.17223145,0.2030518,0.23205921,0.26287958,0.69436467,1.1276628,1.5591478,1.9924458,2.4257438,2.0722163,1.7205015,1.3669738,1.015259,0.66173136,0.59283876,0.52213323,0.45324063,0.3825351,0.31182957,0.2955129,0.27738327,0.25925365,0.24293698,0.22480737,1.0478923,1.8691645,2.6922495,3.5153344,4.3366065,3.7492065,3.1618068,2.5744069,1.987007,1.3996071,1.9543737,2.5091403,3.0657198,3.6204863,4.175253,3.6766882,3.1799364,2.6831846,2.18462,1.6878681,1.5083848,1.3270886,1.1476053,0.968122,0.7868258,1.2944553,1.8020848,2.3097143,2.817344,3.3249733,2.7466383,2.1701162,1.5917811,1.015259,0.43692398,0.37165734,0.30820364,0.24293698,0.17767033,0.11240368,0.5402629,0.968122,1.3941683,1.8220274,2.2498865,2.0432088,1.8347181,1.6280404,1.4195497,1.2128719,0.97718686,0.7433147,0.5076295,0.27194437,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.11240368,0.22480737,0.33721104,0.44961473,0.5620184,0.4949388,0.42785916,0.36077955,0.291887,0.22480737,1.2328146,2.2408218,3.247016,4.255023,5.2630305,10.642091,16.022963,21.402023,26.782896,32.161957,28.530592,24.897415,21.264238,17.632874,13.999697,13.337966,12.674421,12.012691,11.349146,10.687414,10.022058,9.3567,8.693155,8.027799,7.362441,6.1296263,4.896812,3.6658103,2.4329958,1.2001812,1.2545701,1.310772,1.3651608,1.4195497,1.4757515,1.310772,1.1457924,0.9808127,0.81583315,0.6508536,0.52575916,0.40066472,0.2755703,0.15047589,0.025381476,0.8919776,1.7603867,2.6269827,3.4953918,4.361988,3.5225863,2.6831846,1.84197,1.0025684,0.16316663,0.17585737,0.18673515,0.19942589,0.21211663,0.22480737,0.1794833,0.13415924,0.09064813,0.045324065,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.07070554,0.07795739,0.08520924,0.092461094,0.099712946,0.11059072,0.11965553,0.13053331,0.13959812,0.15047589,0.13778515,0.12509441,0.11240368,0.099712946,0.0870222,0.0870222,0.0870222,0.0870222,0.0870222,0.0870222,0.09427405,0.10333887,0.11059072,0.11784257,0.12509441,0.17223145,0.21936847,0.26831847,0.3154555,0.36259252,0.36259252,0.36259252,0.36259252,0.36259252,0.36259252,0.33177215,0.30276474,0.27194437,0.24293698,0.21211663,0.1794833,0.14684997,0.11421664,0.08339628,0.05076295,0.045324065,0.03988518,0.034446288,0.030820364,0.025381476,4.9131284,4.7916603,4.6720047,4.552349,4.4326935,4.313038,4.780782,5.2467136,5.714458,6.1822023,6.6499467,6.6191263,6.590119,6.5592985,6.530291,6.4994707,7.157576,7.8156815,8.471974,9.130079,9.788185,9.40565,9.023115,8.640579,8.258044,7.8755093,7.987913,8.100317,8.212721,8.325124,8.437528,8.138389,7.837437,7.5382986,7.2373466,6.9382076,6.7079616,6.4777155,6.247469,6.017223,5.7869763,5.75253,5.718084,5.6818247,5.6473784,5.612932,6.492219,7.3733187,8.252605,9.131892,10.012992,9.612328,9.211663,8.812811,8.412147,8.013294,8.089439,8.167397,8.245354,8.323311,8.399456,7.8827615,7.364254,6.8475595,6.3308654,5.812358,9.7773075,13.742256,17.707205,21.672155,25.637104,21.184467,16.731833,12.279196,7.8265595,3.3757362,2.6995013,2.0250793,1.3506571,0.6744221,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.04169814,0.08520924,0.12690738,0.17041849,0.21211663,1.3198367,2.427557,3.5352771,4.6429973,5.750717,4.74271,3.7347028,2.7266958,1.7205015,0.7124943,0.56927025,0.42785916,0.28463513,0.14322405,0.0,0.0,0.0,0.0,0.0,0.0,0.11965553,0.23931105,0.36077955,0.48043507,0.6000906,0.5475147,0.4949388,0.44236287,0.38978696,0.33721104,0.77232206,1.2074331,1.6425442,2.077655,2.5127661,2.9641938,3.4174345,3.870675,4.322103,4.7753434,5.5929894,6.4106355,7.228282,8.044115,8.861761,8.609759,8.357758,8.105756,7.851941,7.5999393,7.41683,7.2355337,7.0524244,6.869315,6.688019,7.5401115,8.392203,9.244296,10.098202,10.950294,10.988366,11.024626,11.062697,11.10077,11.137029,11.030065,10.9230995,10.8143215,10.707357,10.600392,10.834265,11.069949,11.3056345,11.539507,11.775192,11.273002,10.770811,10.266808,9.764616,9.262425,9.6504,10.038374,10.424535,10.812509,11.200482,10.890467,10.58045,10.270433,9.960417,9.6504,10.107266,10.564133,11.022813,11.479679,11.938358,12.919171,13.901797,14.884423,15.867048,16.849674,16.92582,17.00015,17.074482,17.150625,17.224958,16.300346,15.375735,14.449312,13.524701,12.60009,13.198368,13.794832,14.39311,14.989574,15.5878525,16.762651,17.937452,19.112251,20.287052,21.461851,22.259554,23.057259,23.854961,24.652666,25.450369,26.949688,28.45082,29.950142,31.449461,32.950596,33.117386,33.28418,33.452785,33.61958,33.788185,32.08944,30.392506,28.695572,26.996826,25.299892,27.772774,30.245655,32.716724,35.1896,37.662483,38.61429,39.56791,40.519714,41.47333,42.425137,43.525604,44.62426,45.724728,46.8252,47.925667,48.0145,48.10515,48.195797,48.284634,48.375282,47.624714,46.87415,46.125393,45.37483,44.62426,39.92506,35.225864,30.52485,25.825651,21.12464,19.672457,18.220274,16.768091,15.314095,13.861912,12.661731,11.463363,10.263181,9.063,7.8628187,7.1466985,6.432391,5.718084,5.0019636,4.2876563,3.720199,3.152742,2.5852847,2.0178273,1.4503701,1.8673514,2.2843328,2.7031271,3.1201086,3.53709,3.4083695,3.2778363,3.147303,3.0167696,2.8880494,2.9478772,3.007705,3.0675328,3.1273603,3.1871881,2.7992141,2.4130533,2.0250793,1.6371052,1.2491312,1.5954071,1.93987,2.2843328,2.6306088,2.9750717,3.7618973,4.550536,5.337362,6.1241875,6.9128265,6.155008,5.3971896,4.6393714,3.8833659,3.1255474,4.933071,6.740595,8.548119,10.355642,12.163166,12.018129,11.873092,11.728055,11.583018,11.437981,10.649343,9.862516,9.07569,8.287052,7.500226,6.717026,5.9356394,5.1524396,4.36924,3.587853,3.290527,2.9932013,2.6958754,2.3967366,2.0994108,2.8608549,3.6204863,4.3801174,5.139749,5.89938,7.3406854,8.780178,10.21967,11.6591625,13.100468,13.45037,13.800271,14.150173,14.500074,14.849977,15.517147,16.184317,16.8533,17.52047,18.187641,17.186886,16.187943,15.187187,14.188245,13.1874895,13.28539,13.383289,13.479377,13.577277,13.675177,13.954373,14.235382,14.514579,14.795588,15.074784,13.519262,11.965553,10.410031,8.854509,7.3008003,7.322556,7.344311,7.36788,7.3896356,7.413204,6.880193,6.347182,5.814171,5.282973,4.749962,4.2223897,3.6948178,3.1672456,2.6396735,2.1121013,1.7168756,1.3216497,0.92823684,0.533011,0.13778515,0.14503701,0.15228885,0.15954071,0.16679256,0.17585737,0.67986095,1.1856775,1.6896812,2.1954978,2.6995013,2.3024626,1.9054236,1.5083848,1.1095331,0.7124943,0.6327239,0.5529536,0.47318324,0.39159992,0.31182957,0.291887,0.27194437,0.2520018,0.23205921,0.21211663,0.7777609,1.3415923,1.9072367,2.472881,3.0367124,2.6251698,2.2118144,1.8002719,1.3869164,0.97537386,1.5083848,2.039583,2.572594,3.105605,3.636803,3.198066,2.7575161,2.3169663,1.8782293,1.4376793,1.2545701,1.0732739,0.8901646,0.7070554,0.52575916,0.9300498,1.3343405,1.7404441,2.1447346,2.5508385,2.1157274,1.6806163,1.2455053,0.8103943,0.37528324,0.3154555,0.25562772,0.19579996,0.13415924,0.07433146,0.48587397,0.89560354,1.305333,1.7150626,2.124792,1.9579996,1.789394,1.6226015,1.455809,1.2872034,1.0352017,0.78319985,0.5293851,0.27738327,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07433146,0.15047589,0.22480737,0.2991388,0.37528324,0.32995918,0.28463513,0.23931105,0.19579996,0.15047589,1.4177368,2.6849976,3.9522583,5.219519,6.48678,13.720501,20.952408,28.184317,35.418037,42.649944,36.0562,29.464268,22.872335,16.280403,9.686659,10.500679,11.312886,12.125093,12.937301,13.749508,12.476809,11.205922,9.933222,8.660522,7.3878226,6.2692246,5.1524396,4.0356545,2.9170568,1.8002719,1.845596,1.889107,1.9344311,1.9797552,2.0250793,1.7150626,1.405046,1.0950294,0.7850128,0.4749962,0.387974,0.2991388,0.21211663,0.12509441,0.038072214,0.8575313,1.6769904,2.4982624,3.3177216,4.137181,3.339477,2.5417736,1.74407,0.9481794,0.15047589,0.16316663,0.17585737,0.18673515,0.19942589,0.21211663,0.17041849,0.12690738,0.08520924,0.04169814,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.06707962,0.072518505,0.07795739,0.08339628,0.0870222,0.10333887,0.11784257,0.13234627,0.14684997,0.16316663,0.15047589,0.13778515,0.12509441,0.11240368,0.099712946,0.099712946,0.099712946,0.099712946,0.099712946,0.099712946,0.10515183,0.11059072,0.11421664,0.11965553,0.12509441,0.16497959,0.20486477,0.24474995,0.28463513,0.3245203,0.3245203,0.3245203,0.3245203,0.3245203,0.3245203,0.3045777,0.28463513,0.26469254,0.24474995,0.22480737,0.19579996,0.16497959,0.13415924,0.10515183,0.07433146,0.06707962,0.059827764,0.052575916,0.045324065,0.038072214,5.612932,5.4533916,5.292038,5.132497,4.972956,4.8116026,5.2648435,5.718084,6.169512,6.622752,7.07418,7.12313,7.170267,7.217404,7.264541,7.311678,7.897265,8.482852,9.066626,9.652213,10.2378,9.728357,9.217102,8.70766,8.198216,7.686961,7.8882003,8.087626,8.287052,8.488291,8.6877165,8.412147,8.138389,7.8628187,7.5872483,7.311678,7.0342946,6.7569118,6.4795284,6.202145,5.924762,5.9447045,5.964647,5.9845896,6.004532,6.0244746,6.9019485,7.7794223,8.656897,9.53437,10.411844,9.849826,9.287807,8.725789,8.161958,7.5999393,7.7195945,7.83925,7.9607186,8.080374,8.200029,7.835624,7.4694057,7.1050005,6.740595,6.3743763,11.256684,16.138992,21.023113,25.905422,30.787731,24.96812,19.14851,13.327088,7.507478,1.6878681,1.3506571,1.0116332,0.6744221,0.33721104,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.052575916,0.10515183,0.15772775,0.21030366,0.26287958,1.0841516,1.9072367,2.7303216,3.5534067,4.3746786,3.589666,2.8046532,2.0196402,1.2346275,0.44961473,0.36077955,0.27013144,0.1794833,0.09064813,0.0,0.0,0.0,0.0,0.0,0.0,0.09789998,0.19579996,0.291887,0.38978696,0.48768693,0.42967212,0.37165734,0.3154555,0.2574407,0.19942589,0.5420758,0.88472575,1.2273756,1.5700256,1.9126755,2.4329958,2.953316,3.4718235,3.9921436,4.512464,5.328297,6.1423173,6.9581504,7.7721705,8.588004,8.192778,7.797552,7.402326,7.0071006,6.6118746,6.4777155,6.341743,6.207584,6.071612,5.9374523,7.170267,8.403082,9.635896,10.866898,12.099712,12.099712,12.099712,12.099712,12.099712,12.099712,11.876718,11.655537,11.432542,11.209548,10.988366,10.979301,10.97205,10.964798,10.957546,10.950294,10.529687,10.110892,9.690285,9.269678,8.8508835,9.336758,9.824444,10.312131,10.799818,11.287505,10.919474,10.553255,10.185224,9.817192,9.449161,9.684846,9.920531,10.154404,10.390089,10.625773,11.947423,13.2690735,14.592536,15.914186,17.237648,17.475147,17.712645,17.950142,18.187641,18.425138,17.174194,15.925063,14.674119,13.424988,12.175857,12.766883,13.359721,13.95256,14.545399,15.138238,16.325727,17.513218,18.700708,19.888199,21.07569,21.791811,22.509743,23.227676,23.94561,24.66173,26.525455,28.387367,30.24928,32.113007,33.97492,34.114517,34.254116,34.395527,34.535126,34.67472,32.669586,30.66445,28.659313,26.654177,24.650852,25.80571,26.960567,28.115423,29.27028,30.425138,32.281612,34.1399,35.998184,37.85466,39.712944,40.887745,42.062546,43.237343,44.412144,45.586945,45.71929,45.851635,45.985794,46.11814,46.25049,46.16165,46.07463,45.98761,45.900585,45.811752,41.237648,36.663544,32.087624,27.511707,22.937603,21.643147,20.34688,19.052423,17.757969,16.4617,14.737573,13.013446,11.287505,9.563377,7.837437,7.0306687,6.2220874,5.4153194,4.606738,3.7999697,3.1853752,2.570781,1.9543737,1.3397794,0.72518504,1.1022812,1.4793775,1.8582866,2.2353828,2.612479,2.8608549,3.1074178,3.3557937,3.6023567,3.8507326,3.4555066,3.0602808,2.665055,2.269829,1.8746033,1.7875811,1.7005589,1.6117238,1.5247015,1.4376793,1.4467441,1.4576219,1.4666867,1.4775645,1.4866294,2.6868105,3.8869917,5.087173,6.2873545,7.4875355,6.6644506,5.8431783,5.0200934,4.1970086,3.3757362,4.76084,6.14413,7.5292335,8.914337,10.29944,10.701918,11.104396,11.506873,11.909351,12.311829,11.486931,10.662033,9.837135,9.012237,8.187339,7.0016613,5.8177967,4.632119,3.4482548,2.2625773,2.1701162,2.077655,1.9851941,1.892733,1.8002719,2.70494,3.6096084,4.514277,5.4207582,6.3254266,7.6198816,8.914337,10.210606,11.50506,12.799516,12.87566,12.949992,13.024323,13.100468,13.174799,14.103036,15.02946,15.957697,16.88412,17.812357,16.73727,15.662184,14.587097,13.512011,12.436923,12.3916,12.348088,12.302764,12.25744,12.212116,12.23931,12.268318,12.295512,12.322706,12.349901,11.184166,10.020245,8.854509,7.690587,6.5248523,6.4178877,6.3091097,6.202145,6.09518,5.9882154,5.4896507,4.992899,4.494334,3.9975824,3.5008307,3.092914,2.6849976,2.277081,1.8691645,1.4630609,1.2019942,0.94274056,0.68167394,0.4224203,0.16316663,0.14684997,0.13234627,0.11784257,0.10333887,0.0870222,0.6653573,1.2418793,1.8202144,2.3967366,2.9750717,2.5327086,2.0903459,1.647983,1.2056202,0.76325727,0.6726091,0.581961,0.49312583,0.40247768,0.31182957,0.29007402,0.26831847,0.24474995,0.2229944,0.19942589,0.5076295,0.81583315,1.1222239,1.4304274,1.7368182,1.49932,1.261822,1.0243238,0.7868258,0.5493277,1.0605831,1.5700256,2.079468,2.5907235,3.100166,2.7176309,2.335096,1.9525607,1.5700256,1.1874905,1.0025684,0.81764615,0.6327239,0.44780177,0.26287958,0.5656443,0.8665961,1.1693609,1.4721256,1.7748904,1.4830034,1.1893034,0.8974165,0.6055295,0.31182957,0.2574407,0.2030518,0.14684997,0.092461094,0.038072214,0.42967212,0.823085,1.214685,1.6080978,1.9996977,1.8727903,1.745883,1.6171626,1.4902552,1.3633479,1.0932164,0.823085,0.5529536,0.28282216,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.16497959,0.14322405,0.11965553,0.09789998,0.07433146,1.6026589,3.1291735,4.6575007,6.185828,7.7123427,16.798912,25.881853,34.968422,44.053177,53.13793,43.583622,34.032932,24.480434,14.927934,5.375434,7.663393,9.949538,12.237497,14.525456,16.811602,14.93156,13.05333,11.173288,9.293246,7.413204,6.4106355,5.408067,4.405499,3.4029307,2.4003625,2.4348087,2.469255,2.5055144,2.5399606,2.5744069,2.1193533,1.6642996,1.209246,0.7541924,0.2991388,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.823085,1.5954071,2.3677292,3.1400511,3.9123733,3.1581807,2.4021754,1.647983,0.8919776,0.13778515,0.15047589,0.16316663,0.17585737,0.18673515,0.19942589,0.15954071,0.11965553,0.07977036,0.03988518,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.065266654,0.06707962,0.07070554,0.072518505,0.07433146,0.09427405,0.11421664,0.13415924,0.15410182,0.17585737,0.16316663,0.15047589,0.13778515,0.12509441,0.11240368,0.11240368,0.11240368,0.11240368,0.11240368,0.11240368,0.11421664,0.11784257,0.11965553,0.12328146,0.12509441,0.15772775,0.19036107,0.2229944,0.25562772,0.28826106,0.28826106,0.28826106,0.28826106,0.28826106,0.28826106,0.27738327,0.26831847,0.2574407,0.24837588,0.2374981,0.21030366,0.18310922,0.15410182,0.12690738,0.099712946,0.09064813,0.07977036,0.07070554,0.059827764,0.05076295,6.3127356,6.11331,5.9120708,5.712645,5.5132194,5.3119802,5.750717,6.187641,6.624565,7.063302,7.500226,7.6253204,7.750415,7.8755093,8.000604,8.125698,8.636953,9.1500225,9.663091,10.174346,10.687414,10.049252,9.412902,8.774739,8.138389,7.500226,7.7866745,8.074935,8.363196,8.649645,8.937905,8.6877165,8.437528,8.187339,7.93715,7.686961,7.362441,7.037921,6.7115874,6.3870673,6.0625467,6.1368785,6.2130227,6.2873545,6.3616858,6.43783,7.311678,8.187339,9.063,9.936848,10.812509,10.087324,9.362139,8.636953,7.911769,7.1883965,7.3497505,7.512917,7.6742706,7.837437,8.000604,7.7866745,7.574558,7.362441,7.1503243,6.9382076,12.737875,18.537542,24.33721,30.136877,35.93836,28.74996,21.563377,14.37498,7.1865835,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06164073,0.12509441,0.18673515,0.25018883,0.31182957,0.85027945,1.3869164,1.9253663,2.4620032,3.000453,2.4366217,1.8746033,1.3125849,0.7505665,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.0,0.0,0.0,0.0,0.0,0.07433146,0.15047589,0.22480737,0.2991388,0.37528324,0.31182957,0.25018883,0.18673515,0.12509441,0.06164073,0.31182957,0.5620184,0.8122072,1.062396,1.3125849,1.8999848,2.4873846,3.0747845,3.6621845,4.249584,5.0617914,5.8758116,6.688019,7.500226,8.312433,7.7757964,7.2373466,6.70071,6.16226,5.6256227,5.5367875,5.4497657,5.3627434,5.275721,5.186886,6.8004227,8.412147,10.025683,11.637406,13.24913,13.212872,13.174799,13.136727,13.100468,13.062395,12.725184,12.387974,12.050762,11.711739,11.374527,11.124338,10.874149,10.625773,10.375585,10.125396,9.788185,9.449161,9.11195,8.774739,8.437528,9.024928,9.612328,10.199727,10.7871275,11.374527,10.950294,10.524248,10.100015,9.675781,9.249735,9.262425,9.275117,9.287807,9.300498,9.313189,10.975676,12.638163,14.300649,15.963136,17.625622,18.024473,18.425138,18.825804,19.224655,19.62532,18.049856,16.474392,14.90074,13.325275,11.74981,12.337211,12.92461,13.512011,14.09941,14.68681,15.8869915,17.087172,18.287354,19.487535,20.687716,21.325878,21.962229,22.600391,23.236742,23.874905,26.09941,28.325727,30.550232,32.77474,34.99924,35.111645,35.225864,35.33827,35.450672,35.563072,33.249733,30.938206,28.624866,26.31334,23.999998,23.836832,23.675478,23.512312,23.349146,23.187792,25.950747,28.71189,31.474844,34.237797,37.00075,38.249886,39.500828,40.74996,42.000904,43.250034,43.42589,43.599937,43.775795,43.94984,44.125698,44.700405,45.275116,45.849823,46.424534,46.99924,42.550232,38.099407,33.6504,29.199575,24.750565,23.612024,22.475298,21.336756,20.20003,19.063301,16.813416,14.561715,12.311829,10.061942,7.8120556,6.9128265,6.011784,5.1125546,4.213325,3.3122826,2.6505513,1.987007,1.3252757,0.66173136,0.0,0.33721104,0.6744221,1.0116332,1.3506571,1.6878681,2.3133402,2.9369993,3.5624714,4.1879435,4.8116026,3.9631362,3.1128569,2.2625773,1.4122978,0.5620184,0.774135,0.9880646,1.2001812,1.4122978,1.6244144,1.2998942,0.97537386,0.6508536,0.3245203,0.0,1.6117238,3.2252605,4.836984,6.450521,8.062244,7.175706,6.2873545,5.4008155,4.512464,3.6241121,4.5867953,5.5494785,6.5121617,7.474845,8.437528,9.38752,10.337513,11.287505,12.237497,13.1874895,12.32452,11.463363,10.600392,9.737422,8.874452,7.28811,5.6999545,4.1117992,2.525457,0.93730164,1.0497054,1.162109,1.2745126,1.3869164,1.49932,2.5508385,3.6005437,4.650249,5.6999545,6.7496595,7.900891,9.050309,10.199727,11.349146,12.500377,12.299138,12.099712,11.900287,11.700861,11.499621,12.687112,13.874602,15.062093,16.249584,17.437075,16.287657,15.138238,13.987006,12.837588,11.6881695,11.499621,11.312886,11.124338,10.937603,10.750868,10.524248,10.29944,10.074633,9.849826,9.625018,8.849071,8.074935,7.3008003,6.5248523,5.750717,5.5132194,5.275721,5.038223,4.800725,4.5632267,4.099108,3.636803,3.1744974,2.712192,2.2498865,1.9616255,1.6751775,1.3869164,1.1004683,0.8122072,0.6871128,0.5620184,0.43692398,0.31182957,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.6508536,1.2998942,1.9507477,2.5997884,3.2506418,2.762955,2.275268,1.7875811,1.2998942,0.8122072,0.7124943,0.61278135,0.51306844,0.41335547,0.31182957,0.28826106,0.26287958,0.2374981,0.21211663,0.18673515,0.2374981,0.28826106,0.33721104,0.387974,0.43692398,0.37528324,0.31182957,0.25018883,0.18673515,0.12509441,0.61278135,1.1004683,1.5881553,2.0758421,2.561716,2.2371957,1.9126755,1.5881553,1.261822,0.93730164,0.7505665,0.5620184,0.37528324,0.18673515,0.0,0.19942589,0.40066472,0.6000906,0.7995165,1.0007553,0.85027945,0.69980353,0.5493277,0.40066472,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.37528324,0.7505665,1.1258497,1.49932,1.8746033,1.7875811,1.7005589,1.6117238,1.5247015,1.4376793,1.1494182,0.8629702,0.5747091,0.28826106,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.7875811,3.5751622,5.3627434,7.1503243,8.937905,19.87551,30.811298,41.750717,52.68832,63.624107,51.111042,38.599785,26.08672,13.575464,1.062396,4.8261065,8.588004,12.349901,16.1118,19.87551,17.388124,14.90074,12.411542,9.924157,7.4367723,6.550234,5.661882,4.7753434,3.8869917,3.000453,3.0258346,3.049403,3.0747845,3.100166,3.1255474,2.525457,1.9253663,1.3252757,0.72518504,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.7868258,1.5120108,2.2371957,2.962381,3.6875658,2.9750717,2.2625773,1.550083,0.8375887,0.12509441,0.13778515,0.15047589,0.16316663,0.17585737,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.0870222,0.11240368,0.13778515,0.16316663,0.18673515,0.17585737,0.16316663,0.15047589,0.13778515,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.15047589,0.17585737,0.19942589,0.22480737,0.25018883,0.25018883,0.25018883,0.25018883,0.25018883,0.25018883,0.25018883,0.25018883,0.25018883,0.25018883,0.25018883,0.22480737,0.19942589,0.17585737,0.15047589,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,5.863121,5.710832,5.5567303,5.4044414,5.2521524,5.0998635,5.580299,6.060734,6.539356,7.019791,7.500226,7.706904,7.915395,8.122072,8.330563,8.537241,8.834567,9.131892,9.429218,9.728357,10.025683,9.56519,9.104698,8.644206,8.185526,7.7250338,7.9226465,8.120259,8.317872,8.515485,8.713099,8.627889,8.54268,8.457471,8.372261,8.287052,7.842876,7.3968873,6.9527116,6.506723,6.0625467,6.209397,6.35806,6.5049095,6.6517596,6.8004227,7.690587,8.580752,9.470917,10.359268,11.249433,10.5695715,9.88971,9.20985,8.529989,7.850128,7.851941,7.855567,7.85738,7.859193,7.8628187,8.470161,9.077503,9.684846,10.292189,10.899531,14.601601,18.305483,22.007553,25.709621,29.411692,23.61565,17.817797,12.019942,6.2220874,0.42423326,0.34083697,0.25562772,0.17041849,0.08520924,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06164073,0.12509441,0.18673515,0.25018883,0.31182957,0.8974165,1.4830034,2.0667772,2.6523643,3.2379513,2.6251698,2.0123885,1.3996071,0.7868258,0.17585737,0.13959812,0.10515183,0.07070554,0.034446288,0.0,0.0,0.0,0.0,0.0,0.0,0.059827764,0.11965553,0.1794833,0.23931105,0.2991388,0.2520018,0.20486477,0.15772775,0.11059072,0.06164073,0.28463513,0.5076295,0.7306239,0.95180535,1.1747998,1.9507477,2.7248828,3.5008307,4.274966,5.049101,5.6074934,6.165886,6.722465,7.2808576,7.837437,7.4422116,7.0469856,6.6517596,6.258347,5.863121,5.6256227,5.388125,5.1506267,4.9131284,4.6756306,6.200332,7.7250338,9.249735,10.774437,12.299138,12.368031,12.43511,12.50219,12.569269,12.638163,12.456866,12.277383,12.097899,11.916603,11.73712,11.809638,11.882156,11.954676,12.027194,12.099712,11.885782,11.67004,11.454298,11.240368,11.024626,11.127964,11.22949,11.332829,11.434355,11.537694,11.262123,10.988366,10.712796,10.437225,10.161655,10.607644,11.05182,11.497808,11.941984,12.387974,13.475751,14.561715,15.649493,16.73727,17.825048,18.122374,18.4197,18.717026,19.01435,19.311678,18.07705,16.842422,15.607795,14.373167,13.136727,13.60991,14.083094,14.554463,15.027647,15.50083,16.764465,18.029913,19.29536,20.560808,21.824444,22.429974,23.035503,23.63922,24.24475,24.850279,26.73576,28.619427,30.504908,32.39039,34.27587,34.3502,34.424534,34.50068,34.57501,34.64934,32.765675,30.880192,28.99471,27.10923,25.225561,24.824896,24.424232,24.025381,23.624716,23.225864,25.584528,27.945005,30.305483,32.664146,35.024624,36.5457,38.06496,39.584225,41.1053,42.624565,42.794983,42.9654,43.13582,43.304424,43.474842,44.31062,45.14458,45.98036,46.81432,47.650097,43.449463,39.25064,35.050007,30.849371,26.65055,25.299892,23.949236,22.600391,21.249735,19.90089,17.730774,15.5606575,13.390542,11.220426,9.050309,8.047741,7.0451727,6.0426044,5.040036,4.0374675,3.7129474,3.386614,3.0620937,2.7375734,2.4130533,2.565342,2.7176309,2.8699198,3.0222087,3.1744974,3.4119956,3.6494937,3.8869917,4.12449,4.361988,3.5806012,2.7974012,2.0142014,1.2328146,0.44961473,1.0551442,1.6606737,2.2643902,2.8699198,3.4754493,2.7992141,2.124792,1.4503701,0.774135,0.099712946,1.6008459,3.100166,4.599486,6.1006193,7.5999393,6.9019485,6.205771,5.5077806,4.8097897,4.1117992,4.900438,5.6872635,6.4759026,7.262728,8.049554,8.814624,9.579695,10.344765,11.109835,11.874905,11.22949,10.585889,9.940474,9.295059,8.649645,7.4277077,6.205771,4.9820213,3.7600844,2.5381477,2.72307,2.907992,3.092914,3.2778363,3.4627585,4.41819,5.371808,6.3272395,7.2826705,8.238102,8.858135,9.4781685,10.098202,10.718235,11.338268,11.030065,10.721861,10.41547,10.107266,9.800876,11.010121,12.219368,13.430427,14.639673,15.850732,14.71763,13.584529,12.45324,11.320138,10.1870365,10.020245,9.851639,9.684846,9.518054,9.349448,9.0956335,8.840006,8.584378,8.330563,8.074935,7.552802,7.0306687,6.506723,5.9845896,5.462456,5.282973,5.101677,4.9221935,4.74271,4.5632267,4.082792,3.6023567,3.1219215,2.6432993,2.1628644,1.8999848,1.6371052,1.3742256,1.1131591,0.85027945,0.7197462,0.58921283,0.4604925,0.32995918,0.19942589,0.17585737,0.15047589,0.12509441,0.099712946,0.07433146,0.80495536,1.5355793,2.2643902,2.9950142,3.7256382,3.4283123,3.1291735,2.8318477,2.5345216,2.2371957,2.0178273,1.7966459,1.5772774,1.357909,1.1367276,1.1022812,1.067835,1.0333886,0.99712944,0.96268314,0.8520924,0.7433147,0.6327239,0.52213323,0.41335547,0.35171473,0.291887,0.23205921,0.17223145,0.11240368,0.5094425,0.90829426,1.305333,1.7023718,2.0994108,1.8292793,1.5591478,1.2908293,1.020698,0.7505665,0.6000906,0.44961473,0.2991388,0.15047589,0.0,0.16679256,0.33539808,0.50219065,0.67079616,0.8375887,0.72337204,0.6073425,0.49312583,0.3770962,0.26287958,0.21030366,0.15772775,0.10515183,0.052575916,0.0,0.3045777,0.6091554,0.9155461,1.2201238,1.5247015,1.4503701,1.3742256,1.2998942,1.2255627,1.1494182,0.922798,0.69436467,0.46774435,0.23931105,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.452183,2.904366,4.358362,5.810545,7.262728,16.274965,25.287203,34.29944,43.313488,52.325726,42.07161,31.82112,21.567003,11.314699,1.062396,4.329355,7.5981264,10.865085,14.132043,17.400814,15.129172,12.859344,10.589515,8.319685,6.049856,5.9483304,5.844991,5.7416525,5.6401267,5.5367875,4.9294453,4.322103,3.7147603,3.1074178,2.5000753,2.1628644,1.8256533,1.4866294,1.1494182,0.8122072,0.9898776,1.167548,1.3452182,1.5228885,1.7005589,1.9670644,2.2353828,2.5018883,2.770207,3.0367124,2.4493124,1.8619126,1.2745126,0.6871128,0.099712946,0.11059072,0.11965553,0.13053331,0.13959812,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.052575916,0.054388877,0.058014803,0.059827764,0.06164073,0.08339628,0.10333887,0.12328146,0.14322405,0.16316663,0.15772775,0.15228885,0.14684997,0.14322405,0.13778515,0.13415924,0.13234627,0.13053331,0.12690738,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.14322405,0.15954071,0.17767033,0.19579996,0.21211663,0.21574254,0.21755551,0.21936847,0.2229944,0.22480737,0.2229944,0.21936847,0.21755551,0.21574254,0.21211663,0.19579996,0.17767033,0.15954071,0.14322405,0.12509441,0.11421664,0.10515183,0.09427405,0.08520924,0.07433146,5.411693,5.3083544,5.2032027,5.0980506,4.992899,4.8877473,5.40988,5.9320135,6.454147,6.978093,7.500226,7.7903004,8.080374,8.370448,8.660522,8.950596,9.03218,9.115576,9.197159,9.280556,9.362139,9.079316,8.798307,8.515485,8.232663,7.949841,8.056806,8.165584,8.272549,8.379513,8.488291,8.568061,8.647832,8.727602,8.807372,8.887142,8.323311,7.757667,7.192023,6.628191,6.0625467,6.281915,6.5030966,6.722465,6.9418335,7.1630154,8.067683,8.972352,9.87702,10.781689,11.6881695,11.05182,10.417283,9.782746,9.14821,8.511859,8.354132,8.198216,8.040489,7.8827615,7.7250338,9.151835,10.58045,12.007251,13.435865,14.862667,16.467138,18.071611,19.677896,21.282368,22.886839,18.479528,14.072216,9.664904,5.2575917,0.85027945,0.67986095,0.5094425,0.34083697,0.17041849,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06164073,0.12509441,0.18673515,0.25018883,0.31182957,0.9445535,1.5772774,2.2100015,2.8427253,3.4754493,2.811905,2.1501737,1.4866294,0.824898,0.16316663,0.13053331,0.09789998,0.065266654,0.032633327,0.0,0.0,0.0,0.0,0.0,0.0,0.045324065,0.09064813,0.13415924,0.1794833,0.22480737,0.19217403,0.15954071,0.12690738,0.09427405,0.06164073,0.2574407,0.45324063,0.64722764,0.8430276,1.0370146,1.9996977,2.962381,3.925064,4.8877473,5.8504305,6.153195,6.454147,6.7569118,7.059676,7.362441,7.1104393,6.8566246,6.604623,6.352621,6.1006193,5.712645,5.3246713,4.936697,4.550536,4.162562,5.600241,7.037921,8.4756,9.91328,11.349146,11.5231905,11.695421,11.867653,12.039885,12.212116,12.19036,12.166792,12.145037,12.123281,12.099712,12.494938,12.890164,13.28539,13.680615,14.075842,13.98338,13.89092,13.796645,13.704185,13.611723,13.229188,12.846653,12.464118,12.083396,11.700861,11.575767,11.450671,11.325577,11.200482,11.075388,11.952863,12.830337,13.70781,14.585284,15.462758,15.975826,16.487082,17.00015,17.513218,18.024473,18.220274,18.41426,18.610062,18.80586,18.999847,18.104244,17.210453,16.31485,15.419247,14.525456,14.882609,15.239763,15.596917,15.955884,16.313038,17.64194,18.972654,20.303368,21.632269,22.962984,23.535881,24.106964,24.67986,25.252756,25.825651,27.370296,28.91494,30.459585,32.004227,33.550686,33.586945,33.625015,33.66309,33.69935,33.73742,32.2798,30.822176,29.364555,27.906933,26.44931,25.812962,25.174799,24.536636,23.900286,23.262123,25.220123,27.178122,29.134308,31.092308,33.05031,34.839703,36.629097,38.420303,40.209698,42.000904,42.165882,42.330864,42.495842,42.660824,42.8258,43.92083,45.01586,46.11089,47.20592,48.299137,44.350502,40.40006,36.44961,32.49917,28.550535,26.98776,25.424988,23.862213,22.29944,20.736666,18.648132,16.557787,14.467442,12.377095,10.28675,9.182655,8.076748,6.972654,5.866747,4.762653,4.7753434,4.788034,4.800725,4.8134155,4.8242936,4.7916603,4.76084,4.7282066,4.695573,4.6629395,4.512464,4.361988,4.213325,4.062849,3.9123733,3.198066,2.4819458,1.7676386,1.0533313,0.33721104,1.3343405,2.333283,3.3304121,4.327542,5.3246713,4.3003473,3.2742105,2.2498865,1.2255627,0.19942589,1.5881553,2.9750717,4.361988,5.750717,7.137634,6.630004,6.1223745,5.614745,5.1071157,4.599486,5.2122674,5.825049,6.43783,7.0506115,7.663393,8.241728,8.821876,9.402024,9.982172,10.56232,10.13446,9.706602,9.280556,8.852696,8.424837,7.567306,6.7097745,5.8522434,4.994712,4.137181,4.3946214,4.652062,4.9095025,5.1669436,5.424384,6.285541,7.1448855,8.00423,8.865387,9.724731,9.815379,9.904215,9.994863,10.085511,10.174346,9.759177,9.345822,8.930654,8.515485,8.100317,9.333132,10.564133,11.7969475,13.029762,14.262577,13.147605,12.032633,10.917661,9.802689,8.6877165,8.540867,8.392203,8.245354,8.096691,7.949841,7.665206,7.380571,7.0941224,6.8094873,6.5248523,6.2547207,5.9845896,5.714458,5.4443264,5.1741953,5.0527267,4.9294453,4.8079767,4.6846952,4.5632267,4.064662,3.5679104,3.0693457,2.572594,2.0758421,1.8383441,1.6008459,1.3633479,1.1258497,0.8883517,0.7523795,0.61822027,0.48224804,0.3480888,0.21211663,0.19942589,0.18673515,0.17585737,0.16316663,0.15047589,0.96087015,1.7694515,2.5798457,3.39024,4.2006345,4.0918565,3.9848917,3.877927,3.7691493,3.6621845,3.3231604,2.9823234,2.6432993,2.3024626,1.9616255,1.9181144,1.8727903,1.8274662,1.7821422,1.7368182,1.4666867,1.1983683,0.92823684,0.65810543,0.387974,0.32995918,0.27194437,0.21574254,0.15772775,0.099712946,0.40791658,0.71430725,1.0225109,1.3307146,1.6371052,1.4231756,1.2074331,0.9916905,0.7777609,0.5620184,0.44961473,0.33721104,0.22480737,0.11240368,0.0,0.13415924,0.27013144,0.40429065,0.5402629,0.6744221,0.5946517,0.5148814,0.43511102,0.35534066,0.2755703,0.21936847,0.16497959,0.11059072,0.054388877,0.0,0.23568514,0.46955732,0.70524246,0.93911463,1.1747998,1.1131591,1.0497054,0.9880646,0.9246109,0.8629702,0.69436467,0.5275721,0.36077955,0.19217403,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.1167849,2.2353828,3.3521678,4.4707656,5.5875506,12.676234,19.763105,26.849976,33.936848,41.02553,33.032177,25.04064,17.047287,9.055748,1.062396,3.834416,6.6082487,9.380268,12.152288,14.924308,12.872034,10.81976,8.767487,6.7152133,4.6629395,5.3446136,6.0281005,6.7097745,7.3932614,8.074935,6.834869,5.5948024,4.3547363,3.1146698,1.8746033,1.8002719,1.7241274,1.649796,1.5754645,1.49932,1.8673514,2.2353828,2.6034143,2.9696326,3.3376641,3.147303,2.956942,2.7683938,2.5780327,2.3876717,1.9253663,1.4630609,1.0007553,0.53663695,0.07433146,0.08339628,0.09064813,0.09789998,0.10515183,0.11240368,0.09064813,0.06707962,0.045324065,0.02175555,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.04169814,0.047137026,0.052575916,0.058014803,0.06164073,0.07795739,0.092461094,0.10696479,0.12328146,0.13778515,0.13959812,0.14322405,0.14503701,0.14684997,0.15047589,0.14503701,0.13959812,0.13415924,0.13053331,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.13415924,0.14503701,0.15410182,0.16497959,0.17585737,0.1794833,0.18492219,0.19036107,0.19579996,0.19942589,0.19579996,0.19036107,0.18492219,0.1794833,0.17585737,0.16497959,0.15410182,0.14503701,0.13415924,0.12509441,0.11784257,0.11059072,0.10333887,0.09427405,0.0870222,4.9620786,4.9058766,4.847862,4.7898474,4.7318325,4.6756306,5.239462,5.805106,6.3707504,6.9345818,7.500226,7.8718834,8.245354,8.617011,8.990481,9.362139,9.229793,9.097446,8.9651,8.832754,8.700407,8.595256,8.490104,8.384952,8.2798,8.174648,8.192778,8.209095,8.227224,8.245354,8.26167,8.508233,8.752983,8.997733,9.242483,9.487233,8.801933,8.116633,7.4331465,6.7478466,6.0625467,6.354434,6.6481338,6.9400206,7.231908,7.5256076,8.444779,9.365765,10.284937,11.204109,12.125093,11.535881,10.944855,10.355642,9.764616,9.175404,8.858135,8.540867,8.221786,7.9045167,7.5872483,9.835322,12.081583,14.329657,16.57773,18.825804,18.332678,17.839552,17.34824,16.855114,16.361988,13.345218,10.328448,7.309865,4.2930956,1.2745126,1.020698,0.7650702,0.5094425,0.25562772,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06164073,0.12509441,0.18673515,0.25018883,0.31182957,0.9916905,1.6733645,2.3532255,3.0330863,3.7129474,3.000453,2.2879589,1.5754645,0.8629702,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.0,0.0,0.0,0.0,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.13234627,0.11421664,0.09789998,0.07977036,0.06164073,0.23024625,0.39703882,0.5656443,0.7324369,0.89922947,2.0504606,3.199879,4.349297,5.5005283,6.6499467,6.697084,6.7442207,6.793171,6.8403077,6.887445,6.776854,6.6680765,6.5574856,6.446895,6.338117,5.7996674,5.2630305,4.7245803,4.1879435,3.6494937,5.0001507,6.350808,7.699652,9.050309,10.399154,10.6783495,10.955733,11.233116,11.510499,11.787883,11.922042,12.058014,12.192173,12.328146,12.462305,13.180238,13.898171,14.614291,15.332225,16.050158,16.079165,16.109985,16.140806,16.169813,16.200634,15.332225,14.465629,13.597219,12.730623,11.862214,11.887595,11.912977,11.938358,11.961927,11.9873085,13.29808,14.607039,15.917811,17.22677,18.537542,18.474089,18.412449,18.350807,18.287354,18.225714,18.318174,18.410635,18.503096,18.595556,18.688019,18.133251,17.576672,17.021906,16.467138,15.912373,16.15531,16.398247,16.63937,16.882307,17.125244,18.519413,19.915394,21.309563,22.705544,24.099712,24.639975,25.180237,25.7205,26.260763,26.799213,28.004833,29.210453,30.41426,31.61988,32.8255,32.8255,32.8255,32.8255,32.8255,32.8255,31.795738,30.764162,29.7344,28.704636,27.674873,26.799213,25.925365,25.049704,24.175856,23.300196,24.855717,26.409426,27.964949,29.52047,31.074179,33.135517,35.19504,37.25457,39.315907,41.37543,41.534973,41.694515,41.855865,42.015408,42.17495,43.529232,44.885326,46.23961,47.595707,48.94999,45.249733,41.549477,37.84922,34.150776,30.45052,28.675629,26.90074,25.124035,23.349146,21.574255,19.565493,17.554916,15.544341,13.535579,11.525003,10.31757,9.110137,7.902704,6.695271,5.487838,5.8377395,6.187641,6.5375433,6.887445,7.2373466,7.019791,6.8022356,6.58468,6.3671246,6.149569,5.612932,5.0744824,4.537845,3.9993954,3.4627585,2.8155308,2.1683033,1.5192627,0.872035,0.22480737,1.6153497,3.004079,4.3946214,5.7851634,7.175706,5.7996674,4.4254417,3.049403,1.6751775,0.2991388,1.5754645,2.8499773,4.12449,5.4008155,6.6753283,6.35806,6.0407915,5.7217097,5.4044414,5.087173,5.52591,5.962834,6.399758,6.836682,7.2754188,7.6706448,8.06587,8.459284,8.854509,9.249735,9.039432,8.829127,8.620637,8.410334,8.200029,7.706904,7.215591,6.722465,6.2293396,5.7380266,6.0679855,6.397945,6.7279043,7.057863,7.3878226,8.152893,8.917963,9.683033,10.448103,11.213174,10.772624,10.332074,9.893337,9.452786,9.012237,8.490104,7.9679704,7.4458375,6.921891,6.399758,7.654328,8.910711,10.165281,11.419851,12.674421,11.5775795,10.480737,9.382081,8.285239,7.1883965,7.059676,6.932769,6.8058615,6.677141,6.550234,6.2347784,5.919323,5.6056805,5.290225,4.974769,4.95664,4.940323,4.9221935,4.9058766,4.8877473,4.8224807,4.7572136,4.691947,4.6266804,4.5632267,4.0483456,3.531651,3.0167696,2.5018883,1.987007,1.7748904,1.5627737,1.3506571,1.1367276,0.9246109,0.7850128,0.64541465,0.5058166,0.36440548,0.22480737,0.22480737,0.22480737,0.22480737,0.22480737,0.22480737,1.114972,2.0051367,2.8953013,3.785466,4.6756306,4.7572136,4.84061,4.9221935,5.0055895,5.087173,4.6266804,4.168001,3.7075086,3.247016,2.7883365,2.7321346,2.6777458,2.6233568,2.5671551,2.5127661,2.0830941,1.651609,1.2219368,0.79226464,0.36259252,0.30820364,0.2520018,0.19761293,0.14322405,0.0870222,0.3045777,0.52213323,0.73968875,0.9572442,1.1747998,1.015259,0.8557183,0.69436467,0.53482395,0.37528324,0.2991388,0.22480737,0.15047589,0.07433146,0.0,0.10333887,0.20486477,0.30820364,0.40972954,0.51306844,0.46774435,0.4224203,0.3770962,0.33177215,0.28826106,0.23024625,0.17223145,0.11421664,0.058014803,0.0,0.16497959,0.32995918,0.4949388,0.65991837,0.824898,0.774135,0.72518504,0.6744221,0.62547207,0.5747091,0.46774435,0.36077955,0.2520018,0.14503701,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.78319985,1.5645868,2.3477864,3.1291735,3.9123733,9.07569,14.237195,19.400513,24.562017,29.725334,23.992746,18.260159,12.527572,6.794984,1.062396,3.339477,5.616558,7.895452,10.172533,12.449615,10.614896,8.780178,6.94546,5.1107416,3.2742105,4.74271,6.209397,7.6778965,9.144584,10.613083,8.740293,6.867502,4.994712,3.1219215,1.2491312,1.4376793,1.6244144,1.8129625,1.9996977,2.1882458,2.7448254,3.303218,3.8597972,4.41819,4.974769,4.327542,3.680314,3.0330863,2.3858588,1.7368182,1.3996071,1.062396,0.72518504,0.387974,0.05076295,0.054388877,0.059827764,0.065266654,0.07070554,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.032633327,0.03988518,0.047137026,0.054388877,0.06164073,0.072518505,0.08339628,0.092461094,0.10333887,0.11240368,0.12328146,0.13234627,0.14322405,0.15228885,0.16316663,0.15410182,0.14684997,0.13959812,0.13234627,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12690738,0.13053331,0.13234627,0.13415924,0.13778515,0.14503701,0.15228885,0.15954071,0.16679256,0.17585737,0.16679256,0.15954071,0.15228885,0.14503701,0.13778515,0.13415924,0.13234627,0.13053331,0.12690738,0.12509441,0.11965553,0.11421664,0.11059072,0.10515183,0.099712946,4.512464,4.503399,4.4925213,4.4816437,4.4725785,4.461701,5.0708566,5.678199,6.285541,6.892884,7.500226,7.95528,8.410334,8.865387,9.32044,9.775495,9.427405,9.079316,8.733041,8.384952,8.036863,8.109382,8.1819,8.254418,8.326937,8.399456,8.326937,8.254418,8.1819,8.109382,8.036863,8.446592,8.858135,9.267865,9.677594,10.087324,9.282369,8.477413,7.6724577,6.867502,6.0625467,6.4269524,6.793171,7.157576,7.5219817,7.8882003,8.821876,9.757364,10.692853,11.628342,12.562017,12.018129,11.472427,10.926725,10.382836,9.837135,9.360326,8.881703,8.404895,7.9280853,7.4494634,10.516996,13.584529,16.652061,19.719595,22.787127,20.198215,17.607492,15.016769,12.427858,9.837135,8.209095,6.582867,4.954827,3.3267863,1.7005589,1.3597219,1.020698,0.67986095,0.34083697,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06164073,0.12509441,0.18673515,0.25018883,0.31182957,1.0406405,1.7676386,2.4946365,3.2216346,3.9504454,3.1871881,2.4257438,1.6624867,0.89922947,0.13778515,0.11059072,0.08339628,0.054388877,0.027194439,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.072518505,0.07070554,0.06707962,0.065266654,0.06164073,0.2030518,0.34264994,0.48224804,0.62184614,0.76325727,2.0994108,3.437377,4.7753434,6.11331,7.4494634,7.2427855,7.0342946,6.827617,6.6191263,6.412449,6.445082,6.4777155,6.510349,6.542982,6.5756154,5.8866897,5.199577,4.512464,3.825351,3.1382382,4.40006,5.661882,6.925517,8.187339,9.449161,9.8316965,10.2142315,10.596766,10.979301,11.361836,11.655537,11.947423,12.23931,12.5330105,12.824898,13.865538,14.904366,15.945006,16.985647,18.024473,18.176764,18.330864,18.483154,18.635443,18.787731,17.43526,16.08279,14.730321,13.377851,12.025381,12.199425,12.375282,12.549327,12.725184,12.899229,14.643299,16.385555,18.127813,19.87007,21.612328,20.974165,20.337814,19.699652,19.063301,18.425138,18.41426,18.405195,18.394318,18.385254,18.374376,18.160446,17.944704,17.730774,17.515032,17.29929,17.428009,17.554916,17.681824,17.810545,17.937452,19.396887,20.858135,22.31757,23.777004,25.238253,25.745882,26.251698,26.759327,27.266956,27.774588,28.63937,29.504152,30.370749,31.235533,32.100315,32.062244,32.02417,31.987911,31.949839,31.911768,31.309864,30.70796,30.104244,29.50234,28.900436,27.787277,26.675932,25.562773,24.449614,23.338266,24.489498,25.642542,26.795588,27.946817,29.099863,31.42952,33.759174,36.090645,38.420303,40.74996,40.905876,41.059975,41.215893,41.36999,41.524094,43.139446,44.754795,46.370144,47.985493,49.60084,46.150776,42.700706,39.25064,35.80057,32.350506,30.361685,28.374678,26.38767,24.400663,22.411844,20.482851,18.552046,16.623055,14.692248,12.763257,11.452485,10.141713,8.832754,7.5219817,6.2130227,6.9001355,7.5872483,8.274362,8.963287,9.6504,9.247922,8.845445,8.442966,8.040489,7.6380115,6.7134004,5.7869763,4.8623657,3.9377546,3.0131438,2.4329958,1.8528478,1.2726997,0.69255173,0.11240368,1.8945459,3.6766882,5.4606433,7.2427855,9.024928,7.3008003,5.57486,3.8507326,2.124792,0.40066472,1.5627737,2.7248828,3.8869917,5.050914,6.2130227,6.0843024,5.957395,5.8304877,5.7017674,5.57486,5.8377395,6.1006193,6.3616858,6.624565,6.887445,7.0977483,7.308052,7.518356,7.7268467,7.93715,7.944402,7.951654,7.9607186,7.9679704,7.9752226,7.8483152,7.7195945,7.592687,7.46578,7.3370595,7.7395372,8.1420145,8.544493,8.94697,9.349448,10.020245,10.689227,11.3600235,12.03082,12.699803,11.729868,10.7599325,9.789998,8.820063,7.850128,7.219217,6.590119,5.959208,5.33011,4.699199,5.977338,7.2554765,8.531802,9.80994,11.088079,10.007553,8.927028,7.8483152,6.7677894,5.6872635,5.580299,5.473334,5.3645563,5.2575917,5.1506267,4.804351,4.459888,4.115425,3.7691493,3.4246864,3.6603715,3.8942437,4.1299286,4.365614,4.599486,4.592234,4.5849824,4.5777307,4.5704784,4.5632267,4.0302157,3.4972048,2.9641938,2.4329958,1.8999848,1.7132497,1.5247015,1.3379664,1.1494182,0.96268314,0.81764615,0.6726091,0.5275721,0.3825351,0.2374981,0.25018883,0.26287958,0.2755703,0.28826106,0.2991388,1.2708868,2.2408218,3.2107568,4.1806917,5.1506267,5.422571,5.6945157,5.9682727,6.240217,6.5121617,5.9320135,5.351866,4.7717175,4.1933823,3.6132345,3.5479677,3.482701,3.4174345,3.3521678,3.2869012,2.6976883,2.1066625,1.5174497,0.92823684,0.33721104,0.28463513,0.23205921,0.1794833,0.12690738,0.07433146,0.2030518,0.32995918,0.45686656,0.5855869,0.7124943,0.6073425,0.50219065,0.39703882,0.291887,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.07070554,0.13959812,0.21030366,0.27919623,0.34990177,0.34083697,0.32995918,0.3208944,0.3100166,0.2991388,0.23931105,0.1794833,0.11965553,0.059827764,0.0,0.09427405,0.19036107,0.28463513,0.38072214,0.4749962,0.43692398,0.40066472,0.36259252,0.3245203,0.28826106,0.23931105,0.19217403,0.14503701,0.09789998,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.44780177,0.89560354,1.3415923,1.789394,2.2371957,5.475147,8.713099,11.949236,15.187187,18.425138,14.951503,11.479679,8.007855,4.5342193,1.062396,2.8445382,4.6266804,6.4106355,8.192778,9.97492,8.357758,6.740595,5.121619,3.5044568,1.887294,4.1408067,6.392506,8.644206,10.897718,13.149418,10.645717,8.140202,5.634688,3.1291735,0.62547207,1.0750868,1.5247015,1.9743162,2.4257438,2.8753586,3.6222992,4.36924,5.1179934,5.864934,6.6118746,5.5077806,4.401873,3.2977788,2.1918716,1.0877775,0.87566096,0.66173136,0.44961473,0.2374981,0.025381476,0.027194439,0.030820364,0.032633327,0.034446288,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.02175555,0.032633327,0.04169814,0.052575916,0.06164073,0.06707962,0.072518505,0.07795739,0.08339628,0.0870222,0.10515183,0.12328146,0.13959812,0.15772775,0.17585737,0.16497959,0.15410182,0.14503701,0.13415924,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.11965553,0.11421664,0.11059072,0.10515183,0.099712946,0.11059072,0.11965553,0.13053331,0.13959812,0.15047589,0.13959812,0.13053331,0.11965553,0.11059072,0.099712946,0.10515183,0.11059072,0.11421664,0.11965553,0.12509441,0.12328146,0.11965553,0.11784257,0.11421664,0.11240368,4.062849,4.099108,4.137181,4.175253,4.213325,4.249584,4.900438,5.5494785,6.200332,6.849373,7.500226,8.036863,8.575313,9.11195,9.6504,10.1870365,9.625018,9.063,8.499168,7.93715,7.3751316,7.6253204,7.8755093,8.125698,8.375887,8.624263,8.46291,8.299743,8.138389,7.9752226,7.8120556,8.386765,8.963287,9.537996,10.112705,10.687414,9.762803,8.838193,7.911769,6.987158,6.0625467,6.4994707,6.9382076,7.3751316,7.8120556,8.2507925,9.200785,10.150778,11.10077,12.050762,13.000754,12.500377,11.999999,11.499621,10.999244,10.500679,9.862516,9.224354,8.588004,7.949841,7.311678,11.200482,15.087475,18.974466,22.863272,26.750263,22.061941,17.375433,12.687112,8.000604,3.3122826,3.0747845,2.8372865,2.5997884,2.3622901,2.124792,1.7005589,1.2745126,0.85027945,0.42423326,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06164073,0.12509441,0.18673515,0.25018883,0.31182957,1.0877775,1.8619126,2.6378605,3.4119956,4.1879435,3.3757362,2.561716,1.7495089,0.93730164,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.17585737,0.28826106,0.40066472,0.51306844,0.62547207,2.1501737,3.6748753,5.199577,6.7242785,8.2507925,7.7866745,7.324369,6.8620634,6.399758,5.9374523,6.11331,6.2873545,6.4632115,6.637256,6.813113,5.975525,5.137936,4.3003473,3.4627585,2.6251698,3.7999697,4.974769,6.149569,7.324369,8.499168,8.9868555,9.474543,9.96223,10.449916,10.937603,11.3872175,11.836833,12.28826,12.737875,13.1874895,14.5508375,15.912373,17.27572,18.637255,20.000603,20.27436,20.54993,20.8255,21.099258,21.374828,19.538298,17.699953,15.861609,14.025079,12.186734,12.513068,12.837588,13.162108,13.486629,13.812962,15.986704,18.16226,20.337814,22.513369,24.68711,23.47424,22.26318,21.050308,19.837437,18.624565,18.512161,18.399757,18.287354,18.17495,18.062546,18.187641,18.312735,18.43783,18.562923,18.688019,18.700708,18.7134,18.724277,18.736969,18.749659,20.27436,21.799063,23.325577,24.850279,26.374979,26.849976,27.324972,27.799969,28.274965,28.74996,29.27572,29.799665,30.325424,30.849371,31.37513,31.300798,31.224655,31.150324,31.074179,30.999847,30.825802,30.649946,30.4759,30.300043,30.124186,28.775343,27.424685,26.07584,24.725183,23.374527,24.125093,24.87566,25.624413,26.374979,27.125546,29.725334,32.325123,34.92491,37.5247,40.12449,40.274963,40.425438,40.574104,40.72458,40.875053,42.749657,44.62426,46.50068,48.375282,50.249886,47.050003,43.850124,40.650246,37.450367,34.25049,32.049553,29.85043,27.649492,25.450369,23.249432,21.40021,19.549175,17.699953,15.850732,13.999697,12.5873995,11.175101,9.762803,8.350506,6.9382076,7.9625316,8.9868555,10.012992,11.037316,12.06164,11.47424,10.88684,10.29944,9.712041,9.12464,7.8120556,6.4994707,5.186886,3.874301,2.561716,2.0504606,1.5373923,1.0243238,0.51306844,0.0,2.175555,4.349297,6.5248523,8.700407,10.874149,8.80012,6.7242785,4.650249,2.5744069,0.50037766,1.550083,2.5997884,3.6494937,4.699199,5.750717,5.812358,5.8758116,5.9374523,6.000906,6.0625467,6.149569,6.2365913,6.3254266,6.412449,6.4994707,6.5248523,6.550234,6.5756154,6.599184,6.624565,6.849373,7.07418,7.3008003,7.5256076,7.750415,7.987913,8.225411,8.46291,8.700407,8.937905,9.412902,9.8878975,10.362894,10.837891,11.312886,11.887595,12.462305,13.037014,13.611723,14.188245,12.687112,11.187792,9.686659,8.187339,6.688019,5.9501433,5.2122674,4.4743915,3.738329,3.000453,4.3003473,5.600241,6.9001355,8.200029,9.499924,8.437528,7.3751316,6.3127356,5.2503395,4.1879435,4.099108,4.0120864,3.925064,3.8380418,3.7492065,3.3757362,3.000453,2.6251698,2.2498865,1.8746033,2.3622901,2.8499773,3.3376641,3.825351,4.313038,4.361988,4.4127507,4.461701,4.512464,4.5632267,4.0120864,3.4627585,2.911618,2.3622901,1.8129625,1.649796,1.4866294,1.3252757,1.162109,1.0007553,0.85027945,0.69980353,0.5493277,0.40066472,0.25018883,0.2755703,0.2991388,0.3245203,0.34990177,0.37528324,1.4249886,2.474694,3.5243993,4.5759177,5.6256227,6.0879283,6.550234,7.0125394,7.474845,7.93715,7.2373466,6.5375433,5.8377395,5.137936,4.4381323,4.361988,4.2876563,4.213325,4.137181,4.062849,3.3122826,2.561716,1.8129625,1.062396,0.31182957,0.26287958,0.21211663,0.16316663,0.11240368,0.06164073,0.099712946,0.13778515,0.17585737,0.21211663,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.0,0.0,0.0,0.0,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.21211663,0.2374981,0.26287958,0.28826106,0.31182957,0.25018883,0.18673515,0.12509441,0.06164073,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.11240368,0.22480737,0.33721104,0.44961473,0.5620184,1.8746033,3.1871881,4.499773,5.812358,7.124943,5.9120708,4.699199,3.48814,2.275268,1.062396,2.3495996,3.636803,4.9258194,6.2130227,7.500226,6.1006193,4.699199,3.299592,1.8999848,0.50037766,3.53709,6.5756154,9.612328,12.650853,15.687565,12.549327,9.412902,6.2746634,3.1382382,0.0,0.7124943,1.4249886,2.137483,2.8499773,3.5624714,4.499773,5.4370747,6.3743763,7.311678,8.2507925,6.688019,5.125245,3.5624714,1.9996977,0.43692398,0.34990177,0.26287958,0.17585737,0.0870222,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.0870222,0.11240368,0.13778515,0.16316663,0.18673515,0.17585737,0.16316663,0.15047589,0.13778515,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,4.249584,4.2930956,4.3347936,4.3783045,4.420003,4.461701,5.0055895,5.5476656,6.089741,6.6318173,7.175706,7.665206,8.154706,8.644206,9.135518,9.625018,9.14821,8.669587,8.192778,7.7141557,7.2373466,7.507478,7.7776093,8.047741,8.317872,8.588004,8.3051815,8.02236,7.7395372,7.456715,7.175706,7.799365,8.424837,9.050309,9.675781,10.29944,9.479981,8.660522,7.83925,7.019791,6.200332,6.834869,7.4694057,8.105756,8.740293,9.374829,10.107266,10.839704,11.57214,12.304577,13.037014,12.407916,11.777005,11.147907,10.516996,9.8878975,9.606889,9.327692,9.046683,8.767487,8.488291,12.092461,15.6966305,19.302612,22.906782,26.512764,21.770054,17.027344,12.284635,7.5419245,2.7992141,2.5798457,2.3604772,2.1392958,1.9199274,1.7005589,1.3597219,1.020698,0.67986095,0.34083697,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07070554,0.13959812,0.21030366,0.27919623,0.34990177,1.2074331,2.0649643,2.9224956,3.780027,4.6375585,3.729264,2.8227828,1.9144884,1.0080072,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0,0.0,0.0,0.0,0.0,0.09064813,0.1794833,0.27013144,0.36077955,0.44961473,0.56020546,0.67079616,0.7795739,0.8901646,1.0007553,1.3071461,1.6153497,1.9217403,2.229944,2.5381477,3.8126602,5.087173,6.3616858,7.6380115,8.912524,8.299743,7.686961,7.07418,6.4632115,5.8504305,6.0480433,6.245656,6.4432693,6.640882,6.836682,6.300045,5.763408,5.224958,4.688321,4.1498713,5.2521524,6.354434,7.456715,8.560809,9.663091,10.012992,10.362894,10.712796,11.062697,11.4126,11.938358,12.462305,12.988064,13.512011,14.037769,15.089288,16.142618,17.194138,18.247469,19.3008,19.50929,19.719595,19.929897,20.140202,20.350506,18.961775,17.57486,16.187943,14.799213,13.412297,13.589968,13.767638,13.945308,14.122978,14.300649,15.970387,17.640125,19.309864,20.979603,22.649342,21.708414,20.765673,19.822933,18.880192,17.937452,17.837738,17.738026,17.638313,17.536787,17.437075,17.870373,18.301857,18.735155,19.166641,19.59994,20.250792,20.899832,21.550686,22.199726,22.85058,24.126905,25.405045,26.683184,27.959509,29.237648,29.382685,29.527721,29.672758,29.817795,29.962833,30.394318,30.827616,31.260914,31.692398,32.125698,32.093063,32.06043,32.027798,31.995163,31.96253,31.750414,31.538298,31.324368,31.112251,30.900135,29.598427,28.294907,26.9932,25.68968,24.387972,25.060581,25.73319,26.4058,27.07841,27.749205,29.721708,31.694212,33.666714,35.639217,37.61172,37.727753,37.84197,37.957996,38.072216,38.188244,40.3076,42.42695,44.548115,46.66747,48.786823,45.93322,43.077805,40.22239,37.36697,34.51337,32.471973,30.43239,28.392807,26.353224,24.311829,22.323008,20.332375,18.341742,16.352922,14.362289,13.1874895,12.012691,10.837891,9.663091,8.488291,9.211663,9.936848,10.662033,11.3872175,12.112403,11.418038,10.721861,10.027496,9.333132,8.636953,7.454902,6.2728505,5.090799,3.9069343,2.7248828,2.179181,1.6352923,1.0895905,0.54570174,0.0,1.9017978,3.8054085,5.7072062,7.610817,9.512614,7.7195945,5.9283876,4.135368,2.3423476,0.5493277,1.5301404,2.5091403,3.489953,4.4707656,5.4497657,5.42801,5.4044414,5.382686,5.3591175,5.337362,5.431636,5.527723,5.621997,5.718084,5.812358,5.8794374,5.9483304,6.01541,6.0824895,6.149569,6.338117,6.5248523,6.7134004,6.9001355,7.0868707,7.2844834,7.4820967,7.6797094,7.877322,8.074935,8.343254,8.609759,8.8780775,9.144584,9.412902,10.002114,10.593141,11.182353,11.773379,12.362592,11.129777,9.896963,8.664148,7.4331465,6.200332,5.710832,5.219519,4.7300196,4.2405195,3.7492065,4.597673,5.4443264,6.2927933,7.1394467,7.987913,7.063302,6.1368785,5.2122674,4.2876563,3.3630457,3.290527,3.2180085,3.1454902,3.0729716,3.000453,2.70494,2.4094272,2.1157274,1.8202144,1.5247015,1.9199274,2.3151531,2.7103791,3.105605,3.5008307,3.673062,3.8452935,4.017525,4.1897564,4.361988,4.1970086,4.0320287,3.8670492,3.7020695,3.53709,3.2343252,2.9333735,2.6306088,2.327844,2.0250793,1.6896812,1.3542831,1.020698,0.6852999,0.34990177,0.6345369,0.91917205,1.2056202,1.4902552,1.7748904,2.617918,3.4591327,4.3021603,5.145188,5.9882154,6.0843024,6.1822023,6.2801023,6.378002,6.474089,6.0770507,5.6800117,5.282973,4.8841214,4.4870825,4.49796,4.507025,4.517903,4.5269675,4.537845,3.7999697,3.0620937,2.324218,1.5881553,0.85027945,0.69073874,0.5293851,0.36984438,0.21030366,0.05076295,0.09427405,0.13959812,0.18492219,0.23024625,0.2755703,0.23024625,0.18492219,0.13959812,0.09427405,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.17585737,0.19942589,0.22480737,0.25018883,0.2755703,0.2229944,0.17041849,0.11784257,0.065266654,0.012690738,0.034446288,0.058014803,0.07977036,0.10333887,0.12509441,0.11784257,0.11059072,0.10333887,0.09427405,0.0870222,0.07977036,0.072518505,0.065266654,0.058014803,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.09064813,0.1794833,0.27013144,0.36077955,0.44961473,1.49932,2.5508385,3.6005437,4.650249,5.6999545,4.76084,3.8199122,2.8807976,1.93987,1.0007553,2.5073273,4.0157123,5.522284,7.0306687,8.537241,6.9092,5.282973,3.6549325,2.0268922,0.40066472,2.8300345,5.2594047,7.690587,10.119957,12.549327,10.040187,7.5292335,5.0200934,2.5091403,0.0,0.6000906,1.2001812,1.8002719,2.4003625,3.000453,3.7945306,4.590421,5.384499,6.1803894,6.9744673,5.6491914,4.325729,3.000453,1.6751775,0.34990177,0.27919623,0.21030366,0.13959812,0.07070554,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.01994259,0.027194439,0.034446288,0.04169814,0.05076295,0.054388877,0.059827764,0.065266654,0.07070554,0.07433146,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.06707962,0.072518505,0.07795739,0.08339628,0.0870222,0.10515183,0.12328146,0.13959812,0.15772775,0.17585737,0.16679256,0.15954071,0.15228885,0.14503701,0.13778515,0.13415924,0.13234627,0.13053331,0.12690738,0.12509441,0.11421664,0.10515183,0.09427405,0.08520924,0.07433146,0.07977036,0.08520924,0.09064813,0.09427405,0.099712946,0.09064813,0.07977036,0.07070554,0.059827764,0.05076295,0.059827764,0.07070554,0.07977036,0.09064813,0.099712946,0.099712946,0.099712946,0.099712946,0.099712946,0.099712946,4.4381323,4.4852695,4.5324063,4.5795436,4.6266804,4.6756306,5.1107416,5.5458527,5.979151,6.414262,6.849373,7.2917356,7.7340984,8.178274,8.620637,9.063,8.669587,8.2779875,7.8845744,7.4929743,7.0995617,7.3896356,7.6797094,7.9697833,8.259857,8.549932,8.147454,7.744976,7.3424983,6.9400206,6.5375433,7.211965,7.8882003,8.562622,9.237044,9.91328,9.197159,8.482852,7.7667317,7.0524244,6.338117,7.170267,8.002417,8.834567,9.666717,10.500679,11.015561,11.530442,12.045323,12.5602045,13.075087,12.3154545,11.555823,10.794379,10.034748,9.275117,9.353074,9.429218,9.507175,9.585134,9.663091,12.984438,16.307598,19.630758,22.952106,26.275267,21.478168,16.679256,11.882156,7.0850577,2.2879589,2.084907,1.8818551,1.6806163,1.4775645,1.2745126,1.020698,0.7650702,0.5094425,0.25562772,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07795739,0.15410182,0.23205921,0.3100166,0.387974,1.3270886,2.268016,3.207131,4.1480584,5.087173,4.0846047,3.0820365,2.079468,1.0768998,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.1794833,0.36077955,0.5402629,0.7197462,0.89922947,1.1077201,1.3143979,1.5228885,1.7295663,1.938057,2.4402475,2.9424384,3.444629,3.9468195,4.4508233,5.475147,6.4994707,7.5256076,8.549932,9.574255,8.812811,8.049554,7.28811,6.5248523,5.7615952,5.9827766,6.202145,6.4233265,6.642695,6.8620634,6.624565,6.3870673,6.149569,5.9120708,5.674573,6.7043357,7.7340984,8.765674,9.795437,10.825199,11.037316,11.249433,11.463363,11.675479,11.887595,12.487686,13.087777,13.687867,14.287958,14.888049,15.62955,16.372866,17.114367,17.857681,18.599184,18.74422,18.889257,19.034294,19.17933,19.324368,18.387066,17.449764,16.512463,15.575162,14.63786,14.666867,14.697688,14.726695,14.757515,14.788336,15.952258,17.117992,18.281914,19.447649,20.613384,19.940775,19.268166,18.595556,17.922949,17.25034,17.163317,17.074482,16.98746,16.900436,16.811602,17.553104,18.292793,19.03248,19.77217,20.511858,21.800875,23.088078,24.375282,25.662485,26.949688,27.979452,29.009214,30.04079,31.070553,32.100315,31.915394,31.73047,31.54555,31.360626,31.175705,31.514729,31.855566,32.194588,32.535427,32.87445,32.885326,32.894394,32.90527,32.914337,32.925213,32.675026,32.424835,32.17465,31.924458,31.674269,30.419699,29.165129,27.910559,26.654177,25.399607,25.994257,26.590723,27.185373,27.780025,28.374678,29.719896,31.065113,32.41033,33.75555,35.10077,35.18054,35.26031,35.34008,35.41985,35.49962,37.865536,40.22964,42.595554,44.95966,47.325577,44.81462,42.30548,39.79453,37.28539,34.774437,32.894394,31.01435,29.134308,27.254267,25.374224,23.245806,21.115576,18.985344,16.855114,14.724882,13.7875805,12.850279,11.912977,10.975676,10.038374,10.462607,10.88684,11.312886,11.73712,12.163166,11.3600235,10.556881,9.755551,8.952409,8.149267,7.0977483,6.0444174,4.992899,3.9395678,2.8880494,2.3097143,1.7331922,1.1548572,0.57833505,0.0,1.6298534,3.2597067,4.88956,6.5194135,8.149267,6.640882,5.130684,3.6204863,2.1102884,0.6000906,1.5101979,2.420305,3.3304121,4.2405195,5.1506267,5.041849,4.934884,4.8279195,4.7191415,4.612177,4.7155156,4.8170414,4.9203806,5.0219064,5.125245,5.235836,5.3446136,5.4552045,5.565795,5.674573,5.825049,5.975525,6.1241875,6.2746634,6.4251394,6.582867,6.740595,6.8983226,7.0542374,7.211965,7.271793,7.3316207,7.3932614,7.453089,7.512917,8.116633,8.722163,9.327692,9.933222,10.536939,9.572442,8.607946,7.6416373,6.677141,5.712645,5.469708,5.2267714,4.985647,4.74271,4.499773,4.894999,5.290225,5.6854506,6.0806766,6.474089,5.6872635,4.900438,4.1117992,3.3249733,2.5381477,2.4801328,2.422118,2.3641033,2.3079014,2.2498865,2.034144,1.8202144,1.6044719,1.3905423,1.1747998,1.4775645,1.7803292,2.0830941,2.3858588,2.6868105,2.9823234,3.2778363,3.5733492,3.8670492,4.162562,4.3819304,4.603112,4.8224807,5.041849,5.2630305,4.8206677,4.3783045,3.9341288,3.491766,3.049403,2.5290828,2.0105755,1.4902552,0.969935,0.44961473,0.99531645,1.5392052,2.084907,2.6306088,3.1744974,3.8108473,4.445384,5.0799212,5.714458,6.350808,6.0824895,5.814171,5.5476656,5.279347,5.0128417,4.9167547,4.8224807,4.7282066,4.632119,4.537845,4.632119,4.7282066,4.8224807,4.9167547,5.0128417,4.2876563,3.5624714,2.8372865,2.1121013,1.3869164,1.1167849,0.8466535,0.57833505,0.30820364,0.038072214,0.09064813,0.14322405,0.19579996,0.24837588,0.2991388,0.25925365,0.21936847,0.1794833,0.13959812,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.13778515,0.16316663,0.18673515,0.21211663,0.2374981,0.19579996,0.15228885,0.11059072,0.06707962,0.025381476,0.045324065,0.065266654,0.08520924,0.10515183,0.12509441,0.13415924,0.14503701,0.15410182,0.16497959,0.17585737,0.14684997,0.11965553,0.092461094,0.065266654,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06707962,0.13415924,0.2030518,0.27013144,0.33721104,1.1258497,1.9126755,2.6995013,3.48814,4.274966,3.6077955,2.9406252,2.2716422,1.6044719,0.93730164,2.665055,4.3928084,6.1205616,7.8483152,9.574255,7.7195945,5.864934,4.0102735,2.1556125,0.2991388,2.1229792,3.9450066,5.767034,7.590874,9.412902,7.5292335,5.6473784,3.7655232,1.8818551,0.0,0.48768693,0.97537386,1.4630609,1.9507477,2.4366217,3.0892882,3.7419548,4.3946214,5.047288,5.6999545,4.612177,3.5243993,2.4366217,1.3506571,0.26287958,0.21030366,0.15772775,0.10515183,0.052575916,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.027194439,0.030820364,0.032633327,0.034446288,0.038072214,0.047137026,0.058014803,0.06707962,0.07795739,0.0870222,0.07433146,0.06164073,0.05076295,0.038072214,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.072518505,0.08339628,0.092461094,0.10333887,0.11240368,0.12328146,0.13234627,0.14322405,0.15228885,0.16316663,0.15954071,0.15772775,0.15410182,0.15228885,0.15047589,0.14503701,0.13959812,0.13415924,0.13053331,0.12509441,0.11784257,0.11059072,0.10333887,0.09427405,0.0870222,0.08520924,0.08339628,0.07977036,0.07795739,0.07433146,0.06707962,0.059827764,0.052575916,0.045324065,0.038072214,0.045324065,0.052575916,0.059827764,0.06707962,0.07433146,0.07433146,0.07433146,0.07433146,0.07433146,0.07433146,4.6248674,4.6774435,4.7300196,4.782595,4.835171,4.8877473,5.2158933,5.542227,5.870373,6.1967063,6.5248523,6.9200783,7.315304,7.71053,8.105756,8.499168,8.192778,7.8845744,7.5781837,7.26998,6.9617763,7.271793,7.5818095,7.891826,8.201842,8.511859,7.989726,7.4675927,6.94546,6.4233265,5.89938,6.624565,7.3497505,8.074935,8.80012,9.525306,8.914337,8.3051815,7.6942134,7.0850577,6.4759026,7.5056653,8.535428,9.56519,10.594954,11.624716,11.922042,12.219368,12.516694,12.815832,13.113158,12.222994,11.332829,10.442664,9.5525,8.662335,9.097446,9.5325575,9.967669,10.40278,10.837891,13.878228,16.916754,19.957092,22.99743,26.03777,21.184467,16.33298,11.479679,6.628191,1.7748904,1.5899682,1.405046,1.2201238,1.0352017,0.85027945,0.67986095,0.5094425,0.34083697,0.17041849,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08520924,0.17041849,0.25562772,0.34083697,0.42423326,1.4467441,2.469255,3.491766,4.514277,5.5367875,4.439945,3.343103,2.2444477,1.1476053,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.27013144,0.5402629,0.8103943,1.0805258,1.3506571,1.6552348,1.9598125,2.2643902,2.570781,2.8753586,3.5733492,4.269527,4.9675174,5.6655083,6.3616858,7.137634,7.911769,8.6877165,9.461852,10.2378,9.325879,8.412147,7.500226,6.588306,5.674573,5.91751,6.1604466,6.4033837,6.644508,6.887445,6.9508986,7.0125394,7.07418,7.137634,7.1992745,8.158332,9.115576,10.07282,11.030065,11.9873085,12.06164,12.137785,12.212116,12.28826,12.362592,13.037014,13.713249,14.387671,15.062093,15.738328,16.169813,16.603111,17.034595,17.467894,17.89938,17.97915,18.060734,18.140503,18.220274,18.300045,17.812357,17.32467,16.836983,16.349297,15.861609,15.74558,15.627737,15.509895,15.392053,15.27421,15.934128,16.59586,17.255777,17.915697,18.575615,18.173138,17.770658,17.368181,16.965704,16.563227,16.487082,16.41275,16.336605,16.262274,16.187943,17.235836,18.281914,19.329807,20.377699,21.425592,23.349146,25.274511,27.199877,29.125244,31.05061,31.831997,32.615196,33.398396,34.179783,34.962982,34.4481,33.93322,33.41834,32.901646,32.386765,32.63514,32.881702,33.130077,33.37664,33.625015,33.677593,33.730167,33.782745,33.83532,33.887897,33.599636,33.313187,33.024925,32.736664,32.45022,31.242785,30.03535,28.827917,27.620485,26.413052,26.929747,27.448254,27.964949,28.481642,29.000149,29.718082,30.434202,31.152136,31.87007,32.588,32.633327,32.676838,32.72216,32.767487,32.81281,35.42166,38.03233,40.642994,43.25185,45.862514,43.697838,41.53316,39.36667,37.201992,35.037315,33.316814,31.598125,29.877623,28.157122,26.43662,24.166792,21.896961,19.627132,17.357304,15.087475,14.387671,13.687867,12.988064,12.28826,11.586644,11.711739,11.836833,11.961927,12.087022,12.212116,11.302009,10.391902,9.481794,8.571687,7.663393,6.740595,5.8177967,4.894999,3.972201,3.049403,2.4402475,1.8292793,1.2201238,0.6091554,0.0,1.357909,2.715818,4.071914,5.429823,6.787732,5.560356,4.3329806,3.105605,1.8782293,0.6508536,1.4902552,2.3296568,3.1708715,4.0102735,4.8496747,4.6575007,4.465327,4.273153,4.079166,3.8869917,3.9975824,4.1081734,4.216951,4.327542,4.4381323,4.590421,4.74271,4.894999,5.047288,5.199577,5.3119802,5.424384,5.5367875,5.6491914,5.763408,5.8794374,5.99728,6.115123,6.2329655,6.350808,6.202145,6.055295,5.906632,5.7597823,5.612932,6.2329655,6.8529987,7.473032,8.093065,8.713099,8.015107,7.317117,6.6191263,5.922949,5.224958,5.230397,5.235836,5.239462,5.2449007,5.2503395,5.1923246,5.1343102,5.0781083,5.0200934,4.9620786,4.313038,3.6621845,3.0131438,2.3622901,1.7132497,1.6697385,1.6280404,1.5845293,1.5428312,1.49932,1.3651608,1.2291887,1.0950294,0.96087015,0.824898,1.0352017,1.2455053,1.455809,1.6642996,1.8746033,2.2933977,2.7103791,3.1273603,3.5443418,3.9631362,4.5668526,5.1723824,5.7779117,6.3816285,6.987158,6.4051967,5.823236,5.239462,4.6575007,4.07554,3.3702974,2.665055,1.9598125,1.2545701,0.5493277,1.3542831,2.1592383,2.9641938,3.7691493,4.574105,5.0019636,5.429823,5.857682,6.285541,6.7134004,6.0806766,5.4479527,4.8152285,4.1825047,3.5497808,3.7582715,3.9649491,4.171627,4.3801174,4.5867953,4.7680917,4.947575,5.127058,5.3083544,5.487838,4.7753434,4.062849,3.350355,2.6378605,1.9253663,1.5446441,1.1657349,0.7850128,0.40429065,0.025381476,0.08520924,0.14503701,0.20486477,0.26469254,0.3245203,0.29007402,0.25562772,0.21936847,0.18492219,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.099712946,0.12509441,0.15047589,0.17585737,0.19942589,0.16679256,0.13415924,0.10333887,0.07070554,0.038072214,0.054388877,0.072518505,0.09064813,0.10696479,0.12509441,0.15228885,0.1794833,0.20667773,0.23568514,0.26287958,0.21574254,0.16679256,0.11965553,0.072518505,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.045324065,0.09064813,0.13415924,0.1794833,0.22480737,0.7505665,1.2745126,1.8002719,2.324218,2.8499773,2.4547513,2.0595255,1.6642996,1.2708868,0.87566096,2.8227828,4.7699046,6.717026,8.664148,10.613083,8.529989,6.446895,4.365614,2.2825198,0.19942589,1.4159238,2.6306088,3.8452935,5.0599785,6.2746634,5.0200934,3.7655232,2.5091403,1.2545701,0.0,0.37528324,0.7505665,1.1258497,1.49932,1.8746033,2.3858588,2.8953013,3.4047437,3.9141862,4.4254417,3.5751622,2.7248828,1.8746033,1.0243238,0.17585737,0.13959812,0.10515183,0.07070554,0.034446288,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.034446288,0.032633327,0.030820364,0.027194439,0.025381476,0.03988518,0.054388877,0.07070554,0.08520924,0.099712946,0.0870222,0.07433146,0.06164073,0.05076295,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.07795739,0.092461094,0.10696479,0.12328146,0.13778515,0.13959812,0.14322405,0.14503701,0.14684997,0.15047589,0.15228885,0.15410182,0.15772775,0.15954071,0.16316663,0.15410182,0.14684997,0.13959812,0.13234627,0.12509441,0.11965553,0.11421664,0.11059072,0.10515183,0.099712946,0.09064813,0.07977036,0.07070554,0.059827764,0.05076295,0.045324065,0.03988518,0.034446288,0.030820364,0.025381476,0.030820364,0.034446288,0.03988518,0.045324065,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,4.8116026,4.8696175,4.9276323,4.985647,5.041849,5.0998635,5.319232,5.540414,5.7597823,5.979151,6.200332,6.546608,6.8946967,7.2427855,7.590874,7.93715,7.7141557,7.4929743,7.26998,7.0469856,6.825804,7.155763,7.4857225,7.8156815,8.145641,8.4756,7.8319983,7.1902094,6.546608,5.904819,5.2630305,6.037165,6.813113,7.5872483,8.363196,9.137331,8.6333275,8.127511,7.6216946,7.117691,6.6118746,7.83925,9.066626,10.2958145,11.5231905,12.750566,12.830337,12.910107,12.989877,13.069647,13.149418,12.130532,11.109835,10.089137,9.070251,8.049554,8.841819,9.634083,10.428161,11.220426,12.012691,14.770206,17.527721,20.285238,23.042755,25.80027,20.89258,15.984891,11.077202,6.169512,1.261822,1.0950294,0.92823684,0.75963134,0.59283876,0.42423326,0.34083697,0.25562772,0.17041849,0.08520924,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.092461094,0.18492219,0.27738327,0.36984438,0.46230546,1.5682126,2.6723068,3.778214,4.882308,5.9882154,4.795286,3.6023567,2.4094272,1.2183108,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.36077955,0.7197462,1.0805258,1.4394923,1.8002719,2.2027495,2.6052272,3.007705,3.4101827,3.8126602,4.704638,5.5966153,6.490406,7.382384,8.274362,8.80012,9.325879,9.849826,10.375585,10.899531,9.837135,8.774739,7.7123427,6.6499467,5.5875506,5.8522434,6.1169357,6.3816285,6.6481338,6.9128265,7.2754188,7.6380115,8.000604,8.363196,8.725789,9.610515,10.49524,11.379966,12.264692,13.149418,13.087777,13.024323,12.962683,12.899229,12.837588,13.588155,14.336908,15.087475,15.838041,16.586794,16.710075,16.833357,16.954826,17.078108,17.199575,17.215893,17.230396,17.2449,17.259403,17.27572,17.237648,17.199575,17.163317,17.125244,17.087172,16.82248,16.557787,16.293095,16.028402,15.761897,15.917811,16.071913,16.227829,16.38193,16.537846,16.405499,16.273151,16.140806,16.006647,15.8743,15.812659,15.749206,15.687565,15.624111,15.56247,16.916754,18.27285,19.627132,20.983229,22.337511,24.89923,27.462757,30.024473,32.588,35.14972,35.684544,36.219368,36.75419,37.29083,37.825653,36.980812,36.13416,35.289318,34.444477,33.599636,33.75555,33.909653,34.065567,34.21967,34.375584,34.469856,34.564133,34.660217,34.754494,34.85058,34.524246,34.199726,33.875206,33.550686,33.224354,32.06587,30.905573,29.745277,28.584982,27.424685,27.865234,28.305784,28.744522,29.185072,29.625622,29.714457,29.805105,29.895754,29.984589,30.075235,30.084301,30.095179,30.104244,30.115122,30.124186,32.979603,35.83502,38.690434,41.54585,44.399452,42.57924,40.760838,38.940624,37.120407,35.300194,33.739235,32.180084,30.619125,29.059977,27.50083,25.08959,22.680162,20.270735,17.859495,15.4500675,14.9877615,14.525456,14.06315,13.600845,13.136727,12.962683,12.786825,12.612781,12.436923,12.262879,11.245807,10.226922,9.20985,8.192778,7.175706,6.3816285,5.5893636,4.797099,4.004834,3.2125697,2.570781,1.9271792,1.2853905,0.6417888,0.0,1.0841516,2.1701162,3.254268,4.3402324,5.424384,4.4798307,3.5352771,2.5907235,1.6443571,0.69980353,1.4703126,2.2408218,3.009518,3.780027,4.550536,4.273153,3.9957695,3.7183862,3.43919,3.1618068,3.2796493,3.397492,3.5153344,3.633177,3.7492065,3.9450066,4.1408067,4.3347936,4.5305934,4.7245803,4.800725,4.8750563,4.949388,5.0255322,5.0998635,5.177821,5.2557783,5.331923,5.40988,5.487838,5.132497,4.7771564,4.421816,4.068288,3.7129474,4.347484,4.9820213,5.618371,6.2529078,6.887445,6.4577727,6.0281005,5.5966153,5.1669436,4.7372713,4.989273,5.243088,5.4950895,5.7470913,6.000906,5.4896507,4.9802084,4.4707656,3.9595103,3.4500678,2.9369993,2.4257438,1.9126755,1.3996071,0.8883517,0.85934424,0.8321498,0.80495536,0.7777609,0.7505665,0.69436467,0.6399758,0.5855869,0.5293851,0.4749962,0.59283876,0.7106813,0.82671094,0.9445535,1.062396,1.6026589,2.1429217,2.6831846,3.2216346,3.7618973,4.751775,5.7416525,6.733343,7.723221,8.713099,7.989726,7.268167,6.544795,5.823236,5.0998635,4.209699,3.3195345,2.42937,1.5392052,0.6508536,1.7150626,2.7792716,3.8452935,4.9095025,5.975525,6.1948934,6.414262,6.635443,6.8548117,7.07418,6.0770507,5.0799212,4.082792,3.0856624,2.08672,2.5979755,3.1074178,3.6168604,4.1281157,4.6375585,4.902251,5.1669436,5.431636,5.6981416,5.962834,5.2630305,4.5632267,3.8616104,3.1618068,2.4620032,1.9725033,1.4830034,0.9916905,0.50219065,0.012690738,0.07977036,0.14684997,0.21574254,0.28282216,0.34990177,0.3208944,0.29007402,0.25925365,0.23024625,0.19942589,0.15954071,0.11965553,0.07977036,0.03988518,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.06164073,0.0870222,0.11240368,0.13778515,0.16316663,0.13959812,0.11784257,0.09427405,0.072518505,0.05076295,0.065266654,0.07977036,0.09427405,0.11059072,0.12509441,0.17041849,0.21574254,0.25925365,0.3045777,0.34990177,0.28282216,0.21574254,0.14684997,0.07977036,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.37528324,0.63816285,0.89922947,1.162109,1.4249886,1.3017071,1.1802386,1.0569572,0.9354887,0.8122072,2.9805105,5.147001,7.315304,9.481794,11.650098,9.340384,7.0306687,4.7191415,2.4094272,0.099712946,0.7070554,1.3143979,1.9217403,2.5290828,3.1382382,2.5091403,1.8818551,1.2545701,0.62728506,0.0,0.26287958,0.52575916,0.7868258,1.0497054,1.3125849,1.6806163,2.0468347,2.4148662,2.7828975,3.149116,2.5381477,1.9253663,1.3125849,0.69980353,0.0870222,0.07070554,0.052575916,0.034446288,0.018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.04169814,0.034446288,0.027194439,0.01994259,0.012690738,0.032633327,0.052575916,0.072518505,0.092461094,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.08339628,0.10333887,0.12328146,0.14322405,0.16316663,0.15772775,0.15228885,0.14684997,0.14322405,0.13778515,0.14503701,0.15228885,0.15954071,0.16679256,0.17585737,0.16497959,0.15410182,0.14503701,0.13415924,0.12509441,0.12328146,0.11965553,0.11784257,0.11421664,0.11240368,0.09427405,0.07795739,0.059827764,0.04169814,0.025381476,0.02175555,0.01994259,0.018129626,0.014503701,0.012690738,0.014503701,0.018129626,0.01994259,0.02175555,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,5.0001507,5.0617914,5.125245,5.186886,5.2503395,5.3119802,5.424384,5.5367875,5.6491914,5.763408,5.8758116,6.1749506,6.474089,6.775041,7.07418,7.3751316,7.2373466,7.0995617,6.9617763,6.825804,6.688019,7.037921,7.3878226,7.7377243,8.087626,8.437528,7.6742706,6.9128265,6.149569,5.388125,4.6248674,5.4497657,6.2746634,7.0995617,7.9244595,8.749357,8.350506,7.949841,7.549176,7.1503243,6.7496595,8.174648,9.599637,11.024626,12.449615,13.874602,13.736817,13.600845,13.46306,13.325275,13.1874895,12.038072,10.88684,9.737422,8.588004,7.4367723,8.588004,9.737422,10.88684,12.038072,13.1874895,15.662184,18.136877,20.613384,23.088078,25.562773,20.600695,15.636803,10.674724,5.712645,0.7505665,0.6000906,0.44961473,0.2991388,0.15047589,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.099712946,0.19942589,0.2991388,0.40066472,0.50037766,1.6878681,2.8753586,4.062849,5.2503395,6.43783,5.1506267,3.8634233,2.5744069,1.2872034,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.44961473,0.89922947,1.3506571,1.8002719,2.2498865,2.7502642,3.2506418,3.7492065,4.249584,4.749962,5.8377395,6.925517,8.013294,9.099259,10.1870365,10.462607,10.738177,11.011934,11.287505,11.563075,10.3502035,9.137331,7.9244595,6.7115874,5.5005283,5.7869763,6.0752378,6.3616858,6.6499467,6.9382076,7.5999393,8.26167,8.925215,9.5869465,10.25049,11.062697,11.874905,12.687112,13.499319,14.313339,14.112101,13.912675,13.713249,13.512011,13.312584,14.137483,14.96238,15.787278,16.612177,17.437075,17.25034,17.06179,16.875055,16.68832,16.499773,16.450823,16.400059,16.349297,16.300346,16.249584,16.66294,17.074482,17.487837,17.89938,18.312735,17.89938,17.487837,17.074482,16.66294,16.249584,15.899682,15.54978,15.199879,14.849977,14.500074,14.63786,14.775645,14.911617,15.049402,15.187187,15.138238,15.087475,15.036712,14.9877615,14.936998,16.599485,18.261972,19.92446,21.586945,23.249432,26.44931,29.64919,32.850883,36.050762,39.25064,39.537086,39.825348,40.111797,40.40006,40.68832,39.511707,38.336906,37.162106,35.98731,34.812508,34.87415,34.937603,34.99924,35.062695,35.124336,35.262123,35.399906,35.537693,35.675476,35.813263,35.450672,35.088078,34.725487,34.362892,34.0003,32.887142,31.775795,30.662636,29.549477,28.438131,28.800724,29.163317,29.52591,29.886688,30.24928,29.712645,29.174194,28.637556,28.099108,27.56247,27.537088,27.511707,27.488138,27.462757,27.437376,30.537542,33.637707,36.737873,39.83804,42.938206,41.462456,39.986702,38.512764,37.037014,35.563072,34.161655,32.762047,31.36244,29.962833,28.563225,26.012386,23.463362,20.912523,18.361685,15.812659,15.5878525,15.363045,15.138238,14.911617,14.68681,14.211814,13.736817,13.261822,12.786825,12.311829,11.187792,10.061942,8.937905,7.8120556,6.688019,6.0244746,5.3627434,4.699199,4.0374675,3.3757362,2.6995013,2.0250793,1.3506571,0.6744221,0.0,0.8122072,1.6244144,2.4366217,3.2506418,4.062849,3.3993049,2.7375734,2.0758421,1.4122978,0.7505665,1.4503701,2.1501737,2.8499773,3.5497808,4.249584,3.8869917,3.5243993,3.1618068,2.7992141,2.4366217,2.561716,2.6868105,2.811905,2.9369993,3.0620937,3.299592,3.53709,3.774588,4.0120864,4.249584,4.2876563,4.325729,4.361988,4.40006,4.4381323,4.4743915,4.512464,4.550536,4.5867953,4.6248674,4.062849,3.5008307,2.9369993,2.374981,1.8129625,2.4620032,3.1128569,3.7618973,4.4127507,5.0617914,4.900438,4.7372713,4.574105,4.4127507,4.249584,4.749962,5.2503395,5.750717,6.249282,6.7496595,5.7869763,4.8242936,3.8616104,2.9007401,1.938057,1.5627737,1.1874905,0.8122072,0.43692398,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.15047589,0.17585737,0.19942589,0.22480737,0.25018883,0.9119202,1.5754645,2.2371957,2.9007401,3.5624714,4.936697,6.3127356,7.686961,9.063,10.437225,9.574255,8.713099,7.850128,6.987158,6.1241875,5.049101,3.975827,2.9007401,1.8256533,0.7505665,2.0758421,3.3993049,4.7245803,6.049856,7.3751316,7.3878226,7.400513,7.413204,7.4258947,7.4367723,6.0752378,4.7118897,3.350355,1.987007,0.62547207,1.4376793,2.2498865,3.0620937,3.874301,4.688321,5.038223,5.388125,5.7380266,6.0879283,6.43783,5.750717,5.0617914,4.3746786,3.6875658,3.000453,2.4003625,1.8002719,1.2001812,0.6000906,0.0,0.07433146,0.15047589,0.22480737,0.2991388,0.37528324,0.34990177,0.3245203,0.2991388,0.2755703,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.18673515,0.25018883,0.31182957,0.37528324,0.43692398,0.34990177,0.26287958,0.17585737,0.0870222,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.15047589,0.2991388,0.44961473,0.6000906,0.7505665,3.1382382,5.524097,7.911769,10.29944,12.687112,10.148965,7.61263,5.0744824,2.5381477,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.15047589,0.2991388,0.44961473,0.6000906,0.7505665,0.97537386,1.2001812,1.4249886,1.649796,1.8746033,1.49932,1.1258497,0.7505665,0.37528324,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.0870222,0.11240368,0.13778515,0.16316663,0.18673515,0.17585737,0.16316663,0.15047589,0.13778515,0.12509441,0.13778515,0.15047589,0.16316663,0.17585737,0.18673515,0.17585737,0.16316663,0.15047589,0.13778515,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,4.900438,5.0074024,5.1143675,5.223145,5.33011,5.4370747,5.375434,5.3119802,5.2503395,5.186886,5.125245,5.524097,5.924762,6.3254266,6.7242785,7.124943,7.179332,7.2355337,7.2899227,7.344311,7.400513,7.5346723,7.6706448,7.804804,7.9407763,8.074935,7.4694057,6.8656893,6.26016,5.65463,5.049101,5.7017674,6.354434,7.0071006,7.6597667,8.312433,8.138389,7.9625316,7.7866745,7.61263,7.4367723,8.747544,10.058316,11.367275,12.678047,13.987006,13.747695,13.508384,13.267261,13.027949,12.786825,11.83502,10.883214,9.929596,8.977791,8.024173,9.492672,10.959359,12.427858,13.894546,15.363045,17.375433,19.387821,21.40021,23.4126,25.424988,20.56806,15.709321,10.852394,5.995467,1.1367276,0.91735905,0.6979906,0.47680917,0.2574407,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.11965553,0.23931105,0.36077955,0.48043507,0.6000906,0.5656443,0.5293851,0.4949388,0.4604925,0.42423326,0.42060733,0.41516843,0.40972954,0.40429065,0.40066472,1.4866294,2.5744069,3.6621845,4.749962,5.8377395,4.6792564,3.5225863,2.3641033,1.2074331,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.8031424,1.6044719,2.4076142,3.2107568,4.0120864,4.465327,4.9167547,5.369995,5.823236,6.2746634,7.2554765,8.234476,9.215289,10.194288,11.175101,11.082641,10.990179,10.897718,10.805257,10.712796,9.684846,8.656897,7.6307597,6.60281,5.57486,5.964647,6.354434,6.7442207,7.135821,7.5256076,8.0858135,8.644206,9.2044115,9.764616,10.324821,11.008308,11.689982,12.371656,13.055143,13.736817,13.651608,13.568212,13.483003,13.397794,13.312584,13.992445,14.672306,15.352167,16.032028,16.71189,16.617615,16.52334,16.427254,16.33298,16.236893,16.177065,16.117237,16.05741,15.9975815,15.937754,16.287657,16.637558,16.98746,17.33736,17.687263,17.400814,17.112555,16.824293,16.537846,16.249584,15.952258,15.654932,15.357606,15.06028,14.762955,14.90074,15.036712,15.174497,15.312282,15.4500675,15.495391,15.540715,15.584227,15.62955,15.674874,16.980207,18.285542,19.590874,20.894394,22.199726,24.817644,27.435562,30.051668,32.669586,35.287502,35.483303,35.67729,35.87309,36.067078,36.26288,35.60477,34.946667,34.290375,33.632267,32.974163,33.309563,33.64496,33.98036,34.315754,34.64934,34.866898,35.084454,35.302006,35.51956,35.737118,35.635593,35.532253,35.43073,35.32739,35.225864,34.194286,33.164524,32.13476,31.105,30.075235,30.410635,30.744219,31.079618,31.415016,31.750414,31.119503,30.490404,29.859493,29.230396,28.599485,28.369238,28.140804,27.910559,27.680313,27.450066,30.167698,32.885326,35.60296,38.32059,41.03822,39.945004,38.851788,37.760384,36.667168,35.575764,34.54056,33.50536,32.47016,31.434958,30.399757,27.395678,24.389786,21.385706,18.379814,15.375735,16.08279,16.789846,17.496902,18.20577,18.912827,17.389936,15.867048,14.34416,12.823084,11.300196,10.388275,9.474543,8.562622,7.650702,6.736969,5.9302006,5.121619,4.314851,3.5080826,2.6995013,2.3024626,1.9054236,1.5083848,1.1095331,0.7124943,1.5428312,2.373168,3.2016919,4.0320287,4.8623657,4.0157123,3.1672456,2.3205922,1.4721256,0.62547207,1.1802386,1.7350051,2.2897718,2.8445382,3.3993049,3.1255474,2.8499773,2.5744069,2.3006494,2.0250793,2.2643902,2.5055144,2.7448254,2.9841363,3.2252605,3.3322253,3.43919,3.5479677,3.6549325,3.7618973,3.8180993,3.872488,3.926877,3.9830787,4.0374675,4.0102735,3.9830787,3.9558845,3.926877,3.8996825,3.4101827,2.9206827,2.42937,1.93987,1.4503701,2.2933977,3.1346123,3.97764,4.8206677,5.661882,5.6927023,5.7217097,5.75253,5.7833505,5.812358,5.859495,5.906632,5.955582,6.002719,6.049856,5.1923246,4.3347936,3.4772623,2.619731,1.7621996,1.4195497,1.0768998,0.73424983,0.39159992,0.05076295,0.15954071,0.27013144,0.38072214,0.4894999,0.6000906,0.56745726,0.53482395,0.50219065,0.46955732,0.43692398,0.44780177,0.45686656,0.46774435,0.47680917,0.48768693,0.9644961,1.4431182,1.9199274,2.3967366,2.8753586,4.0374675,5.199577,6.3616858,7.5256076,8.6877165,8.009668,7.3316207,6.6553855,5.977338,5.2992897,4.441758,3.584227,2.7266958,1.8691645,1.0116332,2.0667772,3.1219215,4.177066,5.23221,6.2873545,6.2293396,6.1731377,6.115123,6.057108,5.999093,4.900438,3.7999697,2.6995013,1.6008459,0.50037766,1.1566701,1.8147756,2.472881,3.1291735,3.787279,4.1806917,4.572292,4.9657044,5.3573046,5.750717,5.1542525,4.559601,3.9649491,3.3702974,2.7756457,2.222692,1.6697385,1.1167849,0.5656443,0.012690738,0.07433146,0.13778515,0.19942589,0.26287958,0.3245203,0.3208944,0.3154555,0.3100166,0.3045777,0.2991388,0.23931105,0.1794833,0.11965553,0.059827764,0.0,0.0,0.0,0.0,0.0,0.0,0.027194439,0.054388877,0.08339628,0.11059072,0.13778515,0.12328146,0.10696479,0.092461094,0.07795739,0.06164073,0.099712946,0.13778515,0.17585737,0.21211663,0.25018883,0.27194437,0.2955129,0.31726846,0.34083697,0.36259252,0.38072214,0.39703882,0.41516843,0.43329805,0.44961473,0.36077955,0.27013144,0.1794833,0.09064813,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.059827764,0.11965553,0.1794833,0.23931105,0.2991388,0.89922947,1.49932,2.0994108,2.6995013,3.299592,2.7792716,2.2607644,1.7404441,1.2201238,0.69980353,2.5907235,4.4798307,6.3707504,8.259857,10.150778,8.147454,6.145943,4.1426196,2.1392958,0.13778515,0.11059072,0.08339628,0.054388877,0.027194439,0.0,0.052575916,0.10515183,0.15772775,0.21030366,0.26287958,0.32995918,0.39703882,0.46411842,0.533011,0.6000906,0.85027945,1.1004683,1.3506571,1.6008459,1.8492218,1.4793775,1.1095331,0.73968875,0.36984438,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.027194439,0.04169814,0.058014803,0.072518505,0.0870222,0.072518505,0.058014803,0.04169814,0.027194439,0.012690738,0.034446288,0.058014803,0.07977036,0.10333887,0.12509441,0.12328146,0.11965553,0.11784257,0.11421664,0.11240368,0.09427405,0.07795739,0.059827764,0.04169814,0.025381476,0.02175555,0.01994259,0.018129626,0.014503701,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.02175555,0.032633327,0.04169814,0.052575916,0.06164073,0.0870222,0.11240368,0.13778515,0.16316663,0.18673515,0.18310922,0.17767033,0.17223145,0.16679256,0.16316663,0.18492219,0.20667773,0.23024625,0.2520018,0.2755703,0.2574407,0.23931105,0.2229944,0.20486477,0.18673515,0.17767033,0.16679256,0.15772775,0.14684997,0.13778515,0.11421664,0.092461094,0.07070554,0.047137026,0.025381476,0.02175555,0.01994259,0.018129626,0.014503701,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,4.800725,4.953014,5.105303,5.2575917,5.40988,5.562169,5.3246713,5.087173,4.8496747,4.612177,4.3746786,4.8750563,5.375434,5.8758116,6.3743763,6.874754,7.12313,7.369693,7.6180687,7.8646317,8.113008,8.033237,7.951654,7.8718834,7.7921133,7.7123427,7.264541,6.816739,6.3707504,5.922949,5.475147,5.955582,6.434204,6.9146395,7.3950744,7.8755093,7.9244595,7.9752226,8.024173,8.074935,8.125698,9.32044,10.515183,11.709926,12.904668,14.09941,13.75676,13.41411,13.073273,12.730623,12.387974,11.631968,10.877775,10.12177,9.367578,8.613385,10.397341,12.183108,13.967064,15.752831,17.536787,19.08687,20.636953,22.187037,23.73712,25.287203,20.535427,15.781839,11.030065,6.2782893,1.5247015,1.2346275,0.9445535,0.6544795,0.36440548,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.23931105,0.48043507,0.7197462,0.96087015,1.2001812,1.1294757,1.0605831,0.9898776,0.91917205,0.85027945,0.73968875,0.630911,0.52032024,0.40972954,0.2991388,1.2872034,2.275268,3.2633326,4.249584,5.237649,4.209699,3.1817493,2.1556125,1.1276628,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0,0.0,0.0,0.0,0.0,1.1548572,2.3097143,3.4645715,4.6194286,5.774286,6.1803894,6.58468,6.9907837,7.3950744,7.799365,8.673213,9.545248,10.417283,11.289318,12.163166,11.702674,11.242181,10.781689,10.323009,9.862516,9.019489,8.178274,7.3352466,6.492219,5.6491914,6.1423173,6.635443,7.1267557,7.6198816,8.113008,8.569874,9.026741,9.48542,9.9422865,10.399154,10.952107,11.50506,12.058014,12.609155,13.162108,13.192928,13.221936,13.252756,13.281764,13.312584,13.847408,14.382232,14.917056,15.45188,15.986704,15.984891,15.983078,15.979452,15.977639,15.975826,15.905121,15.834415,15.765523,15.694818,15.624111,15.912373,16.200634,16.487082,16.775343,17.06179,16.900436,16.73727,16.574104,16.41275,16.249584,16.004833,15.760084,15.515334,15.270584,15.025834,15.161806,15.299591,15.437376,15.575162,15.712947,15.852545,15.992143,16.13174,16.273151,16.41275,17.359118,18.307297,19.255476,20.201841,21.15002,23.184166,25.220123,27.254267,29.290224,31.324368,31.427706,31.529232,31.63257,31.734097,31.837437,31.697838,31.558239,31.416828,31.277231,31.137632,31.744974,32.352318,32.95966,33.567,34.174343,34.471672,34.77081,35.068134,35.36546,35.66279,35.820515,35.97824,36.13416,36.291885,36.44961,35.503246,34.555065,33.606888,32.660522,31.712341,32.020546,32.326935,32.63514,32.943344,33.249733,32.528175,31.804802,31.083244,30.35987,29.638311,29.203201,28.768091,28.33298,27.89787,27.462757,29.797853,32.13295,34.468044,36.80314,39.138237,38.427555,37.716873,37.008007,36.297325,35.586643,34.91766,34.246864,33.57788,32.907085,32.238102,28.777155,25.318022,21.857077,18.397943,14.936998,16.57773,18.216648,19.85738,21.49811,23.137028,20.56806,17.99728,15.428311,12.857531,10.28675,9.5869465,8.887142,8.187339,7.4875355,6.787732,5.8341136,4.882308,3.930503,2.9768846,2.0250793,1.9054236,1.7857682,1.6642996,1.5446441,1.4249886,2.2716422,3.1201086,3.966762,4.8152285,5.661882,4.6303062,3.5969179,2.565342,1.5319533,0.50037766,0.9101072,1.3198367,1.7295663,2.1392958,2.5508385,2.3622901,2.175555,1.987007,1.8002719,1.6117238,1.9670644,2.322405,2.6777458,3.0330863,3.386614,3.3648586,3.343103,3.3195345,3.2977788,3.2742105,3.346729,3.4192474,3.491766,3.5642843,3.636803,3.5443418,3.4518807,3.3594196,3.2669585,3.1744974,2.7575161,2.3405347,1.9217403,1.504759,1.0877775,2.1229792,3.1581807,4.1933823,5.2267714,6.261973,6.484967,6.7079616,6.929143,7.1521373,7.3751316,6.970841,6.5647373,6.1604466,5.754343,5.3500524,4.597673,3.8452935,3.092914,2.3405347,1.5881553,1.2781386,0.968122,0.65810543,0.3480888,0.038072214,0.27013144,0.50219065,0.73424983,0.968122,1.2001812,1.1095331,1.020698,0.9300498,0.83940166,0.7505665,0.7451276,0.73968875,0.73424983,0.7306239,0.72518504,1.017072,1.310772,1.6026589,1.8945459,2.1882458,3.1382382,4.0882306,5.038223,5.9882154,6.9382076,6.445082,5.9519563,5.4606433,4.9675174,4.4743915,3.834416,3.1944401,2.5544643,1.9144884,1.2745126,2.0595255,2.8445382,3.6295512,4.4145637,5.199577,5.0726695,4.945762,4.8170414,4.690134,4.5632267,3.7256382,2.8880494,2.0504606,1.2128719,0.37528324,0.8774739,1.3796645,1.8818551,2.3858588,2.8880494,3.3231604,3.7582715,4.1933823,4.6266804,5.0617914,4.559601,4.0574102,3.5552197,3.053029,2.5508385,2.0450218,1.5392052,1.0352017,0.5293851,0.025381476,0.07433146,0.12509441,0.17585737,0.22480737,0.2755703,0.29007402,0.3045777,0.3208944,0.33539808,0.34990177,0.27919623,0.21030366,0.13959812,0.07070554,0.0,0.0,0.0,0.0,0.0,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.13234627,0.11421664,0.09789998,0.07977036,0.06164073,0.12509441,0.18673515,0.25018883,0.31182957,0.37528324,0.35715362,0.34083697,0.32270733,0.3045777,0.28826106,0.40972954,0.533011,0.6544795,0.7777609,0.89922947,0.7197462,0.5402629,0.36077955,0.1794833,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.11965553,0.23931105,0.36077955,0.48043507,0.6000906,1.8002719,3.000453,4.2006345,5.4008155,6.599184,5.40988,4.220577,3.0294604,1.840157,0.6508536,2.0432088,3.435564,4.8279195,6.2202744,7.61263,6.14413,4.6774435,3.2107568,1.742257,0.2755703,0.21936847,0.16497959,0.11059072,0.054388877,0.0,0.10515183,0.21030366,0.3154555,0.42060733,0.52575916,0.5094425,0.4949388,0.48043507,0.46411842,0.44961473,0.72518504,1.0007553,1.2745126,1.550083,1.8256533,1.4594349,1.0950294,0.7306239,0.36440548,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.04169814,0.059827764,0.07795739,0.09427405,0.11240368,0.09427405,0.07795739,0.059827764,0.04169814,0.025381476,0.045324065,0.065266654,0.08520924,0.10515183,0.12509441,0.13234627,0.13959812,0.14684997,0.15410182,0.16316663,0.13959812,0.11784257,0.09427405,0.072518505,0.05076295,0.045324065,0.03988518,0.034446288,0.030820364,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.032633327,0.03988518,0.047137026,0.054388877,0.06164073,0.0870222,0.11240368,0.13778515,0.16316663,0.18673515,0.19036107,0.19217403,0.19579996,0.19761293,0.19942589,0.23205921,0.26469254,0.29732585,0.32995918,0.36259252,0.34083697,0.31726846,0.2955129,0.27194437,0.25018883,0.23024625,0.21030366,0.19036107,0.17041849,0.15047589,0.13053331,0.11059072,0.09064813,0.07070554,0.05076295,0.045324065,0.03988518,0.034446288,0.030820364,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,4.699199,4.896812,5.0944247,5.292038,5.4896507,5.6872635,5.275721,4.8623657,4.4508233,4.0374675,3.6241121,4.2242026,4.8242936,5.424384,6.0244746,6.624565,7.065115,7.5056653,7.944402,8.384952,8.825501,8.529989,8.234476,7.9407763,7.645263,7.3497505,7.059676,6.7696023,6.4795284,6.189454,5.89938,6.207584,6.5157876,6.8221784,7.130382,7.4367723,7.7123427,7.987913,8.26167,8.537241,8.812811,9.893337,10.97205,12.052575,13.1331005,14.211814,13.767638,13.321649,12.877473,12.433297,11.9873085,11.430729,10.872336,10.315757,9.757364,9.200785,11.302009,13.4050455,15.508082,17.609306,19.712341,20.80012,21.887897,22.975676,24.06164,25.149418,20.502794,15.854358,11.207735,6.5592985,1.9126755,1.551896,1.1929294,0.8321498,0.47318324,0.11240368,0.09064813,0.06707962,0.045324065,0.02175555,0.0,0.36077955,0.7197462,1.0805258,1.4394923,1.8002719,1.69512,1.5899682,1.4848163,1.3796645,1.2745126,1.0605831,0.8448406,0.629098,0.41516843,0.19942589,1.0877775,1.9743162,2.8626678,3.7492065,4.6375585,3.7401419,2.8427253,1.9453088,1.0478923,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.0,0.0,0.0,0.0,0.0,1.5065719,3.0149567,4.5233417,6.0299134,7.5382986,7.895452,8.252605,8.609759,8.966913,9.325879,10.089137,10.854207,11.619277,12.384347,13.149418,12.322706,11.494183,10.667472,9.840761,9.012237,8.354132,7.6978393,7.039734,6.3816285,5.7253356,6.319988,6.9146395,7.509291,8.105756,8.700407,9.055748,9.409276,9.764616,10.119957,10.475298,10.897718,11.320138,11.7425585,12.164979,12.5873995,12.732436,12.877473,13.022511,13.167547,13.312584,13.702372,14.092158,14.481945,14.871732,15.263332,15.352167,15.442815,15.531651,15.622298,15.712947,15.633177,15.553406,15.471823,15.392053,15.312282,15.537089,15.761897,15.986704,16.213324,16.438131,16.400059,16.361988,16.325727,16.287657,16.249584,16.05741,15.865235,15.673061,15.480887,15.2869005,15.4246855,15.56247,15.700256,15.838041,15.975826,16.209698,16.445383,16.679256,16.914942,17.150625,17.73984,18.330864,18.920078,19.50929,20.100317,21.5525,23.004683,24.456865,25.910862,27.363045,27.372108,27.382986,27.392052,27.40293,27.411995,27.790903,28.168,28.545095,28.922192,29.299288,30.180387,31.059675,31.940775,32.82006,33.69935,34.07826,34.455353,34.83245,35.209545,35.586643,36.005436,36.422417,36.8394,37.258194,37.675175,36.81039,35.94561,35.080826,34.21423,33.349445,33.630455,33.909653,34.190662,34.469856,34.750866,33.93503,33.1192,32.30518,31.489347,30.675327,30.03535,29.395376,28.7554,28.115423,27.475449,29.428009,31.38057,33.33313,35.28569,37.23825,36.910107,36.58196,36.255627,35.92748,35.599335,35.294754,34.990177,34.6856,34.379208,34.07463,30.160446,26.244446,22.33026,18.41426,14.500074,17.072668,19.645262,22.217857,24.790451,27.363045,23.744371,20.12751,16.51065,12.891977,9.275117,8.78743,8.299743,7.8120556,7.324369,6.836682,5.7398396,4.6429973,3.5443418,2.4474995,1.3506571,1.5083848,1.6642996,1.8220274,1.9797552,2.137483,3.002266,3.8670492,4.7318325,5.5966153,6.4632115,5.2449007,4.028403,2.810092,1.5917811,0.37528324,0.6399758,0.90466833,1.1693609,1.4358664,1.7005589,1.6008459,1.49932,1.3996071,1.2998942,1.2001812,1.6697385,2.1392958,2.610666,3.0802233,3.5497808,3.397492,3.245203,3.092914,2.9406252,2.7883365,2.8771715,2.9678197,3.056655,3.147303,3.2379513,3.0802233,2.9224956,2.764768,2.6070402,2.4493124,2.1048496,1.7603867,1.4141108,1.0696479,0.72518504,1.9525607,3.1799364,4.407312,5.634688,6.8620634,7.2772317,7.6924005,8.107569,8.5227375,8.937905,8.080374,7.2228427,6.3653116,5.5077806,4.650249,4.0030212,3.3557937,2.7067533,2.0595255,1.4122978,1.1349145,0.8575313,0.58014804,0.30276474,0.025381476,0.38072214,0.73424983,1.0895905,1.4449311,1.8002719,1.651609,1.504759,1.357909,1.209246,1.062396,1.0424535,1.0225109,1.0025684,0.9826257,0.96268314,1.0696479,1.1766127,1.2853905,1.3923552,1.49932,2.2371957,2.9750717,3.7129474,4.4508233,5.186886,4.880495,4.572292,4.265901,3.9576974,3.6494937,3.2270734,2.8046532,2.382233,1.9598125,1.5373923,2.0522738,2.5671551,3.0820365,3.5969179,4.1117992,3.9141862,3.7183862,3.5207734,3.3231604,3.1255474,2.5508385,1.9743162,1.3996071,0.824898,0.25018883,0.5982776,0.9445535,1.2926424,1.6407311,1.987007,2.465629,2.9424384,3.4192474,3.8978696,4.3746786,3.9649491,3.5552197,3.1454902,2.7357605,2.324218,1.8673514,1.4104849,0.95180535,0.4949388,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.22480737,0.25925365,0.2955129,0.32995918,0.36440548,0.40066472,0.3208944,0.23931105,0.15954071,0.07977036,0.0,0.0,0.0,0.0,0.0,0.0,0.032633327,0.065266654,0.09789998,0.13053331,0.16316663,0.14322405,0.12328146,0.10333887,0.08339628,0.06164073,0.15047589,0.2374981,0.3245203,0.41335547,0.50037766,0.44236287,0.38434806,0.32814622,0.27013144,0.21211663,0.4405499,0.6671702,0.89560354,1.1222239,1.3506571,1.0805258,0.8103943,0.5402629,0.27013144,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1794833,0.36077955,0.5402629,0.7197462,0.89922947,2.6995013,4.499773,6.300045,8.100317,9.900589,8.040489,6.1803894,4.3202896,2.4601903,0.6000906,1.4956942,2.3894846,3.2850883,4.1806917,5.0744824,4.1426196,3.2107568,2.277081,1.3452182,0.41335547,0.32995918,0.24837588,0.16497959,0.08339628,0.0,0.15772775,0.3154555,0.47318324,0.629098,0.7868258,0.69073874,0.59283876,0.4949388,0.39703882,0.2991388,0.6000906,0.89922947,1.2001812,1.49932,1.8002719,1.4394923,1.0805258,0.7197462,0.36077955,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.058014803,0.07795739,0.09789998,0.11784257,0.13778515,0.11784257,0.09789998,0.07795739,0.058014803,0.038072214,0.054388877,0.072518505,0.09064813,0.10696479,0.12509441,0.14322405,0.15954071,0.17767033,0.19579996,0.21211663,0.18492219,0.15772775,0.13053331,0.10333887,0.07433146,0.06707962,0.059827764,0.052575916,0.045324065,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.04169814,0.047137026,0.052575916,0.058014803,0.06164073,0.0870222,0.11240368,0.13778515,0.16316663,0.18673515,0.19761293,0.20667773,0.21755551,0.22662032,0.2374981,0.27919623,0.32270733,0.36440548,0.40791658,0.44961473,0.4224203,0.39522585,0.3680314,0.34083697,0.31182957,0.28282216,0.2520018,0.2229944,0.19217403,0.16316663,0.14503701,0.12690738,0.11059072,0.092461094,0.07433146,0.06707962,0.059827764,0.052575916,0.045324065,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,4.599486,4.842423,5.08536,5.328297,5.569421,5.812358,5.224958,4.6375585,4.0501585,3.4627585,2.8753586,3.5751622,4.274966,4.974769,5.674573,6.3743763,7.0071006,7.6398244,8.272549,8.9052725,9.537996,9.026741,8.517298,8.007855,7.4966,6.987158,6.8548117,6.722465,6.590119,6.4577727,6.3254266,6.4595857,6.5955577,6.7297173,6.8656893,6.9998484,7.500226,8.000604,8.499168,8.999546,9.499924,10.46442,11.430729,12.395226,13.359721,14.324218,13.776703,13.229188,12.681673,12.134158,11.586644,11.227677,10.866898,10.507931,10.147152,9.788185,12.206677,14.626982,17.047287,19.467592,21.887897,22.513369,23.137028,23.7625,24.387972,25.011631,20.470161,15.926876,11.385405,6.8421206,2.3006494,1.8691645,1.4394923,1.0098201,0.58014804,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.48043507,0.96087015,1.4394923,1.9199274,2.4003625,2.2607644,2.1193533,1.9797552,1.840157,1.7005589,1.3796645,1.0605831,0.73968875,0.42060733,0.099712946,0.8883517,1.6751775,2.4620032,3.2506418,4.0374675,3.2705846,2.5018883,1.7350051,0.968122,0.19942589,0.15954071,0.11965553,0.07977036,0.03988518,0.0,0.0,0.0,0.0,0.0,0.0,1.8600996,3.720199,5.580299,7.440398,9.300498,9.610515,9.920531,10.230548,10.540565,10.850581,11.506873,12.164979,12.823084,13.479377,14.137483,12.9427395,11.747997,10.553255,9.3567,8.161958,7.690587,7.217404,6.7442207,6.2728505,5.7996674,6.497658,7.1956487,7.891826,8.589817,9.287807,9.539809,9.791811,10.045626,10.297627,10.549629,10.843329,11.135216,11.427103,11.720803,12.012691,12.271944,12.5330105,12.792264,13.05333,13.312584,13.557334,13.802084,14.046834,14.293397,14.538147,14.719443,14.902553,15.085662,15.266958,15.4500675,15.359419,15.270584,15.179935,15.089288,15.000452,15.161806,15.324973,15.488139,15.649493,15.812659,15.899682,15.986704,16.075539,16.162561,16.249584,16.109985,15.970387,15.83079,15.689378,15.54978,15.687565,15.825351,15.963136,16.099108,16.236893,16.566853,16.89681,17.22677,17.55673,17.886688,18.120562,18.352621,18.584679,18.816738,19.050611,19.920834,20.789242,21.659464,22.529686,23.399908,23.318325,23.234928,23.151533,23.069948,22.986553,23.882156,24.77776,25.673363,26.567154,27.462757,28.6158,29.767033,30.920076,32.07312,33.224354,33.683033,34.1399,34.596764,35.055443,35.51231,36.190357,36.866592,37.544643,38.22269,38.900738,38.11754,37.33434,36.55295,35.769753,34.988365,35.240368,35.492367,35.74437,35.998184,36.250187,35.341892,34.43541,33.52712,32.620636,31.712341,30.8675,30.022661,29.17782,28.33298,27.488138,29.058165,30.62819,32.198215,33.76824,35.33827,35.392654,35.447044,35.503246,35.557636,35.612022,35.671852,35.731678,35.79332,35.85315,35.912975,31.541924,27.172684,22.80163,18.43239,14.06315,17.567608,21.072063,24.578333,28.08279,31.587248,26.922495,22.257742,17.592989,12.928236,8.26167,7.987913,7.7123427,7.4367723,7.1630154,6.887445,5.6455655,4.401873,3.159994,1.9181144,0.6744221,1.1095331,1.5446441,1.9797552,2.4148662,2.8499773,3.73289,4.615803,5.4969025,6.379815,7.262728,5.859495,4.458075,3.054842,1.651609,0.25018883,0.36984438,0.4894999,0.6091554,0.7306239,0.85027945,0.8375887,0.824898,0.8122072,0.7995165,0.7868258,1.3724127,1.9579996,2.5417736,3.1273603,3.7129474,3.4301252,3.147303,2.864481,2.5816586,2.3006494,2.4076142,2.514579,2.6233568,2.7303216,2.8372865,2.6142921,2.3931105,2.1701162,1.9471219,1.7241274,1.452183,1.1802386,0.90829426,0.6345369,0.36259252,1.7821422,3.2016919,4.6230545,6.0426044,7.462154,8.069496,8.676839,9.284182,9.893337,10.500679,9.189907,7.8809485,6.5701766,5.2594047,3.9504454,3.4065566,2.864481,2.322405,1.7803292,1.2382535,0.9916905,0.7469406,0.50219065,0.2574407,0.012690738,0.4894999,0.968122,1.4449311,1.9217403,2.4003625,2.1954978,1.9906329,1.7857682,1.5809034,1.3742256,1.3397794,1.305333,1.2708868,1.2346275,1.2001812,1.1222239,1.0442665,0.968122,0.8901646,0.8122072,1.3379664,1.8619126,2.3876717,2.911618,3.437377,3.3140955,3.1926272,3.0693457,2.9478772,2.8245957,2.619731,2.4148662,2.2100015,2.0051367,1.8002719,2.0450218,2.2897718,2.5345216,2.7792716,3.0258346,2.7575161,2.4891977,2.222692,1.9543737,1.6878681,1.3742256,1.062396,0.7505665,0.43692398,0.12509441,0.31726846,0.5094425,0.7016165,0.89560354,1.0877775,1.6080978,2.126605,2.6469254,3.1672456,3.6875658,3.3702974,3.053029,2.7357605,2.4166791,2.0994108,1.6896812,1.2799516,0.87022203,0.4604925,0.05076295,0.07433146,0.099712946,0.12509441,0.15047589,0.17585737,0.23024625,0.28463513,0.34083697,0.39522585,0.44961473,0.36077955,0.27013144,0.1794833,0.09064813,0.0,0.0,0.0,0.0,0.0,0.0,0.034446288,0.07070554,0.10515183,0.13959812,0.17585737,0.15228885,0.13053331,0.10696479,0.08520924,0.06164073,0.17585737,0.28826106,0.40066472,0.51306844,0.62547207,0.5275721,0.42967212,0.33177215,0.23568514,0.13778515,0.46955732,0.8031424,1.1349145,1.4666867,1.8002719,1.4394923,1.0805258,0.7197462,0.36077955,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.23931105,0.48043507,0.7197462,0.96087015,1.2001812,3.6005437,5.999093,8.399456,10.799818,13.200181,10.669285,8.140202,5.6093063,3.0802233,0.5493277,0.9481794,1.3452182,1.742257,2.1392958,2.5381477,2.1392958,1.742257,1.3452182,0.9481794,0.5493277,0.4405499,0.32995918,0.21936847,0.11059072,0.0,0.21030366,0.42060733,0.630911,0.83940166,1.0497054,0.87022203,0.69073874,0.5094425,0.32995918,0.15047589,0.4749962,0.7995165,1.1258497,1.4503701,1.7748904,1.4195497,1.064209,0.7106813,0.35534066,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.072518505,0.09427405,0.11784257,0.13959812,0.16316663,0.13959812,0.11784257,0.09427405,0.072518505,0.05076295,0.065266654,0.07977036,0.09427405,0.11059072,0.12509441,0.15228885,0.1794833,0.20667773,0.23568514,0.26287958,0.23024625,0.19761293,0.16497959,0.13234627,0.099712946,0.09064813,0.07977036,0.07070554,0.059827764,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.052575916,0.054388877,0.058014803,0.059827764,0.06164073,0.0870222,0.11240368,0.13778515,0.16316663,0.18673515,0.20486477,0.2229944,0.23931105,0.2574407,0.2755703,0.32814622,0.38072214,0.43329805,0.48587397,0.53663695,0.5058166,0.47318324,0.4405499,0.40791658,0.37528324,0.33539808,0.2955129,0.25562772,0.21574254,0.17585737,0.15954071,0.14503701,0.13053331,0.11421664,0.099712946,0.09064813,0.07977036,0.07070554,0.059827764,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,4.499773,4.788034,5.0744824,5.3627434,5.6491914,5.9374523,5.1741953,4.4127507,3.6494937,2.8880494,2.124792,2.9243085,3.7256382,4.5251546,5.3246713,6.1241875,6.9490857,7.7757964,8.600695,9.425592,10.25049,9.525306,8.80012,8.074935,7.3497505,6.624565,6.6499467,6.6753283,6.70071,6.7242785,6.7496595,6.7134004,6.6753283,6.637256,6.599184,6.5629244,7.28811,8.013294,8.736667,9.461852,10.1870365,11.037316,11.887595,12.737875,13.588155,14.436621,13.7875805,13.136727,12.487686,11.836833,11.187792,11.024626,10.863272,10.700105,10.536939,10.375585,13.113158,15.850732,18.588305,21.325878,24.06164,24.224806,24.387972,24.549326,24.712494,24.87566,20.437527,15.999394,11.563075,7.124943,2.6868105,2.1882458,1.6878681,1.1874905,0.6871128,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.6000906,1.2001812,1.8002719,2.4003625,3.000453,2.8245957,2.6505513,2.474694,2.3006494,2.124792,1.7005589,1.2745126,0.85027945,0.42423326,0.0,0.6871128,1.3742256,2.0631514,2.7502642,3.437377,2.7992141,2.1628644,1.5247015,0.8883517,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.0,0.0,0.0,0.0,0.0,2.2118144,4.4254417,6.637256,8.8508835,11.062697,11.325577,11.586644,11.849524,12.112403,12.375282,12.92461,13.475751,14.025079,14.574407,15.125546,13.562773,11.999999,10.437225,8.874452,7.311678,7.02523,6.736969,6.450521,6.16226,5.8758116,6.6753283,7.474845,8.274362,9.07569,9.875207,10.025683,10.174346,10.324821,10.475298,10.625773,10.7871275,10.950294,11.111648,11.274815,11.437981,11.813264,12.186734,12.562017,12.937301,13.312584,13.412297,13.512011,13.611723,13.713249,13.812962,14.0867195,14.362289,14.63786,14.911617,15.187187,15.087475,14.9877615,14.888049,14.788336,14.68681,14.788336,14.888049,14.9877615,15.087475,15.187187,15.399304,15.613234,15.825351,16.037468,16.249584,16.162561,16.075539,15.986704,15.899682,15.812659,15.950445,16.08823,16.224201,16.361988,16.499773,16.92582,17.350052,17.774284,18.20033,18.624565,18.49947,18.374376,18.24928,18.124187,18.000906,18.287354,18.575615,18.862062,19.150324,19.436771,19.262728,19.08687,18.912827,18.736969,18.562923,19.975222,21.38752,22.799818,24.212114,25.624413,27.049402,28.47439,29.89938,31.324368,32.749355,33.287807,33.824444,34.362892,34.89953,35.43798,36.375282,37.312584,38.249886,39.187187,40.12449,39.424683,38.72488,38.025078,37.325275,36.62547,36.850277,37.075085,37.299892,37.5247,37.749508,36.750565,35.74981,34.750866,33.75011,32.749355,31.69965,30.649946,29.60024,28.550535,27.50083,28.68832,29.87581,31.063301,32.25079,33.438282,33.875206,34.31213,34.750866,35.18779,35.624714,36.050762,36.474995,36.899227,37.325275,37.749508,32.925213,28.10092,23.274813,18.45052,13.6244135,18.062546,22.500679,26.936998,31.37513,35.813263,30.100618,24.387972,18.675327,12.962683,7.250037,7.1883965,7.124943,7.063302,6.9998484,6.9382076,5.5494785,4.162562,2.7756457,1.3869164,0.0,0.7124943,1.4249886,2.137483,2.8499773,3.5624714,4.461701,5.3627434,6.261973,7.1630154,8.062244,6.4759026,4.8877473,3.299592,1.7132497,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.07433146,0.15047589,0.22480737,0.2991388,0.37528324,1.0750868,1.7748904,2.474694,3.1744974,3.874301,3.4627585,3.049403,2.6378605,2.2245052,1.8129625,1.938057,2.0631514,2.1882458,2.3133402,2.4366217,2.1501737,1.8619126,1.5754645,1.2872034,1.0007553,0.7995165,0.6000906,0.40066472,0.19942589,0.0,1.6117238,3.2252605,4.836984,6.450521,8.062244,8.861761,9.663091,10.462607,11.262123,12.06164,10.29944,8.537241,6.775041,5.0128417,3.2506418,2.811905,2.374981,1.938057,1.49932,1.062396,0.85027945,0.63816285,0.42423326,0.21211663,0.0,0.6000906,1.2001812,1.8002719,2.4003625,3.000453,2.7375734,2.474694,2.2118144,1.9507477,1.6878681,1.6371052,1.5881553,1.5373923,1.4866294,1.4376793,1.1747998,0.9119202,0.6508536,0.387974,0.12509441,0.43692398,0.7505665,1.062396,1.3742256,1.6878681,1.7495089,1.8129625,1.8746033,1.938057,1.9996977,2.0123885,2.0250793,2.03777,2.0504606,2.0631514,2.03777,2.0123885,1.987007,1.9616255,1.938057,1.6008459,1.261822,0.9246109,0.5873999,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.7505665,1.3125849,1.8746033,2.4366217,3.000453,2.7756457,2.5508385,2.324218,2.0994108,1.8746033,1.5120108,1.1494182,0.7868258,0.42423326,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.19942589,0.2755703,0.34990177,0.42423326,0.50037766,0.40066472,0.2991388,0.19942589,0.099712946,0.0,0.0,0.0,0.0,0.0,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.16316663,0.13778515,0.11240368,0.0870222,0.06164073,0.19942589,0.33721104,0.4749962,0.61278135,0.7505665,0.61278135,0.4749962,0.33721104,0.19942589,0.06164073,0.50037766,0.93730164,1.3742256,1.8129625,2.2498865,1.8002719,1.3506571,0.89922947,0.44961473,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.2991388,0.6000906,0.89922947,1.2001812,1.49932,4.499773,7.500226,10.500679,13.499319,16.499773,13.299893,10.100015,6.9001355,3.7002566,0.50037766,0.40066472,0.2991388,0.19942589,0.099712946,0.0,0.13778515,0.2755703,0.41335547,0.5493277,0.6871128,0.5493277,0.41335547,0.2755703,0.13778515,0.0,0.26287958,0.52575916,0.7868258,1.0497054,1.3125849,1.0497054,0.7868258,0.52575916,0.26287958,0.0,0.34990177,0.69980353,1.0497054,1.3996071,1.7495089,1.3996071,1.0497054,0.69980353,0.34990177,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.0870222,0.11240368,0.13778515,0.16316663,0.18673515,0.16316663,0.13778515,0.11240368,0.0870222,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.16316663,0.19942589,0.2374981,0.2755703,0.31182957,0.2755703,0.2374981,0.19942589,0.16316663,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.0870222,0.11240368,0.13778515,0.16316663,0.18673515,0.21211663,0.2374981,0.26287958,0.28826106,0.31182957,0.37528324,0.43692398,0.50037766,0.5620184,0.62547207,0.5873999,0.5493277,0.51306844,0.4749962,0.43692398,0.387974,0.33721104,0.28826106,0.2374981,0.18673515,0.17585737,0.16316663,0.15047589,0.13778515,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,4.5251546,4.74271,4.9602656,5.177821,5.3953767,5.612932,5.0146546,4.41819,3.8199122,3.2216346,2.6251698,3.199879,3.774588,4.349297,4.9258194,5.5005283,6.2801023,7.059676,7.83925,8.620637,9.400211,8.907085,8.415772,7.9226465,7.4295206,6.9382076,6.9055743,6.872941,6.8403077,6.8076744,6.775041,6.813113,6.849373,6.887445,6.925517,6.9617763,7.7340984,8.508233,9.280556,10.052877,10.825199,11.4416065,12.059827,12.678047,13.294455,13.912675,13.318023,12.7233715,12.126906,11.532255,10.937603,11.062697,11.187792,11.312886,11.437981,11.563075,15.147303,18.73153,22.31757,25.901796,29.487837,28.037466,26.587097,25.136726,23.68817,22.237799,18.660824,15.082036,11.50506,7.9280853,4.349297,3.5117085,2.675933,1.8383441,1.0007553,0.16316663,0.1794833,0.19761293,0.21574254,0.23205921,0.25018883,0.69255173,1.1349145,1.5772774,2.0196402,2.4620032,2.3097143,2.1574254,2.0051367,1.8528478,1.7005589,1.5156367,1.3307146,1.1457924,0.96087015,0.774135,1.2418793,1.7096237,2.1773682,2.6451125,3.1128569,2.5308957,1.9471219,1.3651608,0.78319985,0.19942589,0.16316663,0.12509441,0.0870222,0.05076295,0.012690738,0.5148814,1.017072,1.5192627,2.0232663,2.525457,4.177066,5.8304877,7.4820967,9.135518,10.7871275,11.302009,11.81689,12.331772,12.846653,13.363347,13.495693,13.628039,13.760386,13.892733,14.025079,12.732436,11.439794,10.147152,8.854509,7.5618668,7.3950744,7.228282,7.059676,6.892884,6.7242785,7.2917356,7.859193,8.42665,8.994107,9.563377,9.9422865,10.323009,10.701918,11.082641,11.463363,11.789696,12.117842,12.444175,12.772322,13.100468,13.345218,13.589968,13.834718,14.079468,14.324218,14.289771,14.255324,14.220879,14.184619,14.150173,14.293397,14.434808,14.5780325,14.719443,14.862667,14.715817,14.567154,14.420304,14.271642,14.124791,14.255324,14.385859,14.514579,14.645112,14.775645,14.777458,14.779271,14.782897,14.78471,14.788336,14.929747,15.072971,15.214382,15.357606,15.50083,15.749206,15.999394,16.249584,16.499773,16.749962,17.192324,17.634687,18.07705,18.519413,18.961775,18.691645,18.423326,18.153194,17.883062,17.612932,17.939264,18.26741,18.595556,18.92189,19.250036,18.998035,18.74422,18.492218,18.240217,17.988214,19.099562,20.212719,21.325878,22.437225,23.550385,25.412296,27.27421,29.137934,30.999847,32.86176,33.287807,33.71204,34.138084,34.562317,34.988365,35.68998,36.391598,37.095028,37.796642,38.500072,38.157425,37.814774,37.472122,37.129475,36.786823,37.147602,37.508385,37.867348,38.22813,38.587097,37.424988,36.26288,35.10077,33.936848,32.77474,31.770357,30.764162,29.75978,28.7554,27.749205,28.91494,30.080675,31.244596,32.41033,33.574253,34.390087,35.20411,36.01994,36.835773,37.649796,36.922794,36.195797,35.466988,34.73999,34.012993,30.294605,26.578032,22.859646,19.143072,15.4246855,19.482096,23.539507,27.596916,31.654327,35.71174,29.815983,23.918415,18.019035,12.123281,6.2257137,6.3218007,6.4197006,6.5176005,6.6155005,6.7134004,5.4969025,4.2822175,3.0675328,1.8528478,0.63816285,1.261822,1.887294,2.5127661,3.1382382,3.7618973,4.3003473,4.836984,5.375434,5.9120708,6.450521,5.179634,3.9105604,2.6396735,1.3705997,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.059827764,0.11965553,0.1794833,0.23931105,0.2991388,0.8629702,1.4249886,1.987007,2.5508385,3.1128569,2.8028402,2.4928236,2.182807,1.8727903,1.5627737,1.6642996,1.7676386,1.8691645,1.9725033,2.0758421,1.8202144,1.5645868,1.310772,1.0551442,0.7995165,0.6399758,0.48043507,0.3208944,0.15954071,0.0,1.2908293,2.5798457,3.870675,5.1596913,6.450521,7.574558,8.700407,9.824444,10.950294,12.07433,10.681975,9.28962,7.897265,6.5049095,5.1125546,4.519716,3.926877,3.3358512,2.7430124,2.1501737,1.7821422,1.4141108,1.0478923,0.67986095,0.31182957,0.7469406,1.1820517,1.6171626,2.0522738,2.4873846,2.2607644,2.032331,1.8057107,1.5772774,1.3506571,1.3651608,1.3796645,1.3941683,1.4104849,1.4249886,1.214685,1.0043813,0.79589057,0.5855869,0.37528324,0.57833505,0.7795739,0.9826257,1.1856775,1.3869164,1.4304274,1.4721256,1.5156367,1.5573349,1.6008459,1.6117238,1.6244144,1.6371052,1.649796,1.6624867,1.7295663,1.7966459,1.8655385,1.9326181,1.9996977,1.6642996,1.3307146,0.99531645,0.65991837,0.3245203,0.25925365,0.19579996,0.13053331,0.065266654,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.6055295,1.0605831,1.5156367,1.9706904,2.4257438,2.3169663,2.2100015,2.1030366,1.9942589,1.887294,1.5301404,1.1729867,0.81583315,0.45686656,0.099712946,0.099712946,0.099712946,0.099712946,0.099712946,0.099712946,0.16316663,0.22480737,0.28826106,0.34990177,0.41335547,0.32995918,0.24837588,0.16497959,0.08339628,0.0,0.0,0.0,0.0,0.0,0.0,0.032633327,0.065266654,0.09789998,0.13053331,0.16316663,0.14322405,0.12328146,0.10333887,0.08339628,0.06164073,0.18310922,0.30276474,0.4224203,0.5420758,0.66173136,0.6200332,0.57833505,0.53482395,0.49312583,0.44961473,0.726998,1.0043813,1.2817645,1.5591478,1.8383441,1.5899682,1.3434052,1.0950294,0.8466535,0.6000906,0.48587397,0.36984438,0.25562772,0.13959812,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.24293698,0.48587397,0.726998,0.969935,1.2128719,4.4870825,7.763106,11.037316,14.313339,17.58755,14.545399,11.503247,8.459284,5.4171324,2.374981,1.9054236,1.4358664,0.9644961,0.4949388,0.025381476,0.20486477,0.38434806,0.5656443,0.7451276,0.9246109,0.79226464,0.65991837,0.5275721,0.39522585,0.26287958,0.8103943,1.357909,1.9054236,2.4529383,3.000453,2.6070402,2.2154403,1.8220274,1.4304274,1.0370146,1.1095331,1.1820517,1.2545701,1.3270886,1.3996071,1.1204109,0.83940166,0.56020546,0.27919623,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.072518505,0.09427405,0.11784257,0.13959812,0.16316663,0.13959812,0.11784257,0.09427405,0.072518505,0.05076295,0.065266654,0.07977036,0.09427405,0.11059072,0.12509441,0.18673515,0.25018883,0.31182957,0.37528324,0.43692398,0.3825351,0.32814622,0.27194437,0.21755551,0.16316663,0.14503701,0.12690738,0.11059072,0.092461094,0.07433146,0.072518505,0.07070554,0.06707962,0.065266654,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.032633327,0.052575916,0.072518505,0.092461094,0.11240368,0.11421664,0.11784257,0.11965553,0.12328146,0.12509441,0.13234627,0.13959812,0.14684997,0.15410182,0.16316663,0.18492219,0.20667773,0.23024625,0.2520018,0.2755703,0.32995918,0.38434806,0.4405499,0.4949388,0.5493277,0.52575916,0.50037766,0.4749962,0.44961473,0.42423326,0.61459434,0.80495536,0.99531645,1.1856775,1.3742256,1.1457924,0.9155461,0.6852999,0.4550536,0.22480737,0.19942589,0.17585737,0.15047589,0.12509441,0.099712946,0.08520924,0.07070554,0.054388877,0.03988518,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,4.550536,4.6973863,4.844236,4.992899,5.139749,5.2865987,4.855114,4.421816,3.9903307,3.5570326,3.1255474,3.4754493,3.825351,4.175253,4.5251546,4.8750563,5.6093063,6.345369,7.079619,7.8156815,8.549932,8.290678,8.029612,7.7703576,7.509291,7.250037,7.159389,7.0705543,6.979906,6.889258,6.8004227,6.9128265,7.02523,7.137634,7.250037,7.362441,8.1819,9.003172,9.822631,10.642091,11.463363,11.847711,12.232059,12.618219,13.002567,13.386916,12.846653,12.308203,11.7679405,11.227677,10.687414,11.10077,11.512312,11.925668,12.337211,12.750566,17.18326,21.61414,26.046833,30.479527,34.91222,31.850126,28.788033,25.724127,22.662033,19.59994,16.882307,14.164677,11.447045,8.729415,6.011784,4.836984,3.6621845,2.4873846,1.3125849,0.13778515,0.21030366,0.28282216,0.35534066,0.42785916,0.50037766,0.7850128,1.0696479,1.3542831,1.6407311,1.9253663,1.794833,1.6642996,1.5355793,1.405046,1.2745126,1.3307146,1.3851035,1.4394923,1.4956942,1.550083,1.7966459,2.0450218,2.2933977,2.5399606,2.7883365,2.2607644,1.7331922,1.2056202,0.678048,0.15047589,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,1.0297627,2.034144,3.0403383,4.0447197,5.050914,6.1423173,7.2355337,8.326937,9.420154,10.51337,11.280253,12.047136,12.815832,13.582716,14.349599,14.064963,13.780329,13.495693,13.209246,12.92461,11.9021,10.879588,9.857078,8.834567,7.8120556,7.764919,7.7177815,7.6706448,7.6216946,7.574558,7.909956,8.245354,8.580752,8.914337,9.249735,9.860703,10.469859,11.080828,11.689982,12.299138,12.792264,13.28539,13.776703,14.269829,14.762955,14.877171,14.9932,15.107417,15.221634,15.337664,15.167245,14.996826,14.828221,14.657803,14.487384,14.498261,14.507326,14.518205,14.527269,14.538147,14.342347,14.14836,13.95256,13.75676,13.562773,13.722314,13.881854,14.043208,14.202749,14.362289,14.155612,13.947122,13.740443,13.531953,13.325275,13.696932,14.070402,14.4420595,14.81553,15.187187,15.54978,15.912373,16.274965,16.637558,17.00015,17.460642,17.919323,18.379814,18.840307,19.3008,18.885632,18.470463,18.055294,17.640125,17.224958,17.592989,17.959208,18.327238,18.69527,19.063301,18.733343,18.403383,18.071611,17.741652,17.411694,18.225714,19.03792,19.850128,20.662334,21.474543,23.77519,26.074028,28.374678,30.675327,32.974163,33.287807,33.599636,33.913277,34.22511,34.536938,35.00468,35.472427,35.94017,36.407913,36.87566,36.890163,36.904667,36.91917,36.935486,36.94999,37.44493,37.93987,38.434807,38.929745,39.424683,38.099407,36.775948,35.450672,34.125393,32.800117,31.839249,30.880192,29.919321,28.960264,27.999393,29.143373,30.28554,31.427706,32.569874,33.71204,34.90497,36.097897,37.29083,38.481945,39.674873,37.79483,35.914787,34.034748,32.154705,30.274662,27.66581,25.055143,22.444477,19.835623,17.224958,20.901646,24.580147,28.256834,31.935335,35.612022,29.529535,23.447044,17.364555,11.282066,5.199577,5.4570174,5.714458,5.9718986,6.2293396,6.48678,5.4443264,4.401873,3.3594196,2.3169663,1.2745126,1.8129625,2.3495996,2.8880494,3.4246864,3.9631362,4.137181,4.313038,4.4870825,4.6629395,4.836984,3.8851788,2.9333735,1.9797552,1.0279498,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.045324065,0.09064813,0.13415924,0.1794833,0.22480737,0.6508536,1.0750868,1.49932,1.9253663,2.3495996,2.1429217,1.9344311,1.7277533,1.5192627,1.3125849,1.3923552,1.4721256,1.551896,1.6316663,1.7132497,1.4902552,1.2672608,1.0442665,0.823085,0.6000906,0.48043507,0.36077955,0.23931105,0.11965553,0.0,0.968122,1.9344311,2.902553,3.870675,4.836984,6.2873545,7.7377243,9.188094,10.636651,12.087022,11.06451,10.042,9.019489,7.996978,6.9744673,6.2275267,5.480586,4.7318325,3.9848917,3.2379513,2.715818,2.1918716,1.6697385,1.1476053,0.62547207,0.89560354,1.1657349,1.4358664,1.7041848,1.9743162,1.7821422,1.5899682,1.3977941,1.2056202,1.0116332,1.0932164,1.1729867,1.2527572,1.3325275,1.4122978,1.2545701,1.0968424,0.93911463,0.78319985,0.62547207,0.7179332,0.8103943,0.90285534,0.99531645,1.0877775,1.1095331,1.1331016,1.1548572,1.1766127,1.2001812,1.2128719,1.2255627,1.2382535,1.2491312,1.261822,1.4231756,1.5827163,1.742257,1.9017978,2.0631514,1.7295663,1.3977941,1.064209,0.7324369,0.40066472,0.3208944,0.23931105,0.15954071,0.07977036,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.4604925,0.80676836,1.1548572,1.502946,1.8492218,1.8600996,1.8691645,1.8800422,1.889107,1.8999848,1.54827,1.1947423,0.8430276,0.4894999,0.13778515,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.12509441,0.17585737,0.22480737,0.2755703,0.3245203,0.25925365,0.19579996,0.13053331,0.065266654,0.0,0.0,0.0,0.0,0.0,0.0,0.027194439,0.054388877,0.08339628,0.11059072,0.13778515,0.12328146,0.10696479,0.092461094,0.07795739,0.06164073,0.16497959,0.26831847,0.36984438,0.47318324,0.5747091,0.62728506,0.67986095,0.7324369,0.7850128,0.8375887,0.9554313,1.0732739,1.1893034,1.3071461,1.4249886,1.3796645,1.3343405,1.2908293,1.2455053,1.2001812,0.969935,0.73968875,0.5094425,0.27919623,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.18492219,0.36984438,0.55476654,0.73968875,0.9246109,4.4743915,8.024173,11.575767,15.125546,18.675327,15.789091,12.904668,10.020245,7.135821,4.249584,3.4101827,2.570781,1.7295663,0.8901646,0.05076295,0.27194437,0.4949388,0.7179332,0.93911463,1.162109,1.0352017,0.90829426,0.7795739,0.6526665,0.52575916,1.357909,2.1900587,3.0222087,3.8543584,4.688321,4.164375,3.6422417,3.1201086,2.5979755,2.0758421,1.8691645,1.6642996,1.4594349,1.2545701,1.0497054,0.83940166,0.630911,0.42060733,0.21030366,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.058014803,0.07795739,0.09789998,0.11784257,0.13778515,0.11784257,0.09789998,0.07795739,0.058014803,0.038072214,0.054388877,0.072518505,0.09064813,0.10696479,0.12509441,0.21211663,0.2991388,0.387974,0.4749962,0.5620184,0.4894999,0.4169814,0.3444629,0.27194437,0.19942589,0.17767033,0.15410182,0.13234627,0.11059072,0.0870222,0.08339628,0.07795739,0.072518505,0.06707962,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.052575916,0.07977036,0.10696479,0.13415924,0.16316663,0.16679256,0.17223145,0.17767033,0.18310922,0.18673515,0.17767033,0.16679256,0.15772775,0.14684997,0.13778515,0.15772775,0.17767033,0.19761293,0.21755551,0.2374981,0.28463513,0.33177215,0.38072214,0.42785916,0.4749962,0.46230546,0.44961473,0.43692398,0.42423326,0.41335547,0.8430276,1.2726997,1.7023718,2.132044,2.561716,2.1157274,1.6679256,1.2201238,0.77232206,0.3245203,0.28826106,0.25018883,0.21211663,0.17585737,0.13778515,0.11965553,0.10333887,0.08520924,0.06707962,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,4.574105,4.652062,4.7300196,4.8079767,4.8841214,4.9620786,4.695573,4.4272547,4.160749,3.8924308,3.6241121,3.7492065,3.874301,3.9993954,4.12449,4.249584,4.940323,5.6292486,6.319988,7.0107265,7.699652,7.6724577,7.645263,7.6180687,7.590874,7.5618668,7.415017,7.268167,7.119504,6.972654,6.825804,7.0125394,7.1992745,7.3878226,7.574558,7.763106,8.629702,9.498111,10.364707,11.233116,12.099712,12.252001,12.40429,12.558392,12.710681,12.862969,12.377095,11.893035,11.407161,10.9230995,10.437225,11.137029,11.836833,12.536636,13.238253,13.938056,19.217403,24.49675,29.77791,35.05726,40.336605,35.66279,30.987156,26.311525,21.637709,16.962078,15.105604,13.247317,11.390844,9.5325575,7.6742706,6.16226,4.650249,3.1382382,1.6244144,0.11240368,0.23931105,0.3680314,0.4949388,0.62184614,0.7505665,0.8774739,1.0043813,1.1331016,1.260009,1.3869164,1.2799516,1.1729867,1.064209,0.9572442,0.85027945,1.1457924,1.4394923,1.7350051,2.030518,2.324218,2.3532255,2.38042,2.4076142,2.4348087,2.4620032,1.9906329,1.5174497,1.0442665,0.5728962,0.099712946,0.0870222,0.07433146,0.06164073,0.05076295,0.038072214,1.5446441,3.053029,4.559601,6.0679855,7.574558,8.107569,8.640579,9.171778,9.704789,10.2378,11.256684,12.277383,13.29808,14.316965,15.337664,14.634234,13.932617,13.229188,12.527572,11.8241415,11.071762,10.319383,9.567003,8.814624,8.062244,8.134763,8.207282,8.2798,8.352319,8.424837,8.528176,8.629702,8.733041,8.834567,8.937905,9.7773075,10.616709,11.457924,12.297325,13.136727,13.794832,14.452938,15.10923,15.767336,16.425442,16.409124,16.39462,16.380117,16.365614,16.349297,16.04472,15.740141,15.435563,15.129172,14.824595,14.703127,14.579845,14.458377,14.335095,14.211814,13.97069,13.727753,13.484816,13.2418785,13.000754,13.189302,13.379663,13.5700245,13.760386,13.9507475,13.531953,13.114971,12.697989,12.279196,11.862214,12.464118,13.067834,13.669738,14.271642,14.875358,15.350354,15.825351,16.300346,16.775343,17.25034,17.727148,18.20577,18.682579,19.15939,19.63801,19.077805,18.5176,17.957394,17.397188,16.836983,17.2449,17.652817,18.060734,18.466837,18.874754,18.466837,18.060734,17.652817,17.2449,16.836983,17.350052,17.863121,18.374376,18.887444,19.400513,22.138086,24.87566,27.613234,30.350807,33.08838,33.287807,33.487232,33.686657,33.887897,34.087322,34.31938,34.553253,34.785313,35.017372,35.24943,35.622902,35.99456,36.36803,36.739685,37.113155,37.742256,38.373165,39.002266,39.633175,40.26227,38.775642,37.2872,35.80057,34.31213,32.8255,31.909954,30.994408,30.080675,29.165129,28.249582,29.369993,30.490404,31.610815,32.729412,33.849823,35.41985,36.989876,38.559902,40.12993,41.69995,38.666866,35.635593,32.602505,29.56942,26.538147,25.0352,23.532255,22.029308,20.528175,19.025229,22.323008,25.620787,28.916754,32.21453,35.51231,29.2449,22.977488,16.710075,10.442664,4.175253,4.592234,5.009216,5.42801,5.844991,6.261973,5.391751,4.5233417,3.6531196,2.7828975,1.9126755,2.3622901,2.811905,3.2633326,3.7129474,4.162562,3.975827,3.787279,3.6005437,3.4119956,3.2252605,2.5907235,1.9543737,1.3198367,0.6852999,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.43692398,0.72518504,1.0116332,1.2998942,1.5881553,1.4830034,1.3778516,1.2726997,1.167548,1.062396,1.1204109,1.1766127,1.2346275,1.2926424,1.3506571,1.1602961,0.969935,0.7795739,0.58921283,0.40066472,0.3208944,0.23931105,0.15954071,0.07977036,0.0,0.64541465,1.2908293,1.9344311,2.5798457,3.2252605,5.0001507,6.775041,8.549932,10.324821,12.099712,11.447045,10.794379,10.141713,9.490859,8.838193,7.935337,7.0324817,6.1296263,5.2267714,4.325729,3.6476808,2.9696326,2.2915847,1.6153497,0.93730164,1.0424535,1.1476053,1.2527572,1.357909,1.4630609,1.305333,1.1476053,0.9898776,0.8321498,0.6744221,0.8194591,0.9644961,1.1095331,1.2545701,1.3996071,1.2944553,1.1893034,1.0841516,0.9808127,0.87566096,0.8575313,0.83940166,0.823085,0.80495536,0.7868258,0.7904517,0.79226464,0.79589057,0.79770356,0.7995165,0.8122072,0.824898,0.8375887,0.85027945,0.8629702,1.114972,1.3669738,1.6207886,1.8727903,2.124792,1.794833,1.4648738,1.1349145,0.80495536,0.4749962,0.38072214,0.28463513,0.19036107,0.09427405,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.3154555,0.55476654,0.79589057,1.0352017,1.2745126,1.403233,1.5301404,1.6570477,1.7857682,1.9126755,1.5645868,1.2183108,0.87022203,0.52213323,0.17585737,0.15047589,0.12509441,0.099712946,0.07433146,0.05076295,0.0870222,0.12509441,0.16316663,0.19942589,0.2374981,0.19036107,0.14322405,0.09427405,0.047137026,0.0,0.0,0.0,0.0,0.0,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.10333887,0.092461094,0.08339628,0.072518505,0.06164073,0.14684997,0.23205921,0.31726846,0.40247768,0.48768693,0.6345369,0.78319985,0.9300498,1.0768998,1.2255627,1.1820517,1.1403534,1.0968424,1.0551442,1.0116332,1.1693609,1.3270886,1.4848163,1.6425442,1.8002719,1.455809,1.1095331,0.7650702,0.42060733,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.12690738,0.25562772,0.3825351,0.5094425,0.63816285,4.463514,8.287052,12.112403,15.937754,19.763105,17.034595,14.3079,11.579392,8.852696,6.1241875,4.914942,3.7056956,2.4946365,1.2853905,0.07433146,0.34083697,0.6055295,0.87022203,1.1349145,1.3996071,1.2781386,1.1548572,1.0333886,0.9101072,0.7868258,1.9054236,3.0222087,4.1408067,5.2575917,6.3743763,5.7217097,5.0708566,4.41819,3.7655232,3.1128569,2.6306088,2.1483607,1.6642996,1.1820517,0.69980353,0.56020546,0.42060733,0.27919623,0.13959812,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.04169814,0.059827764,0.07795739,0.09427405,0.11240368,0.09427405,0.07795739,0.059827764,0.04169814,0.025381476,0.045324065,0.065266654,0.08520924,0.10515183,0.12509441,0.2374981,0.34990177,0.46230546,0.5747091,0.6871128,0.5982776,0.5076295,0.4169814,0.32814622,0.2374981,0.21030366,0.18310922,0.15410182,0.12690738,0.099712946,0.092461094,0.08520924,0.07795739,0.07070554,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.072518505,0.10696479,0.14322405,0.17767033,0.21211663,0.21936847,0.22662032,0.23568514,0.24293698,0.25018883,0.2229944,0.19579996,0.16679256,0.13959812,0.11240368,0.13053331,0.14684997,0.16497959,0.18310922,0.19942589,0.23931105,0.27919623,0.3208944,0.36077955,0.40066472,0.40066472,0.40066472,0.40066472,0.40066472,0.40066472,1.0696479,1.7404441,2.4094272,3.0802233,3.7492065,3.0856624,2.420305,1.7549478,1.0895905,0.42423326,0.37528324,0.3245203,0.2755703,0.22480737,0.17585737,0.15410182,0.13415924,0.11421664,0.09427405,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,4.599486,4.606738,4.615803,4.6230545,4.6303062,4.6375585,4.5342193,4.4326935,4.329355,4.227829,4.12449,4.024777,3.925064,3.825351,3.7256382,3.6241121,4.269527,4.914942,5.560356,6.205771,6.849373,7.0542374,7.2591023,7.46578,7.6706448,7.8755093,7.6706448,7.46578,7.2591023,7.0542374,6.849373,7.112252,7.3751316,7.6380115,7.900891,8.161958,9.077503,9.99305,10.906783,11.822329,12.737875,12.658105,12.578335,12.496751,12.416981,12.337211,11.907538,11.477866,11.048194,10.616709,10.1870365,11.175101,12.163166,13.149418,14.137483,15.125546,21.251547,27.37936,33.507175,39.634987,45.762802,39.47545,33.18809,26.898926,20.611572,14.324218,13.327088,12.329959,11.332829,10.3357,9.336758,7.4875355,5.638314,3.787279,1.938057,0.0870222,0.27013144,0.45324063,0.6345369,0.81764615,1.0007553,0.969935,0.93911463,0.9101072,0.8792868,0.85027945,0.7650702,0.67986095,0.5946517,0.5094425,0.42423326,0.96087015,1.4956942,2.030518,2.565342,3.100166,2.907992,2.715818,2.521831,2.3296568,2.137483,1.7205015,1.3017071,0.88472575,0.46774435,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,2.0595255,4.070101,6.0806766,8.089439,10.100015,10.07282,10.045626,10.016619,9.989424,9.96223,11.234929,12.507628,13.780329,15.053028,16.325727,15.2053175,14.084907,12.964496,11.844085,10.725487,10.243238,9.759177,9.27693,8.794682,8.312433,8.504607,8.696781,8.890768,9.082943,9.275117,9.144584,9.015862,8.885329,8.754796,8.624263,9.695724,10.765372,11.83502,12.904668,13.974316,14.7974,15.620485,16.441757,17.264843,18.087927,17.94289,17.797853,17.652817,17.50778,17.362743,16.922194,16.481644,16.042906,15.602356,15.161806,14.907991,14.652364,14.396736,14.142921,13.887294,13.597219,13.307145,13.017072,12.726997,12.436923,12.658105,12.877473,13.096842,13.318023,13.537392,12.910107,12.282822,11.655537,11.028252,10.399154,11.233116,12.065266,12.897416,13.729566,14.561715,15.149116,15.738328,16.325727,16.913128,17.500528,17.995466,18.490406,18.985344,19.480284,19.975222,19.26998,18.564737,17.859495,17.154251,16.450823,16.89681,17.344612,17.792416,18.240217,18.688019,18.202145,17.718082,17.23221,16.748148,16.262274,16.474392,16.68832,16.900436,17.112555,17.32467,20.499168,23.675478,26.849976,30.024473,33.200783,33.287807,33.37483,33.46185,33.550686,33.637707,33.635895,33.632267,33.630455,33.62683,33.625015,34.35564,35.084454,35.815075,36.5457,37.27451,38.03958,38.80465,39.56972,40.334793,41.09986,39.450066,37.80027,36.150475,34.50068,32.850883,31.98066,31.110437,30.240215,29.369993,28.499771,29.596615,30.695269,31.792112,32.890766,33.98761,35.93473,37.881855,39.830788,41.77791,43.725033,39.540714,35.354584,31.170265,26.984135,22.799818,22.404593,22.009365,21.61414,21.220728,20.8255,23.742558,26.659615,29.578484,32.49554,35.412598,28.960264,22.50793,16.055597,9.603263,3.149116,3.727451,4.305786,4.882308,5.4606433,6.037165,5.3391747,4.6429973,3.9450066,3.247016,2.5508385,2.911618,3.2742105,3.636803,3.9993954,4.361988,3.8126602,3.2633326,2.712192,2.1628644,1.6117238,1.2944553,0.97718686,0.65991837,0.34264994,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.22480737,0.37528324,0.52575916,0.6744221,0.824898,0.823085,0.8194591,0.81764615,0.81583315,0.8122072,0.8466535,0.88291276,0.91735905,0.95180535,0.9880646,0.83033687,0.6726091,0.5148814,0.35715362,0.19942589,0.15954071,0.11965553,0.07977036,0.03988518,0.0,0.32270733,0.64541465,0.968122,1.2908293,1.6117238,3.7129474,5.812358,7.911769,10.012992,12.112403,11.829581,11.546759,11.26575,10.982927,10.700105,9.643148,8.584378,7.5274205,6.4704633,5.411693,4.5795436,3.7473936,2.9152439,2.0830941,1.2491312,1.1893034,1.1294757,1.0696479,1.0098201,0.9499924,0.82671094,0.70524246,0.581961,0.4604925,0.33721104,0.5475147,0.75781834,0.968122,1.1766127,1.3869164,1.3343405,1.2817645,1.2291887,1.1766127,1.1258497,0.99712944,0.87022203,0.7433147,0.61459434,0.48768693,0.46955732,0.45324063,0.43511102,0.4169814,0.40066472,0.41335547,0.42423326,0.43692398,0.44961473,0.46230546,0.80676836,1.1530442,1.4975071,1.84197,2.1882458,1.8600996,1.5319533,1.2056202,0.8774739,0.5493277,0.4405499,0.32995918,0.21936847,0.11059072,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.17041849,0.30276474,0.43511102,0.56745726,0.69980353,0.9445535,1.1893034,1.4358664,1.6806163,1.9253663,1.5827163,1.2400664,0.8974165,0.55476654,0.21211663,0.17585737,0.13778515,0.099712946,0.06164073,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.0,0.0,0.0,0.0,0.0,0.018129626,0.034446288,0.052575916,0.07070554,0.0870222,0.08339628,0.07795739,0.072518505,0.06707962,0.06164073,0.13053331,0.19761293,0.26469254,0.33177215,0.40066472,0.6417888,0.88472575,1.1276628,1.3705997,1.6117238,1.4104849,1.2074331,1.0043813,0.8031424,0.6000906,0.96087015,1.3198367,1.6806163,2.039583,2.4003625,1.93987,1.4793775,1.020698,0.56020546,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07070554,0.13959812,0.21030366,0.27919623,0.34990177,4.4508233,8.549932,12.650853,16.749962,20.850883,18.280102,15.709321,13.140353,10.5695715,8.000604,6.4197006,4.84061,3.2597067,1.6806163,0.099712946,0.40791658,0.71430725,1.0225109,1.3307146,1.6371052,1.5192627,1.403233,1.2853905,1.167548,1.0497054,2.4529383,3.8543584,5.2575917,6.6608243,8.062244,7.2808576,6.497658,5.714458,4.933071,4.1498713,3.39024,2.6306088,1.8691645,1.1095331,0.34990177,0.27919623,0.21030366,0.13959812,0.07070554,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.027194439,0.04169814,0.058014803,0.072518505,0.0870222,0.072518505,0.058014803,0.04169814,0.027194439,0.012690738,0.034446288,0.058014803,0.07977036,0.10333887,0.12509441,0.26287958,0.40066472,0.53663695,0.6744221,0.8122072,0.70524246,0.5982776,0.4894999,0.3825351,0.2755703,0.24293698,0.21030366,0.17767033,0.14503701,0.11240368,0.10333887,0.092461094,0.08339628,0.072518505,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.092461094,0.13415924,0.17767033,0.21936847,0.26287958,0.27194437,0.28282216,0.291887,0.30276474,0.31182957,0.26831847,0.2229944,0.17767033,0.13234627,0.0870222,0.10333887,0.11784257,0.13234627,0.14684997,0.16316663,0.19579996,0.22662032,0.25925365,0.291887,0.3245203,0.33721104,0.34990177,0.36259252,0.37528324,0.387974,1.2980812,2.2081885,3.1182957,4.02659,4.936697,4.0555973,3.1726844,2.2897718,1.4068589,0.52575916,0.46230546,0.40066472,0.33721104,0.2755703,0.21211663,0.19036107,0.16679256,0.14503701,0.12328146,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,4.6248674,4.5632267,4.499773,4.4381323,4.3746786,4.313038,4.3746786,4.4381323,4.499773,4.5632267,4.6248674,4.3003473,3.975827,3.6494937,3.3249733,3.000453,3.6005437,4.2006345,4.800725,5.4008155,6.000906,6.43783,6.874754,7.311678,7.750415,8.187339,7.9244595,7.663393,7.400513,7.137634,6.874754,7.211965,7.549176,7.8882003,8.225411,8.562622,9.525306,10.487988,11.450671,12.413355,13.374225,13.062395,12.750566,12.436923,12.125093,11.813264,11.437981,11.062697,10.687414,10.312131,9.936848,11.213174,12.487686,13.762199,15.036712,16.313038,23.287504,30.26197,37.23825,44.21272,51.187187,43.28811,35.38722,27.488138,19.587248,11.6881695,11.5503845,11.4126,11.274815,11.137029,10.999244,8.812811,6.624565,4.4381323,2.2498865,0.06164073,0.2991388,0.53663695,0.774135,1.0116332,1.2491312,1.062396,0.87566096,0.6871128,0.50037766,0.31182957,0.25018883,0.18673515,0.12509441,0.06164073,0.0,0.774135,1.550083,2.324218,3.100166,3.874301,3.4627585,3.049403,2.6378605,2.2245052,1.8129625,1.4503701,1.0877775,0.72518504,0.36259252,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,2.5744069,5.087173,7.5999393,10.112705,12.625471,12.038072,11.450671,10.863272,10.275872,9.686659,11.213174,12.737875,14.262577,15.787278,17.31198,15.774588,14.237195,12.699803,11.162411,9.625018,9.412902,9.200785,8.9868555,8.774739,8.562622,8.874452,9.188094,9.499924,9.811753,10.125396,9.762803,9.400211,9.037619,8.675026,8.312433,9.612328,10.912222,12.212116,13.512011,14.811904,15.799969,16.788034,17.774284,18.76235,19.750414,19.474844,19.199274,18.925516,18.649946,18.374376,17.799667,17.224958,16.650248,16.075539,15.50083,15.112856,14.724882,14.336908,13.9507475,13.562773,13.225562,12.888351,12.549327,12.212116,11.874905,12.125093,12.375282,12.625471,12.87566,13.125849,12.28826,11.450671,10.613083,9.775495,8.937905,10.000301,11.062697,12.125093,13.1874895,14.249886,14.94969,15.649493,16.349297,17.050913,17.750717,18.261972,18.77504,19.288109,19.799364,20.312433,19.462152,18.611874,17.761595,16.913128,16.062849,16.550535,17.038223,17.52591,18.011784,18.49947,17.937452,17.375433,16.811602,16.249584,15.687565,15.600543,15.511708,15.4246855,15.337664,15.250641,18.862062,22.475298,26.08672,29.699953,33.313187,33.287807,33.262424,33.23704,33.211662,33.18809,32.950596,32.713097,32.475597,32.238102,32.000603,33.08838,34.174343,35.262123,36.3499,37.437675,38.336906,39.23795,40.13718,41.03822,41.93745,40.12449,38.31334,36.500374,34.687412,32.87445,32.049553,31.224655,30.399757,29.574858,28.74996,29.825047,30.900135,31.975222,33.05031,34.125393,36.44961,38.775642,41.09986,43.42589,45.75011,40.41275,35.075386,29.738026,24.400663,19.063301,19.775795,20.48829,21.200785,21.913279,22.625772,25.162107,27.700254,30.238403,32.77474,35.312885,28.675629,22.038374,15.399304,8.762048,2.124792,2.8626678,3.6005437,4.3384194,5.0744824,5.812358,5.2884116,4.762653,4.2368937,3.7129474,3.1871881,3.4627585,3.738329,4.0120864,4.2876563,4.5632267,3.6494937,2.7375734,1.8256533,0.9119202,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.16316663,0.26287958,0.36259252,0.46230546,0.5620184,0.5747091,0.5873999,0.6000906,0.61278135,0.62547207,0.50037766,0.37528324,0.25018883,0.12509441,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.4257438,4.8496747,7.2754188,9.699349,12.125093,12.212116,12.299138,12.387974,12.474996,12.562017,11.349146,10.138086,8.925215,7.7123427,6.4994707,5.5132194,4.5251546,3.53709,2.5508385,1.5627737,1.3379664,1.1131591,0.8883517,0.66173136,0.43692398,0.34990177,0.26287958,0.17585737,0.0870222,0.0,0.2755703,0.5493277,0.824898,1.1004683,1.3742256,1.3742256,1.3742256,1.3742256,1.3742256,1.3742256,1.1367276,0.89922947,0.66173136,0.42423326,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.50037766,0.93730164,1.3742256,1.8129625,2.2498865,1.9253663,1.6008459,1.2745126,0.9499924,0.62547207,0.50037766,0.37528324,0.25018883,0.12509441,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.48768693,0.85027945,1.2128719,1.5754645,1.938057,1.6008459,1.261822,0.9246109,0.5873999,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.11240368,0.16316663,0.21211663,0.26287958,0.31182957,0.6508536,0.9880646,1.3252757,1.6624867,1.9996977,1.6371052,1.2745126,0.9119202,0.5493277,0.18673515,0.7505665,1.3125849,1.8746033,2.4366217,3.000453,2.4257438,1.8492218,1.2745126,0.69980353,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,4.4381323,8.812811,13.1874895,17.562168,21.936848,19.525606,17.112555,14.699501,12.28826,9.875207,7.9244595,5.975525,4.024777,2.0758421,0.12509441,0.4749962,0.824898,1.1747998,1.5247015,1.8746033,1.7621996,1.649796,1.5373923,1.4249886,1.3125849,3.000453,4.688321,6.3743763,8.062244,9.750113,8.838193,7.9244595,7.0125394,6.1006193,5.186886,4.1498713,3.1128569,2.0758421,1.0370146,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.28826106,0.44961473,0.61278135,0.774135,0.93730164,0.8122072,0.6871128,0.5620184,0.43692398,0.31182957,0.2755703,0.2374981,0.19942589,0.16316663,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.11240368,0.16316663,0.21211663,0.26287958,0.31182957,0.3245203,0.33721104,0.34990177,0.36259252,0.37528324,0.31182957,0.25018883,0.18673515,0.12509441,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.15047589,0.17585737,0.19942589,0.22480737,0.25018883,0.2755703,0.2991388,0.3245203,0.34990177,0.37528324,1.5247015,2.675933,3.825351,4.974769,6.1241875,5.0255322,3.925064,2.8245957,1.7259403,0.62547207,0.5493277,0.4749962,0.40066472,0.3245203,0.25018883,0.22480737,0.19942589,0.17585737,0.15047589,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,4.499773,4.458075,4.4145637,4.3728657,4.329355,4.2876563,4.347484,4.407312,4.4671397,4.5269675,4.5867953,4.2967215,4.006647,3.7183862,3.4283123,3.1382382,3.6476808,4.157123,4.668379,5.177821,5.6872635,6.2782893,6.867502,7.456715,8.047741,8.636953,8.455658,8.272549,8.089439,7.9081426,7.7250338,8.040489,8.354132,8.669587,8.985043,9.300498,10.167094,11.035503,11.9021,12.770509,13.637105,13.234627,12.8321495,12.429671,12.027194,11.624716,11.242181,10.859646,10.477111,10.094576,9.712041,11.379966,13.047892,14.715817,16.38193,18.049856,24.652666,31.255474,37.858284,44.459282,51.06209,43.532856,36.003624,28.472578,20.94153,13.412297,12.5058155,11.597522,10.689227,9.782746,8.874452,7.1104393,5.3446136,3.5806012,1.8147756,0.05076295,0.23931105,0.42967212,0.6200332,0.8103943,1.0007553,0.85027945,0.69980353,0.5493277,0.40066472,0.25018883,0.21755551,0.18492219,0.15228885,0.11965553,0.0870222,0.8557183,1.6226015,2.3894846,3.1581807,3.925064,3.633177,3.339477,3.04759,2.7557032,2.4620032,2.2172532,1.9725033,1.7277533,1.4830034,1.2382535,1.3343405,1.4322405,1.5301404,1.6280404,1.7241274,4.0102735,6.294606,8.580752,10.865085,13.149418,13.134913,13.12041,13.1059065,13.08959,13.075087,14.159238,15.245202,16.329353,17.41532,18.49947,17.029158,15.5606575,14.090345,12.620032,11.14972,10.799818,10.449916,10.100015,9.750113,9.400211,9.6141405,9.829884,10.045626,10.259555,10.475298,10.457169,10.440851,10.422722,10.4045925,10.388275,11.202296,12.018129,12.8321495,13.647983,14.462003,15.411995,16.361988,17.31198,18.261972,19.211964,18.845747,18.477715,18.109684,17.741652,17.375433,16.84786,16.32029,15.792717,15.265145,14.737573,14.534521,14.333282,14.13023,13.927178,13.724127,13.53014,13.33434,13.140353,12.944552,12.750566,12.908294,13.064208,13.221936,13.379663,13.537392,12.699803,11.862214,11.024626,10.1870365,9.349448,10.411844,11.47424,12.536636,13.600845,14.663241,15.339477,16.017525,16.695572,17.371807,18.049856,18.269224,18.490406,18.709774,18.929142,19.150324,18.426952,17.705393,16.982021,16.260462,15.537089,16.289469,17.04185,17.794228,18.54842,19.3008,18.503096,17.705393,16.907688,16.109985,15.312282,15.279649,15.247015,15.214382,15.181748,15.149116,18.987158,22.8252,26.66324,30.49947,34.337513,33.92778,33.51805,33.108322,32.69678,32.287052,32.147453,32.007854,31.868256,31.726845,31.587248,32.994106,34.40278,35.809635,37.218307,38.625168,39.41562,40.204258,40.99471,41.78516,42.575615,40.619427,38.665054,36.71068,34.754494,32.800117,31.949839,31.09956,30.24928,29.400814,28.550535,29.516844,30.484966,31.453089,32.419395,33.38752,35.209545,37.031574,38.855415,40.67744,42.49947,37.80571,33.110134,28.414562,23.720802,19.025229,19.518354,20.009668,20.502794,20.994106,21.487232,23.43254,25.37785,27.323158,29.266655,31.211964,25.38329,19.552801,13.722314,7.891826,2.0631514,2.8499773,3.636803,4.4254417,5.2122674,6.000906,5.331923,4.664753,3.9975824,3.3304121,2.663242,3.009518,3.3576066,3.7056956,4.0519714,4.40006,3.5207734,2.6396735,1.7603867,0.8792868,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.045324065,0.03988518,0.034446288,0.030820364,0.025381476,0.06707962,0.11059072,0.15228885,0.19579996,0.2374981,0.28463513,0.33177215,0.38072214,0.42785916,0.4749962,0.48043507,0.48587397,0.4894999,0.4949388,0.50037766,0.41516843,0.32995918,0.24474995,0.15954071,0.07433146,0.07070554,0.065266654,0.059827764,0.054388877,0.05076295,0.48043507,0.9101072,1.3397794,1.7694515,2.1991236,4.022964,5.844991,7.667019,9.490859,11.312886,11.59027,11.867653,12.145037,12.42242,12.699803,11.579392,10.460794,9.340384,8.219973,7.0995617,5.9302006,4.76084,3.589666,2.420305,1.2491312,1.0768998,0.90466833,0.7324369,0.56020546,0.387974,0.46955732,0.5529536,0.6345369,0.7179332,0.7995165,0.95180535,1.1040943,1.258196,1.4104849,1.5627737,1.6352923,1.7078108,1.7803292,1.8528478,1.9253663,1.7005589,1.4757515,1.2491312,1.0243238,0.7995165,0.6399758,0.48043507,0.3208944,0.15954071,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.4169814,0.7850128,1.1530442,1.5192627,1.887294,1.6298534,1.3724127,1.114972,0.8575313,0.6000906,0.48224804,0.36440548,0.24837588,0.13053331,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.42423326,0.73787576,1.0497054,1.3633479,1.6751775,1.3905423,1.1059072,0.8194591,0.53482395,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.09064813,0.13053331,0.17041849,0.21030366,0.25018883,0.52575916,0.7995165,1.0750868,1.3506571,1.6244144,1.3397794,1.0551442,0.7705091,0.48587397,0.19942589,0.6399758,1.0805258,1.5192627,1.9598125,2.4003625,2.0830941,1.7658255,1.4467441,1.1294757,0.8122072,0.90285534,0.9916905,1.0823387,1.1729867,1.261822,1.0098201,0.75781834,0.5058166,0.2520018,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.73424983,1.4703126,2.2045624,2.9406252,3.6748753,6.8221784,9.969481,13.116784,16.2659,19.413204,17.112555,14.811904,12.513068,10.212419,7.911769,6.677141,5.4425135,4.207886,2.9732587,1.7368182,1.7404441,1.742257,1.745883,1.7476959,1.7495089,3.484514,5.219519,6.9545245,8.689529,10.424535,10.087324,9.750113,9.412902,9.07569,8.736667,7.819308,6.9019485,5.9845896,5.06723,4.1498713,3.3195345,2.4891977,1.6606737,0.83033687,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.065266654,0.06707962,0.07070554,0.072518505,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.03988518,0.07977036,0.11965553,0.15954071,0.19942589,0.36077955,0.52032024,0.67986095,0.83940166,1.0007553,0.8520924,0.70524246,0.55839247,0.40972954,0.26287958,0.23205921,0.2030518,0.17223145,0.14322405,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.3245203,0.5493277,0.774135,1.0007553,1.2255627,1.0823387,0.93911463,0.79770356,0.6544795,0.51306844,0.4405499,0.3680314,0.2955129,0.2229944,0.15047589,0.14322405,0.13415924,0.12690738,0.11965553,0.11240368,0.15228885,0.19217403,0.23205921,0.27194437,0.31182957,0.56927025,0.82671094,1.0841516,1.3415923,1.6008459,2.3169663,3.0348995,3.7528327,4.4707656,5.186886,4.274966,3.3630457,2.4493124,1.5373923,0.62547207,0.55839247,0.4894999,0.4224203,0.35534066,0.28826106,0.25925365,0.23205921,0.20486477,0.17767033,0.15047589,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,4.3746786,4.3529234,4.329355,4.307599,4.2858434,4.262275,4.3202896,4.3783045,4.4345064,4.4925213,4.550536,4.2949085,4.0392804,3.785466,3.529838,3.2742105,3.6948178,4.115425,4.5342193,4.954827,5.375434,6.1169357,6.8602505,7.6017523,8.345067,9.088382,8.985043,8.881703,8.780178,8.676839,8.575313,8.8672,9.1609,9.452786,9.744674,10.038374,10.810696,11.583018,12.35534,13.127662,13.899984,13.406858,12.915545,12.42242,11.929294,11.437981,11.048194,10.658407,10.266808,9.87702,9.487233,11.546759,13.608097,15.667623,17.727148,19.786674,26.017826,32.247166,38.478317,44.707657,50.936996,43.777607,36.618217,29.457016,22.297626,15.138238,13.4594345,11.782444,10.1054535,8.42665,6.7496595,5.408067,4.064662,2.72307,1.3796645,0.038072214,0.1794833,0.32270733,0.46411842,0.6073425,0.7505665,0.63816285,0.52575916,0.41335547,0.2991388,0.18673515,0.18492219,0.18310922,0.1794833,0.17767033,0.17585737,0.9354887,1.69512,2.4547513,3.2143826,3.975827,3.8017826,3.6295512,3.4573197,3.2850883,3.1128569,2.9841363,2.857229,2.7303216,2.6016014,2.474694,2.657803,2.8390994,3.0222087,3.2053177,3.386614,5.4443264,7.502039,9.5597515,11.617464,13.675177,14.231756,14.790149,15.346728,15.905121,16.4617,17.107115,17.75253,18.397943,19.04336,19.68696,18.285542,16.882307,15.4790745,14.077655,12.674421,12.186734,11.700861,11.213174,10.725487,10.2378,10.355642,10.471672,10.589515,10.707357,10.825199,11.153346,11.479679,11.807825,12.134158,12.462305,12.792264,13.122223,13.452183,13.782142,14.112101,15.025834,15.937754,16.849674,17.763407,18.675327,18.214834,17.754343,17.295664,16.83517,16.374678,15.894243,15.415621,14.935185,14.454751,13.974316,13.957999,13.939869,13.92174,13.905423,13.887294,13.834718,13.782142,13.729566,13.67699,13.6244135,13.68968,13.754947,13.820213,13.885481,13.9507475,13.113158,12.27557,11.437981,10.600392,9.762803,10.825199,11.887595,12.949992,14.012388,15.074784,15.729263,16.385555,17.040035,17.694515,18.350807,18.278288,18.20577,18.133251,18.060734,17.988214,17.39175,16.797098,16.202446,15.607795,15.013144,16.030214,17.047287,18.06436,19.083244,20.100317,19.066927,18.035353,17.001963,15.970387,14.936998,14.960567,14.982323,15.005891,15.027647,15.049402,19.112251,23.1751,27.23795,31.300798,35.361835,34.567757,33.771866,32.97779,32.1819,31.387821,31.34431,31.302612,31.2591,31.217403,31.175705,32.901646,34.6294,36.35715,38.084904,39.812656,40.49252,41.17238,41.85224,42.5321,43.211964,41.114365,39.01677,36.91917,34.82157,32.72579,31.850126,30.974466,30.100618,29.224957,28.349297,29.210453,30.069798,30.929142,31.790298,32.649643,33.96948,35.289318,36.609154,37.9308,39.25064,35.196857,31.144884,27.092913,23.03913,18.987158,19.259102,19.53286,19.804804,20.076748,20.350506,21.702974,23.055445,24.407915,25.760386,27.112856,22.09095,17.06723,12.045323,7.021604,1.9996977,2.8372865,3.6748753,4.512464,5.3500524,6.187641,5.377247,4.5668526,3.7582715,2.9478772,2.137483,2.5580902,2.9768846,3.397492,3.8180993,4.2368937,3.39024,2.5417736,1.69512,0.8466535,0.0,0.0,0.0,0.0,0.0,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.09064813,0.07977036,0.07070554,0.059827764,0.05076295,0.12328146,0.19579996,0.26831847,0.34083697,0.41335547,0.40791658,0.40247768,0.39703882,0.39159992,0.387974,0.38434806,0.3825351,0.38072214,0.3770962,0.37528324,0.32995918,0.28463513,0.23931105,0.19579996,0.15047589,0.13959812,0.13053331,0.11965553,0.11059072,0.099712946,0.96087015,1.8202144,2.6795588,3.540716,4.40006,5.620184,6.8403077,8.0604315,9.280556,10.500679,10.968424,11.434355,11.9021,12.3698435,12.837588,11.809638,10.781689,9.755551,8.727602,7.699652,6.347182,4.994712,3.6422417,2.2897718,0.93730164,0.81764615,0.6979906,0.57833505,0.45686656,0.33721104,0.58921283,0.8430276,1.0950294,1.3470312,1.6008459,1.6298534,1.6606737,1.6896812,1.7205015,1.7495089,1.8945459,2.039583,2.18462,2.3296568,2.474694,2.2625773,2.0504606,1.8383441,1.6244144,1.4122978,1.1294757,0.8466535,0.5656443,0.28282216,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.33539808,0.6327239,0.9300498,1.2273756,1.5247015,1.3343405,1.1457924,0.9554313,0.7650702,0.5747091,0.46411842,0.35534066,0.24474995,0.13415924,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.36259252,0.62547207,0.8883517,1.1494182,1.4122978,1.1802386,0.9481794,0.71430725,0.48224804,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.06707962,0.09789998,0.12690738,0.15772775,0.18673515,0.40066472,0.61278135,0.824898,1.0370146,1.2491312,1.0424535,0.83577573,0.62728506,0.42060733,0.21211663,0.5293851,0.8466535,1.1657349,1.4830034,1.8002719,1.7404441,1.6806163,1.6207886,1.5591478,1.49932,1.7041848,1.9108626,2.1157274,2.3205922,2.525457,2.0196402,1.5156367,1.0098201,0.5058166,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.4576219,2.9152439,4.3728657,5.8304877,7.28811,9.208037,11.127964,13.047892,14.967819,16.887747,14.699501,12.513068,10.324821,8.136576,5.9501433,5.429823,4.9095025,4.3891826,3.870675,3.350355,3.005892,2.659616,2.3151531,1.9706904,1.6244144,5.2068286,8.789243,12.373469,15.955884,19.538298,17.174194,14.811904,12.449615,10.087324,7.7250338,6.8022356,5.8794374,4.95664,4.0356545,3.1128569,2.4891977,1.8673514,1.2455053,0.62184614,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.06707962,0.072518505,0.07795739,0.08339628,0.0870222,0.07070554,0.052575916,0.034446288,0.018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.054388877,0.11059072,0.16497959,0.21936847,0.2755703,0.43329805,0.58921283,0.7469406,0.90466833,1.062396,0.8919776,0.72337204,0.5529536,0.3825351,0.21211663,0.19036107,0.16679256,0.14503701,0.12328146,0.099712946,0.0870222,0.07433146,0.06164073,0.05076295,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.027194439,0.054388877,0.08339628,0.11059072,0.13778515,0.53663695,0.93730164,1.3379664,1.7368182,2.137483,1.840157,1.5428312,1.2455053,0.9481794,0.6508536,0.56745726,0.48587397,0.40247768,0.3208944,0.2374981,0.21030366,0.18310922,0.15410182,0.12690738,0.099712946,0.15410182,0.21030366,0.26469254,0.3208944,0.37528324,0.86478317,1.3542831,1.845596,2.335096,2.8245957,3.1092308,3.395679,3.680314,3.9649491,4.249584,3.5243993,2.7992141,2.0758421,1.3506571,0.62547207,0.5656443,0.5058166,0.44417584,0.38434806,0.3245203,0.2955129,0.26469254,0.23568514,0.20486477,0.17585737,0.15047589,0.12509441,0.099712946,0.07433146,0.05076295,4.249584,4.2477713,4.2441454,4.2423325,4.2405195,4.2368937,4.2930956,4.347484,4.401873,4.458075,4.512464,4.2930956,4.071914,3.8525455,3.633177,3.4119956,3.7419548,4.071914,4.401873,4.7318325,5.0617914,5.957395,6.8529987,7.746789,8.642392,9.537996,9.514427,9.492672,9.469104,9.447348,9.425592,9.695724,9.965856,10.234174,10.504305,10.774437,11.452485,12.130532,12.806767,13.484816,14.162864,13.580903,12.9971285,12.415168,11.833207,11.249433,10.852394,10.455356,10.058316,9.659465,9.262425,11.715364,14.168303,16.619429,19.072367,21.525305,27.382986,33.24067,39.09835,44.95422,50.8119,44.022358,37.23281,30.441454,23.65191,16.862366,14.4148655,11.967366,9.519867,7.072367,4.6248674,3.7056956,2.7847104,1.8655385,0.9445535,0.025381476,0.11965553,0.21574254,0.3100166,0.40429065,0.50037766,0.42423326,0.34990177,0.2755703,0.19942589,0.12509441,0.15228885,0.1794833,0.20667773,0.23568514,0.26287958,1.015259,1.7676386,2.520018,3.2723975,4.024777,3.972201,3.919625,3.8670492,3.8144734,3.7618973,3.7528327,3.7419548,3.73289,3.7220123,3.7129474,3.9794528,4.2477713,4.514277,4.782595,5.049101,6.880193,8.709473,10.540565,12.3698435,14.199123,15.330412,16.459887,17.589363,18.720652,19.850128,20.054993,20.259857,20.464722,20.669586,20.87445,19.540112,18.20577,16.869617,15.535276,14.199123,13.575464,12.949992,12.32452,11.700861,11.075388,11.095331,11.115273,11.135216,11.155159,11.175101,11.847711,12.52032,13.192928,13.865538,14.538147,14.382232,14.22813,14.072216,13.918114,13.762199,14.63786,15.511708,16.38737,17.26303,18.136877,17.585737,17.032784,16.47983,15.926876,15.375735,14.942437,14.50914,14.077655,13.644357,13.212872,13.379663,13.548269,13.715062,13.881854,14.05046,14.139296,14.229943,14.320591,14.409427,14.500074,14.47288,14.445685,14.416678,14.389484,14.362289,13.524701,12.687112,11.849524,11.011934,10.174346,11.236742,12.299138,13.363347,14.425743,15.488139,16.120863,16.751774,17.384499,18.017221,18.649946,18.285542,17.919323,17.554916,17.190512,16.824293,16.358362,15.890617,15.422873,14.955129,14.487384,15.769149,17.052727,18.33449,19.618069,20.899832,19.632572,18.36531,17.09805,15.83079,14.561715,14.639673,14.71763,14.795588,14.871732,14.94969,19.237347,23.525002,27.812658,32.100315,36.387974,35.207733,34.027496,32.847256,31.667017,30.486778,30.54298,30.59737,30.651758,30.70796,30.762348,32.809185,34.85783,36.904667,38.953316,41.00015,41.56942,42.140503,42.709774,43.280857,43.850124,41.609303,39.370296,37.129475,34.890465,32.649643,31.750414,30.849371,29.950142,29.049099,28.14987,28.90225,29.654629,30.40701,31.159388,31.911768,32.729412,33.54706,34.364704,35.18235,35.999996,32.589817,29.179632,25.76945,22.359268,18.950897,19.001661,19.054237,19.106813,19.15939,19.211964,19.97341,20.73304,21.492672,22.252302,23.011934,18.796797,14.583471,10.36652,6.153195,1.938057,2.8245957,3.7129474,4.599486,5.487838,6.3743763,5.422571,4.4707656,3.5171473,2.565342,1.6117238,2.1048496,2.5979755,3.0892882,3.5824142,4.07554,3.2597067,2.4456866,1.6298534,0.81583315,0.0,0.0,0.0,0.0,0.0,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.13415924,0.11965553,0.10515183,0.09064813,0.07433146,0.17767033,0.27919623,0.3825351,0.48587397,0.5873999,0.5293851,0.47318324,0.41516843,0.35715362,0.2991388,0.29007402,0.27919623,0.27013144,0.25925365,0.25018883,0.24474995,0.23931105,0.23568514,0.23024625,0.22480737,0.21030366,0.19579996,0.1794833,0.16497959,0.15047589,1.4394923,2.7303216,4.019338,5.3101673,6.599184,7.217404,7.835624,8.452031,9.070251,9.686659,10.344765,11.00287,11.6591625,12.317267,12.975373,12.039885,11.104396,10.17072,9.235231,8.299743,6.7641635,5.230397,3.6948178,2.1592383,0.62547207,0.55839247,0.4894999,0.4224203,0.35534066,0.28826106,0.7106813,1.1331016,1.5555218,1.9779422,2.4003625,2.3079014,2.2154403,2.1229792,2.030518,1.938057,2.1556125,2.373168,2.5907235,2.808279,3.0258346,2.8245957,2.6251698,2.4257438,2.2245052,2.0250793,1.6207886,1.214685,0.8103943,0.40429065,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.2520018,0.48043507,0.7070554,0.9354887,1.162109,1.0406405,0.91735905,0.79589057,0.6726091,0.5493277,0.44780177,0.3444629,0.24293698,0.13959812,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.018129626,0.034446288,0.052575916,0.07070554,0.0870222,0.2991388,0.51306844,0.72518504,0.93730164,1.1494182,0.969935,0.7904517,0.6091554,0.42967212,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.045324065,0.065266654,0.08520924,0.10515183,0.12509441,0.2755703,0.42423326,0.5747091,0.72518504,0.87566096,0.7451276,0.61459434,0.48587397,0.35534066,0.22480737,0.42060733,0.61459434,0.8103943,1.0043813,1.2001812,1.3977941,1.5954071,1.79302,1.9906329,2.1882458,2.5073273,2.8282216,3.147303,3.4681973,3.787279,3.0294604,2.2716422,1.5156367,0.75781834,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.180994,4.360175,6.539356,8.72035,10.899531,11.592083,12.284635,12.977186,13.669738,14.362289,12.28826,10.212419,8.136576,6.0625467,3.9867048,4.1825047,4.3783045,4.572292,4.7680917,4.9620786,4.269527,3.576975,2.8844235,2.1918716,1.49932,6.930956,12.358966,17.790602,23.220425,28.650248,24.262878,19.87551,15.488139,11.10077,6.7134004,5.7851634,4.856927,3.930503,3.002266,2.0758421,1.6606737,1.2455053,0.83033687,0.41516843,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.07070554,0.07795739,0.08520924,0.092461094,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.07070554,0.13959812,0.21030366,0.27919623,0.34990177,0.5058166,0.65991837,0.81583315,0.969935,1.1258497,0.9318628,0.73968875,0.5475147,0.35534066,0.16316663,0.14684997,0.13234627,0.11784257,0.10333887,0.0870222,0.07433146,0.06164073,0.05076295,0.038072214,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.034446288,0.07070554,0.10515183,0.13959812,0.17585737,0.7505665,1.3252757,1.8999848,2.474694,3.049403,2.5979755,2.1447346,1.693307,1.2400664,0.7868258,0.69436467,0.60190356,0.5094425,0.4169814,0.3245203,0.27738327,0.23024625,0.18310922,0.13415924,0.0870222,0.15772775,0.22662032,0.29732585,0.3680314,0.43692398,1.1602961,1.8818551,2.6052272,3.3267863,4.0501585,3.9033084,3.7546456,3.6077955,3.4591327,3.3122826,2.7756457,2.2371957,1.7005589,1.162109,0.62547207,0.5728962,0.52032024,0.46774435,0.41516843,0.36259252,0.32995918,0.29732585,0.26469254,0.23205921,0.19942589,0.17585737,0.15047589,0.12509441,0.099712946,0.07433146,4.12449,4.1426196,4.160749,4.177066,4.195195,4.213325,4.265901,4.3166637,4.36924,4.421816,4.4743915,4.2894692,4.1045475,3.919625,3.7347028,3.5497808,3.7890918,4.0302157,4.269527,4.510651,4.749962,5.7978544,6.8457465,7.891826,8.939718,9.987611,10.045626,10.101828,10.1598425,10.217857,10.275872,10.522435,10.770811,11.017374,11.26575,11.512312,12.094274,12.678047,13.260008,13.8419695,14.425743,13.753134,13.080525,12.407916,11.735307,11.062697,10.658407,10.252303,9.848013,9.441909,9.037619,11.882156,14.726695,17.573046,20.417585,23.262123,28.748148,34.23236,39.718384,45.202595,50.68681,44.26711,37.84741,31.427706,25.008005,18.588305,15.3702965,12.152288,8.934279,5.718084,2.5000753,2.0033236,1.504759,1.0080072,0.5094425,0.012690738,0.059827764,0.10696479,0.15410182,0.2030518,0.25018883,0.21211663,0.17585737,0.13778515,0.099712946,0.06164073,0.11965553,0.17767033,0.23568514,0.291887,0.34990177,1.0950294,1.840157,2.5852847,3.3304121,4.07554,4.1426196,4.209699,4.2767787,4.345671,4.4127507,4.519716,4.6266804,4.7354584,4.842423,4.949388,5.3029156,5.65463,6.008158,6.359873,6.7134004,8.314246,9.916905,11.519565,13.122223,14.724882,16.427254,18.129625,19.831997,21.53437,23.236742,23.002869,22.767183,22.533312,22.297626,22.061941,20.794682,19.52742,18.260159,16.992899,15.725637,14.96238,14.200936,13.437678,12.674421,11.912977,11.83502,11.757062,11.679105,11.602961,11.525003,12.542075,13.559147,14.5780325,15.595104,16.612177,15.9722,15.332225,14.692248,14.052273,13.412297,14.249886,15.087475,15.925063,16.762651,17.60024,16.954826,16.309412,15.66581,15.020395,14.37498,13.990632,13.604471,13.220123,12.835775,12.449615,12.803142,13.154857,13.508384,13.860099,14.211814,14.445685,14.677745,14.909804,15.141864,15.375735,15.254267,15.134612,15.014956,14.895301,14.775645,13.938056,13.100468,12.262879,11.42529,10.587702,11.650098,12.712494,13.77489,14.837286,15.899682,16.51065,17.119806,17.730774,18.33993,18.950897,18.292793,17.634687,16.976582,16.32029,15.662184,15.32316,14.982323,14.643299,14.302462,13.961625,15.509895,17.058165,18.604622,20.152891,21.699348,20.198215,18.69527,17.192324,15.689378,14.188245,14.320591,14.452938,14.585284,14.71763,14.849977,19.36244,23.874905,28.387367,32.899834,37.412296,35.84771,34.283123,32.716724,31.152136,29.58755,29.739838,29.892128,30.044416,30.196705,30.350807,32.716724,35.084454,37.452183,39.819912,42.18764,42.648132,43.10681,43.567303,44.027798,44.48829,42.104244,39.72201,37.33978,34.957546,32.575314,31.650702,30.724277,29.799665,28.875055,27.950443,28.59586,29.23946,29.884874,30.53029,31.175705,31.489347,31.804802,32.12026,32.435715,32.749355,29.982775,27.214382,24.4478,21.679407,18.912827,18.74422,18.577427,18.410635,18.24203,18.075237,18.24203,18.410635,18.577427,18.74422,18.912827,15.504456,12.097899,8.689529,5.282973,1.8746033,2.811905,3.7492065,4.688321,5.6256227,6.5629244,5.467895,4.3728657,3.2778363,2.182807,1.0877775,1.651609,2.2172532,2.7828975,3.346729,3.9123733,3.1291735,2.3477864,1.5645868,0.78319985,0.0,0.0,0.0,0.0,0.0,0.0,0.03988518,0.07977036,0.11965553,0.15954071,0.19942589,0.1794833,0.15954071,0.13959812,0.11965553,0.099712946,0.23205921,0.36440548,0.49675176,0.629098,0.76325727,0.6526665,0.5420758,0.43329805,0.32270733,0.21211663,0.19579996,0.17767033,0.15954071,0.14322405,0.12509441,0.15954071,0.19579996,0.23024625,0.26469254,0.2991388,0.27919623,0.25925365,0.23931105,0.21936847,0.19942589,1.9199274,3.6404288,5.3609304,7.079619,8.80012,8.814624,8.829127,8.845445,8.859948,8.874452,9.7229185,10.5695715,11.418038,12.264692,13.113158,12.270131,11.427103,10.584076,9.742861,8.899834,7.1829576,5.464269,3.7473936,2.030518,0.31182957,0.29732585,0.28282216,0.26831847,0.2520018,0.2374981,0.83033687,1.4231756,2.0142014,2.6070402,3.199879,2.9841363,2.770207,2.5544643,2.3405347,2.124792,2.4148662,2.70494,2.9950142,3.2850883,3.5751622,3.386614,3.199879,3.0131438,2.8245957,2.6378605,2.1102884,1.5827163,1.0551442,0.5275721,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.17041849,0.32814622,0.48587397,0.6417888,0.7995165,0.7451276,0.69073874,0.6345369,0.58014804,0.52575916,0.42967212,0.33539808,0.23931105,0.14503701,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.2374981,0.40066472,0.5620184,0.72518504,0.8883517,0.75963134,0.6327239,0.5058166,0.3770962,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.02175555,0.032633327,0.04169814,0.052575916,0.06164073,0.15047589,0.2374981,0.3245203,0.41335547,0.50037766,0.44780177,0.39522585,0.34264994,0.29007402,0.2374981,0.3100166,0.3825351,0.4550536,0.5275721,0.6000906,1.0551442,1.5101979,1.9652514,2.420305,2.8753586,3.3104696,3.7455807,4.1806917,4.615803,5.050914,4.0392804,3.0294604,2.0196402,1.0098201,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.902553,5.805106,8.70766,11.610212,14.512766,13.9779415,13.443117,12.908294,12.371656,11.836833,9.875207,7.911769,5.9501433,3.9867048,2.0250793,2.9351864,3.8452935,4.7554007,5.6655083,6.5756154,5.5349746,4.494334,3.4555066,2.4148662,1.3742256,8.653271,15.930502,23.207733,30.484966,37.7622,31.349749,24.9373,18.52485,12.112403,5.6999545,4.7680917,3.834416,2.902553,1.9706904,1.0370146,0.83033687,0.62184614,0.41516843,0.20667773,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.072518505,0.08339628,0.092461094,0.10333887,0.11240368,0.09064813,0.06707962,0.045324065,0.02175555,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.08520924,0.17041849,0.25562772,0.34083697,0.42423326,0.57833505,0.7306239,0.88291276,1.0352017,1.1874905,0.97174793,0.75781834,0.5420758,0.32814622,0.11240368,0.10515183,0.09789998,0.09064813,0.08339628,0.07433146,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.04169814,0.08520924,0.12690738,0.17041849,0.21211663,0.96268314,1.7132497,2.4620032,3.2125697,3.9631362,3.3557937,2.7466383,2.1392958,1.5319533,0.9246109,0.823085,0.7197462,0.61822027,0.5148814,0.41335547,0.3444629,0.27738327,0.21030366,0.14322405,0.07433146,0.15954071,0.24474995,0.32995918,0.41516843,0.50037766,1.455809,2.4094272,3.3648586,4.3202896,5.275721,4.695573,4.115425,3.5352771,2.955129,2.374981,2.0250793,1.6751775,1.3252757,0.97537386,0.62547207,0.58014804,0.53482395,0.4894999,0.44417584,0.40066472,0.36440548,0.32995918,0.2955129,0.25925365,0.22480737,0.19942589,0.17585737,0.15047589,0.12509441,0.099712946,3.9993954,4.0374675,4.07554,4.1117992,4.1498713,4.1879435,4.2368937,4.2876563,4.3366065,4.3873696,4.4381323,4.2876563,4.137181,3.9867048,3.8380418,3.6875658,3.8380418,3.9867048,4.137181,4.2876563,4.4381323,5.638314,6.836682,8.036863,9.237044,10.437225,10.57501,10.712796,10.850581,10.988366,11.124338,11.349146,11.575767,11.800573,12.025381,12.250188,12.737875,13.225562,13.713249,14.199123,14.68681,13.925365,13.162108,12.400664,11.637406,10.874149,10.462607,10.049252,9.637709,9.224354,8.812811,12.050762,15.2869005,18.52485,21.762802,25.000753,30.113308,35.22405,40.338417,45.450974,50.561714,44.511856,38.462,32.412144,26.36229,20.312433,16.325727,12.337211,8.350506,4.361988,0.37528324,0.2991388,0.22480737,0.15047589,0.07433146,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0870222,0.17585737,0.26287958,0.34990177,0.43692398,1.1747998,1.9126755,2.6505513,3.386614,4.12449,4.313038,4.499773,4.688321,4.8750563,5.0617914,5.2865987,5.5132194,5.7380266,5.962834,6.187641,6.624565,7.063302,7.500226,7.93715,8.375887,9.750113,11.124338,12.500377,13.874602,15.250641,17.524096,19.799364,22.074633,24.349901,26.625168,25.950747,25.274511,24.60009,23.925667,23.249432,22.049252,20.850883,19.650702,18.45052,17.25034,16.349297,15.4500675,14.5508375,13.649796,12.750566,12.574709,12.400664,12.224807,12.050762,11.874905,13.238253,14.599788,15.963136,17.32467,18.688019,17.562168,16.438131,15.312282,14.188245,13.062395,13.861912,14.663241,15.462758,16.262274,17.06179,16.325727,15.5878525,14.849977,14.112101,13.374225,13.037014,12.699803,12.362592,12.025381,11.6881695,12.224807,12.763257,13.299893,13.838344,14.37498,14.750263,15.125546,15.50083,15.8743,16.249584,16.037468,15.825351,15.613234,15.399304,15.187187,14.349599,13.512011,12.674421,11.836833,10.999244,12.06164,13.125849,14.188245,15.250641,16.313038,16.900436,17.487837,18.075237,18.662638,19.250036,18.300045,17.350052,16.400059,15.4500675,14.500074,14.287958,14.075842,13.861912,13.649796,13.437678,15.250641,17.06179,18.874754,20.687716,22.500679,20.762047,19.025229,17.286598,15.54978,13.812962,13.999697,14.188245,14.37498,14.561715,14.750263,19.487535,24.224806,28.962078,33.69935,38.43662,36.487686,34.536938,32.588,30.637255,28.68832,28.936695,29.186884,29.437073,29.687262,29.93745,32.62426,35.312885,37.999695,40.68832,43.37513,43.725033,44.074932,44.424835,44.77474,45.124638,42.599182,40.07554,37.55008,35.024624,32.49917,31.549175,30.599182,29.64919,28.699198,27.749205,28.287655,28.824291,29.362741,29.89938,30.437828,30.24928,30.062546,29.87581,29.687262,29.500526,27.375734,25.250942,23.124338,20.999546,18.874754,18.48678,18.100618,17.712645,17.32467,16.936697,16.512463,16.08823,15.662184,15.23795,14.811904,12.212116,9.612328,7.0125394,4.4127507,1.8129625,2.7992141,3.787279,4.7753434,5.763408,6.7496595,5.5132194,4.274966,3.0367124,1.8002719,0.5620184,1.2001812,1.8383441,2.474694,3.1128569,3.7492065,3.000453,2.2498865,1.49932,0.7505665,0.0,0.0,0.0,0.0,0.0,0.0,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,0.22480737,0.19942589,0.17585737,0.15047589,0.12509441,0.28826106,0.44961473,0.61278135,0.774135,0.93730164,0.774135,0.61278135,0.44961473,0.28826106,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.07433146,0.15047589,0.22480737,0.2991388,0.37528324,0.34990177,0.3245203,0.2991388,0.2755703,0.25018883,2.4003625,4.550536,6.70071,8.8508835,10.999244,10.411844,9.824444,9.237044,8.649645,8.062244,9.099259,10.138086,11.175101,12.212116,13.24913,12.500377,11.74981,10.999244,10.25049,9.499924,7.5999393,5.6999545,3.7999697,1.8999848,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.9499924,1.7132497,2.474694,3.2379513,3.9993954,3.6621845,3.3249733,2.9877625,2.6505513,2.3133402,2.6741197,3.0367124,3.3993049,3.7618973,4.12449,3.9504454,3.774588,3.6005437,3.4246864,3.2506418,2.5997884,1.9507477,1.2998942,0.6508536,0.0,0.0,0.0,0.0,0.0,0.0,0.0870222,0.17585737,0.26287958,0.34990177,0.43692398,0.44961473,0.46230546,0.4749962,0.48768693,0.50037766,0.41335547,0.3245203,0.2374981,0.15047589,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.17585737,0.28826106,0.40066472,0.51306844,0.62547207,0.5493277,0.4749962,0.40066472,0.3245203,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.15047589,0.17585737,0.19942589,0.22480737,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.7124943,1.4249886,2.137483,2.8499773,3.5624714,4.1117992,4.6629395,5.2122674,5.763408,6.3127356,5.049101,3.787279,2.525457,1.261822,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,3.625925,7.250037,10.875962,14.500074,18.124187,16.361988,14.599788,12.837588,11.075388,9.313189,7.462154,5.612932,3.7618973,1.9126755,0.06164073,1.6878681,3.3122826,4.936697,6.5629244,8.187339,6.8004227,5.411693,4.024777,2.6378605,1.2491312,10.375585,19.500225,28.624866,37.749508,46.87415,38.43662,30.000904,21.561563,13.124036,4.688321,3.7492065,2.811905,1.8746033,0.93730164,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.099712946,0.19942589,0.2991388,0.40066472,0.50037766,0.6508536,0.7995165,0.9499924,1.1004683,1.2491312,1.0116332,0.774135,0.53663695,0.2991388,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,1.1747998,2.0994108,3.0258346,3.9504454,4.8750563,4.1117992,3.350355,2.5870976,1.8256533,1.062396,0.9499924,0.8375887,0.72518504,0.61278135,0.50037766,0.41335547,0.3245203,0.2374981,0.15047589,0.06164073,0.16316663,0.26287958,0.36259252,0.46230546,0.5620184,1.7495089,2.9369993,4.12449,5.3119802,6.4994707,5.487838,4.4743915,3.4627585,2.4493124,1.4376793,1.2745126,1.1131591,0.9499924,0.7868258,0.62547207,0.5873999,0.5493277,0.51306844,0.4749962,0.43692398,0.40066472,0.36259252,0.3245203,0.28826106,0.25018883,0.22480737,0.19942589,0.17585737,0.15047589,0.12509441,3.9123733,4.028403,4.1426196,4.256836,4.3728657,4.4870825,4.49796,4.507025,4.517903,4.5269675,4.537845,4.3982472,4.256836,4.117238,3.97764,3.8380418,4.0501585,4.262275,4.4743915,4.688321,4.900438,6.009971,7.119504,8.23085,9.340384,10.449916,10.636651,10.825199,11.011934,11.200482,11.3872175,11.599335,11.813264,12.025381,12.237497,12.449615,12.919171,13.390542,13.860099,14.329657,14.799213,14.066776,13.33434,12.601903,11.869466,11.137029,10.750868,10.362894,9.97492,9.5869465,9.200785,13.528327,17.854055,22.18341,26.510952,30.836681,34.045624,37.252754,40.459885,43.667015,46.87415,41.09805,35.320137,29.542225,23.764313,17.988214,14.492823,10.997431,7.502039,4.006647,0.51306844,0.40972954,0.30820364,0.20486477,0.10333887,0.0,0.10696479,0.21574254,0.32270733,0.42967212,0.53663695,0.533011,0.5275721,0.52213323,0.5166943,0.51306844,0.55839247,0.60190356,0.64722764,0.69255173,0.73787576,1.4594349,2.182807,2.904366,3.6277382,4.349297,4.3420453,4.3347936,4.327542,4.3202896,4.313038,4.7699046,5.2267714,5.6854506,6.1423173,6.599184,7.262728,7.9244595,8.588004,9.249735,9.91328,10.937603,11.961927,12.988064,14.012388,15.036712,16.965704,18.892883,20.820063,22.747242,24.674421,24.019941,23.365461,22.70917,22.05469,21.40021,20.343254,19.284483,18.227526,17.170568,16.1118,15.4500675,14.788336,14.124791,13.46306,12.799516,12.601903,12.40429,12.206677,12.010877,11.813264,12.935488,14.057712,15.179935,16.30216,17.424383,16.592234,15.760084,14.927934,14.095784,13.261822,13.914488,14.567154,15.219821,15.872487,16.525154,15.781839,15.040338,14.297023,13.555521,12.812206,12.513068,12.212116,11.912977,11.612025,11.312886,11.873092,12.433297,12.99169,13.551895,14.112101,14.400362,14.68681,14.975071,15.263332,15.54978,15.272397,14.995013,14.71763,14.440247,14.162864,13.555521,12.948178,12.340837,11.731681,11.124338,12.32452,13.524701,14.724882,15.925063,17.125244,17.560356,17.995466,18.430578,18.865688,19.3008,18.24203,17.185072,16.128115,15.0693445,14.012388,14.139296,14.268016,14.394923,14.521831,14.650551,16.336605,18.024473,19.712341,21.40021,23.088078,21.57063,20.053179,18.53573,17.01828,15.50083,15.95951,16.420002,16.880495,17.339174,17.799667,21.643147,25.484816,29.328295,33.169964,37.01163,35.18054,33.347633,31.514729,29.681824,27.85073,28.24233,28.635744,29.027344,29.420757,29.812357,32.15833,34.50249,36.848465,39.192627,41.536785,42.02447,42.51216,42.999847,43.487534,43.97522,41.84499,39.71476,37.584526,35.454296,33.32588,31.951653,30.57924,29.206827,27.834415,26.462002,26.795588,27.12736,27.459131,27.792717,28.124489,27.952257,27.780025,27.607794,27.435562,27.26333,24.995316,22.727299,20.459282,18.193079,15.925063,15.852545,15.780026,15.707508,15.63499,15.56247,15.201692,14.842725,14.481945,14.122978,13.762199,11.325577,8.887142,6.450521,4.0120864,1.5754645,2.7974012,4.019338,5.243088,6.4650245,7.686961,6.240217,4.7916603,3.3449159,1.8981718,0.44961473,0.96268314,1.4757515,1.987007,2.5000753,3.0131438,2.4547513,1.8981718,1.3397794,0.78319985,0.22480737,0.32814622,0.42967212,0.533011,0.6345369,0.73787576,0.8774739,1.017072,1.1566701,1.2980812,1.4376793,1.2074331,0.97718686,0.7469406,0.5166943,0.28826106,0.40791658,0.5275721,0.64722764,0.7668832,0.8883517,0.89922947,0.9119202,0.9246109,0.93730164,0.9499924,0.75963134,0.56927025,0.38072214,0.19036107,0.0,0.39703882,0.79589057,1.1929294,1.5899682,1.987007,1.7857682,1.5827163,1.3796645,1.1766127,0.97537386,2.7847104,4.594047,6.4051967,8.214534,10.025683,9.644961,9.264238,8.885329,8.504607,8.125698,9.131892,10.139899,11.147907,12.155914,13.162108,12.329959,11.497808,10.665659,9.8316965,8.999546,7.5382986,6.0752378,4.612177,3.149116,1.6878681,1.6733645,1.6570477,1.6425442,1.6280404,1.6117238,2.0105755,2.4076142,2.8046532,3.2016919,3.6005437,3.2850883,2.9696326,2.6541772,2.3405347,2.0250793,2.3097143,2.5943494,2.8807976,3.1654327,3.4500678,3.3757362,3.299592,3.2252605,3.149116,3.0747845,2.6016014,2.1302311,1.6570477,1.1856775,0.7124943,0.61459434,0.5166943,0.42060733,0.32270733,0.22480737,0.25562772,0.28463513,0.3154555,0.3444629,0.37528324,0.387974,0.40066472,0.41335547,0.42423326,0.43692398,0.36440548,0.291887,0.21936847,0.14684997,0.07433146,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.01994259,0.027194439,0.034446288,0.04169814,0.05076295,0.14322405,0.23568514,0.32814622,0.42060733,0.51306844,0.45686656,0.40247768,0.3480888,0.291887,0.2374981,0.19036107,0.14322405,0.09427405,0.047137026,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.11965553,0.13959812,0.15954071,0.1794833,0.19942589,0.16316663,0.12509441,0.0870222,0.05076295,0.012690738,0.6000906,1.1874905,1.7748904,2.3622901,2.94969,3.491766,4.0356545,4.5777307,5.1198063,5.661882,4.550536,3.437377,2.324218,1.2128719,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,3.1309865,6.26016,9.389333,12.52032,15.649493,14.190058,12.730623,11.269376,9.80994,8.350506,6.7496595,5.1506267,3.5497808,1.9507477,0.34990177,1.6624867,2.9750717,4.2876563,5.600241,6.9128265,5.7416525,4.572292,3.4029307,2.231757,1.062396,8.428463,15.792717,23.156971,30.523039,37.88729,31.587248,25.287203,18.987158,12.687112,6.3870673,5.1107416,3.832603,2.5544643,1.2781386,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.059827764,0.07070554,0.07977036,0.09064813,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.06164073,0.099712946,0.13778515,0.17585737,0.21211663,0.17585737,0.13778515,0.099712946,0.06164073,0.025381476,0.27919623,0.53482395,0.7904517,1.0442665,1.2998942,1.2545701,1.209246,1.1657349,1.1204109,1.0750868,0.87022203,0.6653573,0.4604925,0.25562772,0.05076295,0.052575916,0.054388877,0.058014803,0.059827764,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.059827764,0.11965553,0.1794833,0.23931105,0.2991388,1.2672608,2.2353828,3.2016919,4.169814,5.137936,4.3347936,3.531651,2.7303216,1.9271792,1.1258497,0.9898776,0.8557183,0.7197462,0.5855869,0.44961473,0.5493277,0.6508536,0.7505665,0.85027945,0.9499924,0.98443866,1.020698,1.0551442,1.0895905,1.1258497,1.9851941,2.8445382,3.7056956,4.5650396,5.424384,4.603112,3.780027,2.956942,2.13567,1.3125849,1.167548,1.0225109,0.8774739,0.7324369,0.5873999,0.5475147,0.5076295,0.46774435,0.42785916,0.387974,0.36077955,0.33177215,0.3045777,0.27738327,0.25018883,0.23024625,0.21030366,0.19036107,0.17041849,0.15047589,3.825351,4.017525,4.209699,4.401873,4.59586,4.788034,4.7572136,4.7282066,4.6973863,4.668379,4.6375585,4.507025,4.3783045,4.2477713,4.117238,3.9867048,4.262275,4.537845,4.8134155,5.087173,5.3627434,6.3816285,7.402326,8.423024,9.441909,10.462607,10.700105,10.937603,11.175101,11.4126,11.650098,11.849524,12.050762,12.250188,12.449615,12.650853,13.102281,13.555521,14.006948,14.46019,14.911617,14.210001,13.508384,12.804955,12.103338,11.399909,11.037316,10.674724,10.312131,9.949538,9.5869465,15.004078,20.423023,25.840157,31.257288,36.67442,37.97794,39.279648,40.583168,41.884876,43.18658,37.682426,32.178272,26.672306,21.168152,15.662184,12.659918,9.657652,6.6553855,3.6531196,0.6508536,0.52032024,0.38978696,0.25925365,0.13053331,0.0,0.21574254,0.42967212,0.64541465,0.85934424,1.0750868,1.064209,1.0551442,1.0442665,1.0352017,1.0243238,1.0279498,1.0297627,1.0333886,1.0352017,1.0370146,1.745883,2.4529383,3.159994,3.8670492,4.574105,4.3728657,4.169814,3.966762,3.7655232,3.5624714,4.25321,4.942136,5.632875,6.3218007,7.0125394,7.900891,8.78743,9.675781,10.56232,11.450671,12.125093,12.799516,13.475751,14.150173,14.824595,16.405499,17.984589,19.565493,21.144583,22.725487,22.089136,21.4546,20.820063,20.185526,19.549175,18.635443,17.719896,16.80435,15.890617,14.975071,14.5508375,14.124791,13.700559,13.274512,12.850279,12.63091,12.409729,12.19036,11.969179,11.74981,12.632723,13.515636,14.396736,15.279649,16.162561,15.622298,15.082036,14.541773,14.003323,13.46306,13.967064,14.47288,14.976884,15.4827,15.986704,15.239763,14.492823,13.744069,12.9971285,12.250188,11.9873085,11.724429,11.463363,11.200482,10.937603,11.519565,12.103338,12.685299,13.267261,13.849221,14.05046,14.249886,14.449312,14.650551,14.849977,14.507326,14.164677,13.822026,13.479377,13.136727,12.75963,12.382534,12.005438,11.628342,11.249433,12.5873995,13.925365,15.263332,16.599485,17.937452,18.220274,18.503096,18.78592,19.066927,19.34975,18.185827,17.020092,15.854358,14.690435,13.524701,13.992445,14.46019,14.927934,15.3956785,15.861609,17.424383,18.987158,20.54993,22.112705,23.675478,22.377398,21.079315,19.783049,18.484966,17.186886,17.919323,18.651758,19.384195,20.116632,20.850883,23.796947,26.744823,29.692701,32.64058,35.586643,33.873394,32.15833,30.443268,28.728205,27.013142,27.547966,28.08279,28.617615,29.15244,29.687262,31.690586,33.692097,35.69542,37.69693,39.700256,40.325726,40.949387,41.57486,42.20033,42.8258,41.090797,39.355793,37.620785,35.88578,34.150776,32.35413,30.559298,28.764463,26.969631,25.174799,25.301706,25.430426,25.557333,25.68424,25.812962,25.655233,25.497505,25.339779,25.18205,25.024323,22.614895,20.205467,17.794228,15.384801,12.975373,13.21831,13.4594345,13.702372,13.945308,14.188245,13.892733,13.597219,13.301706,13.008006,12.712494,10.437225,8.161958,5.8866897,3.6132345,1.3379664,2.7955883,4.25321,5.710832,7.166641,8.624263,6.967215,5.3101673,3.6531196,1.9942589,0.33721104,0.72518504,1.1131591,1.49932,1.887294,2.275268,1.9108626,1.5446441,1.1802386,0.81583315,0.44961473,0.6544795,0.85934424,1.064209,1.2708868,1.4757515,1.7041848,1.9344311,2.1646774,2.3949237,2.6251698,2.1900587,1.7549478,1.3198367,0.88472575,0.44961473,0.5275721,0.6055295,0.68167394,0.75963134,0.8375887,1.0243238,1.2128719,1.3996071,1.5881553,1.7748904,1.4195497,1.064209,0.7106813,0.35534066,0.0,0.7197462,1.4394923,2.1592383,2.8807976,3.6005437,3.2198215,2.8409123,2.4601903,2.079468,1.7005589,3.1708715,4.6393714,6.109684,7.5799966,9.050309,8.8780775,8.705847,8.531802,8.3595705,8.187339,9.164526,10.141713,11.120712,12.097899,13.075087,12.15954,11.245807,10.330261,9.414715,8.499168,7.474845,6.450521,5.424384,4.40006,3.3757362,3.3068438,3.2397642,3.1726844,3.105605,3.0367124,3.0693457,3.101979,3.1346123,3.1672456,3.199879,2.907992,2.6142921,2.322405,2.030518,1.7368182,1.9453088,2.1519866,2.3604772,2.5671551,2.7756457,2.7992141,2.8245957,2.8499773,2.8753586,2.9007401,2.6052272,2.3097143,2.0142014,1.7205015,1.4249886,1.2291887,1.0352017,0.83940166,0.64541465,0.44961473,0.4224203,0.39522585,0.3680314,0.34083697,0.31182957,0.3245203,0.33721104,0.34990177,0.36259252,0.37528324,0.31726846,0.25925365,0.2030518,0.14503701,0.0870222,0.07433146,0.06164073,0.05076295,0.038072214,0.025381476,0.027194439,0.030820364,0.032633327,0.034446288,0.038072214,0.11059072,0.18310922,0.25562772,0.32814622,0.40066472,0.36440548,0.32995918,0.2955129,0.25925365,0.22480737,0.1794833,0.13415924,0.09064813,0.045324065,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.09064813,0.10515183,0.11965553,0.13415924,0.15047589,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.48768693,0.9499924,1.4122978,1.8746033,2.3369088,2.8717327,3.4083695,3.9431937,4.478018,5.0128417,4.0501585,3.0874753,2.124792,1.162109,0.19942589,0.15954071,0.11965553,0.07977036,0.03988518,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.6360476,5.2702823,7.9045167,10.540565,13.174799,12.018129,10.859646,9.702975,8.544493,7.3878226,6.037165,4.688321,3.3376641,1.987007,0.63816285,1.6371052,2.6378605,3.636803,4.6375585,5.638314,4.6846952,3.73289,2.7792716,1.8274662,0.87566096,6.4795284,12.085209,17.69089,23.294756,28.900436,24.737875,20.575312,16.41275,12.250188,8.087626,6.4704633,4.853301,3.2343252,1.6171626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.045324065,0.052575916,0.059827764,0.06707962,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.11240368,0.17585737,0.2374981,0.2991388,0.36259252,0.2991388,0.2374981,0.17585737,0.11240368,0.05076295,0.4604925,0.87022203,1.2799516,1.6896812,2.0994108,1.8600996,1.6207886,1.3796645,1.1403534,0.89922947,0.726998,0.55476654,0.3825351,0.21030366,0.038072214,0.04169814,0.047137026,0.052575916,0.058014803,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07070554,0.13959812,0.21030366,0.27919623,0.34990177,1.3597219,2.3695421,3.3793623,4.3891826,5.4008155,4.557788,3.7147603,2.8717327,2.030518,1.1874905,1.0297627,0.872035,0.71430725,0.55839247,0.40066472,0.6871128,0.97537386,1.261822,1.550083,1.8383441,1.8075237,1.7767034,1.7476959,1.7168756,1.6878681,2.220879,2.752077,3.2850883,3.8180993,4.349297,3.7165732,3.0856624,2.4529383,1.8202144,1.1874905,1.0605831,0.9318628,0.80495536,0.678048,0.5493277,0.5076295,0.46411842,0.4224203,0.38072214,0.33721104,0.3208944,0.30276474,0.28463513,0.26831847,0.25018883,0.23568514,0.21936847,0.20486477,0.19036107,0.17585737,3.738329,4.006647,4.2767787,4.5469103,4.8170414,5.087173,5.0182805,4.947575,4.876869,4.8079767,4.7372713,4.6176157,4.49796,4.3783045,4.256836,4.137181,4.4743915,4.8116026,5.1506267,5.487838,5.825049,6.755099,7.6851482,8.615198,9.545248,10.475298,10.761745,11.050007,11.338268,11.624716,11.912977,12.099712,12.28826,12.474996,12.661731,12.850279,13.28539,13.720501,14.155612,14.590723,15.025834,14.353225,13.680615,13.008006,12.335398,11.662788,11.325577,10.988366,10.649343,10.312131,9.97492,16.481644,22.99018,29.4969,36.005436,42.51216,41.910255,41.308353,40.704636,40.102734,39.500828,34.266808,29.034595,23.802385,18.570175,13.337966,10.827013,8.317872,5.806919,3.2977788,0.7868258,0.629098,0.47318324,0.3154555,0.15772775,0.0,0.32270733,0.64541465,0.968122,1.2908293,1.6117238,1.5972201,1.5827163,1.5682126,1.551896,1.5373923,1.4975071,1.4576219,1.4177368,1.3778516,1.3379664,2.030518,2.72307,3.4156215,4.1081734,4.800725,4.401873,4.004834,3.6077955,3.2107568,2.811905,3.7347028,4.6575007,5.580299,6.5030966,7.4258947,8.537241,9.6504,10.761745,11.874905,12.988064,13.312584,13.637105,13.961625,14.287958,14.612478,15.845293,17.078108,18.310923,19.541924,20.774738,20.160145,19.54555,18.929142,18.314548,17.699953,16.927631,16.15531,15.382988,14.610665,13.838344,13.649796,13.46306,13.274512,13.087777,12.899229,12.658105,12.415168,12.172231,11.929294,11.6881695,12.329959,12.971747,13.615349,14.257137,14.90074,14.652364,14.405801,14.157425,13.910862,13.662486,14.01964,14.376793,14.73576,15.092914,15.4500675,14.697688,13.945308,13.192928,12.440549,11.6881695,11.463363,11.236742,11.011934,10.7871275,10.56232,11.16785,11.773379,12.377095,12.982625,13.588155,13.700559,13.812962,13.925365,14.037769,14.150173,13.742256,13.33434,12.928236,12.52032,12.112403,11.965553,11.81689,11.67004,11.5231905,11.374527,12.850279,14.324218,15.799969,17.27572,18.749659,18.880192,19.010725,19.139446,19.26998,19.400513,18.127813,16.855114,15.582414,14.309713,13.037014,13.845595,14.652364,15.459132,16.267714,17.074482,18.512161,19.94984,21.38752,22.8252,24.262878,23.184166,22.107265,21.030367,19.951653,18.874754,19.879135,20.885328,21.88971,22.89409,23.900286,25.952559,28.004833,30.057106,32.10938,34.161655,32.564434,30.967215,29.369993,27.772774,26.175554,26.85179,27.529837,28.207886,28.884119,29.562168,31.222841,32.881702,34.542377,36.20305,37.86191,38.625168,39.386612,40.149868,40.913128,41.674572,40.334793,38.99501,37.65523,36.315453,34.975674,32.75842,30.539354,28.322102,26.104849,23.887594,23.809637,23.73168,23.655537,23.577578,23.49962,23.35821,23.214987,23.071762,22.930351,22.787127,20.234476,17.681824,15.129172,12.578335,10.025683,10.582263,11.1406555,11.697234,12.255627,12.812206,12.581961,12.351714,12.123281,11.893035,11.662788,9.550687,7.4367723,5.3246713,3.2125697,1.1004683,2.7919624,4.4852695,6.1767635,7.8700705,9.563377,7.6942134,5.826862,3.9595103,2.0921588,0.22480737,0.48768693,0.7505665,1.0116332,1.2745126,1.5373923,1.3651608,1.1929294,1.020698,0.8466535,0.6744221,0.9826257,1.2908293,1.5972201,1.9054236,2.2118144,2.5327086,2.8517902,3.1726844,3.491766,3.8126602,3.1726844,2.5327086,1.892733,1.2527572,0.61278135,0.64722764,0.68167394,0.7179332,0.7523795,0.7868258,1.1494182,1.5120108,1.8746033,2.2371957,2.5997884,2.079468,1.5591478,1.0406405,0.52032024,0.0,1.0424535,2.084907,3.1273603,4.169814,5.2122674,4.655688,4.0972953,3.540716,2.9823234,2.4257438,3.5552197,4.6846952,5.814171,6.94546,8.074935,8.109382,8.145641,8.180087,8.214534,8.2507925,9.197159,10.145339,11.091705,12.039885,12.988064,11.989121,10.991992,9.994863,8.997733,8.000604,7.413204,6.825804,6.2365913,5.6491914,5.0617914,4.942136,4.8224807,4.702825,4.5831695,4.461701,4.1299286,3.7981565,3.4645715,3.1327994,2.7992141,2.5290828,2.2607644,1.9906329,1.7205015,1.4503701,1.5809034,1.7096237,1.840157,1.9706904,2.0994108,2.2245052,2.3495996,2.474694,2.5997884,2.7248828,2.6070402,2.4891977,2.373168,2.2553256,2.137483,1.845596,1.551896,1.260009,0.968122,0.6744221,0.58921283,0.5058166,0.42060733,0.33539808,0.25018883,0.26287958,0.2755703,0.28826106,0.2991388,0.31182957,0.27013144,0.22662032,0.18492219,0.14322405,0.099712946,0.0870222,0.07433146,0.06164073,0.05076295,0.038072214,0.034446288,0.032633327,0.030820364,0.027194439,0.025381476,0.07795739,0.13053331,0.18310922,0.23568514,0.28826106,0.27194437,0.2574407,0.24293698,0.22662032,0.21211663,0.17041849,0.12690738,0.08520924,0.04169814,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.059827764,0.07070554,0.07977036,0.09064813,0.099712946,0.0870222,0.07433146,0.06164073,0.05076295,0.038072214,0.37528324,0.7124943,1.0497054,1.3869164,1.7241274,2.2516994,2.7792716,3.3068438,3.834416,4.361988,3.5497808,2.7375734,1.9253663,1.1131591,0.2991388,0.23931105,0.1794833,0.11965553,0.059827764,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.1392958,4.2804046,6.4197006,8.560809,10.700105,9.844387,8.990481,8.134763,7.2808576,6.4251394,5.3246713,4.2242026,3.1255474,2.0250793,0.9246109,1.6117238,2.3006494,2.9877625,3.6748753,4.361988,3.6277382,2.8916752,2.1574254,1.4231756,0.6871128,4.5324063,8.3777,12.222994,16.068287,19.911768,17.886688,15.863422,13.838344,11.813264,9.788185,7.8301854,5.8721857,3.9141862,1.9579996,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.030820364,0.034446288,0.03988518,0.045324065,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.16316663,0.25018883,0.33721104,0.42423326,0.51306844,0.42423326,0.33721104,0.25018883,0.16316663,0.07433146,0.6399758,1.2056202,1.7694515,2.335096,2.9007401,2.465629,2.030518,1.5954071,1.1602961,0.72518504,0.5855869,0.44417584,0.3045777,0.16497959,0.025381476,0.032633327,0.03988518,0.047137026,0.054388877,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07977036,0.15954071,0.23931105,0.3208944,0.40066472,1.452183,2.5055144,3.5570326,4.610364,5.661882,4.780782,3.8978696,3.0149567,2.132044,1.2491312,1.0696479,0.8901646,0.7106813,0.5293851,0.34990177,0.824898,1.2998942,1.7748904,2.2498865,2.7248828,2.6306088,2.5345216,2.4402475,2.3441606,2.2498865,2.4547513,2.659616,2.864481,3.0693457,3.2742105,2.8318477,2.3894846,1.9471219,1.504759,1.062396,0.95180535,0.8430276,0.7324369,0.62184614,0.51306844,0.46774435,0.4224203,0.3770962,0.33177215,0.28826106,0.27919623,0.27194437,0.26469254,0.2574407,0.25018883,0.23931105,0.23024625,0.21936847,0.21030366,0.19942589,3.6494937,3.9975824,4.345671,4.691947,5.040036,5.388125,5.277534,5.1669436,5.0581656,4.947575,4.836984,4.7282066,4.6176157,4.507025,4.3982472,4.2876563,4.688321,5.087173,5.487838,5.8866897,6.2873545,7.1267557,7.9679704,8.807372,9.646774,10.487988,10.825199,11.162411,11.499621,11.836833,12.175857,12.349901,12.525759,12.699803,12.87566,13.049705,13.466686,13.885481,14.302462,14.719443,15.138238,14.494636,13.852847,13.209246,12.567456,11.925668,11.612025,11.300196,10.988366,10.674724,10.362894,17.959208,25.557333,33.15546,40.753586,48.3499,45.84257,43.335243,40.82792,38.32059,35.813263,30.852997,25.89273,20.932467,15.9722,11.011934,8.994107,6.978093,4.9602656,2.9424384,0.9246109,0.73968875,0.55476654,0.36984438,0.18492219,0.0,0.42967212,0.85934424,1.2908293,1.7205015,2.1501737,2.1302311,2.1102884,2.0903459,2.0704033,2.0504606,1.9670644,1.8854811,1.8020848,1.7205015,1.6371052,2.3151531,2.9932013,3.6694362,4.347484,5.0255322,4.4326935,3.8398547,3.247016,2.6541772,2.0631514,3.2180085,4.3728657,5.527723,6.68258,7.837437,9.175404,10.51337,11.849524,13.1874895,14.525456,14.500074,14.474693,14.449312,14.425743,14.400362,15.285088,16.169813,17.054539,17.939264,18.825804,18.22934,17.634687,17.040035,16.445383,15.850732,15.219821,14.590723,13.959812,13.330714,12.699803,12.750566,12.799516,12.850279,12.899229,12.949992,12.685299,12.420607,12.154101,11.889409,11.624716,12.027194,12.429671,12.8321495,13.234627,13.637105,13.682428,13.727753,13.773077,13.8184,13.861912,14.072216,14.282519,14.492823,14.703127,14.911617,14.155612,13.397794,12.639976,11.882156,11.124338,10.937603,10.750868,10.56232,10.375585,10.1870365,10.8143215,11.4416065,12.070704,12.697989,13.325275,13.3506565,13.374225,13.399607,13.424988,13.45037,12.977186,12.5058155,12.032633,11.559449,11.088079,11.169662,11.253058,11.334642,11.418038,11.499621,13.113158,14.724882,16.338419,17.950142,19.561867,19.540112,19.518354,19.494787,19.473032,19.449463,18.069798,16.690134,15.310469,13.930804,12.549327,13.696932,14.844538,15.992143,17.139748,18.287354,19.59994,20.912523,22.22511,23.537693,24.850279,23.992746,23.135216,22.277683,21.420153,20.562622,21.84076,23.117086,24.395224,25.673363,26.949688,28.108171,29.264841,30.423325,31.579996,32.736664,31.257288,29.77791,28.29672,26.817343,25.337965,26.157425,26.976883,27.798155,28.617615,29.437073,30.755096,32.07312,33.38933,34.707355,36.02538,36.92461,37.825653,38.72488,39.62411,40.525154,39.5806,38.63423,37.68968,36.745125,35.80057,33.1609,30.519413,27.879738,25.240065,22.600391,22.31757,22.034748,21.751925,21.469103,21.188093,21.059374,20.932467,20.80556,20.676838,20.54993,17.85587,15.159993,12.464118,9.770056,7.07418,7.948028,8.820063,9.692098,10.564133,11.437981,11.273002,11.108022,10.943042,10.778063,10.613083,8.662335,6.7134004,4.762653,2.811905,0.8629702,2.7901495,4.7173285,6.644508,8.571687,10.500679,8.423024,6.345369,4.267714,2.1900587,0.11240368,0.25018883,0.387974,0.52575916,0.66173136,0.7995165,0.8194591,0.83940166,0.85934424,0.8792868,0.89922947,1.310772,1.7205015,2.1302311,2.5399606,2.94969,3.3594196,3.7691493,4.1806917,4.590421,5.0001507,4.15531,3.3104696,2.465629,1.6207886,0.774135,0.7668832,0.75963134,0.7523795,0.7451276,0.73787576,1.2745126,1.8129625,2.3495996,2.8880494,3.4246864,2.7393866,2.0558996,1.3705997,0.6852999,0.0,1.3651608,2.7303216,4.0954823,5.4606433,6.825804,6.089741,5.3554916,4.6194286,3.8851788,3.149116,3.9395678,4.7300196,5.520471,6.3091097,7.0995617,7.3424983,7.5854354,7.8283725,8.069496,8.312433,9.229793,10.147152,11.06451,11.98187,12.899229,11.820516,10.73999,9.659465,8.580752,7.500226,7.3497505,7.1992745,7.0506115,6.9001355,6.7496595,6.5774283,6.4051967,6.2329655,6.060734,5.8866897,5.1905117,4.4925213,3.7945306,3.0983531,2.4003625,2.1519866,1.9054236,1.6570477,1.4104849,1.162109,1.214685,1.2672608,1.3198367,1.3724127,1.4249886,1.649796,1.8746033,2.0994108,2.324218,2.5508385,2.610666,2.6704938,2.7303216,2.7901495,2.8499773,2.4601903,2.0704033,1.6806163,1.2908293,0.89922947,0.75781834,0.61459434,0.47318324,0.32995918,0.18673515,0.19942589,0.21211663,0.22480737,0.2374981,0.25018883,0.2229944,0.19579996,0.16679256,0.13959812,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.05076295,0.04169814,0.034446288,0.027194439,0.01994259,0.012690738,0.045324065,0.07795739,0.11059072,0.14322405,0.17585737,0.1794833,0.18492219,0.19036107,0.19579996,0.19942589,0.15954071,0.11965553,0.07977036,0.03988518,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.030820364,0.034446288,0.03988518,0.045324065,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.26287958,0.4749962,0.6871128,0.89922947,1.1131591,1.6316663,2.1519866,2.6723068,3.1926272,3.7129474,3.049403,2.3876717,1.7241274,1.062396,0.40066472,0.3208944,0.23931105,0.15954071,0.07977036,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.6443571,3.290527,4.934884,6.5792413,8.225411,7.6724577,7.119504,6.5683637,6.01541,5.462456,4.612177,3.7618973,2.911618,2.0631514,1.2128719,1.5881553,1.9616255,2.3369088,2.712192,3.0874753,2.570781,2.0522738,1.5355793,1.017072,0.50037766,2.5852847,4.670192,6.755099,8.840006,10.924912,11.037316,11.14972,11.262123,11.374527,11.486931,9.189907,6.892884,4.594047,2.2970235,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.014503701,0.018129626,0.01994259,0.02175555,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.21211663,0.3245203,0.43692398,0.5493277,0.66173136,0.5493277,0.43692398,0.3245203,0.21211663,0.099712946,0.8194591,1.5392052,2.2607644,2.9805105,3.7002566,3.0693457,2.4402475,1.8093367,1.1802386,0.5493277,0.44236287,0.33539808,0.22662032,0.11965553,0.012690738,0.02175555,0.032633327,0.04169814,0.052575916,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.09064813,0.1794833,0.27013144,0.36077955,0.44961473,1.5446441,2.6396735,3.7347028,4.8297324,5.924762,5.0019636,4.079166,3.1581807,2.2353828,1.3125849,1.1095331,0.90829426,0.70524246,0.50219065,0.2991388,0.96268314,1.6244144,2.2879589,2.94969,3.6132345,3.4518807,3.29234,3.1327994,2.9732587,2.811905,2.6904364,2.5671551,2.4456866,2.322405,2.1991236,1.9471219,1.69512,1.4431182,1.1893034,0.93730164,0.8448406,0.7523795,0.65991837,0.56745726,0.4749962,0.42785916,0.38072214,0.33177215,0.28463513,0.2374981,0.23931105,0.24293698,0.24474995,0.24837588,0.25018883,0.24474995,0.23931105,0.23568514,0.23024625,0.22480737,3.5624714,3.9867048,4.4127507,4.836984,5.2630305,5.6872635,5.5367875,5.388125,5.237649,5.087173,4.936697,4.836984,4.7372713,4.6375585,4.537845,4.4381323,4.900438,5.3627434,5.825049,6.2873545,6.7496595,7.500226,8.2507925,8.999546,9.750113,10.500679,10.88684,11.274815,11.662788,12.050762,12.436923,12.60009,12.763257,12.92461,13.087777,13.24913,13.649796,14.05046,14.449312,14.849977,15.250641,14.63786,14.025079,13.412297,12.799516,12.186734,11.900287,11.612025,11.325577,11.037316,10.750868,19.436771,28.124489,36.812206,45.499924,54.187637,49.774887,45.362137,40.949387,36.536636,32.125698,27.437376,22.750868,18.062546,13.374225,8.6877165,7.1630154,5.638314,4.1117992,2.5870976,1.062396,0.85027945,0.63816285,0.42423326,0.21211663,0.0,0.53663695,1.0750868,1.6117238,2.1501737,2.6868105,2.663242,2.6378605,2.612479,2.5870976,2.561716,2.4366217,2.3133402,2.1882458,2.0631514,1.938057,2.5997884,3.2633326,3.925064,4.5867953,5.2503395,4.461701,3.6748753,2.8880494,2.0994108,1.3125849,2.6995013,4.0882306,5.475147,6.8620634,8.2507925,9.811753,11.374527,12.937301,14.500074,16.062849,15.687565,15.312282,14.936998,14.561715,14.188245,14.724882,15.263332,15.799969,16.336605,16.875055,16.300346,15.725637,15.149116,14.574407,13.999697,13.512011,13.024323,12.536636,12.050762,11.563075,11.849524,12.137785,12.4242325,12.712494,13.000754,12.712494,12.4242325,12.137785,11.849524,11.563075,11.724429,11.887595,12.050762,12.212116,12.375282,12.712494,13.049705,13.386916,13.724127,14.06315,14.124791,14.188245,14.249886,14.313339,14.37498,13.611723,12.850279,12.087022,11.325577,10.56232,10.411844,10.263181,10.112705,9.96223,9.811753,10.462607,11.111648,11.762501,12.413355,13.062395,13.000754,12.937301,12.87566,12.812206,12.750566,12.212116,11.675479,11.137029,10.600392,10.061942,10.375585,10.687414,10.999244,11.312886,11.624716,13.374225,15.125546,16.875055,18.624565,20.375887,20.20003,20.024172,19.850128,19.67427,19.500225,18.011784,16.525154,15.036712,13.550082,12.06164,13.550082,15.036712,16.525154,18.011784,19.500225,20.687716,21.875206,23.062696,24.250187,25.437677,24.799515,24.163166,23.525002,22.886839,22.25049,23.800573,25.350657,26.90074,28.45082,30.000904,30.26197,30.52485,30.787731,31.05061,31.311676,29.950142,28.586794,27.22526,25.861912,24.500376,25.46306,26.425743,27.388426,28.349297,29.31198,30.287354,31.262726,32.238102,33.211662,34.187035,35.225864,36.26288,37.299892,38.336906,39.375732,38.824593,38.275265,37.724125,37.174797,36.62547,33.563377,30.49947,27.437376,24.375282,21.313189,20.8255,20.337814,19.850128,19.36244,18.874754,18.76235,18.649946,18.537542,18.425138,18.312735,15.475449,12.638163,9.799063,6.9617763,4.12449,5.3119802,6.4994707,7.686961,8.874452,10.061942,9.96223,9.862516,9.762803,9.663091,9.563377,7.7757964,5.9882154,4.2006345,2.4130533,0.62547207,2.7883365,4.949388,7.112252,9.275117,11.437981,9.1500225,6.8620634,4.574105,2.2879589,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.2755703,0.48768693,0.69980353,0.9119202,1.1258497,1.6371052,2.1501737,2.663242,3.1744974,3.6875658,4.1879435,4.688321,5.186886,5.6872635,6.187641,5.137936,4.0882306,3.0367124,1.987007,0.93730164,0.8883517,0.8375887,0.7868258,0.73787576,0.6871128,1.3996071,2.1121013,2.8245957,3.53709,4.249584,3.3993049,2.5508385,1.7005589,0.85027945,0.0,1.6878681,3.3757362,5.0617914,6.7496595,8.437528,7.5256076,6.6118746,5.6999545,4.788034,3.874301,4.325729,4.7753434,5.224958,5.674573,6.1241875,6.5756154,7.02523,7.474845,7.9244595,8.375887,9.262425,10.150778,11.037316,11.925668,12.812206,11.650098,10.487988,9.324066,8.161958,6.9998484,7.28811,7.574558,7.8628187,8.149267,8.437528,8.212721,7.987913,7.763106,7.5382986,7.311678,6.249282,5.186886,4.12449,3.0620937,1.9996977,1.7748904,1.550083,1.3252757,1.1004683,0.87566096,0.85027945,0.824898,0.7995165,0.774135,0.7505665,1.0750868,1.3996071,1.7241274,2.0504606,2.374981,2.612479,2.8499773,3.0874753,3.3249733,3.5624714,3.0747845,2.5870976,2.0994108,1.6117238,1.1258497,0.9246109,0.72518504,0.52575916,0.3245203,0.12509441,0.13778515,0.15047589,0.16316663,0.17585737,0.18673515,0.17585737,0.16316663,0.15047589,0.13778515,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.0870222,0.11240368,0.13778515,0.16316663,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.15047589,0.2374981,0.3245203,0.41335547,0.50037766,1.0116332,1.5247015,2.03777,2.5508385,3.0620937,2.5508385,2.03777,1.5247015,1.0116332,0.50037766,0.40066472,0.2991388,0.19942589,0.099712946,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.1494182,2.3006494,3.4500678,4.599486,5.750717,5.5005283,5.2503395,5.0001507,4.749962,4.499773,3.8996825,3.299592,2.6995013,2.0994108,1.49932,1.5627737,1.6244144,1.6878681,1.7495089,1.8129625,1.5120108,1.2128719,0.9119202,0.61278135,0.31182957,0.63816285,0.96268314,1.2872034,1.6117238,1.938057,4.1879435,6.43783,8.6877165,10.937603,13.1874895,10.549629,7.911769,5.275721,2.6378605,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.26287958,0.40066472,0.53663695,0.6744221,0.8122072,0.6744221,0.53663695,0.40066472,0.26287958,0.12509441,1.0007553,1.8746033,2.7502642,3.6241121,4.499773,3.6748753,2.8499773,2.0250793,1.2001812,0.37528324,0.2991388,0.22480737,0.15047589,0.07433146,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.099712946,0.19942589,0.2991388,0.40066472,0.50037766,1.6371052,2.7756457,3.9123733,5.049101,6.187641,5.224958,4.262275,3.299592,2.3369088,1.3742256,1.1494182,0.9246109,0.69980353,0.4749962,0.25018883,1.1004683,1.9507477,2.7992141,3.6494937,4.499773,4.274966,4.0501585,3.825351,3.6005437,3.3757362,2.9243085,2.474694,2.0250793,1.5754645,1.1258497,1.062396,1.0007553,0.93730164,0.87566096,0.8122072,0.73787576,0.66173136,0.5873999,0.51306844,0.43692398,0.387974,0.33721104,0.28826106,0.2374981,0.18673515,0.19942589,0.21211663,0.22480737,0.2374981,0.25018883,0.25018883,0.25018883,0.25018883,0.25018883,0.25018883,3.5751622,3.9957695,4.4145637,4.835171,5.2557783,5.674573,5.4969025,5.319232,5.143375,4.9657044,4.788034,4.7916603,4.797099,4.802538,4.8079767,4.8116026,5.1651306,5.516845,5.870373,6.2220874,6.5756154,7.3298078,8.0858135,8.840006,9.594198,10.3502035,10.930351,11.510499,12.090648,12.670795,13.24913,13.363347,13.475751,13.588155,13.700559,13.812962,14.066776,14.322405,14.5780325,14.831847,15.087475,14.369541,13.653421,12.935488,12.217555,11.499621,11.628342,11.755249,11.882156,12.010877,12.137785,21.07569,30.011782,38.949688,47.887592,56.8255,51.480885,46.13446,40.789845,35.445232,30.100618,25.945307,21.789997,17.634687,13.479377,9.325879,7.6307597,5.9356394,4.2405195,2.5453994,0.85027945,0.67986095,0.5094425,0.34083697,0.17041849,0.0,0.43692398,0.87566096,1.3125849,1.7495089,2.1882458,2.1701162,2.1519866,2.13567,2.1175404,2.0994108,1.9942589,1.889107,1.7857682,1.6806163,1.5754645,2.1519866,2.7303216,3.3068438,3.8851788,4.461701,3.870675,3.2778363,2.6849976,2.0921588,1.49932,3.0675328,4.6357455,6.202145,7.7703576,9.336758,10.500679,11.662788,12.824898,13.987006,15.149116,14.7683935,14.385859,14.003323,13.620788,13.238253,13.617162,13.997884,14.376793,14.757515,15.138238,14.964193,14.791962,14.61973,14.447499,14.275268,13.68968,13.1059065,12.52032,11.934732,11.349146,11.662788,11.974618,12.28826,12.60009,12.91192,12.552953,12.192173,11.833207,11.472427,11.111648,11.234929,11.358211,11.479679,11.602961,11.724429,12.059827,12.395226,12.730623,13.064208,13.399607,13.394168,13.390542,13.385102,13.379663,13.374225,12.774135,12.175857,11.575767,10.975676,10.375585,10.20698,10.040187,9.873394,9.704789,9.537996,10.05469,10.573197,11.089892,11.608399,12.125093,12.090648,12.054388,12.019942,11.985496,11.949236,11.546759,11.144281,10.741803,10.339326,9.936848,10.154404,10.371959,10.589515,10.80707,11.024626,12.60009,14.175554,15.749206,17.32467,18.900135,18.742407,18.584679,18.426952,18.269224,18.11331,16.771717,15.431937,14.092158,12.752378,11.4126,12.835775,14.257137,15.680313,17.101677,18.52485,19.667019,20.809185,21.953163,23.095331,24.237497,23.760687,23.282066,22.805256,22.326633,21.849825,23.209547,24.56927,25.930803,27.290525,28.650248,29.0074,29.364555,29.721708,30.080675,30.437828,29.243086,28.048344,26.85179,25.657047,24.462305,25.385101,26.3079,27.230698,28.151684,29.07448,29.984589,30.894695,31.804802,32.71491,33.625015,34.596764,35.570328,36.542072,37.515636,38.48738,38.03233,37.577274,37.122223,36.667168,36.212116,33.11195,30.011782,26.911617,23.813263,20.713097,19.822933,18.932768,18.042604,17.15244,16.262274,16.287657,16.313038,16.336605,16.361988,16.38737,13.852847,11.318325,8.781991,6.247469,3.7129474,5.177821,6.642695,8.107569,9.572442,11.037316,10.674724,10.312131,9.949538,9.5869465,9.224354,7.5854354,5.9447045,4.305786,2.665055,1.0243238,2.9968271,4.9693303,6.9418335,8.914337,10.88684,8.892582,6.8983226,4.902251,2.907992,0.9119202,0.73968875,0.56745726,0.39522585,0.2229944,0.05076295,0.21936847,0.38978696,0.56020546,0.7306239,0.89922947,1.5120108,2.124792,2.7375734,3.350355,3.9631362,4.327542,4.691947,5.0581656,5.422571,5.7869763,4.9076896,4.028403,3.147303,2.268016,1.3869164,1.3325275,1.2781386,1.2219368,1.167548,1.1131591,1.5700256,2.0268922,2.4855716,2.9424384,3.3993049,2.9478772,2.4946365,2.0432088,1.5899682,1.1367276,2.3876717,3.636803,4.8877473,6.1368785,7.3878226,6.5375433,5.6872635,4.836984,3.9867048,3.1382382,3.491766,3.8471067,4.2024474,4.557788,4.9131284,5.5458527,6.1767635,6.8094873,7.4422116,8.074935,8.885329,9.695724,10.504305,11.314699,12.125093,11.062697,10.000301,8.937905,7.8755093,6.813113,7.5799966,8.34688,9.115576,9.882459,10.649343,10.174346,9.699349,9.224354,8.749357,8.274362,8.02236,7.7703576,7.518356,7.264541,7.0125394,6.3127356,5.612932,4.9131284,4.213325,3.5117085,2.9297476,2.3477864,1.7658255,1.1820517,0.6000906,0.8629702,1.1258497,1.3869164,1.649796,1.9126755,2.1701162,2.427557,2.6849976,2.9424384,3.199879,2.7430124,2.2843328,1.8274662,1.3705997,0.9119202,0.7505665,0.5873999,0.42423326,0.26287958,0.099712946,0.12690738,0.15410182,0.18310922,0.21030366,0.2374981,0.23205921,0.22662032,0.2229944,0.21755551,0.21211663,0.1794833,0.14684997,0.11421664,0.08339628,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.072518505,0.09427405,0.11784257,0.13959812,0.16316663,0.13053331,0.09789998,0.065266654,0.032633327,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.11965553,0.19036107,0.25925365,0.32995918,0.40066472,0.8103943,1.2201238,1.6298534,2.039583,2.4493124,2.039583,1.6298534,1.2201238,0.8103943,0.40066472,0.3245203,0.25018883,0.17585737,0.099712946,0.025381476,0.5293851,1.0352017,1.5392052,2.0450218,2.5508385,2.0631514,1.5754645,1.0877775,0.6000906,0.11240368,1.017072,1.9217403,2.8282216,3.73289,4.6375585,5.125245,5.612932,6.1006193,6.588306,7.07418,6.096993,5.1198063,4.1426196,3.1654327,2.1882458,2.039583,1.892733,1.745883,1.5972201,1.4503701,1.2491312,1.0497054,0.85027945,0.6508536,0.44961473,0.8919776,1.3343405,1.7767034,2.220879,2.663242,4.6393714,6.6173134,8.595256,10.573197,12.549327,10.127209,7.705091,5.282973,2.8608549,0.43692398,0.34990177,0.26287958,0.17585737,0.0870222,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.052575916,0.06707962,0.08339628,0.09789998,0.11240368,0.2574407,0.40247768,0.5475147,0.69255173,0.8375887,0.726998,0.61822027,0.5076295,0.39703882,0.28826106,0.968122,1.647983,2.327844,3.007705,3.6875658,3.0131438,2.3369088,1.6624867,0.9880646,0.31182957,0.25018883,0.18673515,0.12509441,0.06164073,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.01994259,0.027194439,0.034446288,0.04169814,0.05076295,0.64722764,1.2455053,1.84197,2.4402475,3.0367124,3.489953,3.9431937,4.3946214,4.847862,5.2992897,4.4798307,3.6603715,2.8390994,2.0196402,1.2001812,1.0333886,0.86478317,0.6979906,0.5293851,0.36259252,1.0352017,1.7078108,2.38042,3.053029,3.7256382,3.5570326,3.39024,3.2216346,3.054842,2.8880494,2.514579,2.1429217,1.7694515,1.3977941,1.0243238,0.96268314,0.89922947,0.8375887,0.774135,0.7124943,0.6399758,0.56745726,0.4949388,0.4224203,0.34990177,0.5420758,0.73424983,0.92823684,1.1204109,1.3125849,1.5156367,1.7168756,1.9199274,2.1229792,2.324218,2.1882458,2.0504606,1.9126755,1.7748904,1.6371052,3.587853,4.0030212,4.41819,4.8333583,5.2467136,5.661882,5.4570174,5.2521524,5.047288,4.842423,4.6375585,4.748149,4.856927,4.9675174,5.0781083,5.186886,5.429823,5.67276,5.915697,6.156821,6.399758,7.159389,7.9208336,8.680465,9.440096,10.199727,10.97205,11.744371,12.516694,13.290829,14.06315,14.124791,14.188245,14.249886,14.313339,14.37498,14.485571,14.594349,14.70494,14.81553,14.924308,14.103036,13.279951,12.456866,11.635593,10.812509,11.354585,11.896661,12.440549,12.982625,13.524701,22.712795,31.899076,41.08717,50.275265,59.46336,53.18507,46.908592,40.630306,34.352016,28.075539,24.45324,20.83094,17.206827,13.584529,9.96223,8.096691,6.2329655,4.367427,2.5018883,0.63816285,0.5094425,0.3825351,0.25562772,0.12690738,0.0,0.33721104,0.6744221,1.0116332,1.3506571,1.6878681,1.6769904,1.6679256,1.6570477,1.647983,1.6371052,1.551896,1.4666867,1.3832904,1.2980812,1.2128719,1.7041848,2.1973107,2.6904364,3.1817493,3.6748753,3.2778363,2.8807976,2.4819458,2.084907,1.6878681,3.435564,5.18326,6.930956,8.676839,10.424535,11.187792,11.949236,12.712494,13.475751,14.237195,13.847408,13.457622,13.067834,12.678047,12.28826,12.509441,12.732436,12.955431,13.176612,13.399607,13.629852,13.860099,14.090345,14.320591,14.5508375,13.867351,13.185677,12.50219,11.820516,11.137029,11.47424,11.813264,12.1504755,12.487686,12.824898,12.393413,11.9601145,11.526816,11.095331,10.662033,10.745429,10.827013,10.910409,10.991992,11.075388,11.407161,11.740746,12.072517,12.40429,12.737875,12.665357,12.592838,12.52032,12.447801,12.375282,11.938358,11.499621,11.062697,10.625773,10.1870365,10.002114,9.817192,9.63227,9.447348,9.262425,9.646774,10.032935,10.417283,10.801631,11.187792,11.18054,11.173288,11.164224,11.156972,11.14972,10.883214,10.614896,10.348391,10.080072,9.811753,9.935035,10.058316,10.179785,10.303066,10.424535,11.8241415,13.225562,14.625169,16.024776,17.424383,17.284784,17.145187,17.005589,16.864178,16.72458,15.531651,14.340534,13.147605,11.954676,10.761745,12.119655,13.477564,14.835473,16.193382,17.549479,18.648132,19.744976,20.841818,21.940474,23.037315,22.720047,22.402779,22.08551,21.768242,21.44916,22.620335,23.789696,24.960869,26.13023,27.299591,27.75283,28.204258,28.6575,29.11074,29.562168,28.534218,27.508081,26.480131,25.45218,24.424232,25.307144,26.190058,27.07297,27.955883,28.836983,29.681824,30.526665,31.373318,32.21816,33.063,33.96948,34.877773,35.784256,36.69255,37.600845,37.240063,36.879284,36.520317,36.15954,35.80057,32.662334,29.52591,26.38767,23.249432,20.113007,18.820364,17.527721,16.23508,14.942437,13.649796,13.812962,13.974316,14.137483,14.300649,14.462003,12.230246,9.9966755,7.764919,5.5331616,3.299592,5.041849,6.784106,8.528176,10.270433,12.012691,11.3872175,10.761745,10.138086,9.512614,8.887142,7.3950744,5.903006,4.409125,2.9170568,1.4249886,3.207131,4.989273,6.773228,8.55537,10.337513,8.63514,6.932769,5.230397,3.5280252,1.8256533,1.4666867,1.1095331,0.7523795,0.39522585,0.038072214,0.16497959,0.291887,0.42060733,0.5475147,0.6744221,1.3869164,2.0994108,2.811905,3.5243993,4.2368937,4.4671397,4.6973863,4.9276323,5.1578784,5.388125,4.6774435,3.966762,3.2578938,2.5472124,1.8383441,1.7767034,1.7168756,1.6570477,1.5972201,1.5373923,1.7404441,1.9416829,2.1447346,2.3477864,2.5508385,2.4946365,2.4402475,2.3858588,2.3296568,2.275268,3.0874753,3.8996825,4.7118897,5.52591,6.338117,5.5494785,4.762653,3.975827,3.1871881,2.4003625,2.659616,2.9206827,3.1799364,3.43919,3.7002566,4.514277,5.33011,6.14413,6.9599633,7.7757964,8.508233,9.24067,9.973107,10.705544,11.437981,10.475298,9.512614,8.549932,7.5872483,6.624565,7.8718834,9.119202,10.368333,11.615651,12.862969,12.137785,11.4126,10.687414,9.96223,9.237044,9.795437,10.352016,10.910409,11.466989,12.025381,10.850581,9.675781,8.499168,7.324369,6.149569,5.009216,3.870675,2.7303216,1.5899682,0.44961473,0.6508536,0.85027945,1.0497054,1.2491312,1.4503701,1.7277533,2.0051367,2.2825198,2.5599031,2.8372865,2.4094272,1.983381,1.5555218,1.1276628,0.69980353,0.5747091,0.44961473,0.3245203,0.19942589,0.07433146,0.11784257,0.15954071,0.2030518,0.24474995,0.28826106,0.29007402,0.291887,0.2955129,0.29732585,0.2991388,0.24837588,0.19579996,0.14322405,0.09064813,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.058014803,0.07795739,0.09789998,0.11784257,0.13778515,0.11059072,0.08339628,0.054388877,0.027194439,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.09064813,0.14322405,0.19579996,0.24837588,0.2991388,0.6073425,0.9155461,1.2219368,1.5301404,1.8383441,1.5301404,1.2219368,0.9155461,0.6073425,0.2991388,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,1.0605831,2.0704033,3.0802233,4.0900435,5.0998635,4.12449,3.150929,2.175555,1.2001812,0.22480737,0.88472575,1.5446441,2.2045624,2.864481,3.5243993,4.749962,5.975525,7.1992745,8.424837,9.6504,8.294304,6.9400206,5.5857377,4.229642,2.8753586,2.518205,2.1592383,1.8020848,1.4449311,1.0877775,0.9880646,0.8883517,0.7868258,0.6871128,0.5873999,1.1476053,1.7078108,2.268016,2.8282216,3.386614,5.092612,6.796797,8.502794,10.20698,11.912977,9.704789,7.498413,5.290225,3.0820365,0.87566096,0.69980353,0.52575916,0.34990177,0.17585737,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.07977036,0.08520924,0.09064813,0.09427405,0.099712946,0.2520018,0.40429065,0.55839247,0.7106813,0.8629702,0.7795739,0.6979906,0.61459434,0.533011,0.44961473,0.9354887,1.4195497,1.9054236,2.3894846,2.8753586,2.3495996,1.8256533,1.2998942,0.774135,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.03988518,0.054388877,0.07070554,0.08520924,0.099712946,1.1947423,2.2897718,3.3848011,4.4798307,5.57486,5.3428006,5.1107416,4.876869,4.64481,4.4127507,3.7347028,3.056655,2.38042,1.7023718,1.0243238,0.9155461,0.80495536,0.69436467,0.5855869,0.4749962,0.969935,1.4648738,1.9598125,2.4547513,2.94969,2.8390994,2.7303216,2.619731,2.5091403,2.4003625,2.1048496,1.8093367,1.5156367,1.2201238,0.9246109,0.8629702,0.7995165,0.73787576,0.6744221,0.61278135,0.5420758,0.47318324,0.40247768,0.33177215,0.26287958,0.6979906,1.1331016,1.5682126,2.0033236,2.4366217,2.8300345,3.2234476,3.6150475,4.006647,4.40006,4.12449,3.8507326,3.5751622,3.299592,3.0258346,3.6005437,4.0102735,4.420003,4.8297324,5.239462,5.6491914,5.4171324,5.185073,4.953014,4.7191415,4.4870825,4.702825,4.9167547,5.132497,5.3482394,5.562169,5.6945157,5.826862,5.959208,6.093367,6.2257137,6.9907837,7.755854,8.520925,9.284182,10.049252,11.015561,11.980057,12.944552,13.910862,14.875358,14.888049,14.90074,14.911617,14.924308,14.936998,14.902553,14.868106,14.831847,14.7974,14.762955,13.834718,12.908294,11.980057,11.05182,10.125396,11.082641,12.039885,12.9971285,13.954373,14.911617,24.349901,33.78637,43.224655,52.662937,62.099407,54.889256,47.680916,40.468952,33.260612,26.050459,22.959358,19.87007,16.78078,13.68968,10.600392,8.564435,6.530291,4.494334,2.4601903,0.42423326,0.34083697,0.25562772,0.17041849,0.08520924,0.0,0.2374981,0.4749962,0.7124943,0.9499924,1.1874905,1.1856775,1.1820517,1.1802386,1.1766127,1.1747998,1.1095331,1.0442665,0.9808127,0.9155461,0.85027945,1.258196,1.6642996,2.0722163,2.4801328,2.8880494,2.6849976,2.4819458,2.280707,2.077655,1.8746033,3.8017826,5.730775,7.6579537,9.585134,11.512312,11.874905,12.237497,12.60009,12.962683,13.325275,12.928236,12.529385,12.132345,11.735307,11.338268,11.401722,11.466989,11.532255,11.597522,11.662788,12.295512,12.928236,13.559147,14.191871,14.824595,14.045021,13.265448,12.485873,11.704487,10.924912,11.287505,11.650098,12.012691,12.375282,12.737875,12.232059,11.728055,11.222239,10.718235,10.212419,10.254116,10.297627,10.339326,10.382836,10.424535,10.754494,11.084454,11.4144125,11.744371,12.07433,11.934732,11.795135,11.655537,11.514126,11.374527,11.10077,10.825199,10.549629,10.275872,10.000301,9.79725,9.594198,9.39296,9.189907,8.9868555,9.24067,9.492672,9.744674,9.9966755,10.25049,10.270433,10.290376,10.310318,10.330261,10.3502035,10.217857,10.085511,9.953164,9.820818,9.686659,9.715667,9.742861,9.770056,9.79725,9.824444,11.050007,12.27557,13.499319,14.724882,15.950445,15.827164,15.705695,15.582414,15.459132,15.337664,14.293397,13.247317,12.203052,11.156972,10.112705,11.405348,12.697989,13.990632,15.283275,16.574104,17.627436,18.680767,19.732285,20.785616,21.837133,21.679407,21.521679,21.365765,21.208036,21.050308,22.029308,23.01012,23.990934,24.969934,25.950747,26.49826,27.045776,27.59329,28.140804,28.68832,27.827162,26.96782,26.10666,25.247316,24.387972,25.229187,26.072214,26.915243,27.75827,28.599485,29.38087,30.160446,30.94002,31.719593,32.49917,33.342194,34.185223,35.02825,35.869465,36.712494,36.4478,36.183105,35.916603,35.65191,35.38722,32.21272,29.038221,25.861912,22.687414,19.512917,17.817797,16.122677,14.427556,12.732436,11.037316,11.338268,11.637406,11.938358,12.237497,12.536636,10.607644,8.676839,6.7478466,4.8170414,2.8880494,4.9076896,6.92733,8.94697,10.968424,12.988064,12.099712,11.213174,10.324821,9.438283,8.549932,7.2047133,5.859495,4.514277,3.1708715,1.8256533,3.4174345,5.009216,6.60281,8.194591,9.788185,8.3777,6.967215,5.5567303,4.1480584,2.7375734,2.1954978,1.651609,1.1095331,0.56745726,0.025381476,0.11059072,0.19579996,0.27919623,0.36440548,0.44961473,1.261822,2.0758421,2.8880494,3.7002566,4.512464,4.606738,4.702825,4.797099,4.893186,4.98746,4.4471974,3.9069343,3.3666716,2.8282216,2.2879589,2.222692,2.1574254,2.0921588,2.0268922,1.9616255,1.9108626,1.8582866,1.8057107,1.7531348,1.7005589,2.0432088,2.3858588,2.7266958,3.0693457,3.4119956,3.787279,4.162562,4.537845,4.9131284,5.2884116,4.5632267,3.8380418,3.1128569,2.3876717,1.6624867,1.8274662,1.9924458,2.1574254,2.322405,2.4873846,3.484514,4.4816437,5.480586,6.4777155,7.474845,8.129324,8.785617,9.440096,10.094576,10.750868,9.8878975,9.024928,8.161958,7.3008003,6.43783,8.165584,9.893337,11.619277,13.347031,15.074784,14.09941,13.125849,12.1504755,11.175101,10.199727,11.566701,12.935488,14.302462,15.6694355,17.038223,15.386614,13.736817,12.087022,10.437225,8.78743,7.0904965,5.391751,3.6948178,1.9978848,0.2991388,0.43692398,0.5747091,0.7124943,0.85027945,0.9880646,1.2853905,1.5827163,1.8800422,2.1773682,2.474694,2.077655,1.6806163,1.2817645,0.88472575,0.48768693,0.40066472,0.31182957,0.22480737,0.13778515,0.05076295,0.10696479,0.16497959,0.2229944,0.27919623,0.33721104,0.3480888,0.35715362,0.3680314,0.3770962,0.387974,0.3154555,0.24293698,0.17041849,0.09789998,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.04169814,0.059827764,0.07795739,0.09427405,0.11240368,0.09064813,0.06707962,0.045324065,0.02175555,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.059827764,0.09427405,0.13053331,0.16497959,0.19942589,0.40429065,0.6091554,0.81583315,1.020698,1.2255627,1.020698,0.81583315,0.6091554,0.40429065,0.19942589,0.17585737,0.15047589,0.12509441,0.099712946,0.07433146,1.5899682,3.105605,4.6194286,6.1350656,7.650702,6.187641,4.7245803,3.2633326,1.8002719,0.33721104,0.7523795,1.167548,1.5827163,1.9978848,2.4130533,4.3746786,6.338117,8.299743,10.263181,12.224807,10.491614,8.760235,7.027043,5.295664,3.5624714,2.9950142,2.427557,1.8600996,1.2926424,0.72518504,0.72518504,0.72518504,0.72518504,0.72518504,0.72518504,1.403233,2.079468,2.7575161,3.435564,4.1117992,5.5458527,6.978093,8.410334,9.842574,11.274815,9.282369,7.2899227,5.297477,3.3050308,1.3125849,1.0497054,0.7868258,0.52575916,0.26287958,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.10696479,0.10333887,0.09789998,0.092461094,0.0870222,0.24837588,0.40791658,0.56745726,0.726998,0.8883517,0.8321498,0.7777609,0.72337204,0.6671702,0.61278135,0.90285534,1.1929294,1.4830034,1.7730774,2.0631514,1.6878681,1.3125849,0.93730164,0.5620184,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.059827764,0.08339628,0.10515183,0.12690738,0.15047589,1.742257,3.3358512,4.9276323,6.5194135,8.113008,7.1956487,6.2764764,5.3591175,4.441758,3.5243993,2.9895754,2.4547513,1.9199274,1.3851035,0.85027945,0.79770356,0.7451276,0.69255173,0.6399758,0.5873999,0.90466833,1.2219368,1.5392052,1.8582866,2.175555,2.1229792,2.0704033,2.0178273,1.9652514,1.9126755,1.69512,1.4775645,1.260009,1.0424535,0.824898,0.76325727,0.69980353,0.63816285,0.5747091,0.51306844,0.44417584,0.3770962,0.3100166,0.24293698,0.17585737,0.8520924,1.5301404,2.2081885,2.8844235,3.5624714,4.1444325,4.7282066,5.3101673,5.8921285,6.474089,6.0625467,5.6491914,5.237649,4.8242936,4.4127507,3.6132345,4.017525,4.421816,4.8279195,5.23221,5.638314,5.377247,5.1179934,4.856927,4.597673,4.3366065,4.6575007,4.9783955,5.297477,5.618371,5.9374523,5.959208,5.9827766,6.004532,6.0281005,6.049856,6.8203654,7.590874,8.3595705,9.130079,9.900589,11.057259,12.215742,13.372412,14.530895,15.687565,15.649493,15.613234,15.575162,15.537089,15.50083,15.319533,15.140051,14.960567,14.779271,14.599788,13.568212,12.534823,11.503247,10.469859,9.438283,10.810696,12.183108,13.555521,14.927934,16.300346,25.987005,35.675476,45.362137,55.05061,64.73727,56.595253,48.45324,40.30941,32.167397,24.025381,21.46729,18.9092,16.352922,13.794832,11.236742,9.03218,6.827617,4.6230545,2.4166791,0.21211663,0.17041849,0.12690738,0.08520924,0.04169814,0.0,0.13778515,0.2755703,0.41335547,0.5493277,0.6871128,0.69255173,0.6979906,0.7016165,0.7070554,0.7124943,0.6671702,0.62184614,0.57833505,0.533011,0.48768693,0.8103943,1.1331016,1.455809,1.7767034,2.0994108,2.0921588,2.084907,2.077655,2.0704033,2.0631514,4.169814,6.2782893,8.384952,10.493427,12.60009,12.562017,12.525759,12.487686,12.449615,12.413355,12.007251,11.602961,11.1968565,10.792566,10.388275,10.2958145,10.203354,10.109079,10.016619,9.924157,10.959359,11.99456,13.029762,14.064963,15.100165,14.222692,13.345218,12.467744,11.59027,10.712796,11.10077,11.486931,11.874905,12.262879,12.650853,12.072517,11.494183,10.917661,10.339326,9.762803,9.764616,9.768243,9.770056,9.771869,9.775495,10.101828,10.429974,10.75812,11.084454,11.4126,11.204109,10.997431,10.790753,10.582263,10.375585,10.263181,10.150778,10.038374,9.924157,9.811753,9.592385,9.373016,9.151835,8.9324665,8.713099,8.832754,8.952409,9.072064,9.19172,9.313189,9.360326,9.407463,9.4546,9.501737,9.550687,9.5525,9.554313,9.557939,9.5597515,9.563377,9.494485,9.427405,9.360326,9.293246,9.224354,10.275872,11.325577,12.375282,13.424988,14.474693,14.369541,14.26439,14.159238,14.054086,13.9507475,13.05333,12.155914,11.256684,10.359268,9.461852,10.689227,11.916603,13.145792,14.373167,15.600543,16.606737,17.614744,18.622751,19.630758,20.636953,20.64058,20.642391,20.644205,20.647831,20.649643,21.440096,22.230547,23.019186,23.809637,24.60009,25.241879,25.885479,26.52727,27.17087,27.812658,27.120108,26.427555,25.735004,25.042452,24.349901,25.153044,25.954372,26.757515,27.560658,28.361986,29.078106,29.792414,30.506721,31.222841,31.93715,32.71491,33.492672,34.27043,35.04819,35.824142,35.655537,35.485115,35.314697,35.14428,34.975674,31.763105,28.550535,25.337965,22.125395,18.912827,16.815228,14.71763,12.620032,10.522435,8.424837,8.861761,9.300498,9.737422,10.174346,10.613083,8.985043,7.3570023,5.730775,4.102734,2.474694,4.7717175,7.0705543,9.367578,11.664601,13.961625,12.812206,11.662788,10.51337,9.362139,8.212721,7.0143523,5.8177967,4.6194286,3.4228733,2.2245052,3.6277382,5.029158,6.432391,7.835624,9.237044,8.120259,7.0016613,5.8848767,4.7680917,3.6494937,2.9224956,2.1954978,1.4666867,0.73968875,0.012690738,0.054388877,0.09789998,0.13959812,0.18310922,0.22480737,1.1367276,2.0504606,2.962381,3.874301,4.788034,4.748149,4.708264,4.668379,4.6266804,4.5867953,4.216951,3.8471067,3.4772623,3.1074178,2.7375734,2.666868,2.5979755,2.5272698,2.4583774,2.3876717,2.079468,1.7730774,1.4648738,1.1566701,0.85027945,1.5899682,2.3296568,3.0693457,3.8108473,4.550536,4.4870825,4.4254417,4.361988,4.3003473,4.2368937,3.5751622,2.911618,2.2498865,1.5881553,0.9246109,0.99531645,1.064209,1.1349145,1.2056202,1.2745126,2.4547513,3.63499,4.8152285,5.995467,7.175706,7.752228,8.330563,8.907085,9.48542,10.061942,9.300498,8.537241,7.7757964,7.0125394,6.249282,8.457471,10.665659,12.872034,15.080223,17.288412,16.062849,14.837286,13.611723,12.387974,11.162411,13.339779,15.517147,17.694515,19.871883,22.049252,19.92446,17.799667,15.674874,13.550082,11.42529,9.169965,6.9146395,4.6593137,2.4058013,0.15047589,0.22480737,0.2991388,0.37528324,0.44961473,0.52575916,0.8430276,1.1602961,1.4775645,1.794833,2.1121013,1.74407,1.3778516,1.0098201,0.6417888,0.2755703,0.22480737,0.17585737,0.12509441,0.07433146,0.025381476,0.09789998,0.17041849,0.24293698,0.3154555,0.387974,0.40429065,0.4224203,0.4405499,0.45686656,0.4749962,0.3825351,0.29007402,0.19761293,0.10515183,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.027194439,0.04169814,0.058014803,0.072518505,0.0870222,0.07070554,0.052575916,0.034446288,0.018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.030820364,0.047137026,0.065266654,0.08339628,0.099712946,0.2030518,0.3045777,0.40791658,0.5094425,0.61278135,0.5094425,0.40791658,0.3045777,0.2030518,0.099712946,0.099712946,0.099712946,0.099712946,0.099712946,0.099712946,2.1193533,4.1408067,6.1604466,8.180087,10.199727,8.2507925,6.300045,4.349297,2.4003625,0.44961473,0.6200332,0.7904517,0.96087015,1.1294757,1.2998942,3.9993954,6.70071,9.400211,12.099712,14.799213,12.690738,10.58045,8.470161,6.359873,4.249584,3.4718235,2.6958754,1.9181144,1.1403534,0.36259252,0.46230546,0.5620184,0.66173136,0.76325727,0.8629702,1.6570477,2.4529383,3.247016,4.0429068,4.836984,5.99728,7.157576,8.317872,9.4781685,10.636651,8.859948,7.083245,5.3047285,3.5280252,1.7495089,1.3996071,1.0497054,0.69980353,0.34990177,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.13415924,0.11965553,0.10515183,0.09064813,0.07433146,0.24293698,0.40972954,0.57833505,0.7451276,0.9119202,0.88472575,0.8575313,0.83033687,0.8031424,0.774135,0.87022203,0.9644961,1.0605831,1.1548572,1.2491312,1.0243238,0.7995165,0.5747091,0.34990177,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.07977036,0.11059072,0.13959812,0.17041849,0.19942589,2.2897718,4.3801174,6.4704633,8.560809,10.649343,9.046683,7.4440246,5.8431783,4.2405195,2.6378605,2.2444477,1.8528478,1.4594349,1.067835,0.6744221,0.67986095,0.6852999,0.69073874,0.69436467,0.69980353,0.83940166,0.9808127,1.1204109,1.260009,1.3996071,1.405046,1.4104849,1.4141108,1.4195497,1.4249886,1.2853905,1.1457924,1.0043813,0.86478317,0.72518504,0.66173136,0.6000906,0.53663695,0.4749962,0.41335547,0.3480888,0.28282216,0.21755551,0.15228885,0.0870222,1.0080072,1.9271792,2.8481643,3.7673361,4.688321,5.4606433,6.2329655,7.0052876,7.7776093,8.549932,8.000604,7.4494634,6.9001355,6.350808,5.7996674,3.6241121,4.024777,4.4254417,4.8242936,5.224958,5.6256227,5.337362,5.050914,4.762653,4.4743915,4.1879435,4.612177,5.038223,5.462456,5.8866897,6.3127356,6.2257137,6.1368785,6.049856,5.962834,5.8758116,6.6499467,7.424082,8.200029,8.974165,9.750113,11.10077,12.449615,13.800271,15.149116,16.499773,16.41275,16.325727,16.236893,16.14987,16.062849,15.738328,15.411995,15.087475,14.762955,14.436621,13.299893,12.163166,11.024626,9.8878975,8.749357,10.536939,12.32452,14.112101,15.899682,17.687263,27.624111,37.56277,47.49962,57.438282,67.37513,58.29944,49.22556,40.149868,31.074179,22.000301,19.975222,17.950142,15.925063,13.899984,11.874905,9.499924,7.124943,4.749962,2.374981,0.0,0.0,0.0,0.0,0.0,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.19942589,0.21211663,0.22480737,0.2374981,0.25018883,0.22480737,0.19942589,0.17585737,0.15047589,0.12509441,0.36259252,0.6000906,0.8375887,1.0750868,1.3125849,1.49932,1.6878681,1.8746033,2.0631514,2.2498865,4.537845,6.825804,9.11195,11.399909,13.687867,13.24913,12.812206,12.375282,11.938358,11.499621,11.088079,10.674724,10.263181,9.849826,9.438283,9.188094,8.937905,8.6877165,8.437528,8.187339,9.625018,11.062697,12.500377,13.938056,15.375735,14.400362,13.424988,12.449615,11.47424,10.500679,10.912222,11.325577,11.73712,12.1504755,12.562017,11.912977,11.262123,10.613083,9.96223,9.313189,9.275117,9.237044,9.200785,9.162713,9.12464,9.449161,9.775495,10.100015,10.424535,10.750868,10.475298,10.199727,9.924157,9.6504,9.374829,9.425592,9.474543,9.525306,9.574255,9.625018,9.38752,9.1500225,8.912524,8.675026,8.437528,8.424837,8.412147,8.399456,8.386765,8.375887,8.450218,8.52455,8.600695,8.675026,8.749357,8.887142,9.024928,9.162713,9.300498,9.438283,9.275117,9.11195,8.950596,8.78743,8.624263,9.499924,10.375585,11.249433,12.125093,13.000754,12.91192,12.824898,12.737875,12.650853,12.562017,11.813264,11.062697,10.312131,9.563377,8.812811,9.97492,11.137029,12.299138,13.46306,14.625169,15.5878525,16.550535,17.513218,18.475903,19.436771,19.59994,19.763105,19.92446,20.087626,20.250792,20.850883,21.44916,22.049252,22.649342,23.249432,23.987309,24.725183,25.46306,26.199121,26.936998,26.413052,25.887293,25.363346,24.837587,24.311829,25.075085,25.838343,26.599787,27.363045,28.124489,28.775343,29.424383,30.075235,30.724277,31.37513,32.087624,32.800117,33.512615,34.22511,34.937603,34.86327,34.787125,34.712795,34.63665,34.562317,31.311676,28.062847,24.812206,21.561563,18.312735,15.812659,13.312584,10.812509,8.312433,5.812358,6.3870673,6.9617763,7.5382986,8.113008,8.6877165,7.362441,6.037165,4.7118897,3.386614,2.0631514,4.6375585,7.211965,9.788185,12.362592,14.936998,13.524701,12.112403,10.700105,9.287807,7.8755093,6.825804,5.774286,4.7245803,3.6748753,2.6251698,3.8380418,5.049101,6.261973,7.474845,8.6877165,7.8628187,7.037921,6.2130227,5.388125,4.5632267,3.6494937,2.7375734,1.8256533,0.9119202,0.0,0.0,0.0,0.0,0.0,0.0,1.0116332,2.0250793,3.0367124,4.0501585,5.0617914,4.8877473,4.7118897,4.537845,4.361988,4.1879435,3.9867048,3.787279,3.587853,3.386614,3.1871881,3.1128569,3.0367124,2.962381,2.8880494,2.811905,2.2498865,1.6878681,1.1258497,0.5620184,0.0,1.1367276,2.275268,3.4119956,4.550536,5.6872635,5.186886,4.688321,4.1879435,3.6875658,3.1871881,2.5870976,1.987007,1.3869164,0.7868258,0.18673515,0.16316663,0.13778515,0.11240368,0.0870222,0.06164073,1.4249886,2.7883365,4.1498713,5.5132194,6.874754,7.3751316,7.8755093,8.375887,8.874452,9.374829,8.713099,8.049554,7.3878226,6.7242785,6.0625467,8.749357,11.437981,14.124791,16.813416,19.500225,18.024473,16.550535,15.074784,13.600845,12.125093,15.112856,18.100618,21.08838,24.07433,27.062092,24.462305,21.862516,19.262728,16.66294,14.06315,11.249433,8.437528,5.6256227,2.811905,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.40066472,0.73787576,1.0750868,1.4122978,1.7495089,1.4122978,1.0750868,0.73787576,0.40066472,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0870222,0.17585737,0.26287958,0.34990177,0.43692398,0.46230546,0.48768693,0.51306844,0.53663695,0.5620184,0.44961473,0.33721104,0.22480737,0.11240368,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,2.6505513,5.1741953,7.699652,10.225109,12.750566,10.312131,7.8755093,5.4370747,3.000453,0.5620184,0.48768693,0.41335547,0.33721104,0.26287958,0.18673515,3.625925,7.061489,10.500679,13.938056,17.375433,14.888049,12.400664,9.91328,7.424082,4.936697,3.9504454,2.962381,1.9743162,0.9880646,0.0,0.19942589,0.40066472,0.6000906,0.7995165,1.0007553,1.9126755,2.8245957,3.738329,4.650249,5.562169,6.450521,7.3370595,8.225411,9.11195,10.000301,8.437528,6.874754,5.3119802,3.7492065,2.1882458,1.7495089,1.3125849,0.87566096,0.43692398,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.16316663,0.13778515,0.11240368,0.0870222,0.06164073,0.2374981,0.41335547,0.5873999,0.76325727,0.93730164,0.93730164,0.93730164,0.93730164,0.93730164,0.93730164,0.8375887,0.73787576,0.63816285,0.53663695,0.43692398,0.36259252,0.28826106,0.21211663,0.13778515,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.099712946,0.13778515,0.17585737,0.21211663,0.25018883,2.8372865,5.426197,8.013294,10.600392,13.1874895,10.899531,8.611572,6.3254266,4.0374675,1.7495089,1.49932,1.2491312,1.0007553,0.7505665,0.50037766,0.5620184,0.62547207,0.6871128,0.7505665,0.8122072,0.774135,0.73787576,0.69980353,0.66173136,0.62547207,0.6871128,0.7505665,0.8122072,0.87566096,0.93730164,0.87566096,0.8122072,0.7505665,0.6871128,0.62547207,0.5620184,0.50037766,0.43692398,0.37528324,0.31182957,0.25018883,0.18673515,0.12509441,0.06164073,0.0,1.162109,2.326031,3.48814,4.650249,5.812358,6.775041,7.7377243,8.700407,9.663091,10.625773,9.936848,9.249735,8.562622,7.8755093,7.1883965,3.7129474,4.004834,4.2967215,4.590421,4.882308,5.1741953,5.0146546,4.855114,4.695573,4.5342193,4.3746786,4.9802084,5.5857377,6.189454,6.794984,7.400513,7.324369,7.250037,7.175706,7.0995617,7.02523,7.5781837,8.129324,8.682278,9.235231,9.788185,10.98474,12.183108,13.379663,14.5780325,15.774588,15.747393,15.720199,15.693004,15.66581,15.636803,15.531651,15.428311,15.32316,15.218008,15.112856,13.954373,12.797703,11.63922,10.48255,9.325879,12.31908,15.314095,18.310923,21.305937,24.299137,31.525606,38.750263,45.97492,53.199574,60.42423,52.06466,43.70509,35.34552,26.984135,18.624565,16.80979,14.995013,13.180238,11.365462,9.550687,7.6398244,5.730775,3.8199122,1.9108626,0.0,0.058014803,0.11421664,0.17223145,0.23024625,0.28826106,0.25925365,0.23205921,0.20486477,0.17767033,0.15047589,0.16316663,0.17585737,0.18673515,0.19942589,0.21211663,0.24837588,0.28282216,0.31726846,0.35171473,0.387974,0.52213323,0.65810543,0.79226464,0.92823684,1.062396,1.5446441,2.0268922,2.5091403,2.9932013,3.4754493,5.524097,7.574558,9.625018,11.675479,13.724127,13.234627,12.745127,12.255627,11.764315,11.274815,10.89228,10.509744,10.127209,9.744674,9.362139,9.349448,9.336758,9.325879,9.313189,9.300498,10.194288,11.089892,11.985496,12.879286,13.77489,12.9971285,12.219368,11.4416065,10.665659,9.8878975,10.4045925,10.9230995,11.439794,11.958302,12.474996,11.735307,10.995618,10.254116,9.514427,8.774739,8.700407,8.624263,8.549932,8.4756,8.399456,8.780178,9.159087,9.539809,9.920531,10.29944,10.00574,9.710228,9.414715,9.119202,8.825501,8.9651,9.104698,9.244296,9.385707,9.525306,9.28962,9.055748,8.820063,8.584378,8.350506,8.3777,8.404895,8.432089,8.459284,8.488291,8.557183,8.627889,8.696781,8.767487,8.838193,9.102885,9.367578,9.63227,9.896963,10.161655,10.014805,9.867955,9.719293,9.572442,9.425592,10.234174,11.044568,11.854962,12.665357,13.475751,13.67699,13.880041,14.083094,14.284332,14.487384,13.589968,12.692551,11.795135,10.897718,10.000301,10.991992,11.985496,12.977186,13.97069,14.96238,15.854358,16.748148,17.640125,18.532103,19.425894,19.739536,20.054993,20.370447,20.685904,20.999546,21.432844,21.864328,22.297626,22.729113,23.16241,24.126905,25.093216,26.05771,27.022207,27.986704,27.515333,27.04215,26.57078,26.097597,25.624413,26.046833,26.469254,26.891674,27.315907,27.738327,28.024776,28.313036,28.599485,28.887745,29.174194,29.61293,30.049854,30.486778,30.925516,31.36244,31.69965,32.03686,32.375885,32.713097,33.05031,30.015408,26.980509,23.94561,20.910711,17.87581,15.319533,12.76507,10.210606,7.654328,5.0998635,5.714458,6.3308654,6.94546,7.560054,8.174648,7.230095,6.285541,5.3391747,4.3946214,3.4500678,5.7217097,7.995165,10.266808,12.540262,14.811904,13.347031,11.882156,10.417283,8.952409,7.4875355,6.5719895,5.658256,4.74271,3.827164,2.911618,4.070101,5.2267714,6.3852544,7.5419245,8.700407,8.1148205,7.5292335,6.94546,6.359873,5.774286,4.6194286,3.4645715,2.3097143,1.1548572,0.0,0.032633327,0.065266654,0.09789998,0.13053331,0.16316663,1.0406405,1.9181144,2.7955883,3.673062,4.550536,4.358362,4.164375,3.972201,3.780027,3.587853,3.53709,3.48814,3.437377,3.386614,3.3376641,3.1581807,2.9768846,2.7974012,2.617918,2.4366217,2.521831,2.6070402,2.6922495,2.7774587,2.8626678,4.6393714,6.4178877,8.194591,9.973107,11.74981,10.040187,8.330563,6.6191263,4.9095025,3.199879,2.6251698,2.0504606,1.4757515,0.89922947,0.3245203,0.65991837,0.99531645,1.3307146,1.6642996,1.9996977,3.3104696,4.6194286,5.9302006,7.2391596,8.549932,9.084756,9.619579,10.154404,10.689227,11.225864,10.419096,9.6141405,8.809185,8.00423,7.1992745,9.131892,11.06451,12.9971285,14.929747,16.862366,15.656745,14.452938,13.247317,12.0416975,10.837891,13.075087,15.312282,17.549479,19.786674,22.025682,20.740292,19.4549,18.169512,16.88412,15.600543,12.714307,9.829884,6.94546,4.059223,1.1747998,0.9499924,0.72518504,0.50037766,0.2755703,0.05076295,0.3208944,0.58921283,0.85934424,1.1294757,1.3996071,1.1331016,0.86478317,0.5982776,0.32995918,0.06164073,0.052575916,0.04169814,0.032633327,0.02175555,0.012690738,0.08520924,0.15772775,0.23024625,0.30276474,0.37528324,0.39522585,0.41516843,0.43511102,0.4550536,0.4749962,0.38072214,0.28463513,0.19036107,0.09427405,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.027194439,0.054388877,0.08339628,0.11059072,0.13778515,2.1501737,4.162562,6.1749506,8.187339,10.199727,8.24898,6.300045,4.349297,2.4003625,0.44961473,0.38978696,0.32995918,0.27013144,0.21030366,0.15047589,2.9007401,5.6491914,8.399456,11.14972,13.899984,11.909351,9.920531,7.9298983,5.9392653,3.9504454,3.1744974,2.4003625,1.6244144,0.85027945,0.07433146,0.21936847,0.36440548,0.5094425,0.6544795,0.7995165,2.9678197,5.1343102,7.3026133,9.470917,11.637406,11.777005,11.918416,12.058014,12.197612,12.337211,10.252303,8.167397,6.0824895,3.9975824,1.9126755,1.5301404,1.1476053,0.7650702,0.3825351,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.09427405,0.19036107,0.28463513,0.38072214,0.4749962,0.39159992,0.3100166,0.22662032,0.14503701,0.06164073,0.21574254,0.3680314,0.52032024,0.6726091,0.824898,1.0478923,1.2708868,1.4920682,1.7150626,1.938057,1.6226015,1.3071461,0.9916905,0.678048,0.36259252,0.2991388,0.2374981,0.17585737,0.11240368,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.052575916,0.092461094,0.13234627,0.17223145,0.21211663,0.72337204,1.2328146,1.742257,2.2516994,2.762955,4.847862,6.932769,9.017676,11.102583,13.1874895,10.832452,8.477413,6.1223745,3.7673361,1.4122978,1.209246,1.0080072,0.80495536,0.60190356,0.40066472,0.44961473,0.50037766,0.5493277,0.6000906,0.6508536,0.6200332,0.58921283,0.56020546,0.5293851,0.50037766,0.5493277,0.6000906,0.6508536,0.69980353,0.7505665,0.69980353,0.6508536,0.6000906,0.5493277,0.50037766,0.44961473,0.40066472,0.34990177,0.2991388,0.25018883,0.25925365,0.27013144,0.27919623,0.29007402,0.2991388,1.5845293,2.8699198,4.15531,5.4407005,6.7242785,7.3751316,8.025986,8.675026,9.324066,9.97492,9.474543,8.974165,8.4756,7.9752226,7.474845,3.7999697,3.9848917,4.169814,4.3547363,4.539658,4.7245803,4.691947,4.6593137,4.6266804,4.59586,4.5632267,5.3482394,6.1332526,6.9182653,7.703278,8.488291,8.424837,8.363196,8.299743,8.238102,8.174648,8.504607,8.834567,9.164526,9.494485,9.824444,10.870523,11.91479,12.96087,14.005136,15.049402,15.082036,15.114669,15.147303,15.179935,15.212569,15.326786,15.442815,15.557032,15.673061,15.787278,14.610665,13.43224,12.255627,11.077202,9.900589,14.103036,18.305483,22.50793,26.710379,30.912825,35.42529,39.93775,44.45022,48.96268,53.475143,45.82988,38.184616,30.539354,22.89409,15.250641,13.644357,12.039885,10.435412,8.829127,7.224656,5.7797246,4.3347936,2.8898623,1.4449311,0.0,0.11421664,0.23024625,0.3444629,0.4604925,0.5747091,0.48224804,0.38978696,0.29732585,0.20486477,0.11240368,0.12509441,0.13778515,0.15047589,0.16316663,0.17585737,0.27013144,0.36440548,0.4604925,0.55476654,0.6508536,0.68167394,0.71430725,0.7469406,0.7795739,0.8122072,1.5899682,2.3677292,3.1454902,3.923251,4.699199,6.5121617,8.325124,10.138086,11.949236,13.762199,13.220123,12.678047,12.134158,11.592083,11.050007,10.698292,10.344765,9.99305,9.639522,9.287807,9.512614,9.737422,9.96223,10.1870365,10.411844,10.765372,11.117086,11.470614,11.822329,12.175857,11.595709,11.015561,10.435412,9.855265,9.275117,9.896963,10.520622,11.142468,11.764315,12.387974,11.557636,10.7273,9.896963,9.066626,8.238102,8.125698,8.013294,7.900891,7.7866745,7.6742706,8.109382,8.544493,8.979604,9.414715,9.849826,9.53437,9.220728,8.9052725,8.589817,8.274362,8.504607,8.734854,8.9651,9.195346,9.425592,9.19172,8.9596615,8.727602,8.495543,8.26167,8.330563,8.397643,8.464723,8.531802,8.600695,8.664148,8.729415,8.794682,8.859948,8.925215,9.316814,9.710228,10.101828,10.49524,10.88684,10.754494,10.622148,10.489801,10.357455,10.225109,10.970237,11.715364,12.460492,13.20562,13.9507475,14.4420595,14.935185,15.428311,15.919624,16.41275,15.366671,14.322405,13.278138,12.232059,11.187792,12.010877,12.8321495,13.655234,14.478319,15.299591,16.122677,16.94576,17.767033,18.590118,19.413204,19.879135,20.34688,20.814623,21.282368,21.750113,22.014805,22.279497,22.54419,22.810696,23.075388,24.268316,25.459433,26.652363,27.845293,29.038221,28.617615,28.197006,27.778214,27.357605,26.936998,27.020395,27.101978,27.185373,27.266956,27.350353,27.27421,27.199877,27.125546,27.049402,26.97507,27.138237,27.299591,27.462757,27.624111,27.787277,28.537844,29.286598,30.037165,30.787731,31.538298,28.717327,25.89817,23.0772,20.258043,17.437075,14.828221,12.217555,9.606889,6.9980354,4.3873696,5.041849,5.6981416,6.352621,7.0071006,7.663393,7.0977483,6.532104,5.9682727,5.4026284,4.836984,6.8076744,8.776552,10.747242,12.717933,14.68681,13.16936,11.651911,10.13446,8.617011,7.0995617,6.319988,5.540414,4.76084,3.9794528,3.199879,4.3021603,5.4044414,6.506723,7.610817,8.713099,8.366822,8.02236,7.6778965,7.3316207,6.987158,5.5893636,4.1933823,2.7955883,1.3977941,0.0,0.065266654,0.13053331,0.19579996,0.25925365,0.3245203,1.067835,1.8093367,2.5526514,3.294153,4.0374675,3.827164,3.6168604,3.4083695,3.198066,2.9877625,3.0874753,3.1871881,3.2869012,3.386614,3.48814,3.2016919,2.9170568,2.6324217,2.3477864,2.0631514,2.7955883,3.5280252,4.2604623,4.992899,5.7253356,8.1420145,10.560507,12.977186,15.3956785,17.812357,14.891675,11.972805,9.052122,6.1332526,3.2125697,2.663242,2.1121013,1.5627737,1.0116332,0.46230546,1.1566701,1.8528478,2.5472124,3.24339,3.9377546,5.195951,6.452334,7.71053,8.966913,10.225109,10.794379,11.365462,11.934732,12.5058155,13.075087,12.126906,11.18054,10.232361,9.284182,8.337815,9.514427,10.692853,11.869466,13.047892,14.224504,13.290829,12.35534,11.419851,10.484363,9.550687,11.037316,12.525759,14.012388,15.50083,16.98746,17.01828,17.047287,17.078108,17.107115,17.137936,14.17918,11.222239,8.265296,5.3083544,2.3495996,1.887294,1.4249886,0.96268314,0.50037766,0.038072214,0.23931105,0.44236287,0.64541465,0.8466535,1.0497054,0.8520924,0.6544795,0.45686656,0.25925365,0.06164073,0.054388877,0.047137026,0.03988518,0.032633327,0.025381476,0.08339628,0.13959812,0.19761293,0.25562772,0.31182957,0.32814622,0.34264994,0.35715362,0.37165734,0.387974,0.3100166,0.23205921,0.15410182,0.07795739,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,1.649796,3.149116,4.650249,6.149569,7.650702,6.187641,4.7245803,3.2633326,1.8002719,0.33721104,0.291887,0.24837588,0.2030518,0.15772775,0.11240368,2.175555,4.2368937,6.300045,8.363196,10.424535,8.9324665,7.440398,5.9483304,4.454449,2.962381,2.4003625,1.8383441,1.2745126,0.7124943,0.15047589,0.23931105,0.32995918,0.42060733,0.5094425,0.6000906,4.022964,7.4440246,10.866898,14.289771,17.712645,17.105303,16.49796,15.890617,15.283275,14.674119,12.067079,9.460039,6.8529987,4.2441454,1.6371052,1.310772,0.9826257,0.6544795,0.32814622,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.15228885,0.3045777,0.45686656,0.6091554,0.76325727,0.62184614,0.48224804,0.34264994,0.2030518,0.06164073,0.19217403,0.32270733,0.45324063,0.581961,0.7124943,1.1566701,1.6026589,2.0468347,2.4928236,2.9369993,2.4076142,1.8782293,1.3470312,0.81764615,0.28826106,0.2374981,0.18673515,0.13778515,0.0870222,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.092461094,0.15954071,0.22662032,0.2955129,0.36259252,1.3452182,2.327844,3.3104696,4.2930956,5.275721,6.8584375,8.439341,10.022058,11.6047735,13.1874895,10.765372,8.341441,5.919323,3.4972048,1.0750868,0.91917205,0.7650702,0.6091554,0.4550536,0.2991388,0.33721104,0.37528324,0.41335547,0.44961473,0.48768693,0.46411842,0.44236287,0.42060733,0.39703882,0.37528324,0.41335547,0.44961473,0.48768693,0.52575916,0.5620184,0.52575916,0.48768693,0.44961473,0.41335547,0.37528324,0.33721104,0.2991388,0.26287958,0.22480737,0.18673515,0.27013144,0.35171473,0.43511102,0.5166943,0.6000906,2.0069497,3.4156215,4.8224807,6.2293396,7.6380115,7.9752226,8.312433,8.649645,8.9868555,9.325879,9.012237,8.700407,8.386765,8.074935,7.763106,3.8869917,3.9649491,4.0429068,4.120864,4.1970086,4.274966,4.36924,4.465327,4.559601,4.655688,4.749962,5.714458,6.680767,7.645263,8.609759,9.574255,9.525306,9.474543,9.425592,9.374829,9.325879,9.432844,9.539809,9.646774,9.755551,9.862516,10.754494,11.648285,12.540262,13.43224,14.324218,14.416678,14.50914,14.601601,14.695875,14.788336,15.121921,15.457319,15.792717,16.128115,16.4617,15.265145,14.066776,12.870221,11.671853,10.475298,15.885179,21.29506,26.704939,32.11482,37.5247,39.32497,41.125244,42.925514,44.72579,46.524246,39.595104,32.66596,25.735004,18.804049,11.874905,10.480737,9.084756,7.690587,6.294606,4.900438,3.919625,2.9406252,1.9598125,0.9808127,0.0,0.17223145,0.3444629,0.5166943,0.69073874,0.8629702,0.70524246,0.5475147,0.38978696,0.23205921,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.13778515,0.291887,0.44780177,0.60190356,0.75781834,0.9119202,0.8430276,0.77232206,0.7016165,0.6327239,0.5620184,1.6352923,2.7067533,3.780027,4.853301,5.924762,7.500226,9.07569,10.649343,12.224807,13.800271,13.20562,12.609155,12.0145035,11.419851,10.825199,10.502492,10.179785,9.857078,9.53437,9.211663,9.675781,10.138086,10.600392,11.062697,11.525003,11.334642,11.144281,10.955733,10.765372,10.57501,10.192475,9.80994,9.427405,9.04487,8.662335,9.389333,10.118144,10.845142,11.57214,12.299138,11.379966,10.460794,9.539809,8.620637,7.699652,7.549176,7.400513,7.250037,7.0995617,6.9508986,7.440398,7.9298983,8.419398,8.910711,9.400211,9.064813,8.729415,8.39583,8.0604315,7.7250338,8.044115,8.365009,8.685904,9.004985,9.325879,9.0956335,8.865387,8.63514,8.404895,8.174648,8.281613,8.39039,8.497355,8.604321,8.713099,8.772926,8.832754,8.892582,8.952409,9.012237,9.5325575,10.052877,10.573197,11.091705,11.612025,11.494183,11.378153,11.26031,11.142468,11.024626,11.704487,12.384347,13.064208,13.745882,14.425743,15.20713,15.99033,16.771717,17.554916,18.338116,17.145187,15.952258,14.759329,13.568212,12.375282,13.027949,13.680615,14.333282,14.984136,15.636803,16.389181,17.143373,17.895754,18.648132,19.400513,20.020546,20.64058,21.260612,21.880646,22.500679,22.596766,22.694666,22.792566,22.890465,22.988365,24.407915,25.827465,27.247015,28.668377,30.087927,29.719896,29.351864,28.985645,28.617615,28.249582,27.992142,27.734701,27.47726,27.21982,26.96238,26.525455,26.08672,25.649796,25.212872,24.774134,24.66173,24.549326,24.436922,24.324518,24.212114,25.374224,26.538147,27.700254,28.862364,30.024473,27.419247,24.815832,22.210604,19.605377,17.00015,14.335095,11.67004,9.004985,6.33993,3.6748753,4.36924,5.0654173,5.7597823,6.454147,7.1503243,6.965402,6.78048,6.5955577,6.4106355,6.2257137,7.891826,9.5597515,11.227677,12.895603,14.561715,12.99169,11.421664,9.851639,8.281613,6.7134004,6.0679855,5.422571,4.7771564,4.1317415,3.48814,4.5342193,5.582112,6.630004,7.6778965,8.725789,8.620637,8.515485,8.410334,8.3051815,8.200029,6.5592985,4.9203806,3.2796493,1.6407311,0.0,0.09789998,0.19579996,0.291887,0.38978696,0.48768693,1.0950294,1.7023718,2.3097143,2.9170568,3.5243993,3.2977788,3.0693457,2.8427253,2.6142921,2.3876717,2.6378605,2.8880494,3.1382382,3.386614,3.636803,3.247016,2.857229,2.467442,2.077655,1.6878681,3.0675328,4.4471974,5.826862,7.208339,8.588004,11.644659,14.703127,17.75978,20.818249,23.874905,19.744976,15.6150465,11.485118,7.3551893,3.2252605,2.6995013,2.175555,1.649796,1.1258497,0.6000906,1.6552348,2.7103791,3.7655232,4.8206677,5.8758116,7.079619,8.285239,9.490859,10.694666,11.900287,12.5058155,13.109532,13.715062,14.320591,14.924308,13.834718,12.745127,11.655537,10.564133,9.474543,9.896963,10.319383,10.741803,11.164224,11.586644,10.9230995,10.257742,9.592385,8.927028,8.26167,8.999546,9.737422,10.475298,11.213174,11.949236,13.294455,14.639673,15.984891,17.330109,18.675327,15.644054,12.6145935,9.585134,6.5556726,3.5243993,2.8245957,2.124792,1.4249886,0.72518504,0.025381476,0.15954071,0.2955129,0.42967212,0.5656443,0.69980353,0.5728962,0.44417584,0.31726846,0.19036107,0.06164073,0.058014803,0.052575916,0.047137026,0.04169814,0.038072214,0.07977036,0.12328146,0.16497959,0.20667773,0.25018883,0.25925365,0.27013144,0.27919623,0.29007402,0.2991388,0.23931105,0.1794833,0.11965553,0.059827764,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.032633327,0.065266654,0.09789998,0.13053331,0.16316663,1.1494182,2.137483,3.1255474,4.1117992,5.0998635,4.12449,3.150929,2.175555,1.2001812,0.22480737,0.19579996,0.16497959,0.13415924,0.10515183,0.07433146,1.4503701,2.8245957,4.2006345,5.57486,6.9508986,5.955582,4.9602656,3.9649491,2.9696326,1.9743162,1.6244144,1.2745126,0.9246109,0.5747091,0.22480737,0.25925365,0.2955129,0.32995918,0.36440548,0.40066472,5.0781083,9.755551,14.432995,19.11044,23.787882,22.431786,21.077503,19.72322,18.367125,17.01284,13.881854,10.752681,7.6216946,4.4925213,1.3633479,1.0895905,0.81764615,0.54570174,0.27194437,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.21030366,0.42060733,0.630911,0.83940166,1.0497054,0.8520924,0.6544795,0.45686656,0.25925365,0.06164073,0.17041849,0.27738327,0.38434806,0.49312583,0.6000906,1.2672608,1.9344311,2.6034143,3.2705846,3.9377546,3.1926272,2.4474995,1.7023718,0.9572442,0.21211663,0.17585737,0.13778515,0.099712946,0.06164073,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.13234627,0.22662032,0.32270733,0.4169814,0.51306844,1.9670644,3.4228733,4.876869,6.3326783,7.7866745,8.8672,9.947725,11.028252,12.106964,13.1874895,10.696479,8.207282,5.718084,3.2270734,0.73787576,0.629098,0.52213323,0.41516843,0.30820364,0.19942589,0.22480737,0.25018883,0.2755703,0.2991388,0.3245203,0.3100166,0.2955129,0.27919623,0.26469254,0.25018883,0.2755703,0.2991388,0.3245203,0.34990177,0.37528324,0.34990177,0.3245203,0.2991388,0.2755703,0.25018883,0.22480737,0.19942589,0.17585737,0.15047589,0.12509441,0.27919623,0.43511102,0.58921283,0.7451276,0.89922947,2.42937,3.9595103,5.4896507,7.019791,8.549932,8.575313,8.600695,8.624263,8.649645,8.675026,8.549932,8.424837,8.299743,8.174648,8.049554,3.975827,3.9450066,3.9141862,3.8851788,3.8543584,3.825351,4.0483456,4.269527,4.4925213,4.7155156,4.936697,6.0824895,7.228282,8.372261,9.518054,10.662033,10.625773,10.587702,10.549629,10.51337,10.475298,10.359268,10.245051,10.130835,10.014805,9.900589,10.640278,11.379966,12.119655,12.859344,13.600845,13.753134,13.905423,14.057712,14.210001,14.362289,14.917056,15.471823,16.028402,16.583168,17.137936,15.919624,14.703127,13.484816,12.268318,11.050007,17.66732,24.284634,30.901947,37.521072,44.138386,43.224655,42.312733,41.400814,40.48708,39.57516,33.360325,27.145489,20.92884,14.7140045,8.499168,7.315304,6.1296263,4.945762,3.7600844,2.5744069,2.0595255,1.5446441,1.0297627,0.5148814,0.0,0.23024625,0.4604925,0.69073874,0.91917205,1.1494182,0.92823684,0.70524246,0.48224804,0.25925365,0.038072214,0.05076295,0.06164073,0.07433146,0.0870222,0.099712946,0.3154555,0.5293851,0.7451276,0.96087015,1.1747998,1.0025684,0.83033687,0.65810543,0.48587397,0.31182957,1.6806163,3.04759,4.4145637,5.7833505,7.1503243,8.488291,9.824444,11.162411,12.500377,13.838344,13.189302,12.542075,11.894848,11.24762,10.600392,10.306692,10.014805,9.7229185,9.429218,9.137331,9.837135,10.536939,11.236742,11.938358,12.638163,11.9057255,11.173288,10.440851,9.706602,8.974165,8.789243,8.604321,8.419398,8.234476,8.049554,8.881703,9.715667,10.547816,11.379966,12.212116,11.202296,10.192475,9.182655,8.172835,7.1630154,6.9744673,6.787732,6.599184,6.412449,6.2257137,6.7696023,7.315304,7.859193,8.404895,8.950596,8.595256,8.239915,7.8845744,7.5292335,7.175706,7.5854354,7.995165,8.404895,8.814624,9.224354,8.997733,8.7693,8.54268,8.314246,8.087626,8.234476,8.383139,8.529989,8.676839,8.825501,8.87989,8.934279,8.990481,9.04487,9.099259,9.7483,10.395528,11.042755,11.689982,12.337211,12.235684,12.132345,12.03082,11.927481,11.8241415,12.440549,13.055143,13.669738,14.284332,14.90074,15.9722,17.045475,18.116936,19.190208,20.26167,18.92189,17.582111,16.242332,14.902553,13.562773,14.045021,14.527269,15.009518,15.491765,15.975826,16.6575,17.339174,18.022661,18.704334,19.387821,20.160145,20.932467,21.704788,22.47711,23.249432,23.18054,23.109835,23.03913,22.970236,22.89953,24.547514,26.195496,27.841667,29.489649,31.137632,30.822176,30.506721,30.193079,29.877623,29.562168,28.965704,28.367426,27.769148,27.172684,26.574406,25.774889,24.975372,24.175856,23.374527,22.57501,22.187037,21.800875,21.4129,21.024927,20.636953,22.212418,23.787882,25.363346,26.936998,28.512463,26.122978,23.73168,21.342196,18.952711,16.563227,13.8419695,11.122525,8.403082,5.6818247,2.962381,3.6966307,4.4326935,5.1669436,5.903006,6.637256,6.833056,7.027043,7.2228427,7.41683,7.61263,8.977791,10.342952,11.708113,13.073273,14.436621,12.815832,11.193231,9.570629,7.948028,6.3254266,5.814171,5.3047285,4.795286,4.2858434,3.774588,4.7680917,5.7597823,6.7532854,7.744976,8.736667,8.872639,9.006798,9.142771,9.27693,9.412902,7.5292335,5.6473784,3.7655232,1.8818551,0.0,0.13053331,0.25925365,0.38978696,0.52032024,0.6508536,1.1222239,1.5954071,2.0667772,2.5399606,3.0131438,2.7683938,2.521831,2.277081,2.032331,1.7875811,2.1882458,2.5870976,2.9877625,3.386614,3.787279,3.29234,2.7974012,2.3024626,1.8075237,1.3125849,3.339477,5.368182,7.3950744,9.421967,11.450671,15.147303,18.845747,22.542377,26.24082,29.93745,24.596464,19.257288,13.918114,8.577126,3.2379513,2.7375734,2.2371957,1.7368182,1.2382535,0.73787576,2.1519866,3.5679104,4.9820213,6.397945,7.8120556,8.9651,10.118144,11.269376,12.42242,13.575464,14.21544,14.855415,15.495391,16.135366,16.775343,15.542528,14.309713,13.0769,11.845898,10.613083,10.279498,9.947725,9.6141405,9.282369,8.950596,8.55537,8.160145,7.764919,7.369693,6.9744673,6.9617763,6.9490857,6.9382076,6.925517,6.9128265,9.572442,12.232059,14.891675,17.553104,20.212719,17.108929,14.006948,10.90497,7.802991,4.699199,3.7618973,2.8245957,1.887294,0.9499924,0.012690738,0.07977036,0.14684997,0.21574254,0.28282216,0.34990177,0.291887,0.23568514,0.17767033,0.11965553,0.06164073,0.059827764,0.058014803,0.054388877,0.052575916,0.05076295,0.07795739,0.10515183,0.13234627,0.15954071,0.18673515,0.19217403,0.19761293,0.2030518,0.20667773,0.21211663,0.17041849,0.12690738,0.08520924,0.04169814,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.034446288,0.07070554,0.10515183,0.13959812,0.17585737,0.6508536,1.1258497,1.6008459,2.0758421,2.5508385,2.0631514,1.5754645,1.0877775,0.6000906,0.11240368,0.09789998,0.08339628,0.06707962,0.052575916,0.038072214,0.72518504,1.4122978,2.0994108,2.7883365,3.4754493,2.9768846,2.4801328,1.9815681,1.4848163,0.9880646,0.85027945,0.7124943,0.5747091,0.43692398,0.2991388,0.27919623,0.25925365,0.23931105,0.21936847,0.19942589,6.1332526,12.065266,17.99728,23.929293,29.86312,27.760082,25.657047,23.555822,21.452785,19.34975,15.6966305,12.045323,8.392203,4.7390842,1.0877775,0.87022203,0.6526665,0.43511102,0.21755551,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.26831847,0.53482395,0.8031424,1.0696479,1.3379664,1.0823387,0.82671094,0.5728962,0.31726846,0.06164073,0.14684997,0.23205921,0.31726846,0.40247768,0.48768693,1.3778516,2.268016,3.1581807,4.0483456,4.936697,3.97764,3.0167696,2.0577126,1.0968424,0.13778515,0.11240368,0.0870222,0.06164073,0.038072214,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.17223145,0.2955129,0.4169814,0.5402629,0.66173136,2.5907235,4.517903,6.445082,8.372261,10.29944,10.877775,11.454298,12.032633,12.609155,13.1874895,10.629399,8.071309,5.5150323,2.956942,0.40066472,0.34083697,0.27919623,0.21936847,0.15954071,0.099712946,0.11240368,0.12509441,0.13778515,0.15047589,0.16316663,0.15410182,0.14684997,0.13959812,0.13234627,0.12509441,0.13778515,0.15047589,0.16316663,0.17585737,0.18673515,0.17585737,0.16316663,0.15047589,0.13778515,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.29007402,0.5166943,0.7451276,0.97174793,1.2001812,2.8517902,4.505212,6.156821,7.8102427,9.461852,9.175404,8.887142,8.600695,8.312433,8.024173,8.087626,8.149267,8.212721,8.274362,8.337815,4.062849,3.925064,3.787279,3.6494937,3.5117085,3.3757362,3.7256382,4.07554,4.4254417,4.7753434,5.125245,6.450521,7.7757964,9.099259,10.424535,11.74981,11.724429,11.700861,11.675479,11.650098,11.624716,11.287505,10.950294,10.613083,10.275872,9.936848,10.524248,11.111648,11.700861,12.28826,12.87566,13.087777,13.299893,13.512011,13.724127,13.938056,14.712192,15.488139,16.262274,17.038223,17.812357,16.575916,15.337664,14.09941,12.862969,11.624716,19.449463,27.27421,35.10077,42.925514,50.750263,47.124336,43.500225,39.8743,36.250187,32.62426,27.125546,21.625017,16.124489,10.625773,5.125245,4.1498713,3.1744974,2.1991236,1.2255627,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.28826106,0.5747091,0.8629702,1.1494182,1.4376793,1.1494182,0.8629702,0.5747091,0.28826106,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.33721104,0.61278135,0.8883517,1.162109,1.4376793,1.162109,0.8883517,0.61278135,0.33721104,0.06164073,1.7241274,3.386614,5.050914,6.7134004,8.375887,9.474543,10.57501,11.675479,12.774135,13.874602,13.174799,12.474996,11.775192,11.075388,10.375585,10.112705,9.849826,9.5869465,9.325879,9.063,10.000301,10.937603,11.874905,12.812206,13.749508,12.474996,11.200482,9.924157,8.649645,7.3751316,7.3878226,7.400513,7.413204,7.4258947,7.4367723,8.375887,9.313189,10.25049,11.187792,12.125093,11.024626,9.924157,8.825501,7.7250338,6.624565,6.399758,6.1749506,5.9501433,5.7253356,5.5005283,6.1006193,6.70071,7.3008003,7.900891,8.499168,8.125698,7.750415,7.3751316,6.9998484,6.624565,7.124943,7.6253204,8.125698,8.624263,9.12464,8.899834,8.675026,8.450218,8.225411,8.000604,8.187339,8.375887,8.562622,8.749357,8.937905,8.9868555,9.037619,9.088382,9.137331,9.188094,9.96223,10.738177,11.512312,12.28826,13.062395,12.975373,12.888351,12.799516,12.712494,12.625471,13.174799,13.724127,14.275268,14.824595,15.375735,16.73727,18.100618,19.462152,20.8255,22.187037,20.700407,19.211964,17.725336,16.236893,14.750263,15.062093,15.375735,15.687565,15.999394,16.313038,16.92582,17.536787,18.149569,18.76235,19.375132,20.299742,21.224354,22.150776,23.075388,23.999998,23.7625,23.525002,23.287504,23.050007,22.812508,24.68711,26.561714,28.438131,30.312735,32.187336,31.924458,31.663391,31.400513,31.137632,30.874752,29.93745,29.000149,28.062847,27.125546,26.188244,25.024323,23.862213,22.700104,21.537996,20.375887,19.712341,19.050611,18.387066,17.725336,17.06179,19.050611,21.037619,23.024624,25.011631,27.000452,24.824896,22.649342,20.4756,18.300045,16.124489,13.3506565,10.57501,7.799365,5.0255322,2.2498865,3.0258346,3.7999697,4.5759177,5.3500524,6.1241875,6.70071,7.2754188,7.850128,8.424837,8.999546,10.061942,11.124338,12.186734,13.24913,14.313339,12.638163,10.962985,9.287807,7.61263,5.9374523,5.562169,5.186886,4.8116026,4.4381323,4.062849,5.0001507,5.9374523,6.874754,7.8120556,8.749357,9.12464,9.499924,9.875207,10.25049,10.625773,8.499168,6.3743763,4.249584,2.124792,0.0,0.16316663,0.3245203,0.48768693,0.6508536,0.8122072,1.1494182,1.4866294,1.8256533,2.1628644,2.5000753,2.2371957,1.9743162,1.7132497,1.4503701,1.1874905,1.7368182,2.2879589,2.8372865,3.386614,3.9377546,3.3376641,2.7375734,2.137483,1.5373923,0.93730164,3.6132345,6.2873545,8.963287,11.637406,14.313339,18.649946,22.986553,27.324972,31.663391,35.999996,29.449764,22.89953,16.349297,9.799063,3.2506418,2.7756457,2.3006494,1.8256533,1.3506571,0.87566096,2.6505513,4.4254417,6.200332,7.9752226,9.750113,10.850581,11.949236,13.049705,14.150173,15.250641,15.925063,16.599485,17.27572,17.950142,18.624565,17.25034,15.8743,14.500074,13.125849,11.74981,10.662033,9.574255,8.488291,7.400513,6.3127356,6.187641,6.0625467,5.9374523,5.812358,5.6872635,4.9258194,4.162562,3.3993049,2.6378605,1.8746033,5.8504305,9.824444,13.800271,17.774284,21.750113,18.575615,15.399304,12.224807,9.050309,5.8758116,4.699199,3.5243993,2.3495996,1.1747998,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07433146,0.15047589,0.22480737,0.2991388,0.37528324,0.2991388,0.22480737,0.15047589,0.07433146,0.0,7.1883965,14.37498,21.563377,28.74996,35.93836,33.086567,30.238403,27.386612,24.536636,21.686659,17.511406,13.337966,9.162713,4.98746,0.8122072,0.6508536,0.48768693,0.3245203,0.16316663,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.3245203,0.6508536,0.97537386,1.2998942,1.6244144,1.3125849,1.0007553,0.6871128,0.37528324,0.06164073,0.12509441,0.18673515,0.25018883,0.31182957,0.37528324,1.4884423,2.5997884,3.7129474,4.8242936,5.9374523,4.762653,3.587853,2.4130533,1.2382535,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.21211663,0.36259252,0.51306844,0.66173136,0.8122072,3.2125697,5.612932,8.013294,10.411844,12.812206,12.888351,12.962683,13.037014,13.113158,13.1874895,10.56232,7.93715,5.3119802,2.6868105,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.2991388,0.6000906,0.89922947,1.2001812,1.49932,3.2742105,5.050914,6.825804,8.600695,10.375585,9.775495,9.175404,8.575313,7.9752226,7.3751316,7.6253204,7.8755093,8.125698,8.375887,8.624263,4.099108,4.0519714,4.004834,3.9576974,3.9105604,3.8616104,4.137181,4.4127507,4.688321,4.9620786,5.237649,6.5701766,7.902704,9.235231,10.567759,11.900287,12.059827,12.219368,12.380721,12.540262,12.699803,12.328146,11.954676,11.583018,11.209548,10.837891,11.184166,11.532255,11.880343,12.22662,12.574709,12.855718,13.134913,13.41411,13.695119,13.974316,14.828221,15.680313,16.532406,17.384499,18.238403,16.936697,15.636803,14.336908,13.037014,11.73712,19.948027,28.157122,36.36803,44.577126,52.788033,48.600086,44.412144,40.2242,36.03807,31.850126,26.376793,20.905272,15.431937,9.960417,4.4870825,3.8144734,3.141864,2.469255,1.7966459,1.1258497,1.0932164,1.0605831,1.0279498,0.99531645,0.96268314,1.1222239,1.2817645,1.4431182,1.6026589,1.7621996,1.4141108,1.067835,0.7197462,0.37165734,0.025381476,0.030820364,0.034446288,0.03988518,0.045324065,0.05076295,0.27738327,0.5058166,0.7324369,0.96087015,1.1874905,1.162109,1.1367276,1.1131591,1.0877775,1.062396,2.3006494,3.53709,4.7753434,6.011784,7.250037,8.716724,10.185224,11.651911,13.12041,14.587097,14.084907,13.582716,13.080525,12.578335,12.07433,11.6047735,11.135216,10.665659,10.194288,9.724731,10.246864,10.770811,11.292944,11.815077,12.337211,11.225864,10.112705,8.999546,7.8882003,6.775041,6.9055743,7.0342946,7.1648283,7.2953615,7.4258947,8.056806,8.689529,9.322253,9.954978,10.587702,9.663091,8.736667,7.8120556,6.887445,5.962834,5.7470913,5.5331616,5.317419,5.101677,4.8877473,5.9374523,6.987158,8.036863,9.088382,10.138086,9.333132,8.528176,7.723221,6.9182653,6.11331,6.630004,7.1466985,7.665206,8.1819,8.700407,8.488291,8.274362,8.062244,7.850128,7.6380115,7.607191,7.5781837,7.5473633,7.518356,7.4875355,7.6706448,7.851941,8.03505,8.21816,8.399456,9.1500225,9.900589,10.649343,11.399909,12.1504755,12.119655,12.090648,12.059827,12.03082,11.999999,12.6417885,13.28539,13.927178,14.57078,15.212569,16.507025,17.803293,19.097748,20.392202,21.686659,20.397642,19.106813,17.817797,16.526966,15.23795,15.674874,16.1118,16.550535,16.98746,17.424383,18.04079,18.655384,19.26998,19.884573,20.499168,21.052122,21.605076,22.15803,22.70917,23.262123,23.24218,23.222239,23.202295,23.182352,23.16241,24.837587,26.512764,28.187943,29.86312,31.538298,31.066927,30.59737,30.127811,29.658255,29.186884,28.151684,27.118294,26.083092,25.047892,24.01269,22.799818,21.586945,20.374073,19.163015,17.950142,17.462456,16.97477,16.487082,15.999394,15.511708,17.29929,19.08687,20.87445,22.662033,24.449614,22.580448,20.70947,18.840307,16.96933,15.100165,12.692551,10.284937,7.877322,5.469708,3.0620937,3.975827,4.8877473,5.7996674,6.7134004,7.6253204,8.39039,9.155461,9.920531,10.685601,11.450671,11.760688,12.070704,12.380721,12.690738,13.000754,11.539507,10.080072,8.620637,7.159389,5.6999545,5.3428006,4.985647,4.6266804,4.269527,3.9123733,4.7227674,5.5331616,6.341743,7.1521373,7.9625316,8.479226,8.997733,9.514427,10.032935,10.549629,8.439341,6.3308654,4.220577,2.1102884,0.0,0.13053331,0.25925365,0.38978696,0.52032024,0.6508536,0.9644961,1.2799516,1.5954071,1.9108626,2.2245052,2.0105755,1.794833,1.5790904,1.3651608,1.1494182,1.6896812,2.229944,2.770207,3.3104696,3.8507326,3.2306993,2.610666,1.9906329,1.3705997,0.7505665,4.071914,7.3950744,10.718235,14.039582,17.362743,19.837437,22.31213,24.786825,27.26333,29.738026,24.697989,19.657953,14.617917,9.577881,4.537845,4.1299286,3.7220123,3.3140955,2.907992,2.5000753,4.17344,5.844991,7.518356,9.189907,10.863272,11.744371,12.627284,13.510198,14.39311,15.27421,15.464571,15.654932,15.845293,16.035654,16.224201,15.027647,13.829279,12.632723,11.434355,10.2378,9.626831,9.017676,8.406708,7.797552,7.1883965,7.039734,6.892884,6.7442207,6.5973706,6.450521,5.678199,4.9058766,4.1317415,3.3594196,2.5870976,5.600241,8.611572,11.624716,14.63786,17.64919,15.06028,12.469557,9.880646,7.2899227,4.699199,3.7600844,2.819157,1.8800422,0.93911463,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.052575916,0.054388877,0.058014803,0.059827764,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.12690738,0.13053331,0.13234627,0.13415924,0.13778515,0.11421664,0.092461094,0.07070554,0.047137026,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.030820364,0.034446288,0.03988518,0.045324065,0.05076295,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.09789998,0.08339628,0.06707962,0.052575916,0.038072214,0.032633327,0.027194439,0.02175555,0.018129626,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.027194439,0.054388877,0.08339628,0.11059072,0.13778515,0.13959812,0.14322405,0.14503701,0.14684997,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.6726091,1.3452182,2.0178273,2.6904364,3.3630457,3.0421512,2.72307,2.4021754,2.0830941,1.7621996,1.4104849,1.0569572,0.70524246,0.35171473,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.07977036,0.13415924,0.19036107,0.24474995,0.2991388,0.75781834,1.214685,1.6733645,2.1302311,2.5870976,7.893639,13.196554,18.503096,23.807825,29.112553,27.05484,24.997128,22.939415,20.881702,18.825804,15.189,11.555823,7.9190207,4.2858434,0.6508536,0.52032024,0.38978696,0.25925365,0.13053331,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.1349145,2.269829,3.4047437,4.539658,5.674573,4.550536,3.4246864,2.3006494,1.1747998,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,0.2991388,1.5555218,2.810092,4.064662,5.319232,6.5756154,5.2865987,3.9993954,2.712192,1.4249886,0.13778515,0.11240368,0.0870222,0.06164073,0.038072214,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.70342946,1.3415923,1.983381,2.6233568,3.2633326,3.48814,3.7129474,3.9377546,4.162562,4.3873696,6.697084,9.006798,11.318325,13.628039,15.937754,14.891675,13.847408,12.803142,11.757062,10.712796,8.580752,6.446895,4.314851,2.182807,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.25562772,0.49675176,0.73968875,0.9826257,1.2255627,2.7176309,4.209699,5.7017674,7.1956487,8.6877165,8.406708,8.127511,7.8483152,7.567306,7.28811,7.474845,7.663393,7.850128,8.036863,8.225411,4.137181,4.1806917,4.2223897,4.265901,4.307599,4.349297,4.550536,4.749962,4.949388,5.1506267,5.3500524,6.6898317,8.029612,9.3693905,10.70917,12.050762,12.395226,12.739688,13.084151,13.430427,13.77489,13.366973,12.96087,12.552953,12.145037,11.73712,11.845898,11.952863,12.059827,12.166792,12.27557,12.621845,12.969934,13.318023,13.664299,14.012388,14.942437,15.872487,16.802538,17.732588,18.662638,17.29929,15.937754,14.574407,13.212872,11.849524,20.444778,29.040035,37.635292,46.230545,54.8258,50.07584,45.32588,40.574104,35.824142,31.074179,25.629852,20.185526,14.739386,9.295059,3.8507326,3.4808881,3.1092308,2.7393866,2.3695421,1.9996977,1.9851941,1.9706904,1.9543737,1.93987,1.9253663,1.9579996,1.9906329,2.0232663,2.0558996,2.08672,1.6806163,1.2726997,0.86478317,0.45686656,0.05076295,0.047137026,0.045324065,0.04169814,0.03988518,0.038072214,0.21755551,0.39703882,0.57833505,0.75781834,0.93730164,1.162109,1.3869164,1.6117238,1.8383441,2.0631514,2.8753586,3.6875658,4.499773,5.3119802,6.1241875,7.9607186,9.795437,11.630155,13.464873,15.299591,14.995013,14.690435,14.385859,14.079468,13.77489,13.096842,12.420607,11.7425585,11.06451,10.388275,10.49524,10.602205,10.70917,10.817947,10.924912,9.97492,9.024928,8.074935,7.124943,6.1749506,6.4233265,6.6698895,6.9182653,7.1648283,7.413204,7.7395372,8.067683,8.39583,8.722163,9.050309,8.299743,7.549176,6.8004227,6.049856,5.2992897,5.0944247,4.88956,4.6846952,4.4798307,4.274966,5.774286,7.2754188,8.774739,10.275872,11.775192,10.540565,9.305937,8.069496,6.834869,5.600241,6.1350656,6.6698895,7.2047133,7.7395372,8.274362,8.074935,7.8755093,7.6742706,7.474845,7.2754188,7.027043,6.78048,6.532104,6.285541,6.037165,6.352621,6.6680765,6.981719,7.2971745,7.61263,8.337815,9.063,9.788185,10.51337,11.236742,11.26575,11.292944,11.320138,11.347333,11.374527,12.11059,12.84484,13.580903,14.315152,15.049402,16.276777,17.504154,18.733343,19.960718,21.188093,20.094877,19.001661,17.910257,16.817041,15.725637,16.287657,16.849674,17.411694,17.975525,18.537542,19.155762,19.77217,20.39039,21.006798,21.625017,21.8045,21.985798,22.165281,22.344765,22.524246,22.72186,22.919474,23.117086,23.3147,23.512312,24.988064,26.462002,27.937754,29.411692,30.887444,30.209396,29.533161,28.855112,28.177065,27.50083,26.367727,25.234627,24.103338,22.970236,21.837133,20.575312,19.311678,18.049856,16.788034,15.524399,15.212569,14.90074,14.587097,14.275268,13.961625,15.54978,17.137936,18.724277,20.312433,21.900587,20.334188,18.769602,17.205015,15.640429,14.075842,12.034446,9.994863,7.95528,5.915697,3.874301,4.9258194,5.975525,7.02523,8.074935,9.12464,10.080072,11.035503,11.990934,12.944552,13.899984,13.457622,13.015259,12.572895,12.130532,11.6881695,10.442664,9.197159,7.951654,6.7079616,5.462456,5.121619,4.782595,4.441758,4.102734,3.7618973,4.445384,5.127058,5.810545,6.492219,7.175706,7.835624,8.495543,9.155461,9.815379,10.475298,8.379513,6.285541,4.1897564,2.0957847,0.0,0.09789998,0.19579996,0.291887,0.38978696,0.48768693,0.7795739,1.0732739,1.3651608,1.6570477,1.9507477,1.7821422,1.6153497,1.4467441,1.2799516,1.1131591,1.6425442,2.1719291,2.7031271,3.2325122,3.7618973,3.1219215,2.4819458,1.84197,1.2019942,0.5620184,4.5324063,8.502794,12.473183,16.441757,20.412146,21.024927,21.637709,22.25049,22.863272,23.47424,19.9444,16.414564,12.884725,9.354887,5.825049,5.484212,5.145188,4.804351,4.465327,4.12449,5.6945157,7.264541,8.834567,10.4045925,11.974618,12.639976,13.305332,13.97069,14.634234,15.299591,15.004078,14.710379,14.4148655,14.119352,13.825653,12.804955,11.784257,10.765372,9.744674,8.725789,8.59163,8.459284,8.326937,8.194591,8.062244,7.891826,7.723221,7.552802,7.382384,7.211965,6.430578,5.6473784,4.8641787,4.082792,3.299592,5.3500524,7.400513,9.449161,11.499621,13.550082,11.544946,9.539809,7.5346723,5.529536,3.5243993,2.819157,2.1157274,1.4104849,0.70524246,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.04169814,0.047137026,0.052575916,0.058014803,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.13053331,0.13415924,0.13959812,0.14503701,0.15047589,0.13053331,0.11059072,0.09064813,0.07070554,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.059827764,0.07070554,0.07977036,0.09064813,0.099712946,0.11240368,0.12509441,0.13778515,0.15047589,0.16316663,0.14503701,0.12690738,0.11059072,0.092461094,0.07433146,0.065266654,0.054388877,0.045324065,0.034446288,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.054388877,0.11059072,0.16497959,0.21936847,0.2755703,0.24293698,0.21030366,0.17767033,0.14503701,0.11240368,0.09064813,0.06707962,0.045324065,0.02175555,0.0,1.3452182,2.6904364,4.0356545,5.3808727,6.7242785,6.0843024,5.4443264,4.804351,4.164375,3.5243993,2.819157,2.1157274,1.4104849,0.70524246,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.08520924,0.11965553,0.15410182,0.19036107,0.22480737,1.214685,2.2045624,3.1944401,4.1843176,5.1741953,8.597069,12.019942,15.442815,18.865688,22.286749,21.023113,19.757666,18.492218,17.22677,15.963136,12.866595,9.771869,6.677141,3.5824142,0.48768693,0.38978696,0.291887,0.19579996,0.09789998,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.9453088,3.8906176,5.8359265,7.7794223,9.724731,7.7866745,5.8504305,3.9123733,1.9743162,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.22480737,1.6226015,3.0203958,4.41819,5.814171,7.211965,5.812358,4.4127507,3.0131438,1.6117238,0.21211663,0.17585737,0.13778515,0.099712946,0.06164073,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,1.3923552,2.659616,3.926877,5.1941376,6.4632115,6.7623506,7.063302,7.362441,7.663393,7.9625316,10.183411,12.402477,14.623356,16.842422,19.063301,16.89681,14.732134,12.567456,10.40278,8.238102,6.5973706,4.95664,3.3177216,1.6769904,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.21030366,0.39522585,0.58014804,0.7650702,0.9499924,2.1592383,3.3702974,4.5795436,5.7906027,6.9998484,7.039734,7.079619,7.119504,7.159389,7.1992745,7.324369,7.4494634,7.574558,7.699652,7.8247466,4.175253,4.307599,4.439945,4.572292,4.704638,4.836984,4.9620786,5.087173,5.2122674,5.337362,5.462456,6.8094873,8.158332,9.5053625,10.852394,12.199425,12.730623,13.260008,13.789393,14.320591,14.849977,14.407614,13.965251,13.522888,13.080525,12.638163,12.5058155,12.371656,12.23931,12.106964,11.974618,12.389787,12.804955,13.220123,13.635292,14.05046,15.056654,16.064661,17.072668,18.080675,19.08687,17.661882,16.236893,14.811904,13.386916,11.961927,20.94153,29.922947,38.90255,47.882156,56.86176,51.549778,46.237797,40.924004,35.612022,30.300043,24.882912,19.465778,14.046834,8.629702,3.2125697,3.1454902,3.0765975,3.009518,2.9424384,2.8753586,2.8771715,2.8807976,2.8826106,2.8844235,2.8880494,2.7919624,2.6976883,2.6016014,2.5073273,2.4130533,1.9453088,1.4775645,1.0098201,0.5420758,0.07433146,0.065266654,0.054388877,0.045324065,0.034446288,0.025381476,0.15772775,0.29007402,0.4224203,0.55476654,0.6871128,1.162109,1.6371052,2.1121013,2.5870976,3.0620937,3.4500678,3.8380418,4.2242026,4.612177,5.0001507,7.2029004,9.40565,11.608399,13.809336,16.012085,15.905121,15.798156,15.689378,15.582414,15.475449,14.590723,13.704185,12.819458,11.934732,11.050007,10.741803,10.435412,10.127209,9.820818,9.512614,8.725789,7.93715,7.1503243,6.3616858,5.57486,5.9392653,6.305484,6.6698895,7.0342946,7.400513,7.422269,7.4458375,7.4675927,7.4893484,7.512917,6.9382076,6.3616858,5.7869763,5.2122674,4.6375585,4.441758,4.2477713,4.0519714,3.8579843,3.6621845,5.612932,7.5618668,9.512614,11.463363,13.412297,11.747997,10.081885,8.417585,6.7532854,5.087173,5.6401267,6.19308,6.7442207,7.2971745,7.850128,7.663393,7.474845,7.28811,7.0995617,6.9128265,6.446895,5.9827766,5.516845,5.0527267,4.5867953,5.034597,5.482399,5.9302006,6.378002,6.825804,7.5256076,8.225411,8.925215,9.625018,10.324821,10.410031,10.49524,10.58045,10.665659,10.750868,11.5775795,12.40429,13.232814,14.059525,14.888049,16.048346,17.206827,18.367125,19.52742,20.687716,19.792112,18.898321,18.002718,17.107115,16.213324,16.900436,17.58755,18.274662,18.961775,19.650702,20.270735,20.890768,21.510801,22.130835,22.750868,22.55688,22.364706,22.172533,21.980358,21.788185,22.203352,22.616709,23.031878,23.447044,23.862213,25.136726,26.413052,27.687565,28.962078,30.238403,29.351864,28.467138,27.582413,26.697687,25.812962,24.581959,23.352772,22.121769,20.89258,19.663393,18.350807,17.038223,15.725637,14.413053,13.100468,12.962683,12.824898,12.687112,12.549327,12.413355,13.800271,15.187187,16.575916,17.962833,19.34975,18.08974,16.829731,15.569723,14.309713,13.049705,11.378153,9.704789,8.033237,6.359873,4.688321,5.8758116,7.063302,8.2507925,9.438283,10.625773,11.769753,12.915545,14.059525,15.2053175,16.349297,15.154554,13.959812,12.76507,11.570327,10.375585,9.345822,8.314246,7.2844834,6.2547207,5.224958,4.902251,4.5795436,4.256836,3.9341288,3.6132345,4.168001,4.7227674,5.277534,5.8323007,6.3870673,7.1902094,7.993352,8.794682,9.597824,10.399154,8.319685,6.240217,4.160749,2.079468,0.0,0.065266654,0.13053331,0.19579996,0.25925365,0.3245203,0.5946517,0.86478317,1.1349145,1.405046,1.6751775,1.5555218,1.4358664,1.3143979,1.1947423,1.0750868,1.5954071,2.1157274,2.6342347,3.1545548,3.6748753,3.0149567,2.3550384,1.69512,1.0352017,0.37528324,4.992899,9.610515,14.22813,18.845747,23.463362,22.212418,20.963285,19.712341,18.463211,17.212267,15.192626,13.172986,11.153346,9.131892,7.112252,6.8403077,6.5683637,6.294606,6.0226617,5.750717,7.217404,8.684091,10.152591,11.619277,13.087777,13.535579,13.98338,14.429369,14.877171,15.324973,14.545399,13.765825,12.984438,12.2048645,11.42529,10.582263,9.739235,8.898021,8.054993,7.211965,7.558241,7.902704,8.247167,8.59163,8.937905,8.745731,8.551744,8.3595705,8.167397,7.9752226,7.1829576,6.390693,5.5966153,4.804351,4.0120864,5.0998635,6.187641,7.2754188,8.363196,9.449161,8.029612,6.6100616,5.1905117,3.7691493,2.3495996,1.8800422,1.4104849,0.93911463,0.46955732,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.032633327,0.03988518,0.047137026,0.054388877,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.13234627,0.13959812,0.14684997,0.15410182,0.16316663,0.14503701,0.12690738,0.11059072,0.092461094,0.07433146,0.07433146,0.07433146,0.07433146,0.07433146,0.07433146,0.09064813,0.10515183,0.11965553,0.13415924,0.15047589,0.16316663,0.17585737,0.18673515,0.19942589,0.21211663,0.19217403,0.17223145,0.15228885,0.13234627,0.11240368,0.09789998,0.08339628,0.06707962,0.052575916,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08339628,0.16497959,0.24837588,0.32995918,0.41335547,0.3444629,0.27738327,0.21030366,0.14322405,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,2.0178273,4.0356545,6.051669,8.069496,10.087324,9.128266,8.167397,7.208339,6.247469,5.2865987,4.229642,3.1726844,2.1157274,1.0569572,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.09064813,0.10515183,0.11965553,0.13415924,0.15047589,1.6733645,3.1944401,4.7173285,6.240217,7.763106,9.302311,10.843329,12.382534,13.92174,15.462758,14.989574,14.518205,14.045021,13.571837,13.100468,10.54419,7.989726,5.4352617,2.8807976,0.3245203,0.25925365,0.19579996,0.13053331,0.065266654,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.7557032,5.5095935,8.265296,11.019187,13.77489,11.024626,8.274362,5.524097,2.7756457,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.15047589,1.6896812,3.2306993,4.7699046,6.3091097,7.850128,6.338117,4.8242936,3.3122826,1.8002719,0.28826106,0.2374981,0.18673515,0.13778515,0.0870222,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,2.0830941,3.97764,5.8721857,7.7667317,9.663091,10.038374,10.411844,10.7871275,11.162411,11.537694,13.667925,15.798156,17.928387,20.056805,22.187037,18.901947,15.616859,12.331772,9.048496,5.763408,4.615803,3.4681973,2.3205922,1.1729867,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.16497959,0.291887,0.42060733,0.5475147,0.6744221,1.6026589,2.5308957,3.4573197,4.3855567,5.3119802,5.67276,6.0317264,6.392506,6.7532854,7.112252,7.175706,7.2373466,7.3008003,7.362441,7.4258947,4.213325,4.4345064,4.6575007,4.880495,5.101677,5.3246713,5.375434,5.424384,5.475147,5.52591,5.57486,6.929143,8.285239,9.639522,10.995618,12.349901,13.064208,13.780329,14.494636,15.210756,15.925063,15.448255,14.969632,14.492823,14.014201,13.537392,13.165734,12.792264,12.420607,12.047136,11.675479,12.157727,12.639976,13.122223,13.604471,14.0867195,15.172684,16.256836,17.3428,18.426952,19.512917,18.024473,16.537846,15.049402,13.562773,12.07433,21.440096,30.804047,40.16981,49.535576,58.89953,53.025528,47.14972,41.27572,35.399906,29.524096,24.135971,18.746033,13.354282,7.9643445,2.5744069,2.810092,3.045777,3.2796493,3.5153344,3.7492065,3.7691493,3.7909048,3.8108473,3.83079,3.8507326,3.6277382,3.4047437,3.1817493,2.960568,2.7375734,2.2100015,1.6824293,1.1548572,0.62728506,0.099712946,0.08339628,0.065266654,0.047137026,0.030820364,0.012690738,0.09789998,0.18310922,0.26831847,0.35171473,0.43692398,1.162109,1.887294,2.612479,3.3376641,4.062849,4.024777,3.9867048,3.9504454,3.9123733,3.874301,6.445082,9.01405,11.584831,14.155612,16.72458,16.815228,16.905876,16.99471,17.08536,17.174194,16.08279,14.989574,13.898171,12.804955,11.711739,10.990179,10.266808,9.545248,8.821876,8.100317,7.474845,6.849373,6.2257137,5.600241,4.974769,5.4570174,5.9392653,6.4233265,6.9055743,7.3878226,7.1050005,6.8221784,6.539356,6.258347,5.975525,5.57486,5.1741953,4.7753434,4.3746786,3.975827,3.7890918,3.6041696,3.4192474,3.2343252,3.049403,5.4497657,7.850128,10.25049,12.650853,15.049402,12.955431,10.859646,8.765674,6.6698895,4.574105,5.145188,5.714458,6.285541,6.8548117,7.4258947,7.250037,7.07418,6.9001355,6.7242785,6.550234,5.866747,5.185073,4.501586,3.8199122,3.1382382,3.7165732,4.2967215,4.876869,5.4570174,6.037165,6.7115874,7.3878226,8.062244,8.736667,9.412902,9.554313,9.697536,9.840761,9.982172,10.125396,11.044568,11.965553,12.884725,13.80571,14.724882,15.818098,16.909502,18.002718,19.094122,20.187338,19.489347,18.79317,18.095179,17.397188,16.699198,17.513218,18.325426,19.137632,19.94984,20.762047,21.385706,22.007553,22.629398,23.253057,23.874905,23.30926,22.745428,22.179785,21.61414,21.050308,21.683033,22.315756,22.946667,23.579391,24.212114,25.287203,26.36229,27.437376,28.512463,29.58755,28.494333,27.40293,26.309713,25.21831,24.125093,22.798004,21.470917,20.142014,18.814926,17.487837,16.124489,14.762955,13.399607,12.038072,10.674724,10.712796,10.750868,10.7871275,10.825199,10.863272,12.050762,13.238253,14.425743,15.613234,16.800724,15.845293,14.889862,13.93443,12.980812,12.025381,10.720048,9.414715,8.109382,6.8058615,5.5005283,6.825804,8.149267,9.474543,10.799818,12.125093,13.4594345,14.795588,16.129929,17.464268,18.800423,16.8533,14.904366,12.957244,11.010121,9.063,8.247167,7.4331465,6.6173134,5.803293,4.98746,4.6828823,4.3783045,4.071914,3.7673361,3.4627585,3.8906176,4.3166637,4.744523,5.1723824,5.600241,6.544795,7.4893484,8.435715,9.380268,10.324821,8.259857,6.1948934,4.1299286,2.0649643,0.0,0.032633327,0.065266654,0.09789998,0.13053331,0.16316663,0.40972954,0.65810543,0.90466833,1.1530442,1.3996071,1.3270886,1.2545701,1.1820517,1.1095331,1.0370146,1.54827,2.0577126,2.5671551,3.0784104,3.587853,2.907992,2.228131,1.54827,0.8665961,0.18673515,5.4533916,10.718235,15.983078,21.247921,26.512764,23.399908,20.287052,17.174194,14.06315,10.950294,10.439038,9.929596,9.420154,8.910711,8.399456,8.194591,7.989726,7.7848616,7.5799966,7.3751316,8.740293,10.1054535,11.470614,12.835775,14.199123,14.429369,14.6596155,14.889862,15.120108,15.350354,14.084907,12.819458,11.555823,10.290376,9.024928,8.3595705,7.6942134,7.0306687,6.3653116,5.6999545,6.5230393,7.344311,8.167397,8.990481,9.811753,9.597824,9.382081,9.168152,8.952409,8.736667,7.935337,7.132195,6.3308654,5.527723,4.7245803,4.8496747,4.974769,5.0998635,5.224958,5.3500524,4.514277,3.680314,2.8445382,2.0105755,1.1747998,0.93911463,0.70524246,0.46955732,0.23568514,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.02175555,0.032633327,0.04169814,0.052575916,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.13415924,0.14503701,0.15410182,0.16497959,0.17585737,0.15954071,0.14503701,0.13053331,0.11421664,0.099712946,0.099712946,0.099712946,0.099712946,0.099712946,0.099712946,0.11965553,0.13959812,0.15954071,0.1794833,0.19942589,0.21211663,0.22480737,0.2374981,0.25018883,0.26287958,0.23931105,0.21755551,0.19579996,0.17223145,0.15047589,0.13053331,0.11059072,0.09064813,0.07070554,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.11059072,0.21936847,0.32995918,0.4405499,0.5493277,0.44780177,0.3444629,0.24293698,0.13959812,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,2.6904364,5.37906,8.069496,10.7599325,13.45037,12.170418,10.890467,9.610515,8.330563,7.0506115,5.6401267,4.229642,2.819157,1.4104849,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.09427405,0.09064813,0.08520924,0.07977036,0.07433146,2.1302311,4.1843176,6.240217,8.294304,10.3502035,10.007553,9.664904,9.322253,8.979604,8.636953,8.957849,9.27693,9.597824,9.916905,10.2378,8.221786,6.207584,4.1915693,2.1773682,0.16316663,0.13053331,0.09789998,0.065266654,0.032633327,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,3.5660975,7.130382,10.694666,14.25895,17.825048,14.262577,10.700105,7.137634,3.5751622,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.07433146,1.7567607,3.43919,5.123432,6.8040485,8.488291,6.8620634,5.237649,3.6132345,1.987007,0.36259252,0.2991388,0.2374981,0.17585737,0.11240368,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,2.7720199,5.295664,7.817495,10.339326,12.862969,13.312584,13.762199,14.211814,14.663241,15.112856,17.15244,19.192022,21.233418,23.273,25.312584,20.907085,16.501585,12.097899,7.6924005,3.2869012,2.6324217,1.9779422,1.3216497,0.6671702,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.11965553,0.19036107,0.25925365,0.32995918,0.40066472,1.0442665,1.6896812,2.335096,2.9805105,3.6241121,4.305786,4.985647,5.6655083,6.345369,7.02523,7.02523,7.02523,7.02523,7.02523,7.02523,4.249584,4.5632267,4.8750563,5.186886,5.5005283,5.812358,5.7869763,5.7615952,5.7380266,5.712645,5.6872635,7.0506115,8.412147,9.775495,11.137029,12.500377,13.399607,14.300649,15.199879,16.100922,17.00015,16.487082,15.975826,15.462758,14.94969,14.436621,13.825653,13.212872,12.60009,11.9873085,11.374527,11.925668,12.474996,13.024323,13.575464,14.124791,15.2869005,16.450823,17.612932,18.77504,19.93715,18.387066,16.836983,15.2869005,13.736817,12.186734,21.936848,31.68696,41.437073,51.187187,60.937298,54.49947,48.06345,41.62562,35.18779,28.74996,23.387217,18.024473,12.661731,7.3008003,1.938057,2.474694,3.0131438,3.5497808,4.0882306,4.6248674,4.6629395,4.699199,4.7372713,4.7753434,4.8116026,4.461701,4.1117992,3.7618973,3.4119956,3.0620937,2.474694,1.887294,1.2998942,0.7124943,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,1.162109,2.137483,3.1128569,4.0882306,5.0617914,4.599486,4.137181,3.6748753,3.2125697,2.7502642,5.6872635,8.624263,11.563075,14.500074,17.437075,17.725336,18.011784,18.300045,18.588305,18.874754,17.57486,16.274965,14.975071,13.675177,12.375282,11.236742,10.100015,8.963287,7.8247466,6.688019,6.2257137,5.763408,5.2992897,4.836984,4.3746786,4.974769,5.57486,6.1749506,6.775041,7.3751316,6.787732,6.200332,5.612932,5.0255322,4.4381323,4.213325,3.9867048,3.7618973,3.53709,3.3122826,3.1382382,2.962381,2.7883365,2.612479,2.4366217,5.2865987,8.136576,10.988366,13.838344,16.68832,14.162864,11.637406,9.11195,6.588306,4.062849,4.650249,5.237649,5.825049,6.412449,6.9998484,6.836682,6.6753283,6.5121617,6.350808,6.187641,5.2884116,4.3873696,3.48814,2.5870976,1.6878681,2.4003625,3.1128569,3.825351,4.537845,5.2503395,5.89938,6.550234,7.1992745,7.850128,8.499168,8.700407,8.899834,9.099259,9.300498,9.499924,10.51337,11.525003,12.536636,13.550082,14.561715,15.5878525,16.612177,17.638313,18.662638,19.68696,19.188396,18.688019,18.187641,17.687263,17.186886,18.124187,19.063301,20.000603,20.937904,21.875206,22.500679,23.124338,23.74981,24.375282,25.000753,24.06164,23.124338,22.187037,21.249735,20.312433,21.162712,22.01299,22.863272,23.711737,24.562017,25.437677,26.31334,27.187187,28.062847,28.936695,27.6368,26.336908,25.037014,23.73712,22.437225,21.012236,19.587248,18.16226,16.73727,15.312282,13.899984,12.487686,11.075388,9.663091,8.2507925,8.46291,8.675026,8.887142,9.099259,9.313189,10.29944,11.287505,12.27557,13.261822,14.249886,13.600845,12.949992,12.299138,11.650098,10.999244,10.061942,9.12464,8.187339,7.250037,6.3127356,7.7757964,9.237044,10.700105,12.163166,13.6244135,15.149116,16.67563,18.20033,19.725033,21.249735,18.550234,15.850732,13.149418,10.449916,7.750415,7.1503243,6.550234,5.9501433,5.3500524,4.749962,4.461701,4.175253,3.8869917,3.6005437,3.3122826,3.6132345,3.9123733,4.213325,4.512464,4.8116026,5.89938,6.987158,8.074935,9.162713,10.25049,8.200029,6.149569,4.099108,2.0504606,0.0,0.0,0.0,0.0,0.0,0.0,0.22480737,0.44961473,0.6744221,0.89922947,1.1258497,1.1004683,1.0750868,1.0497054,1.0243238,1.0007553,1.49932,1.9996977,2.5000753,3.000453,3.5008307,2.7992141,2.0994108,1.3996071,0.69980353,0.0,5.9120708,11.8241415,17.738026,23.650097,29.562168,24.587399,19.612629,14.63786,9.663091,4.688321,5.6872635,6.688019,7.686961,8.6877165,9.686659,9.550687,9.412902,9.275117,9.137331,8.999546,10.263181,11.525003,12.786825,14.05046,15.312282,15.324973,15.337664,15.350354,15.363045,15.375735,13.6244135,11.874905,10.125396,8.374074,6.624565,6.1368785,5.6491914,5.163317,4.6756306,4.1879435,5.487838,6.787732,8.087626,9.38752,10.687414,10.449916,10.212419,9.97492,9.737422,9.499924,8.6877165,7.8755093,7.063302,6.249282,5.4370747,4.599486,3.7618973,2.9243085,2.08672,1.2491312,1.0007553,0.7505665,0.50037766,0.25018883,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.13778515,0.15047589,0.16316663,0.17585737,0.18673515,0.17585737,0.16316663,0.15047589,0.13778515,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.15047589,0.17585737,0.19942589,0.22480737,0.25018883,0.26287958,0.2755703,0.28826106,0.2991388,0.31182957,0.28826106,0.26287958,0.2374981,0.21211663,0.18673515,0.16316663,0.13778515,0.11240368,0.0870222,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13778515,0.2755703,0.41335547,0.5493277,0.6871128,0.5493277,0.41335547,0.2755703,0.13778515,0.0,0.0,0.0,0.0,0.0,0.0,3.3630457,6.7242785,10.087324,13.45037,16.811602,15.212569,13.611723,12.012691,10.411844,8.812811,7.0506115,5.2884116,3.5243993,1.7621996,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,2.5870976,5.1741953,7.763106,10.3502035,12.937301,10.712796,8.488291,6.261973,4.0374675,1.8129625,2.9243085,4.0374675,5.1506267,6.261973,7.3751316,5.89938,4.4254417,2.94969,1.4757515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,4.3746786,8.749357,13.125849,17.500528,21.875206,17.500528,13.125849,8.749357,4.3746786,0.0,0.0,0.0,0.0,0.0,0.0,1.8256533,3.6494937,5.475147,7.2989874,9.12464,7.3878226,5.6491914,3.9123733,2.175555,0.43692398,0.36259252,0.28826106,0.21211663,0.13778515,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.06164073,0.12509441,0.18673515,0.25018883,0.31182957,3.4627585,6.6118746,9.762803,12.91192,16.062849,16.586794,17.112555,17.638313,18.16226,18.688019,20.636953,22.5877,24.538448,26.487383,28.438131,22.912222,17.38631,11.862214,6.338117,0.8122072,0.6508536,0.48768693,0.3245203,0.16316663,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.48768693,0.85027945,1.2128719,1.5754645,1.938057,2.9369993,3.9377546,4.936697,5.9374523,6.9382076,6.874754,6.813113,6.7496595,6.688019,6.624565,3.9867048,4.36924,4.751775,5.1343102,5.516845,5.89938,5.8903155,5.8794374,5.870373,5.859495,5.8504305,7.3424983,8.834567,10.328448,11.820516,13.312584,14.150173,14.9877615,15.825351,16.66294,17.500528,17.143373,16.784407,16.427254,16.0701,15.712947,14.762955,13.812962,12.862969,11.912977,10.962985,11.514126,12.067079,12.620032,13.172986,13.724127,14.4148655,15.105604,15.79453,16.48527,17.174194,17.007402,16.840609,16.672005,16.50521,16.338419,25.062395,33.78637,42.51216,51.23795,59.961926,52.933067,45.9024,38.87173,31.842875,24.812206,20.450218,16.08823,11.724429,7.362441,3.000453,3.1708715,3.339477,3.5098956,3.680314,3.8507326,3.9431937,4.0356545,4.1281157,4.220577,4.313038,3.9450066,3.576975,3.2107568,2.8427253,2.474694,1.9996977,1.5247015,1.0497054,0.5747091,0.099712946,0.17585737,0.25018883,0.3245203,0.40066472,0.4749962,0.40972954,0.3444629,0.27919623,0.21574254,0.15047589,0.9445535,1.7404441,2.5345216,3.3304121,4.12449,3.7528327,3.3793623,3.007705,2.6342347,2.2625773,5.573047,8.881703,12.192173,15.502643,18.813112,20.258043,21.702974,23.147905,24.592838,26.03777,23.684544,21.33313,18.979906,16.62668,14.275268,13.035201,11.795135,10.555068,9.3150015,8.074935,7.6706448,7.264541,6.8602505,6.454147,6.049856,6.506723,6.965402,7.422269,7.8791356,8.337815,7.5818095,6.827617,6.071612,5.317419,4.5632267,4.2876563,4.0120864,3.738329,3.4627585,3.1871881,3.3358512,3.482701,3.6295512,3.778214,3.925064,6.298232,8.669587,11.042755,13.415923,15.787278,13.470312,11.153346,8.834567,6.5176005,4.2006345,4.9221935,5.6455655,6.3671246,7.0904965,7.8120556,7.4857225,7.157576,6.82943,6.5030966,6.1749506,5.3119802,4.4508233,3.587853,2.7248828,1.8619126,2.4003625,2.9369993,3.4754493,4.0120864,4.550536,5.2521524,5.955582,6.6571984,7.360628,8.062244,8.238102,8.412147,8.588004,8.762048,8.937905,9.762803,10.587702,11.4126,12.237497,13.062395,14.122978,15.181748,16.242332,17.302916,18.361685,18.220274,18.07705,17.935638,17.792416,17.64919,18.57924,19.50929,20.43934,21.36939,22.29944,22.66022,23.019186,23.379965,23.740746,24.099712,23.347332,22.594954,21.842573,21.090193,20.337814,21.07569,21.811752,22.54963,23.287504,24.025381,24.560204,25.095028,25.629852,26.164677,26.6995,25.374224,24.050762,22.725487,21.40021,20.074934,18.869314,17.665508,16.459887,15.254267,14.05046,12.888351,11.724429,10.56232,9.400211,8.238102,8.42665,8.617011,8.807372,8.997733,9.188094,10.375585,11.563075,12.750566,13.938056,15.125546,14.692248,14.260764,13.827466,13.394168,12.962683,12.010877,11.057259,10.1054535,9.151835,8.200029,9.304124,10.410031,11.515939,12.620032,13.724127,15.161806,16.599485,18.037165,19.474844,20.912523,18.142317,15.372109,12.601903,9.8316965,7.063302,6.5756154,6.0879283,5.600241,5.1125546,4.6248674,4.229642,3.834416,3.43919,3.045777,2.6505513,3.2143826,3.780027,4.345671,4.9095025,5.475147,6.294606,7.115878,7.935337,8.754796,9.574255,7.8646317,6.155008,4.445384,2.7357605,1.0243238,0.8901646,0.7541924,0.6200332,0.48587397,0.34990177,0.5293851,0.7106813,0.8901646,1.0696479,1.2491312,1.214685,1.1802386,1.1457924,1.1095331,1.0750868,1.4775645,1.8800422,2.2825198,2.6849976,3.0874753,2.715818,2.3423476,1.9706904,1.5972201,1.2255627,5.7960415,10.364707,14.935185,19.505665,24.07433,20.13295,16.189756,12.246562,8.3051815,4.361988,5.219519,6.0770507,6.9345818,7.7921133,8.649645,8.7693,8.890768,9.010424,9.130079,9.249735,10.306692,11.365462,12.42242,13.479377,14.538147,14.501887,14.467442,14.432995,14.396736,14.362289,12.670795,10.9774885,9.284182,7.592687,5.89938,5.732588,5.565795,5.3971896,5.230397,5.0617914,5.9483304,6.833056,7.7177815,8.602508,9.487233,9.316814,9.14821,8.977791,8.807372,8.636953,8.049554,7.462154,6.874754,6.2873545,5.6999545,4.9095025,4.120864,3.3304121,2.5399606,1.7495089,1.3996071,1.0497054,0.69980353,0.34990177,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12328146,0.13234627,0.14322405,0.15228885,0.16316663,0.16497959,0.16679256,0.17041849,0.17223145,0.17585737,0.15954071,0.14503701,0.13053331,0.11421664,0.099712946,0.14503701,0.19036107,0.23568514,0.27919623,0.3245203,0.40247768,0.48043507,0.55839247,0.6345369,0.7124943,0.7850128,0.8575313,0.9300498,1.0025684,1.0750868,1.0696479,1.064209,1.0605831,1.0551442,1.0497054,0.94274056,0.83577573,0.726998,0.6200332,0.51306844,0.41335547,0.31182957,0.21211663,0.11240368,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.018129626,0.02175555,0.027194439,0.032633327,0.038072214,0.045324065,0.052575916,0.059827764,0.06707962,0.07433146,0.17041849,0.26469254,0.36077955,0.4550536,0.5493277,0.5076295,0.46411842,0.4224203,0.38072214,0.33721104,0.2755703,0.21211663,0.15047589,0.0870222,0.025381476,4.1426196,8.259857,12.377095,16.494333,20.613384,17.89938,15.187187,12.474996,9.762803,7.0506115,5.7470913,4.445384,3.141864,1.840157,0.53663695,0.44961473,0.36259252,0.2755703,0.18673515,0.099712946,0.09789998,0.09427405,0.092461094,0.09064813,0.0870222,2.913431,5.7380266,8.562622,11.3872175,14.211814,11.999999,9.788185,7.574558,5.3627434,3.149116,3.8996825,4.650249,5.4008155,6.149569,6.9001355,5.520471,4.1408067,2.759329,1.3796645,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,3.6222992,7.2445984,10.866898,14.489197,18.11331,14.489197,10.866898,7.2445984,3.6222992,0.0,0.0,0.0,0.0,0.0,0.0,1.7495089,3.5008307,5.2503395,6.9998484,8.749357,7.400513,6.049856,4.699199,3.350355,1.9996977,1.6117238,1.2255627,0.8375887,0.44961473,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.11059072,0.21936847,0.32995918,0.4405499,0.5493277,3.3304121,6.109684,8.890768,11.67004,14.449312,14.911617,15.375735,15.838041,16.300346,16.762651,18.07705,19.393261,20.707659,22.022057,23.338266,18.800423,14.262577,9.724731,5.186886,0.6508536,0.52032024,0.38978696,0.25925365,0.13053331,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.12690738,0.20486477,0.28282216,0.36077955,0.43692398,1.0333886,1.6280404,2.222692,2.817344,3.4119956,3.8416677,4.273153,4.702825,5.132497,5.562169,5.661882,5.763408,5.863121,5.962834,6.0625467,3.7256382,4.177066,4.6303062,5.081734,5.5349746,5.9882154,5.9918413,5.99728,6.002719,6.008158,6.011784,7.6343856,9.256987,10.879588,12.50219,14.124791,14.90074,15.674874,16.450823,17.224958,18.000906,17.797853,17.5948,17.39175,17.190512,16.98746,15.700256,14.413053,13.125849,11.836833,10.549629,11.104396,11.6591625,12.215742,12.770509,13.325275,13.54283,13.760386,13.9779415,14.195497,14.413053,15.627737,16.842422,18.057108,19.271791,20.48829,28.187943,35.887596,43.587246,51.2869,58.988365,51.364857,43.74316,36.11965,28.49796,20.87445,17.513218,14.150173,10.7871275,7.424082,4.062849,3.8652363,3.6676233,3.4700103,3.2723975,3.0747845,3.2216346,3.3702974,3.5171473,3.6658103,3.8126602,3.4283123,3.0421512,2.657803,2.2716422,1.887294,1.5247015,1.162109,0.7995165,0.43692398,0.07433146,0.25018883,0.42423326,0.6000906,0.774135,0.9499924,0.78319985,0.61459434,0.44780177,0.27919623,0.11240368,0.726998,1.3415923,1.9579996,2.572594,3.1871881,2.904366,2.6233568,2.3405347,2.0577126,1.7748904,5.4570174,9.139144,12.823084,16.50521,20.187338,22.790752,25.392353,27.995768,30.59737,33.200783,29.794228,26.389482,22.98474,19.579996,16.175253,14.831847,13.490254,12.14685,10.805257,9.461852,9.115576,8.767487,8.419398,8.073122,7.7250338,8.040489,8.354132,8.669587,8.985043,9.300498,8.3777,7.454902,6.532104,5.6093063,4.688321,4.361988,4.0374675,3.7129474,3.386614,3.0620937,3.531651,4.0030212,4.4725785,4.942136,5.411693,7.308052,9.202598,11.097144,12.99169,14.888049,12.7777605,10.667472,8.557183,6.446895,4.3366065,5.1941376,6.051669,6.9092,7.7667317,8.624263,8.13295,7.6398244,7.1466985,6.6553855,6.16226,5.337362,4.512464,3.6875658,2.8626678,2.03777,2.4003625,2.762955,3.1255474,3.48814,3.8507326,4.604925,5.3591175,6.115123,6.869315,7.6253204,7.7757964,7.9244595,8.074935,8.225411,8.375887,9.012237,9.6504,10.28675,10.924912,11.563075,12.658105,13.753134,14.848164,15.9431925,17.038223,17.252151,17.467894,17.681824,17.897566,18.11331,19.034294,19.957092,20.87989,21.802689,22.725487,22.81976,22.915848,23.01012,23.104395,23.200481,22.633024,22.065567,21.49811,20.930653,20.363195,20.986855,21.612328,22.237799,22.863272,23.48693,23.68273,23.876717,24.072517,24.268316,24.462305,23.111647,21.762802,20.412146,19.063301,17.712645,16.728207,15.741954,14.757515,13.773077,12.786825,11.874905,10.962985,10.049252,9.137331,8.225411,8.392203,8.560809,8.727602,8.894395,9.063,10.449916,11.836833,13.225562,14.612478,15.999394,15.785465,15.569723,15.355793,15.140051,14.924308,13.957999,12.989877,12.021755,11.055446,10.087324,10.834265,11.583018,12.329959,13.0769,13.825653,15.174497,16.525154,17.87581,19.224655,20.575312,17.7344,14.895301,12.054388,9.215289,6.3743763,6.000906,5.6256227,5.2503395,4.8750563,4.499773,3.9975824,3.4953918,2.9932013,2.4891977,1.987007,2.817344,3.6476808,4.478018,5.3083544,6.1368785,6.6898317,7.2427855,7.795739,8.34688,8.899834,7.5292335,6.1604466,4.7898474,3.4192474,2.0504606,1.7803292,1.5101979,1.2400664,0.969935,0.69980353,0.83577573,0.969935,1.1059072,1.2400664,1.3742256,1.3307146,1.2853905,1.2400664,1.1947423,1.1494182,1.455809,1.7603867,2.0649643,2.3695421,2.6741197,2.6306088,2.5852847,2.5399606,2.4946365,2.4493124,5.678199,8.9052725,12.132345,15.359419,18.588305,15.676687,12.766883,9.857078,6.947273,4.0374675,4.751775,5.467895,6.1822023,6.8983226,7.61263,7.989726,8.366822,8.745731,9.122828,9.499924,10.352016,11.204109,12.058014,12.910107,13.762199,13.680615,13.597219,13.515636,13.43224,13.3506565,11.715364,10.080072,8.444779,6.8094873,5.1741953,5.328297,5.480586,5.632875,5.7851634,5.9374523,6.4070096,6.87838,7.3479376,7.817495,8.287052,8.185526,8.082188,7.9806614,7.877322,7.7757964,7.413204,7.0506115,6.688019,6.3254266,5.962834,5.219519,4.478018,3.7347028,2.9932013,2.2498865,1.8002719,1.3506571,0.89922947,0.44961473,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.05076295,0.06164073,0.07433146,0.0870222,0.099712946,0.10696479,0.11421664,0.12328146,0.13053331,0.13778515,0.15410182,0.17223145,0.19036107,0.20667773,0.22480737,0.19579996,0.16497959,0.13415924,0.10515183,0.07433146,0.13959812,0.20486477,0.27013144,0.33539808,0.40066472,0.5420758,0.6852999,0.82671094,0.969935,1.1131591,1.2817645,1.452183,1.6226015,1.79302,1.9616255,1.9779422,1.9924458,2.0069497,2.0232663,2.03777,1.8347181,1.6316663,1.4304274,1.2273756,1.0243238,0.824898,0.62547207,0.42423326,0.22480737,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.034446288,0.045324065,0.054388877,0.065266654,0.07433146,0.09064813,0.10515183,0.11965553,0.13415924,0.15047589,0.2030518,0.25562772,0.30820364,0.36077955,0.41335547,0.46411842,0.5166943,0.56927025,0.62184614,0.6744221,0.5493277,0.42423326,0.2991388,0.17585737,0.05076295,4.9221935,9.795437,14.666867,19.540112,24.413355,20.588003,16.762651,12.937301,9.11195,5.2865987,4.445384,3.6023567,2.759329,1.9181144,1.0750868,0.87566096,0.6744221,0.4749962,0.2755703,0.07433146,0.09427405,0.11421664,0.13415924,0.15410182,0.17585737,3.2379513,6.300045,9.362139,12.4242325,15.488139,13.287203,11.088079,8.887142,6.688019,4.4870825,4.8750563,5.2630305,5.6491914,6.037165,6.4251394,5.139749,3.8543584,2.570781,1.2853905,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.8699198,5.7398396,8.609759,11.479679,14.349599,11.479679,8.609759,5.7398396,2.8699198,0.0,0.0,0.0,0.0,0.0,0.0,1.6751775,3.350355,5.0255322,6.70071,8.375887,7.413204,6.450521,5.487838,4.5251546,3.5624714,2.8626678,2.1628644,1.4630609,0.76325727,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.15772775,0.3154555,0.47318324,0.629098,0.7868258,3.198066,5.6074934,8.01692,10.428161,12.837588,13.238253,13.637105,14.037769,14.436621,14.837286,15.517147,16.197008,16.87687,17.55673,18.236591,14.68681,11.137029,7.5872483,4.0374675,0.48768693,0.38978696,0.291887,0.19579996,0.09789998,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.1794833,0.32270733,0.46411842,0.6073425,0.7505665,1.5772774,2.4058013,3.2325122,4.059223,4.8877473,4.748149,4.606738,4.4671397,4.327542,4.1879435,4.4508233,4.7118897,4.974769,5.237649,5.5005283,3.4627585,3.9848917,4.507025,5.029158,5.5531044,6.0752378,6.09518,6.115123,6.1350656,6.155008,6.1749506,7.9280853,9.679407,11.432542,13.185677,14.936998,15.649493,16.361988,17.074482,17.786976,18.49947,18.452333,18.405195,18.358059,18.309109,18.261972,16.637558,15.013144,13.386916,11.762501,10.138086,10.694666,11.253058,11.809638,12.368031,12.92461,12.670795,12.415168,12.15954,11.9057255,11.650098,14.248073,16.844234,19.442211,22.040186,24.63816,31.311676,37.987003,44.662334,51.33766,58.01299,49.79846,41.58211,33.367577,25.153044,16.936697,14.574407,12.212116,9.849826,7.4875355,5.125245,4.559601,3.9957695,3.4301252,2.864481,2.3006494,2.5018883,2.70494,2.907992,3.1092308,3.3122826,2.909805,2.5073273,2.1048496,1.7023718,1.2998942,1.0497054,0.7995165,0.5493277,0.2991388,0.05076295,0.3245203,0.6000906,0.87566096,1.1494182,1.4249886,1.1548572,0.88472575,0.61459434,0.3444629,0.07433146,0.5094425,0.9445535,1.3796645,1.8147756,2.2498865,2.0577126,1.8655385,1.6733645,1.4793775,1.2872034,5.3428006,9.396585,13.452183,17.50778,21.563377,25.321648,29.081734,32.841816,36.601902,40.361984,35.905724,31.447649,26.989574,22.533312,18.075237,16.630306,15.185374,13.740443,12.295512,10.850581,10.560507,10.270433,9.980359,9.690285,9.400211,9.572442,9.744674,9.916905,10.089137,10.263181,9.171778,8.082188,6.9925966,5.903006,4.8116026,4.4381323,4.062849,3.6875658,3.3122826,2.9369993,3.729264,4.5233417,5.315606,6.107871,6.9001355,8.317872,9.735609,11.153346,12.569269,13.987006,12.085209,10.183411,8.2798,6.378002,4.4743915,5.467895,6.4595857,7.453089,8.444779,9.438283,8.780178,8.122072,7.46578,6.8076744,6.149569,5.3627434,4.5759177,3.787279,3.000453,2.2118144,2.4003625,2.5870976,2.7756457,2.962381,3.149116,3.9576974,4.764466,5.573047,6.379815,7.1883965,7.311678,7.4367723,7.5618668,7.686961,7.8120556,8.26167,8.713099,9.162713,9.612328,10.061942,11.193231,12.322706,13.452183,14.581658,15.712947,16.285843,16.856926,17.429823,18.002718,18.575615,19.489347,20.404894,21.32044,22.234173,23.14972,22.979301,22.810696,22.640276,22.469858,22.29944,21.916904,21.53437,21.151834,20.769299,20.386765,20.899832,21.4129,21.924156,22.437225,22.950293,22.805256,22.66022,22.515182,22.370146,22.22511,20.850883,19.474844,18.100618,16.72458,15.350354,14.585284,13.820213,13.055143,12.290073,11.525003,10.863272,10.199727,9.537996,8.874452,8.212721,8.357758,8.502794,8.647832,8.792869,8.937905,10.524248,12.112403,13.700559,15.2869005,16.875055,16.87687,16.880495,16.882307,16.88412,16.887747,15.905121,14.922495,13.939869,12.957244,11.974618,12.364405,12.754191,13.145792,13.535579,13.925365,15.187187,16.450823,17.712645,18.974466,20.238102,17.328297,14.418491,11.506873,8.597069,5.6872635,5.424384,5.163317,4.900438,4.6375585,4.3746786,3.7655232,3.1545548,2.5453994,1.9344311,1.3252757,2.420305,3.5153344,4.610364,5.7053933,6.8004227,7.0850577,7.369693,7.654328,7.9407763,8.225411,7.1956487,6.165886,5.1343102,4.1045475,3.0747845,2.6704938,2.2643902,1.8600996,1.455809,1.0497054,1.1403534,1.2291887,1.3198367,1.4104849,1.49932,1.4449311,1.3905423,1.3343405,1.2799516,1.2255627,1.4322405,1.6407311,1.8474089,2.0558996,2.2625773,2.5453994,2.8282216,3.1092308,3.392053,3.6748753,5.560356,7.4458375,9.329506,11.214987,13.100468,11.222239,9.345822,7.4675927,5.5893636,3.7129474,4.2858434,4.856927,5.429823,6.002719,6.5756154,7.210152,7.844689,8.479226,9.115576,9.750113,10.397341,11.044568,11.691795,12.340837,12.988064,12.857531,12.726997,12.598277,12.467744,12.337211,10.7599325,9.182655,7.605378,6.0281005,4.4508233,4.9221935,5.3953767,5.866747,6.33993,6.813113,6.867502,6.921891,6.978093,7.0324817,7.0868707,7.0524244,7.017978,6.981719,6.947273,6.9128265,6.775041,6.637256,6.4994707,6.3616858,6.2257137,5.529536,4.835171,4.1408067,3.444629,2.7502642,2.1991236,1.649796,1.1004683,0.5493277,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.038072214,0.05076295,0.06164073,0.07433146,0.0870222,0.092461094,0.09789998,0.10333887,0.10696479,0.11240368,0.14503701,0.17767033,0.21030366,0.24293698,0.2755703,0.23024625,0.18492219,0.13959812,0.09427405,0.05076295,0.13415924,0.21936847,0.3045777,0.38978696,0.4749962,0.68167394,0.8901646,1.0968424,1.305333,1.5120108,1.7803292,2.0468347,2.3151531,2.5816586,2.8499773,2.8844235,2.9206827,2.955129,2.9895754,3.0258346,2.7266958,2.42937,2.132044,1.8347181,1.5373923,1.2382535,0.93730164,0.63816285,0.33721104,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.052575916,0.06707962,0.08339628,0.09789998,0.11240368,0.13415924,0.15772775,0.1794833,0.2030518,0.22480737,0.23568514,0.24474995,0.25562772,0.26469254,0.2755703,0.4224203,0.56927025,0.7179332,0.86478317,1.0116332,0.824898,0.63816285,0.44961473,0.26287958,0.07433146,5.7035804,11.329204,16.958452,22.585888,28.213324,23.274813,18.338116,13.399607,8.46291,3.5243993,3.141864,2.759329,2.3767939,1.9942589,1.6117238,1.2998942,0.9880646,0.6744221,0.36259252,0.05076295,0.092461094,0.13415924,0.17767033,0.21936847,0.26287958,3.5624714,6.8620634,10.163468,13.46306,16.762651,14.574407,12.387974,10.199727,8.013294,5.825049,5.8504305,5.8758116,5.89938,5.924762,5.9501433,4.759027,3.5697234,2.38042,1.1893034,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.1175404,4.2350807,6.352621,8.470161,10.587702,8.470161,6.352621,4.2350807,2.1175404,0.0,0.0,0.0,0.0,0.0,0.0,1.6008459,3.199879,4.800725,6.399758,8.000604,7.424082,6.849373,6.2746634,5.6999545,5.125245,4.1117992,3.100166,2.08672,1.0750868,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.20486477,0.40972954,0.61459434,0.8194591,1.0243238,3.0657198,5.105303,7.1448855,9.184468,11.225864,11.563075,11.900287,12.237497,12.574709,12.91192,12.957244,13.002567,13.047892,13.093216,13.136727,10.57501,8.011481,5.4497657,2.8880494,0.3245203,0.25925365,0.19579996,0.13053331,0.065266654,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.23205921,0.4405499,0.64722764,0.8557183,1.062396,2.1229792,3.1817493,4.2423325,5.3029156,6.3616858,5.6528172,4.942136,4.233268,3.5225863,2.811905,3.2379513,3.6621845,4.0882306,4.512464,4.936697,3.199879,3.7927177,4.3855567,4.9783955,5.569421,6.16226,6.1967063,6.2329655,6.2674117,6.301858,6.338117,8.219973,10.101828,11.985496,13.867351,15.749206,16.400059,17.0491,17.699953,18.350807,18.999847,19.106813,19.21559,19.322556,19.42952,19.538298,17.57486,15.613234,13.649796,11.6881695,9.724731,10.284937,10.845142,11.405348,11.965553,12.525759,11.7969475,11.069949,10.342952,9.6141405,8.887142,12.866595,16.84786,20.827314,24.806767,28.788033,34.437225,40.08823,45.73742,51.388424,57.037617,48.230244,39.42287,30.6155,21.808126,13.000754,11.637406,10.275872,8.912524,7.549176,6.187641,5.2557783,4.322103,3.39024,2.4583774,1.5247015,1.7821422,2.039583,2.2970235,2.5544643,2.811905,2.3931105,1.9725033,1.551896,1.1331016,0.7124943,0.5747091,0.43692398,0.2991388,0.16316663,0.025381476,0.40066472,0.774135,1.1494182,1.5247015,1.8999848,1.5283275,1.1548572,0.78319985,0.40972954,0.038072214,0.291887,0.5475147,0.8031424,1.0569572,1.3125849,1.209246,1.1077201,1.0043813,0.90285534,0.7995165,5.2267714,9.654026,14.083094,18.510347,22.937603,27.854357,32.772926,37.68968,42.608246,47.525,42.015408,36.505814,30.994408,25.484816,19.975222,18.426952,16.880495,15.332225,13.785768,12.237497,12.005438,11.773379,11.539507,11.307447,11.075388,11.104396,11.135216,11.164224,11.195044,11.225864,9.967669,8.709473,7.453089,6.1948934,4.936697,4.512464,4.0882306,3.6621845,3.2379513,2.811905,3.926877,5.041849,6.156821,7.271793,8.386765,9.327692,10.266808,11.207735,12.14685,13.087777,11.392657,9.697536,8.002417,6.3072968,4.612177,5.7398396,6.867502,7.995165,9.122828,10.25049,9.427405,8.604321,7.783048,6.9599633,6.1368785,5.388125,4.6375585,3.8869917,3.1382382,2.3876717,2.4003625,2.4130533,2.4257438,2.4366217,2.4493124,3.3104696,4.169814,5.029158,5.8903155,6.7496595,6.849373,6.9490857,7.0506115,7.1503243,7.250037,7.512917,7.7757964,8.036863,8.299743,8.562622,9.728357,10.89228,12.058014,13.221936,14.387671,15.31772,16.24777,17.17782,18.10787,19.03792,19.9444,20.852695,21.759176,22.66747,23.575766,23.140654,22.705544,22.270432,21.835321,21.40021,21.202597,21.004984,20.807371,20.609758,20.412146,20.81281,21.211662,21.612328,22.01299,22.411844,21.927782,21.441908,20.957848,20.471973,19.987913,18.588305,17.186886,15.787278,14.387671,12.988064,12.442362,11.896661,11.352772,10.80707,10.263181,9.849826,9.438283,9.024928,8.613385,8.200029,8.323311,8.444779,8.568061,8.689529,8.812811,10.600392,12.387974,14.175554,15.963136,17.750717,17.970085,18.189453,18.410635,18.630003,18.849373,17.852243,16.855114,15.857984,14.860854,13.861912,13.894546,13.927178,13.959812,13.992445,14.025079,15.199879,16.374678,17.549479,18.724277,19.90089,16.92038,13.939869,10.959359,7.9806614,5.0001507,4.8496747,4.699199,4.550536,4.40006,4.249584,3.531651,2.8155308,2.0975976,1.3796645,0.66173136,2.0232663,3.3829882,4.74271,6.1024323,7.462154,7.4802837,7.4966,7.51473,7.5328593,7.549176,6.8602505,6.169512,5.480586,4.7898474,4.100921,3.5606585,3.0203958,2.4801328,1.93987,1.3996071,1.4449311,1.4902552,1.5355793,1.5809034,1.6244144,1.5591478,1.4956942,1.4304274,1.3651608,1.2998942,1.4104849,1.5192627,1.6298534,1.7404441,1.8492218,2.4601903,3.0693457,3.680314,4.2894692,4.900438,5.4425135,5.9845896,6.526665,7.0705543,7.61263,6.7677894,5.922949,5.0781083,4.233268,3.386614,3.8180993,4.2477713,4.6774435,5.1071157,5.5367875,6.430578,7.322556,8.214534,9.108324,10.000301,10.442664,10.885027,11.327391,11.769753,12.212116,12.034446,11.856775,11.679105,11.503247,11.325577,9.804502,8.285239,6.7641635,5.2449007,3.7256382,4.517903,5.3101673,6.1024323,6.8946967,7.686961,7.327995,6.967215,6.6082487,6.247469,5.8866897,5.919323,5.9519563,5.9845896,6.017223,6.049856,6.1368785,6.2257137,6.3127356,6.399758,6.48678,5.8395524,5.1923246,4.5450974,3.8978696,3.2506418,2.5997884,1.9507477,1.2998942,0.6508536,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.07433146,0.07795739,0.07977036,0.08339628,0.08520924,0.0870222,0.13415924,0.18310922,0.23024625,0.27738327,0.3245203,0.26469254,0.20486477,0.14503701,0.08520924,0.025381476,0.13053331,0.23568514,0.34083697,0.44417584,0.5493277,0.823085,1.0950294,1.3669738,1.6407311,1.9126755,2.277081,2.6432993,3.007705,3.3721104,3.738329,3.7927177,3.8471067,3.9033084,3.9576974,4.0120864,3.6204863,3.2270734,2.8354735,2.4420607,2.0504606,1.649796,1.2491312,0.85027945,0.44961473,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.07070554,0.09064813,0.11059072,0.13053331,0.15047589,0.1794833,0.21030366,0.23931105,0.27013144,0.2991388,0.26831847,0.23568514,0.2030518,0.17041849,0.13778515,0.38072214,0.62184614,0.86478317,1.1077201,1.3506571,1.1004683,0.85027945,0.6000906,0.34990177,0.099712946,6.4831543,12.864782,19.248224,25.629852,32.013294,25.961624,19.913582,13.861912,7.8120556,1.7621996,1.840157,1.9181144,1.9942589,2.0722163,2.1501737,1.7241274,1.2998942,0.87566096,0.44961473,0.025381476,0.09064813,0.15410182,0.21936847,0.28463513,0.34990177,3.8869917,7.424082,10.962985,14.500074,18.037165,15.861609,13.687867,11.512312,9.336758,7.1630154,6.825804,6.48678,6.149569,5.812358,5.475147,4.3801174,3.2850883,2.1900587,1.0950294,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.3651608,2.7303216,4.0954823,5.4606433,6.825804,5.4606433,4.0954823,2.7303216,1.3651608,0.0,0.0,0.0,0.0,0.0,0.0,1.5247015,3.049403,4.5759177,6.1006193,7.6253204,7.4367723,7.250037,7.063302,6.874754,6.688019,5.3627434,4.0374675,2.712192,1.3869164,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.2520018,0.5058166,0.75781834,1.0098201,1.261822,2.9333735,4.603112,6.2728505,7.9425893,9.612328,9.8878975,10.161655,10.437225,10.712796,10.988366,10.397341,9.808127,9.217102,8.627889,8.036863,6.4632115,4.8877473,3.3122826,1.7368182,0.16316663,0.13053331,0.09789998,0.065266654,0.032633327,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.28463513,0.55839247,0.83033687,1.1022812,1.3742256,2.666868,3.9595103,5.2521524,6.544795,7.837437,6.5574856,5.277534,3.9975824,2.7176309,1.4376793,2.0250793,2.612479,3.199879,3.787279,4.3746786,2.9369993,3.6005437,4.262275,4.9258194,5.5875506,6.249282,6.300045,6.350808,6.399758,6.450521,6.4994707,8.511859,10.524248,12.538449,14.5508375,16.563227,17.150625,17.738026,18.325426,18.912827,19.500225,19.763105,20.024172,20.287052,20.54993,20.81281,18.512161,16.213324,13.912675,11.612025,9.313189,9.875207,10.437225,10.999244,11.563075,12.125093,10.924912,9.724731,8.52455,7.324369,6.1241875,11.486931,16.849674,22.212418,27.575161,32.937904,37.56277,42.18764,46.812508,51.437374,56.06224,46.66203,37.263634,27.861609,18.463211,9.063,8.700407,8.337815,7.9752226,7.61263,7.250037,5.9501433,4.650249,3.350355,2.0504606,0.7505665,1.062396,1.3742256,1.6878681,1.9996977,2.3133402,1.8746033,1.4376793,1.0007553,0.5620184,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.4749962,0.9499924,1.4249886,1.8999848,2.374981,1.8999848,1.4249886,0.9499924,0.4749962,0.0,0.07433146,0.15047589,0.22480737,0.2991388,0.37528324,0.36259252,0.34990177,0.33721104,0.3245203,0.31182957,5.1125546,9.911467,14.712192,19.512917,24.311829,30.387066,36.462303,42.53754,48.612778,54.688015,48.12509,41.56217,34.99924,28.438131,21.875206,20.22541,18.575615,16.92582,15.27421,13.6244135,13.45037,13.274512,13.100468,12.92461,12.750566,12.638163,12.525759,12.413355,12.299138,12.186734,10.761745,9.336758,7.911769,6.48678,5.0617914,4.5867953,4.1117992,3.636803,3.1618068,2.6868105,4.12449,5.562169,6.9998484,8.437528,9.875207,10.337513,10.799818,11.262123,11.724429,12.186734,10.700105,9.211663,7.7250338,6.2365913,4.749962,6.011784,7.2754188,8.537241,9.800876,11.062697,10.074633,9.088382,8.100317,7.112252,6.1241875,5.411693,4.699199,3.9867048,3.2742105,2.561716,2.4003625,2.2371957,2.0758421,1.9126755,1.7495089,2.663242,3.5751622,4.4870825,5.4008155,6.3127356,6.3870673,6.4632115,6.5375433,6.6118746,6.688019,6.7623506,6.836682,6.9128265,6.987158,7.063302,8.26167,9.461852,10.662033,11.862214,13.062395,14.349599,15.636803,16.92582,18.213022,19.500225,20.399454,21.300497,22.199726,23.100769,23.999998,23.300196,22.600391,21.900587,21.200785,20.499168,20.48829,20.4756,20.462908,20.450218,20.437527,20.725788,21.012236,21.300497,21.586945,21.875206,21.050308,20.22541,19.400513,18.575615,17.750717,16.325727,14.90074,13.475751,12.050762,10.625773,10.29944,9.97492,9.6504,9.325879,8.999546,8.838193,8.675026,8.511859,8.350506,8.187339,8.287052,8.386765,8.488291,8.588004,8.6877165,10.674724,12.661731,14.650551,16.637558,18.624565,19.063301,19.500225,19.93715,20.375887,20.81281,19.799364,18.787731,17.774284,16.762651,15.749206,15.4246855,15.100165,14.775645,14.449312,14.124791,15.212569,16.300346,17.388124,18.475903,19.561867,16.512463,13.46306,10.411844,7.362441,4.313038,4.274966,4.2368937,4.2006345,4.162562,4.12449,3.299592,2.474694,1.649796,0.824898,0.0,1.6244144,3.2506418,4.8750563,6.4994707,8.125698,7.8755093,7.6253204,7.3751316,7.124943,6.874754,6.5248523,6.1749506,5.825049,5.475147,5.125245,4.4508233,3.774588,3.100166,2.4257438,1.7495089,1.7495089,1.7495089,1.7495089,1.7495089,1.7495089,1.6751775,1.6008459,1.5247015,1.4503701,1.3742256,1.3869164,1.3996071,1.4122978,1.4249886,1.4376793,2.374981,3.3122826,4.249584,5.186886,6.1241875,5.3246713,4.5251546,3.7256382,2.9243085,2.124792,2.3133402,2.5000753,2.6868105,2.8753586,3.0620937,3.350355,3.636803,3.925064,4.213325,4.499773,5.6491914,6.8004227,7.949841,9.099259,10.25049,10.487988,10.725487,10.962985,11.200482,11.437981,11.213174,10.988366,10.761745,10.536939,10.312131,8.849071,7.3878226,5.924762,4.461701,3.000453,4.1117992,5.224958,6.338117,7.4494634,8.562622,7.7866745,7.0125394,6.2365913,5.462456,4.688321,4.788034,4.8877473,4.98746,5.087173,5.186886,5.5005283,5.812358,6.1241875,6.43783,6.7496595,6.149569,5.5494785,4.949388,4.349297,3.7492065,3.000453,2.2498865,1.49932,0.7505665,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.12509441,0.18673515,0.25018883,0.31182957,0.37528324,0.2991388,0.22480737,0.15047589,0.07433146,0.0,0.12509441,0.25018883,0.37528324,0.50037766,0.62547207,0.96268314,1.2998942,1.6371052,1.9743162,2.3133402,2.7756457,3.2379513,3.7002566,4.162562,4.6248674,4.699199,4.7753434,4.8496747,4.9258194,5.0001507,4.512464,4.024777,3.53709,3.049403,2.561716,2.0631514,1.5627737,1.062396,0.5620184,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.0870222,0.11240368,0.13778515,0.16316663,0.18673515,0.22480737,0.26287958,0.2991388,0.33721104,0.37528324,0.2991388,0.22480737,0.15047589,0.07433146,0.0,0.33721104,0.6744221,1.0116332,1.3506571,1.6878681,1.3742256,1.062396,0.7505665,0.43692398,0.12509441,7.262728,14.400362,21.537996,28.675629,35.813263,28.650248,21.487232,14.324218,7.1630154,0.0,0.53663695,1.0750868,1.6117238,2.1501737,2.6868105,2.1501737,1.6117238,1.0750868,0.53663695,0.0,0.0870222,0.17585737,0.26287958,0.34990177,0.43692398,4.213325,7.987913,11.762501,15.537089,19.311678,17.150625,14.9877615,12.824898,10.662033,8.499168,7.799365,7.0995617,6.399758,5.6999545,5.0001507,3.9993954,3.000453,1.9996977,1.0007553,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.61278135,1.2255627,1.8383441,2.4493124,3.0620937,2.4493124,1.8383441,1.2255627,0.61278135,0.0,0.0,0.0,0.0,0.0,0.0,1.4503701,2.9007401,4.349297,5.7996674,7.250037,7.4494634,7.650702,7.850128,8.049554,8.2507925,6.6118746,4.974769,3.3376641,1.7005589,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.2991388,0.6000906,0.89922947,1.2001812,1.49932,2.7992141,4.099108,5.4008155,6.70071,8.000604,8.212721,8.424837,8.636953,8.8508835,9.063,7.837437,6.6118746,5.388125,4.162562,2.9369993,2.3495996,1.7621996,1.1747998,0.5873999,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.33721104,0.6744221,1.0116332,1.3506571,1.6878681,3.2125697,4.7372713,6.261973,7.7866745,9.313189,7.462154,5.612932,3.7618973,1.9126755,0.06164073,0.8122072,1.5627737,2.3133402,3.0620937,3.8126602,2.8372865,3.5280252,4.216951,4.9076896,5.5966153,6.2873545,6.472276,6.6571984,6.8421206,7.027043,7.211965,9.14821,11.082641,13.017072,14.953316,16.887747,17.380873,17.872185,18.36531,18.856625,19.34975,19.360628,19.369692,19.38057,19.389635,19.400513,17.304728,15.210756,13.114971,11.019187,8.925215,9.731983,10.540565,11.347333,12.155914,12.962683,11.680918,10.397341,9.115576,7.8319983,6.550234,13.716875,20.885328,28.05197,35.220425,42.387066,43.84469,45.302307,46.75993,48.217552,49.675175,41.27753,32.87989,24.482246,16.084604,7.686961,7.309865,6.932769,6.5556726,6.1767635,5.7996674,4.7753434,3.7492065,2.7248828,1.7005589,0.6744221,1.1657349,1.6552348,2.1447346,2.6342347,3.1255474,2.8681068,2.610666,2.3532255,2.0957847,1.8383441,1.4902552,1.1421664,0.79589057,0.44780177,0.099712946,0.5855869,1.0696479,1.5555218,2.039583,2.525457,2.0196402,1.5156367,1.0098201,0.5058166,0.0,0.072518505,0.14503701,0.21755551,0.29007402,0.36259252,0.46411842,0.56745726,0.67079616,0.77232206,0.87566096,5.1125546,9.349448,13.588155,17.825048,22.061941,27.520773,32.97779,38.434807,43.891823,49.350655,43.647076,37.94531,32.241726,26.539959,20.838192,19.393261,17.94833,16.501585,15.056654,13.611723,13.575464,13.537392,13.499319,13.46306,13.424988,13.225562,13.024323,12.824898,12.625471,12.4242325,11.035503,9.644961,8.254418,6.8656893,5.475147,4.9657044,4.454449,3.9450066,3.435564,2.9243085,4.1933823,5.4606433,6.7279043,7.995165,9.262425,9.652213,10.042,10.431787,10.823386,11.213174,9.965856,8.716724,7.4694057,6.2220874,4.974769,6.33993,7.705091,9.070251,10.435412,11.800573,10.830639,9.860703,8.890768,7.9208336,6.9508986,6.1296263,5.3101673,4.4907084,3.6694362,2.8499773,2.7266958,2.6052272,2.4819458,2.3604772,2.2371957,3.159994,4.082792,5.0055895,5.9283876,6.849373,6.887445,6.925517,6.9617763,6.9998484,7.037921,7.0506115,7.063302,7.07418,7.0868707,7.0995617,8.200029,9.300498,10.399154,11.499621,12.60009,14.045021,15.489952,16.934883,18.379814,19.824745,20.540867,21.255173,21.96948,22.6856,23.399908,22.600391,21.800875,20.999546,20.20003,19.400513,19.420456,19.440397,19.46034,19.480284,19.500225,19.610817,19.719595,19.830185,19.940775,20.049553,19.36788,18.684393,18.002718,17.319231,16.637558,15.198066,13.75676,12.317267,10.877775,9.438283,9.256987,9.077503,8.898021,8.716724,8.537241,8.410334,8.281613,8.154706,8.027799,7.900891,8.01692,8.134763,8.252605,8.370448,8.488291,10.48255,12.476809,14.47288,16.467138,18.463211,18.628191,18.79317,18.958149,19.123129,19.288109,18.446894,17.607492,16.768091,15.926876,15.087475,14.889862,14.692248,14.494636,14.297023,14.09941,15.179935,16.260462,17.339174,18.4197,19.500225,16.33298,13.165734,9.9966755,6.82943,3.6621845,3.832603,4.0030212,4.171627,4.3420453,4.512464,3.6096084,2.7067533,1.8057107,0.90285534,0.0,1.4467441,2.8953013,4.3420453,5.7906027,7.2373466,7.112252,6.987158,6.8620634,6.736969,6.6118746,6.249282,5.8866897,5.524097,5.163317,4.800725,4.2423325,3.6857529,3.1273603,2.570781,2.0123885,1.892733,1.7730774,1.651609,1.5319533,1.4122978,1.9217403,2.4329958,2.9424384,3.4518807,3.9631362,3.832603,3.7020695,3.5733492,3.442816,3.3122826,4.2223897,5.132497,6.0426044,6.9527116,7.8628187,6.7677894,5.67276,4.5777307,3.482701,2.3876717,2.4529383,2.518205,2.5816586,2.6469254,2.712192,3.2669585,3.8217251,4.3783045,4.933071,5.487838,6.4668374,7.4476504,8.42665,9.407463,10.388275,10.866898,11.347333,11.827768,12.308203,12.786825,12.215742,11.642846,11.069949,10.497053,9.924157,8.54268,7.159389,5.7779117,4.3946214,3.0131438,4.077353,5.141562,6.207584,7.271793,8.337815,7.567306,6.796797,6.0281005,5.2575917,4.4870825,4.572292,4.6575007,4.74271,4.8279195,4.9131284,5.163317,5.411693,5.661882,5.9120708,6.16226,5.5331616,4.902251,4.273153,3.6422417,3.0131438,2.810092,2.6070402,2.4058013,2.2027495,1.9996977,1.6044719,1.209246,0.81583315,0.42060733,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.052575916,0.054388877,0.058014803,0.059827764,0.06164073,0.11240368,0.16316663,0.21211663,0.26287958,0.31182957,0.2520018,0.19217403,0.13234627,0.072518505,0.012690738,0.11240368,0.21211663,0.31182957,0.41335547,0.51306844,1.1022812,1.693307,2.2825198,2.8717327,3.4627585,3.825351,4.1879435,4.550536,4.9131284,5.275721,5.2503395,5.224958,5.199577,5.1741953,5.1506267,4.7300196,4.309412,3.8906176,3.4700103,3.049403,2.6741197,2.3006494,1.9253663,1.550083,1.1747998,0.9445535,0.71430725,0.48587397,0.25562772,0.025381476,0.02175555,0.01994259,0.018129626,0.014503701,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.02175555,0.032633327,0.04169814,0.052575916,0.06164073,0.06707962,0.072518505,0.07795739,0.08339628,0.0870222,0.10696479,0.12690738,0.14684997,0.16679256,0.18673515,0.22480737,0.26287958,0.2991388,0.33721104,0.37528324,0.33539808,0.2955129,0.25562772,0.21574254,0.17585737,0.41335547,0.6508536,0.8883517,1.1258497,1.3633479,1.1131591,0.8629702,0.61278135,0.36259252,0.11240368,6.198519,12.282822,18.367125,24.45324,30.537542,24.49675,18.457771,12.416981,6.378002,0.33721104,0.9354887,1.5319533,2.1302311,2.7266958,3.3249733,2.6704938,2.0142014,1.3597219,0.70524246,0.05076295,0.11784257,0.18492219,0.2520018,0.3208944,0.387974,3.680314,6.972654,10.264994,13.557334,16.849674,15.0421505,13.234627,11.427103,9.619579,7.8120556,7.135821,6.4577727,5.7797246,5.101677,4.4254417,3.540716,2.6541772,1.7694515,0.88472575,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.4894999,0.9808127,1.4703126,1.9598125,2.4493124,1.9815681,1.5156367,1.0478923,0.58014804,0.11240368,0.31182957,0.51306844,0.7124943,0.9119202,1.1131591,2.4094272,3.7075086,5.0055895,6.301858,7.5999393,7.835624,8.069496,8.3051815,8.540867,8.774739,7.0306687,5.2847857,3.540716,1.794833,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.38072214,0.75963134,1.1403534,1.5192627,1.8999848,2.864481,3.83079,4.795286,5.7597823,6.7242785,7.132195,7.5401115,7.948028,8.354132,8.762048,7.4929743,6.2220874,4.953014,3.682127,2.4130533,1.9326181,1.452183,0.97174793,0.49312583,0.012690738,0.014503701,0.018129626,0.01994259,0.02175555,0.025381476,0.030820364,0.034446288,0.03988518,0.045324065,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.291887,0.5855869,0.8774739,1.1693609,1.4630609,3.054842,4.648436,6.240217,7.8319983,9.425592,7.5781837,5.728962,3.881553,2.035957,0.18673515,0.81764615,1.4467441,2.077655,2.7067533,3.3376641,2.7375734,3.4555066,4.171627,4.88956,5.6074934,6.3254266,6.644508,6.965402,7.2844834,7.605378,7.9244595,9.782746,11.63922,13.497506,15.355793,17.212267,17.609306,18.008158,18.405195,18.802235,19.199274,18.958149,18.715212,18.472277,18.22934,17.988214,16.097294,14.208188,12.317267,10.428161,8.537241,9.590572,10.642091,11.695421,12.74694,13.800271,12.43511,11.069949,9.704789,8.339628,6.9744673,15.946819,24.91917,33.893337,42.86569,51.83804,50.128414,48.416977,46.707355,44.99773,43.28811,35.893032,28.49796,21.102884,13.70781,6.3127356,5.919323,5.527723,5.1343102,4.74271,4.349297,3.6005437,2.8499773,2.0994108,1.3506571,0.6000906,1.2672608,1.9344311,2.6034143,3.2705846,3.9377546,3.8597972,3.7818398,3.7056956,3.6277382,3.5497808,2.8807976,2.2100015,1.5392052,0.87022203,0.19942589,0.69436467,1.1893034,1.6842422,2.179181,2.6741197,2.1392958,1.6044719,1.0696479,0.53482395,0.0,0.07070554,0.13959812,0.21030366,0.27919623,0.34990177,0.56745726,0.7850128,1.0025684,1.2201238,1.4376793,5.1125546,8.78743,12.462305,16.13718,19.812056,24.652666,29.491463,34.332073,39.172684,44.013294,39.170868,34.328445,29.484211,24.641787,19.799364,18.559298,17.319231,16.079165,14.839099,13.600845,13.700559,13.800271,13.899984,13.999697,14.09941,13.812962,13.524701,13.238253,12.949992,12.661731,11.307447,9.953164,8.597069,7.2427855,5.8866897,5.3428006,4.797099,4.25321,3.7075086,3.1618068,4.2604623,5.3573046,6.454147,7.552802,8.649645,8.966913,9.284182,9.603263,9.920531,10.2378,9.229793,8.221786,7.215591,6.207584,5.199577,6.6680765,8.134763,9.603263,11.069949,12.536636,11.584831,10.633025,9.679407,8.727602,7.7757964,6.8475595,5.919323,4.992899,4.064662,3.1382382,3.054842,2.9732587,2.8898623,2.808279,2.7248828,3.6567454,4.590421,5.522284,6.454147,7.3878226,7.3878226,7.3878226,7.3878226,7.3878226,7.3878226,7.3370595,7.28811,7.2373466,7.1883965,7.137634,8.138389,9.137331,10.138086,11.137029,12.137785,13.740443,15.343102,16.94576,18.54842,20.149265,20.680464,21.209848,21.739235,22.270432,22.799818,21.900587,20.999546,20.100317,19.199274,18.300045,18.352621,18.405195,18.457771,18.510347,18.562923,18.495844,18.426952,18.359873,18.292793,18.225714,17.68545,17.145187,16.604925,16.064661,15.524399,14.070402,12.6145935,11.160598,9.704789,8.2507925,8.214534,8.180087,8.145641,8.109382,8.074935,7.9824743,7.890013,7.797552,7.705091,7.61263,7.746789,7.8827615,8.01692,8.152893,8.287052,10.290376,12.291886,14.29521,16.29672,18.300045,18.193079,18.084301,17.977337,17.870373,17.761595,17.094423,16.427254,15.760084,15.092914,14.425743,14.355038,14.284332,14.21544,14.144734,14.075842,15.147303,16.220575,17.292038,18.36531,19.436771,16.151684,12.868408,9.581508,6.298232,3.0131438,3.39024,3.7673361,4.1444325,4.5233417,4.900438,3.919625,2.9406252,1.9598125,0.9808127,0.0,1.2690738,2.5399606,3.8108473,5.0799212,6.350808,6.350808,6.350808,6.350808,6.350808,6.350808,5.975525,5.600241,5.224958,4.8496747,4.4743915,4.0356545,3.5951047,3.1545548,2.715818,2.275268,2.034144,1.794833,1.5555218,1.3143979,1.0750868,2.1701162,3.2651455,4.360175,5.4552045,6.550234,6.2782893,6.004532,5.732588,5.4606433,5.186886,6.069799,6.9527116,7.835624,8.716724,9.599637,8.209095,6.8203654,5.429823,4.0392804,2.6505513,2.5925364,2.5345216,2.47832,2.420305,2.3622901,3.1853752,4.006647,4.8297324,5.6528172,6.4759026,7.2844834,8.094878,8.9052725,9.715667,10.524248,11.24762,11.969179,12.692551,13.415923,14.137483,13.21831,12.297325,11.378153,10.457169,9.537996,8.234476,6.932769,5.6292486,4.327542,3.0258346,4.0429068,5.0599785,6.0770507,7.0941224,8.113008,7.3479376,6.582867,5.8177967,5.0527267,4.2876563,4.358362,4.4272547,4.49796,4.5668526,4.6375585,4.8242936,5.0128417,5.199577,5.388125,5.57486,4.914942,4.255023,3.5951047,2.9351864,2.275268,2.619731,2.9641938,3.3104696,3.6549325,3.9993954,3.2107568,2.420305,1.6298534,0.83940166,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.04169814,0.047137026,0.052575916,0.058014803,0.06164073,0.099712946,0.13778515,0.17585737,0.21211663,0.25018883,0.20486477,0.15954071,0.11421664,0.07070554,0.025381476,0.099712946,0.17585737,0.25018883,0.3245203,0.40066472,1.2418793,2.084907,2.9279346,3.7691493,4.612177,4.8750563,5.137936,5.4008155,5.661882,5.924762,5.7996674,5.674573,5.5494785,5.424384,5.2992897,4.947575,4.59586,4.2423325,3.8906176,3.53709,3.2869012,3.0367124,2.7883365,2.5381477,2.2879589,1.840157,1.3923552,0.9445535,0.49675176,0.05076295,0.045324065,0.03988518,0.034446288,0.030820364,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.032633327,0.03988518,0.047137026,0.054388877,0.06164073,0.072518505,0.08339628,0.092461094,0.10333887,0.11240368,0.12690738,0.14322405,0.15772775,0.17223145,0.18673515,0.22480737,0.26287958,0.2991388,0.33721104,0.37528324,0.36984438,0.36440548,0.36077955,0.35534066,0.34990177,0.48768693,0.62547207,0.76325727,0.89922947,1.0370146,0.85027945,0.66173136,0.4749962,0.28826106,0.099712946,5.132497,10.165281,15.198066,20.23085,25.26182,20.345066,15.428311,10.509744,5.5929894,0.6744221,1.3325275,1.9906329,2.6469254,3.3050308,3.9631362,3.1908143,2.4166791,1.6443571,0.872035,0.099712946,0.14684997,0.19579996,0.24293698,0.29007402,0.33721104,3.147303,5.957395,8.767487,11.5775795,14.387671,12.935488,11.483305,10.029309,8.577126,7.124943,6.4704633,5.814171,5.1596913,4.505212,3.8507326,3.0802233,2.3097143,1.5392052,0.7705091,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.3680314,0.73424983,1.1022812,1.4703126,1.8383441,1.5156367,1.1929294,0.87022203,0.5475147,0.22480737,0.62547207,1.0243238,1.4249886,1.8256533,2.2245052,3.3702974,4.514277,5.660069,6.8040485,7.949841,8.219973,8.490104,8.760235,9.030367,9.300498,7.4476504,5.5948024,3.7419548,1.8909199,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.4604925,0.91917205,1.3796645,1.840157,2.3006494,2.9297476,3.5606585,4.1897564,4.8206677,5.4497657,6.051669,6.6553855,7.2572894,7.859193,8.46291,7.1466985,5.8323007,4.517903,3.2016919,1.887294,1.5156367,1.1421664,0.7705091,0.39703882,0.025381476,0.030820364,0.034446288,0.03988518,0.045324065,0.05076295,0.047137026,0.045324065,0.04169814,0.03988518,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.24837588,0.4949388,0.7433147,0.9898776,1.2382535,2.8971143,4.557788,6.2166486,7.877322,9.537996,7.6924005,5.846804,4.0030212,2.1574254,0.31182957,0.823085,1.3325275,1.84197,2.3532255,2.8626678,2.6378605,3.3829882,4.1281157,4.8732433,5.618371,6.3616858,6.816739,7.271793,7.7268467,8.1819,8.636953,10.417283,12.197612,13.9779415,15.758271,17.536787,17.839552,18.142317,18.445082,18.747847,19.050611,18.555672,18.060734,17.565794,17.070856,16.575916,14.889862,13.20562,11.519565,9.835322,8.149267,9.447348,10.745429,12.0416975,13.339779,14.63786,13.189302,11.7425585,10.2958145,8.847258,7.400513,18.176764,28.954826,39.732887,50.510952,61.2872,56.41033,51.533463,46.654778,41.77791,36.899227,30.508533,24.116028,17.721708,11.329204,4.936697,4.5305934,4.122677,3.7147603,3.3068438,2.9007401,2.4257438,1.9507477,1.4757515,1.0007553,0.52575916,1.3705997,2.2154403,3.0602808,3.9051213,4.749962,4.853301,4.954827,5.0581656,5.1596913,5.2630305,4.269527,3.2778363,2.2843328,1.2926424,0.2991388,0.80495536,1.310772,1.8147756,2.3205922,2.8245957,2.2607644,1.69512,1.1294757,0.5656443,0.0,0.06707962,0.13415924,0.2030518,0.27013144,0.33721104,0.67079616,1.0025684,1.3343405,1.6679256,1.9996977,5.1125546,8.225411,11.338268,14.449312,17.562168,21.78456,26.006948,30.229338,34.45173,38.67593,34.692852,30.709774,26.726694,22.745428,18.76235,17.727148,16.691946,15.656745,14.623356,13.588155,13.825653,14.06315,14.300649,14.538147,14.775645,14.400362,14.025079,13.649796,13.274512,12.899229,11.579392,10.259555,8.939718,7.6198816,6.300045,5.719897,5.139749,4.559601,3.9794528,3.3993049,4.327542,5.2557783,6.1822023,7.1104393,8.036863,8.281613,8.528176,8.772926,9.017676,9.262425,8.495543,7.7268467,6.9599633,6.19308,5.424384,6.9944096,8.564435,10.13446,11.704487,13.274512,12.340837,11.405348,10.469859,9.53437,8.600695,7.5654926,6.530291,5.4950895,4.459888,3.4246864,3.3829882,3.339477,3.2977788,3.254268,3.2125697,4.15531,5.0980506,6.0407915,6.981719,7.9244595,7.8882003,7.850128,7.8120556,7.7757964,7.7377243,7.6253204,7.512917,7.400513,7.28811,7.175706,8.074935,8.974165,9.875207,10.774437,11.675479,13.435865,15.194439,16.954826,18.715212,20.4756,20.820063,21.164526,21.510801,21.855265,22.199726,21.200785,20.20003,19.199274,18.20033,17.199575,17.284784,17.369995,17.455204,17.540413,17.625622,17.380873,17.13431,16.889559,16.64481,16.400059,16.003021,15.604169,15.20713,14.810091,14.413053,12.9427395,11.472427,10.002114,8.531802,7.063302,7.17208,7.2826705,7.3932614,7.502039,7.61263,7.554615,7.4966,7.440398,7.382384,7.324369,7.476658,7.6307597,7.783048,7.935337,8.087626,10.098202,12.106964,14.117539,16.128115,18.136877,17.757969,17.377247,16.998337,16.617615,16.236893,15.741954,15.247015,14.752076,14.257137,13.762199,13.820213,13.878228,13.93443,13.992445,14.05046,15.114669,16.18069,17.2449,18.310923,19.375132,15.9722,12.569269,9.168152,5.765221,2.3622901,2.9478772,3.531651,4.117238,4.702825,5.2865987,4.229642,3.1726844,2.1157274,1.0569572,0.0,1.0932164,2.18462,3.2778363,4.36924,5.462456,5.5875506,5.712645,5.8377395,5.962834,6.0879283,5.6999545,5.3119802,4.9258194,4.537845,4.1498713,3.827164,3.5044568,3.1817493,2.8608549,2.5381477,2.1773682,1.8184015,1.4576219,1.0968424,0.73787576,2.4166791,4.0972953,5.7779117,7.456715,9.137331,8.722163,8.306994,7.891826,7.476658,7.063302,7.9172077,8.772926,9.626831,10.48255,11.338268,9.652213,7.9679704,6.281915,4.597673,2.911618,2.7321346,2.5526514,2.373168,2.1918716,2.0123885,3.101979,4.1915693,5.282973,6.3725634,7.462154,8.10213,8.7421055,9.382081,10.022058,10.662033,11.628342,12.592838,13.557334,14.521831,15.488139,14.219066,12.951805,11.684544,10.417283,9.1500225,7.9280853,6.7043357,5.482399,4.2604623,3.0367124,4.00846,4.976582,5.9483304,6.9182653,7.8882003,7.1267557,6.3671246,5.6074934,4.847862,4.0882306,4.1426196,4.1970086,4.25321,4.307599,4.361988,4.4870825,4.612177,4.7372713,4.8623657,4.98746,4.2967215,3.6077955,2.9170568,2.228131,1.5373923,2.42937,3.3231604,4.215138,5.1071157,5.999093,4.8152285,3.6295512,2.4456866,1.260009,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.032633327,0.03988518,0.047137026,0.054388877,0.06164073,0.0870222,0.11240368,0.13778515,0.16316663,0.18673515,0.15772775,0.12690738,0.09789998,0.06707962,0.038072214,0.0870222,0.13778515,0.18673515,0.2374981,0.28826106,1.3832904,2.47832,3.5733492,4.668379,5.7615952,5.924762,6.0879283,6.249282,6.412449,6.5756154,6.350808,6.1241875,5.89938,5.674573,5.4497657,5.1651306,4.880495,4.59586,4.309412,4.024777,3.8996825,3.774588,3.6494937,3.5243993,3.3993049,2.7357605,2.0704033,1.405046,0.73968875,0.07433146,0.06707962,0.059827764,0.052575916,0.045324065,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.04169814,0.047137026,0.052575916,0.058014803,0.06164073,0.07795739,0.092461094,0.10696479,0.12328146,0.13778515,0.14684997,0.15772775,0.16679256,0.17767033,0.18673515,0.22480737,0.26287958,0.2991388,0.33721104,0.37528324,0.40429065,0.43511102,0.46411842,0.4949388,0.52575916,0.5620184,0.6000906,0.63816285,0.6744221,0.7124943,0.5873999,0.46230546,0.33721104,0.21211663,0.0870222,4.068288,8.047741,12.027194,16.00846,19.987913,16.191568,12.397038,8.602508,4.8079767,1.0116332,1.7295663,2.4474995,3.1654327,3.8833659,4.599486,3.7093215,2.819157,1.9308052,1.0406405,0.15047589,0.17767033,0.20486477,0.23205921,0.25925365,0.28826106,2.6142921,4.942136,7.26998,9.597824,11.925668,10.827013,9.73017,8.6333275,7.5346723,6.43783,5.805106,5.1723824,4.539658,3.9069343,3.2742105,2.619731,1.9652514,1.310772,0.6544795,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.24474995,0.4894999,0.73424983,0.9808127,1.2255627,1.0478923,0.87022203,0.69255173,0.5148814,0.33721104,0.93730164,1.5373923,2.137483,2.7375734,3.3376641,4.329355,5.3228583,6.3145485,7.308052,8.299743,8.604321,8.910711,9.215289,9.519867,9.824444,7.8646317,5.904819,3.9450066,1.9851941,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.5402629,1.0805258,1.6207886,2.1592383,2.6995013,2.9950142,3.290527,3.584227,3.87974,4.175253,4.972956,5.77066,6.5683637,7.364254,8.161958,6.8022356,5.4425135,4.082792,2.72307,1.3633479,1.0968424,0.8321498,0.56745726,0.30276474,0.038072214,0.045324065,0.052575916,0.059827764,0.06707962,0.07433146,0.065266654,0.054388877,0.045324065,0.034446288,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.2030518,0.40429065,0.6073425,0.8103943,1.0116332,2.7393866,4.4671397,6.1948934,7.9226465,9.6504,7.806617,5.964647,4.122677,2.280707,0.43692398,0.82671094,1.2183108,1.6080978,1.9978848,2.3876717,2.5381477,3.3104696,4.082792,4.855114,5.6274357,6.399758,6.9907837,7.5799966,8.1692095,8.760235,9.349448,11.05182,12.754191,14.458377,16.160748,17.863121,18.069798,18.278288,18.484966,18.691645,18.900135,18.153194,17.40444,16.6575,15.91056,15.161806,13.682428,12.203052,10.721861,9.242483,7.763106,9.304124,10.846955,12.389787,13.932617,15.475449,13.945308,12.415168,10.885027,9.354887,7.8247466,20.406708,32.99048,45.57244,58.15621,70.738174,62.692245,54.648132,46.602203,38.558086,30.51216,25.122223,19.732285,14.342347,8.952409,3.5624714,3.1400511,2.7176309,2.2952106,1.8727903,1.4503701,1.2491312,1.0497054,0.85027945,0.6508536,0.44961473,1.4721256,2.4946365,3.5171473,4.539658,5.562169,5.844991,6.1278133,6.4106355,6.6916447,6.9744673,5.660069,4.345671,3.0294604,1.7150626,0.40066472,0.9155461,1.4304274,1.9453088,2.4601903,2.9750717,2.38042,1.7857682,1.1893034,0.5946517,0.0,0.065266654,0.13053331,0.19579996,0.25925365,0.3245203,0.77232206,1.2201238,1.6679256,2.1157274,2.561716,5.1125546,7.66158,10.212419,12.763257,15.312282,18.918264,22.522434,26.128416,29.732586,33.336758,30.214834,27.092913,23.96918,20.847258,17.725336,16.894999,16.064661,15.234324,14.405801,13.575464,13.9507475,14.324218,14.699501,15.074784,15.4500675,14.9877615,14.525456,14.06315,13.600845,13.136727,11.853149,10.567759,9.282369,7.996978,6.7134004,6.096993,5.482399,4.8678045,4.25321,3.636803,4.3946214,5.1524396,5.910258,6.6680765,7.4258947,7.5981264,7.7703576,7.9425893,8.1148205,8.287052,7.75948,7.231908,6.7043357,6.1767635,5.6491914,7.322556,8.994107,10.667472,12.340837,14.012388,13.095029,12.17767,11.26031,10.342952,9.425592,8.283426,7.1394467,5.99728,4.855114,3.7129474,3.7093215,3.7075086,3.7056956,3.7020695,3.7002566,4.652062,5.6056805,6.5574856,7.509291,8.46291,8.386765,8.312433,8.238102,8.161958,8.087626,7.911769,7.7377243,7.5618668,7.3878226,7.211965,8.013294,8.812811,9.612328,10.411844,11.213174,13.129475,15.047589,16.965704,18.882006,20.80012,20.95966,21.119202,21.280556,21.440096,21.599636,20.499168,19.400513,18.300045,17.199575,16.099108,16.21695,16.334793,16.452635,16.570478,16.68832,16.264088,15.841667,15.419247,14.996826,14.574407,14.320591,14.064963,13.809336,13.555521,13.299893,11.815077,10.330261,8.845445,7.360628,5.8758116,6.1296263,6.3852544,6.640882,6.8946967,7.1503243,7.1267557,7.1050005,7.083245,7.059676,7.037921,7.208339,7.3769445,7.5473633,7.7177815,7.8882003,9.904215,11.922042,13.939869,15.957697,17.975525,17.322857,16.67019,16.017525,15.364858,14.712192,14.389484,14.066776,13.744069,13.423175,13.100468,13.28539,13.470312,13.655234,13.840157,14.025079,15.082036,16.140806,17.197763,18.25472,19.311678,15.792717,12.271944,8.752983,5.23221,1.7132497,2.5055144,3.2977788,4.0900435,4.882308,5.674573,4.539658,3.4047437,2.269829,1.1349145,0.0,0.9155461,1.8292793,2.7448254,3.6603715,4.574105,4.8242936,5.0744824,5.3246713,5.57486,5.825049,5.424384,5.0255322,4.6248674,4.2242026,3.825351,3.6204863,3.4156215,3.2107568,3.005892,2.7992141,2.3205922,1.840157,1.3597219,0.8792868,0.40066472,2.665055,4.9294453,7.1956487,9.460039,11.724429,11.16785,10.609457,10.052877,9.494485,8.937905,9.764616,10.593141,11.419851,12.248375,13.075087,11.095331,9.115576,7.135821,5.1542525,3.1744974,2.8717327,2.570781,2.268016,1.9652514,1.6624867,3.0203958,4.3783045,5.7344007,7.0923095,8.450218,8.919776,9.389333,9.860703,10.330261,10.799818,12.007251,13.2146845,14.422117,15.62955,16.836983,15.221634,13.608097,11.992747,10.377398,8.762048,7.6198816,6.4777155,5.335549,4.1933823,3.049403,3.972201,4.894999,5.8177967,6.740595,7.663393,6.9073873,6.153195,5.3971896,4.6429973,3.8869917,3.926877,3.966762,4.006647,4.0483456,4.0882306,4.1498713,4.213325,4.274966,4.3366065,4.40006,3.680314,2.960568,2.2408218,1.5192627,0.7995165,2.2408218,3.680314,5.1198063,6.5592985,8.000604,6.4197006,4.84061,3.2597067,1.6806163,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.02175555,0.032633327,0.04169814,0.052575916,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.11059072,0.09427405,0.07977036,0.065266654,0.05076295,0.07433146,0.099712946,0.12509441,0.15047589,0.17585737,1.5228885,2.8699198,4.216951,5.565795,6.9128265,6.9744673,7.037921,7.0995617,7.1630154,7.224656,6.9001355,6.5756154,6.249282,5.924762,5.600241,5.382686,5.1651306,4.947575,4.7300196,4.512464,4.512464,4.512464,4.512464,4.512464,4.512464,3.6295512,2.7466383,1.8655385,0.9826257,0.099712946,0.09064813,0.07977036,0.07070554,0.059827764,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.052575916,0.054388877,0.058014803,0.059827764,0.06164073,0.08339628,0.10333887,0.12328146,0.14322405,0.16316663,0.16679256,0.17223145,0.17767033,0.18310922,0.18673515,0.22480737,0.26287958,0.2991388,0.33721104,0.37528324,0.4405499,0.5058166,0.56927025,0.6345369,0.69980353,0.63816285,0.5747091,0.51306844,0.44961473,0.387974,0.3245203,0.26287958,0.19942589,0.13778515,0.07433146,3.002266,5.9302006,8.858135,11.784257,14.712192,12.039885,9.367578,6.695271,4.022964,1.3506571,2.128418,2.904366,3.682127,4.459888,5.237649,4.229642,3.2216346,2.2154403,1.2074331,0.19942589,0.20667773,0.21574254,0.2229944,0.23024625,0.2374981,2.0830941,3.926877,5.772473,7.6180687,9.461852,8.72035,7.9770355,7.2355337,6.492219,5.750717,5.139749,4.5305934,3.919625,3.3104696,2.6995013,2.1592383,1.6207886,1.0805258,0.5402629,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.12328146,0.24474995,0.3680314,0.4894999,0.61278135,0.58014804,0.5475147,0.5148814,0.48224804,0.44961473,1.2509441,2.0504606,2.8499773,3.6494937,4.4508233,5.290225,6.1296263,6.970841,7.8102427,8.649645,8.990481,9.329506,9.670342,10.009366,10.3502035,8.281613,6.2148356,4.1480584,2.079468,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.6200332,1.2400664,1.8600996,2.4801328,3.100166,3.0602808,3.0203958,2.9805105,2.9406252,2.9007401,3.8924308,4.8841214,5.8776245,6.869315,7.8628187,6.4577727,5.0527267,3.6476808,2.2426348,0.8375887,0.67986095,0.52213323,0.36440548,0.20667773,0.05076295,0.059827764,0.07070554,0.07977036,0.09064813,0.099712946,0.08339628,0.065266654,0.047137026,0.030820364,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.15772775,0.3154555,0.47318324,0.629098,0.7868258,2.5834718,4.3783045,6.1731377,7.9679704,9.762803,7.9226465,6.0824895,4.2423325,2.4021754,0.5620184,0.8321498,1.1022812,1.3724127,1.6425442,1.9126755,2.4366217,3.2379513,4.0374675,4.836984,5.638314,6.43783,7.1630154,7.8882003,8.613385,9.336758,10.061942,11.6881695,13.312584,14.936998,16.563227,18.187641,18.300045,18.412449,18.52485,18.637255,18.749659,17.750717,16.749962,15.749206,14.750263,13.749508,12.474996,11.200482,9.924157,8.649645,7.3751316,9.162713,10.950294,12.737875,14.525456,16.313038,14.699501,13.087777,11.47424,9.862516,8.2507925,22.63665,37.024323,51.413807,65.79967,80.18733,68.975975,57.762802,46.549625,35.336452,24.125093,19.737724,15.350354,10.962985,6.5756154,2.1882458,1.7495089,1.3125849,0.87566096,0.43692398,0.0,0.07433146,0.15047589,0.22480737,0.2991388,0.37528324,1.5754645,2.7756457,3.975827,5.1741953,6.3743763,6.836682,7.3008003,7.763106,8.225411,8.6877165,7.0506115,5.411693,3.774588,2.137483,0.50037766,1.0243238,1.550083,2.0758421,2.5997884,3.1255474,2.5000753,1.8746033,1.2491312,0.62547207,0.0,0.06164073,0.12509441,0.18673515,0.25018883,0.31182957,0.87566096,1.4376793,1.9996977,2.561716,3.1255474,5.1125546,7.0995617,9.088382,11.075388,13.062395,16.050158,19.03792,22.025682,25.013445,27.999393,25.736816,23.47424,21.211662,18.949085,16.68832,16.062849,15.437376,14.811904,14.188245,13.562773,14.075842,14.587097,15.100165,15.613234,16.124489,15.575162,15.025834,14.474693,13.925365,13.374225,12.125093,10.874149,9.625018,8.375887,7.124943,6.4759026,5.825049,5.1741953,4.5251546,3.874301,4.461701,5.049101,5.638314,6.2257137,6.813113,6.9128265,7.0125394,7.112252,7.211965,7.311678,7.02523,6.736969,6.450521,6.16226,5.8758116,7.650702,9.425592,11.200482,12.975373,14.750263,13.849221,12.949992,12.050762,11.14972,10.25049,8.999546,7.750415,6.4994707,5.2503395,3.9993954,4.0374675,4.07554,4.1117992,4.1498713,4.1879435,5.1506267,6.11331,7.07418,8.036863,8.999546,8.887142,8.774739,8.662335,8.549932,8.437528,8.200029,7.9625316,7.7250338,7.4875355,7.250037,7.949841,8.649645,9.349448,10.049252,10.750868,12.824898,14.90074,16.97477,19.050611,21.12464,21.099258,21.07569,21.050308,21.024927,20.999546,19.799364,18.599184,17.400814,16.200634,15.000452,15.149116,15.299591,15.4500675,15.600543,15.749206,15.149116,14.5508375,13.9507475,13.3506565,12.750566,12.638163,12.525759,12.413355,12.299138,12.186734,10.687414,9.188094,7.686961,6.187641,4.688321,5.087173,5.487838,5.8866897,6.2873545,6.688019,6.70071,6.7134004,6.7242785,6.736969,6.7496595,6.9382076,7.124943,7.311678,7.500226,7.686961,9.712041,11.73712,13.762199,15.787278,17.812357,16.887747,15.963136,15.036712,14.112101,13.1874895,13.037014,12.888351,12.737875,12.5873995,12.436923,12.750566,13.062395,13.374225,13.687867,13.999697,15.049402,16.099108,17.150625,18.20033,19.250036,15.613234,11.974618,8.337815,4.699199,1.062396,2.0631514,3.0620937,4.062849,5.0617914,6.0625467,4.8496747,3.636803,2.4257438,1.2128719,0.0,0.73787576,1.4757515,2.2118144,2.94969,3.6875658,4.062849,4.4381323,4.8134155,5.186886,5.562169,5.1506267,4.7372713,4.325729,3.9123733,3.5008307,3.4119956,3.3249733,3.2379513,3.149116,3.0620937,2.4620032,1.8619126,1.261822,0.66173136,0.06164073,2.911618,5.7615952,8.613385,11.463363,14.313339,13.611723,12.91192,12.212116,11.512312,10.812509,11.612025,12.413355,13.212872,14.012388,14.811904,12.536636,10.263181,7.987913,5.712645,3.437377,3.0131438,2.5870976,2.1628644,1.7368182,1.3125849,2.9369993,4.5632267,6.187641,7.8120556,9.438283,9.737422,10.038374,10.337513,10.636651,10.937603,12.387974,13.838344,15.2869005,16.73727,18.187641,16.224201,14.262577,12.299138,10.337513,8.375887,7.311678,6.249282,5.186886,4.12449,3.0620937,3.9377546,4.8116026,5.6872635,6.5629244,7.4367723,6.688019,5.9374523,5.186886,4.4381323,3.6875658,3.7129474,3.738329,3.7618973,3.787279,3.8126602,3.8126602,3.8126602,3.8126602,3.8126602,3.8126602,3.0620937,2.3133402,1.5627737,0.8122072,0.06164073,2.0504606,4.0374675,6.0244746,8.013294,10.000301,8.024173,6.049856,4.07554,2.0994108,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,1.6624867,3.2633326,4.8623657,6.4632115,8.062244,8.024173,7.987913,7.949841,7.911769,7.8755093,7.4494634,7.02523,6.599184,6.1749506,5.750717,5.600241,5.4497657,5.2992897,5.1506267,5.0001507,5.125245,5.2503395,5.375434,5.5005283,5.6256227,4.5251546,3.4246864,2.324218,1.2255627,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.0870222,0.11240368,0.13778515,0.16316663,0.18673515,0.18673515,0.18673515,0.18673515,0.18673515,0.18673515,0.22480737,0.26287958,0.2991388,0.33721104,0.37528324,0.4749962,0.5747091,0.6744221,0.774135,0.87566096,0.7124943,0.5493277,0.387974,0.22480737,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,1.938057,3.8126602,5.6872635,7.5618668,9.438283,7.8882003,6.338117,4.788034,3.2379513,1.6878681,2.525457,3.3630457,4.2006345,5.038223,5.8758116,4.749962,3.625925,2.5000753,1.3742256,0.25018883,0.2374981,0.22480737,0.21211663,0.19942589,0.18673515,1.550083,2.911618,4.274966,5.638314,6.9998484,6.6118746,6.2257137,5.8377395,5.4497657,5.0617914,4.4743915,3.8869917,3.299592,2.712192,2.124792,1.7005589,1.2745126,0.85027945,0.42423326,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.11240368,0.22480737,0.33721104,0.44961473,0.5620184,1.5627737,2.561716,3.5624714,4.5632267,5.562169,6.249282,6.9382076,7.6253204,8.312433,8.999546,9.374829,9.750113,10.125396,10.500679,10.874149,8.700407,6.5248523,4.349297,2.175555,0.0,0.0,0.0,0.0,0.0,0.0,0.69980353,1.3996071,2.0994108,2.7992141,3.5008307,3.1255474,2.7502642,2.374981,1.9996977,1.6244144,2.811905,3.9993954,5.186886,6.3743763,7.5618668,6.11331,4.6629395,3.2125697,1.7621996,0.31182957,0.26287958,0.21211663,0.16316663,0.11240368,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.11240368,0.22480737,0.33721104,0.44961473,0.5620184,2.4257438,4.2876563,6.149569,8.011481,9.875207,8.036863,6.200332,4.361988,2.525457,0.6871128,0.8375887,0.9880646,1.1367276,1.2872034,1.4376793,2.4130533,3.149116,3.8869917,4.6248674,5.3627434,6.1006193,6.755099,7.409578,8.06587,8.72035,9.374829,10.877775,12.380721,13.881854,15.384801,16.887747,17.192324,17.496902,17.803293,18.10787,18.412449,17.375433,16.338419,15.299591,14.262577,13.225562,12.348088,11.470614,10.593141,9.715667,8.838193,10.520622,12.203052,13.885481,15.567909,17.25034,16.236893,15.22526,14.211814,13.200181,12.186734,25.34159,38.49645,51.65312,64.807976,77.96283,66.49222,55.023415,43.5528,32.082188,20.613384,16.92582,13.238253,9.550687,5.863121,2.175555,1.84197,1.5101979,1.1766127,0.8448406,0.51306844,0.5747091,0.63816285,0.69980353,0.76325727,0.824898,2.030518,3.2343252,4.439945,5.6455655,6.849373,6.872941,6.8946967,6.9182653,6.9400206,6.9617763,5.6491914,4.3384194,3.0258346,1.7132497,0.40066472,0.8194591,1.2400664,1.6606737,2.079468,2.5000753,1.9996977,1.49932,1.0007553,0.50037766,0.0,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,0.7650702,1.2799516,1.794833,2.3097143,2.8245957,4.615803,6.4051967,8.194591,9.985798,11.775192,14.4692545,17.16513,19.859192,22.555067,25.24913,23.494183,21.739235,19.984287,18.22934,16.474392,16.042906,15.609608,15.1781225,14.744824,14.313339,14.449312,14.587097,14.724882,14.862667,15.000452,14.559902,14.119352,13.680615,13.240066,12.799516,11.526816,10.255929,8.98323,7.71053,6.43783,5.89938,5.3627434,4.8242936,4.2876563,3.7492065,4.273153,4.795286,5.317419,5.8395524,6.3616858,6.530291,6.697084,6.8656893,7.0324817,7.1992745,6.8983226,6.5955577,6.2927933,5.9900284,5.6872635,7.2591023,8.832754,10.4045925,11.978244,13.550082,12.826711,12.105151,11.381779,10.66022,9.936848,8.7421055,7.5473633,6.352621,5.1578784,3.9631362,4.0918565,4.2223897,4.3529234,4.4816437,4.612177,5.3482394,6.0824895,6.816739,7.552802,8.287052,8.1819,8.076748,7.9715962,7.8682575,7.763106,7.8755093,7.987913,8.100317,8.212721,8.325124,8.577126,8.829127,9.082943,9.334945,9.5869465,11.525003,13.46306,15.399304,17.33736,19.275417,19.750414,20.22541,20.700407,21.175404,21.650398,20.19459,18.740595,17.284784,15.83079,14.37498,14.632421,14.889862,15.147303,15.404743,15.662184,15.045776,14.427556,13.809336,13.192928,12.574709,12.650853,12.725184,12.799516,12.87566,12.949992,11.445232,9.940474,8.435715,6.929143,5.424384,5.5567303,5.6908894,5.823236,5.955582,6.0879283,6.1368785,6.187641,6.2384043,6.2873545,6.338117,6.688019,7.037921,7.3878226,7.7377243,8.087626,9.7229185,11.358211,12.99169,14.626982,16.262274,15.352167,14.4420595,13.531953,12.621845,11.711739,11.9329195,12.152288,12.371656,12.592838,12.812206,13.647983,14.481945,15.31772,16.151684,16.98746,17.371807,17.757969,18.142317,18.526665,18.912827,15.852545,12.792264,9.731983,6.6717024,3.6132345,3.975827,4.3366065,4.699199,5.0617914,5.424384,4.604925,3.785466,2.9641938,2.1447346,1.3252757,1.7404441,2.1556125,2.570781,2.9841363,3.3993049,3.6458678,3.8906176,4.135368,4.3801174,4.6248674,4.421816,4.220577,4.017525,3.8144734,3.6132345,3.6404288,3.6676233,3.6948178,3.7220123,3.7492065,3.2397642,2.7303216,2.220879,1.7096237,1.2001812,3.2506418,5.2992897,7.3497505,9.400211,11.450671,10.890467,10.330261,9.770056,9.20985,8.649645,9.804502,10.959359,12.114216,13.270886,14.425743,12.302764,10.179785,8.056806,5.9356394,3.8126602,3.3231604,2.8318477,2.3423476,1.8528478,1.3633479,2.6922495,4.022964,5.351866,6.68258,8.013294,8.760235,9.507175,10.254116,11.00287,11.74981,12.413355,13.075087,13.736817,14.400362,15.062093,13.424988,11.787883,10.150778,8.511859,6.874754,6.1767635,5.480586,4.782595,4.0846047,3.386614,3.9957695,4.603112,5.2104545,5.8177967,6.4251394,5.730775,5.034597,4.3402324,3.6458678,2.94969,2.9750717,3.000453,3.0258346,3.049403,3.0747845,3.6603715,4.2441454,4.8297324,5.4153194,6.000906,4.936697,3.874301,2.811905,1.7495089,0.6871128,2.1683033,3.6476808,5.127058,6.6082487,8.087626,6.510349,4.933071,3.3557937,1.7767034,0.19942589,0.15954071,0.11965553,0.07977036,0.03988518,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.12328146,0.18310922,0.24293698,0.30276474,0.36259252,0.2991388,0.2374981,0.17585737,0.11240368,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,1.4830034,2.9152439,4.347484,5.7797246,7.211965,7.2772317,7.3424983,7.407765,7.473032,7.5382986,7.2917356,7.0469856,6.8022356,6.5574856,6.3127356,6.2130227,6.11331,6.011784,5.9120708,5.812358,5.864934,5.91751,5.9700856,6.0226617,6.0752378,4.972956,3.870675,2.7665808,1.6642996,0.5620184,0.52575916,0.48768693,0.44961473,0.41335547,0.37528324,0.33539808,0.2955129,0.25562772,0.21574254,0.17585737,0.15954071,0.14503701,0.13053331,0.11421664,0.099712946,0.09789998,0.09427405,0.092461094,0.09064813,0.0870222,0.10515183,0.12328146,0.13959812,0.15772775,0.17585737,0.17223145,0.17041849,0.16679256,0.16497959,0.16316663,0.19217403,0.2229944,0.2520018,0.28282216,0.31182957,0.39703882,0.48224804,0.56745726,0.6526665,0.73787576,0.6073425,0.47680917,0.3480888,0.21755551,0.0870222,0.16497959,0.24293698,0.3208944,0.39703882,0.4749962,1.892733,3.3104696,4.7282066,6.14413,7.5618668,6.3707504,5.177821,3.9848917,2.7919624,1.6008459,2.4493124,3.299592,4.1498713,5.0001507,5.8504305,4.7227674,3.5951047,2.467442,1.3397794,0.21211663,0.2229944,0.23205921,0.24293698,0.2520018,0.26287958,1.3307146,2.3967366,3.4645715,4.5324063,5.600241,5.3029156,5.0055895,4.708264,4.409125,4.1117992,3.6295512,3.147303,2.665055,2.182807,1.7005589,1.3633479,1.0243238,0.6871128,0.34990177,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.04169814,0.034446288,0.027194439,0.01994259,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.09064813,0.1794833,0.27013144,0.36077955,0.44961473,1.3252757,2.1991236,3.0747845,3.9504454,4.8242936,5.3228583,5.81961,6.3181744,6.814926,7.311678,7.6797094,8.047741,8.415772,8.781991,9.1500225,7.3497505,5.5494785,3.7492065,1.9507477,0.15047589,0.12328146,0.09427405,0.06707962,0.03988518,0.012690738,0.59283876,1.1729867,1.7531348,2.333283,2.911618,2.7266958,2.5417736,2.3568513,2.1719291,1.987007,2.9243085,3.8616104,4.800725,5.7380266,6.6753283,5.4570174,4.2405195,3.0222087,1.8057107,0.5873999,0.48224804,0.3770962,0.27194437,0.16679256,0.06164073,0.07070554,0.07795739,0.08520924,0.092461094,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.10333887,0.20486477,0.30820364,0.40972954,0.51306844,1.9978848,3.482701,4.9675174,6.452334,7.93715,6.4632115,4.98746,3.5117085,2.03777,0.5620184,0.69255173,0.823085,0.95180535,1.0823387,1.2128719,2.3876717,3.0620937,3.738329,4.4127507,5.087173,5.7615952,6.347182,6.932769,7.518356,8.10213,8.6877165,10.067381,11.447045,12.826711,14.208188,15.5878525,16.084604,16.583168,17.07992,17.576672,18.075237,17.00015,15.925063,14.849977,13.77489,12.699803,12.219368,11.740746,11.26031,10.779876,10.29944,11.876718,13.455809,15.033086,16.610363,18.187641,17.774284,17.362743,16.949387,16.537846,16.124489,28.046532,39.970387,51.89243,63.81447,75.73833,64.01027,52.282215,40.55416,28.827917,17.099863,14.112101,11.124338,8.136576,5.1506267,2.1628644,1.9344311,1.7078108,1.4793775,1.2527572,1.0243238,1.0750868,1.1258497,1.1747998,1.2255627,1.2745126,2.4855716,3.6948178,4.9058766,6.115123,7.324369,6.9073873,6.490406,6.071612,5.65463,5.237649,4.249584,3.2633326,2.275268,1.2872034,0.2991388,0.61459434,0.9300498,1.2455053,1.5591478,1.8746033,1.49932,1.1258497,0.7505665,0.37528324,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.6544795,1.1222239,1.5899682,2.0577126,2.525457,4.117238,5.710832,7.3026133,8.894395,10.487988,12.890164,15.292339,17.694515,20.096691,22.500679,21.25336,20.004229,18.75691,17.509592,16.262274,16.022963,15.781839,15.542528,15.303217,15.062093,14.824595,14.587097,14.349599,14.112101,13.874602,13.544643,13.2146845,12.884725,12.554766,12.224807,10.930351,9.635896,8.339628,7.0451727,5.750717,5.3246713,4.900438,4.4743915,4.0501585,3.6241121,4.082792,4.539658,4.9983377,5.4552045,5.9120708,6.147756,6.3816285,6.6173134,6.8529987,7.0868707,6.7696023,6.452334,6.1350656,5.8177967,5.5005283,6.869315,8.239915,9.610515,10.979301,12.349901,11.804199,11.26031,10.714609,10.17072,9.625018,8.484665,7.344311,6.205771,5.0654173,3.925064,4.1480584,4.36924,4.592234,4.8152285,5.038223,5.5458527,6.051669,6.5592985,7.066928,7.574558,7.476658,7.380571,7.2826705,7.1847706,7.0868707,7.549176,8.013294,8.4756,8.937905,9.400211,9.2044115,9.010424,8.814624,8.620637,8.424837,10.225109,12.025381,13.825653,15.624111,17.424383,18.399757,19.375132,20.350506,21.325878,22.29944,20.589815,18.880192,17.170568,15.459132,13.749508,14.115726,14.480132,14.844538,15.210756,15.575162,14.940624,14.304275,13.669738,13.035201,12.400664,12.661731,12.92461,13.1874895,13.45037,13.713249,12.203052,10.692853,9.182655,7.6724577,6.16226,6.0281005,5.8921285,5.7579694,5.621997,5.487838,5.57486,5.661882,5.750717,5.8377395,5.924762,6.43783,6.9490857,7.462154,7.9752226,8.488291,9.731983,10.9774885,12.222994,13.466686,14.712192,13.8184,12.922797,12.027194,11.13159,10.2378,10.827013,11.418038,12.007251,12.598277,13.1874895,14.545399,15.903308,17.259403,18.617313,19.975222,19.694212,19.415016,19.13582,18.85481,18.575615,16.091856,13.60991,11.127964,8.644206,6.16226,5.8866897,5.612932,5.337362,5.0617914,4.788034,4.360175,3.9323158,3.5044568,3.0765975,2.6505513,2.7430124,2.8354735,2.9279346,3.0203958,3.1128569,3.2270734,3.343103,3.4573197,3.5733492,3.6875658,3.6948178,3.7020695,3.7093215,3.7183862,3.7256382,3.8670492,4.0102735,4.1516843,4.2949085,4.4381323,4.017525,3.5969179,3.1781235,2.7575161,2.3369088,3.587853,4.836984,6.0879283,7.3370595,8.588004,8.167397,7.746789,7.327995,6.9073873,6.48678,7.996978,9.507175,11.017374,12.527572,14.037769,12.067079,10.098202,8.127511,6.156821,4.1879435,3.633177,3.0784104,2.521831,1.9670644,1.4122978,2.4474995,3.482701,4.517903,5.5531044,6.588306,7.783048,8.977791,10.172533,11.367275,12.562017,12.436923,12.311829,12.186734,12.06164,11.938358,10.625773,9.313189,8.000604,6.688019,5.375434,5.041849,4.710077,4.3783045,4.0447197,3.7129474,4.0519714,4.3928084,4.7318325,5.0726695,5.411693,4.7717175,4.1317415,3.491766,2.8517902,2.2118144,2.2371957,2.2625773,2.2879589,2.3133402,2.3369088,3.5080826,4.6774435,5.846804,7.017978,8.187339,6.813113,5.4370747,4.062849,2.6868105,1.3125849,2.2843328,3.2578938,4.229642,5.2032027,6.1749506,4.994712,3.8144734,2.6342347,1.455809,0.2755703,0.21936847,0.16497959,0.11059072,0.054388877,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.18310922,0.30276474,0.4224203,0.5420758,0.66173136,0.53663695,0.41335547,0.28826106,0.16316663,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,1.3017071,2.5671551,3.832603,5.0980506,6.3616858,6.530291,6.697084,6.8656893,7.0324817,7.1992745,7.135821,7.0705543,7.0052876,6.9400206,6.874754,6.825804,6.775041,6.7242785,6.6753283,6.624565,6.604623,6.58468,6.5647373,6.544795,6.5248523,5.4207582,4.314851,3.2107568,2.1048496,1.0007553,0.93730164,0.87566096,0.8122072,0.7505665,0.6871128,0.6073425,0.5275721,0.44780177,0.3680314,0.28826106,0.2574407,0.22662032,0.19761293,0.16679256,0.13778515,0.13234627,0.12690738,0.12328146,0.11784257,0.11240368,0.12328146,0.13234627,0.14322405,0.15228885,0.16316663,0.15772775,0.15228885,0.14684997,0.14322405,0.13778515,0.15954071,0.18310922,0.20486477,0.22662032,0.25018883,0.3208944,0.38978696,0.4604925,0.5293851,0.6000906,0.50219065,0.40429065,0.30820364,0.21030366,0.11240368,0.26831847,0.4224203,0.57833505,0.7324369,0.8883517,1.8474089,2.808279,3.7673361,4.7282066,5.6872635,4.853301,4.017525,3.1817493,2.3477864,1.5120108,2.374981,3.2379513,4.100921,4.9620786,5.825049,4.695573,3.5642843,2.4348087,1.305333,0.17585737,0.20667773,0.23931105,0.27194437,0.3045777,0.33721104,1.1095331,1.8818551,2.6541772,3.4283123,4.2006345,3.9921436,3.785466,3.576975,3.3702974,3.1618068,2.7847104,2.4076142,2.030518,1.651609,1.2745126,1.0243238,0.774135,0.52575916,0.2755703,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.099712946,0.099712946,0.099712946,0.099712946,0.099712946,0.08520924,0.07070554,0.054388877,0.03988518,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.06707962,0.13415924,0.2030518,0.27013144,0.33721104,1.0877775,1.8383441,2.5870976,3.3376641,4.0882306,4.3946214,4.702825,5.009216,5.317419,5.6256227,5.9845896,6.345369,6.7043357,7.065115,7.424082,5.999093,4.5759177,3.149116,1.7259403,0.2991388,0.24474995,0.19036107,0.13415924,0.07977036,0.025381476,0.48587397,0.9445535,1.405046,1.8655385,2.324218,2.3296568,2.335096,2.3405347,2.3441606,2.3495996,3.0367124,3.7256382,4.4127507,5.0998635,5.7869763,4.802538,3.8180993,2.8318477,1.8474089,0.8629702,0.7016165,0.5420758,0.3825351,0.2229944,0.06164073,0.065266654,0.06707962,0.07070554,0.072518505,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.092461094,0.18492219,0.27738327,0.36984438,0.46230546,1.5700256,2.6777458,3.785466,4.893186,5.999093,4.8877473,3.774588,2.663242,1.550083,0.43692398,0.5475147,0.65810543,0.7668832,0.8774739,0.9880646,2.3622901,2.9750717,3.587853,4.2006345,4.8134155,5.424384,5.9392653,6.454147,6.970841,7.4857225,8.000604,9.256987,10.515183,11.773379,13.029762,14.287958,14.976884,15.667623,16.358362,17.047287,17.738026,16.624866,15.511708,14.400362,13.287203,12.175857,12.092461,12.010877,11.927481,11.845898,11.762501,13.234627,14.706753,16.18069,17.652817,19.124943,19.311678,19.500225,19.68696,19.87551,20.062244,30.75147,41.442513,52.133553,62.82278,73.51201,61.528324,49.542828,37.55733,25.571836,13.588155,11.300196,9.012237,6.7242785,4.4381323,2.1501737,2.0268922,1.9054236,1.7821422,1.6606737,1.5373923,1.5754645,1.6117238,1.649796,1.6878681,1.7241274,2.9406252,4.15531,5.369995,6.58468,7.799365,6.9418335,6.0843024,5.2267714,4.36924,3.5117085,2.8499773,2.1882458,1.5247015,0.8629702,0.19942589,0.40972954,0.6200332,0.83033687,1.0406405,1.2491312,1.0007553,0.7505665,0.50037766,0.25018883,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.54570174,0.9644961,1.3851035,1.8057107,2.2245052,3.6204863,5.0146546,6.4106355,7.804804,9.200785,11.30926,13.419549,15.529838,17.640125,19.750414,19.010725,18.269224,17.529535,16.789846,16.050158,16.003021,15.955884,15.906934,15.859797,15.812659,15.199879,14.587097,13.974316,13.363347,12.750566,12.529385,12.310016,12.090648,11.869466,11.650098,10.332074,9.015862,7.6978393,6.379815,5.0617914,4.749962,4.4381323,4.12449,3.8126602,3.5008307,3.8924308,4.2858434,4.6774435,5.0708566,5.462456,5.765221,6.0679855,6.3707504,6.6717024,6.9744673,6.642695,6.3091097,5.977338,5.6455655,5.3119802,6.4795284,7.647076,8.814624,9.982172,11.14972,10.781689,10.41547,10.047439,9.679407,9.313189,8.227224,7.1430726,6.057108,4.972956,3.8869917,4.2024474,4.517903,4.8333583,5.147001,5.462456,5.7416525,6.0226617,6.301858,6.582867,6.8620634,6.773228,6.68258,6.591932,6.5030966,6.412449,7.224656,8.036863,8.8508835,9.663091,10.475298,9.8316965,9.189907,8.548119,7.9045167,7.262728,8.925215,10.587702,12.250188,13.912675,15.575162,17.0491,18.52485,20.000603,21.474543,22.950293,20.985043,19.01979,17.054539,15.089288,13.125849,13.597219,14.070402,14.541773,15.014956,15.488139,14.835473,14.182806,13.53014,12.877473,12.224807,12.674421,13.125849,13.575464,14.025079,14.474693,12.96087,11.445232,9.929596,8.415772,6.9001355,6.497658,6.09518,5.6927023,5.290225,4.8877473,5.0128417,5.137936,5.2630305,5.388125,5.5132194,6.187641,6.8620634,7.5382986,8.212721,8.887142,9.742861,10.596766,11.452485,12.308203,13.162108,12.282822,11.401722,10.522435,9.643148,8.762048,9.7229185,10.681975,11.642846,12.601903,13.562773,15.442815,17.322857,19.2029,21.082941,22.962984,22.016617,21.072063,20.12751,19.182957,18.238403,16.33298,14.427556,12.522133,10.616709,8.713099,7.799365,6.887445,5.975525,5.0617914,4.1498713,4.115425,4.079166,4.0447197,4.0102735,3.975827,3.7455807,3.5153344,3.2850883,3.054842,2.8245957,2.810092,2.7955883,2.7792716,2.764768,2.7502642,2.9678197,3.1853752,3.4029307,3.6204863,3.8380418,4.0954823,4.3529234,4.610364,4.8678045,5.125245,4.795286,4.465327,4.135368,3.8054085,3.4754493,3.925064,4.3746786,4.8242936,5.275721,5.7253356,5.4443264,5.1651306,4.8841214,4.604925,4.325729,6.189454,8.054993,9.920531,11.784257,13.649796,11.833207,10.014805,8.198216,6.379815,4.5632267,3.9431937,3.3231604,2.7031271,2.0830941,1.4630609,2.2027495,2.9424384,3.682127,4.421816,5.163317,6.8058615,8.446592,10.09095,11.731681,13.374225,12.462305,11.5503845,10.636651,9.724731,8.812811,7.8247466,6.836682,5.8504305,4.8623657,3.874301,3.9069343,3.9395678,3.972201,4.004834,4.0374675,4.1099863,4.1825047,4.255023,4.327542,4.40006,3.8144734,3.2306993,2.6451125,2.0595255,1.4757515,1.49932,1.5247015,1.550083,1.5754645,1.6008459,3.3557937,5.1107416,6.8656893,8.620637,10.375585,8.6877165,6.9998484,5.3119802,3.6241121,1.938057,2.4021754,2.8681068,3.3322253,3.7981565,4.262275,3.4790752,2.6976883,1.9144884,1.1331016,0.34990177,0.27919623,0.21030366,0.13959812,0.07070554,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.24293698,0.4224203,0.60190356,0.78319985,0.96268314,0.774135,0.5873999,0.40066472,0.21211663,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,1.1222239,2.2190661,3.3177216,4.4145637,5.5132194,5.7833505,6.051669,6.3218007,6.591932,6.8620634,6.978093,7.0923095,7.208339,7.322556,7.4367723,7.4367723,7.4367723,7.4367723,7.4367723,7.4367723,7.344311,7.25185,7.159389,7.066928,6.9744673,5.866747,4.76084,3.6531196,2.5453994,1.4376793,1.3506571,1.261822,1.1747998,1.0877775,1.0007553,0.8792868,0.75963134,0.6399758,0.52032024,0.40066472,0.35534066,0.3100166,0.26469254,0.21936847,0.17585737,0.16679256,0.15954071,0.15228885,0.14503701,0.13778515,0.13959812,0.14322405,0.14503701,0.14684997,0.15047589,0.14322405,0.13415924,0.12690738,0.11965553,0.11240368,0.12690738,0.14322405,0.15772775,0.17223145,0.18673515,0.24293698,0.29732585,0.35171473,0.40791658,0.46230546,0.39703882,0.33177215,0.26831847,0.2030518,0.13778515,0.36984438,0.60190356,0.83577573,1.067835,1.2998942,1.8020848,2.3042755,2.808279,3.3104696,3.8126602,3.3358512,2.857229,2.38042,1.9017978,1.4249886,2.3006494,3.1744974,4.0501585,4.9258194,5.7996674,4.666566,3.5352771,2.4021754,1.2708868,0.13778515,0.19217403,0.24837588,0.30276474,0.35715362,0.41335547,0.8901646,1.3669738,1.845596,2.322405,2.7992141,2.6831846,2.565342,2.4474995,2.3296568,2.2118144,1.93987,1.6679256,1.3941683,1.1222239,0.85027945,0.6871128,0.52575916,0.36259252,0.19942589,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.15047589,0.15047589,0.15047589,0.15047589,0.15047589,0.12690738,0.10515183,0.08339628,0.059827764,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.045324065,0.09064813,0.13415924,0.1794833,0.22480737,0.85027945,1.4757515,2.0994108,2.7248828,3.350355,3.4681973,3.584227,3.7020695,3.8199122,3.9377546,4.2894692,4.6429973,4.994712,5.3482394,5.6999545,4.650249,3.6005437,2.5508385,1.49932,0.44961473,0.3680314,0.28463513,0.2030518,0.11965553,0.038072214,0.3770962,0.7179332,1.0569572,1.3977941,1.7368182,1.9326181,2.126605,2.322405,2.518205,2.712192,3.150929,3.587853,4.024777,4.461701,4.900438,4.1480584,3.395679,2.6432993,1.8909199,1.1367276,0.922798,0.7070554,0.49312583,0.27738327,0.06164073,0.059827764,0.058014803,0.054388877,0.052575916,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08339628,0.16497959,0.24837588,0.32995918,0.41335547,1.1421664,1.8727903,2.6034143,3.3322253,4.062849,3.3122826,2.561716,1.8129625,1.062396,0.31182957,0.40247768,0.49312583,0.581961,0.6726091,0.76325727,2.3369088,2.8880494,3.437377,3.9867048,4.537845,5.087173,5.5331616,5.977338,6.4233265,6.867502,7.311678,8.446592,9.583321,10.718235,11.853149,12.988064,13.8691635,14.752076,15.63499,16.517902,17.400814,16.249584,15.100165,13.9507475,12.799516,11.650098,11.965553,12.279196,12.594651,12.910107,13.225562,14.592536,15.95951,17.328297,18.69527,20.062244,20.850883,21.637709,22.424534,23.213173,23.999998,33.458225,42.91464,52.372864,61.829277,71.2875,59.044567,46.803444,34.558693,22.31757,10.074633,8.488291,6.9001355,5.3119802,3.7256382,2.137483,2.1193533,2.1030366,2.084907,2.0667772,2.0504606,2.0758421,2.0994108,2.124792,2.1501737,2.175555,3.395679,4.615803,5.8359265,7.0542374,8.274362,6.978093,5.6800117,4.3819304,3.0856624,1.7875811,1.4503701,1.1131591,0.774135,0.43692398,0.099712946,0.20486477,0.3100166,0.41516843,0.52032024,0.62547207,0.50037766,0.37528324,0.25018883,0.12509441,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.43511102,0.80676836,1.1802386,1.551896,1.9253663,3.1219215,4.3202896,5.516845,6.7152133,7.911769,9.73017,11.546759,13.36516,15.181748,17.00015,16.768091,16.534218,16.30216,16.0701,15.838041,15.983078,16.128115,16.273151,16.41819,16.563227,15.575162,14.587097,13.600845,12.612781,11.624716,11.514126,11.405348,11.294757,11.184166,11.075388,9.735609,8.39583,7.0542374,5.714458,4.3746786,4.175253,3.975827,3.774588,3.5751622,3.3757362,3.7020695,4.0302157,4.358362,4.6846952,5.0128417,5.382686,5.75253,6.1223745,6.492219,6.8620634,6.5157876,6.167699,5.81961,5.473334,5.125245,6.089741,7.0542374,8.020547,8.985043,9.949538,9.759177,9.570629,9.380268,9.189907,8.999546,7.9697833,6.9400206,5.910258,4.880495,3.8507326,4.256836,4.664753,5.0726695,5.480586,5.8866897,5.9392653,5.9918413,6.0444174,6.096993,6.149569,6.0679855,5.9845896,5.903006,5.81961,5.7380266,6.9001355,8.062244,9.224354,10.388275,11.5503845,10.460794,9.3693905,8.2798,7.1902094,6.1006193,7.6253204,9.1500225,10.674724,12.199425,13.724127,15.700256,17.674572,19.650702,21.625017,23.599335,21.380268,19.15939,16.940323,14.719443,12.500377,13.080525,13.660673,14.240821,14.819156,15.399304,14.730321,14.059525,13.390542,12.719746,12.050762,12.687112,13.325275,13.961625,14.599788,15.23795,13.716875,12.197612,10.6783495,9.157274,7.6380115,6.967215,6.298232,5.6274357,4.95664,4.2876563,4.4508233,4.612177,4.7753434,4.936697,5.0998635,5.9374523,6.775041,7.61263,8.450218,9.287807,9.751925,10.217857,10.681975,11.147907,11.612025,10.747242,9.882459,9.017676,8.152893,7.28811,8.617011,9.947725,11.27844,12.607342,13.938056,16.34023,18.742407,21.144583,23.546759,25.950747,24.340836,22.730925,21.119202,19.50929,17.89938,16.57229,15.245202,13.918114,12.589212,11.262123,9.712041,8.161958,6.6118746,5.0617914,3.5117085,3.870675,4.227829,4.5849824,4.942136,5.2992897,4.748149,4.195195,3.6422417,3.0892882,2.5381477,2.3931105,2.2480736,2.1030366,1.9579996,1.8129625,2.2408218,2.666868,3.094727,3.5225863,3.9504454,4.322103,4.695573,5.06723,5.4407005,5.812358,5.573047,5.331923,5.092612,4.853301,4.612177,4.262275,3.9123733,3.5624714,3.2125697,2.8626678,2.72307,2.5816586,2.4420607,2.3024626,2.1628644,4.3819304,6.60281,8.821876,11.042755,13.261822,11.597522,9.933222,8.267109,6.60281,4.936697,4.25321,3.5679104,2.8826106,2.1973107,1.5120108,1.9579996,2.4021754,2.8481643,3.29234,3.738329,5.826862,7.9172077,10.007553,12.097899,14.188245,12.487686,10.7871275,9.086569,7.3878226,5.6872635,5.0255322,4.361988,3.7002566,3.0367124,2.374981,2.7720199,3.1708715,3.5679104,3.9649491,4.361988,4.168001,3.972201,3.778214,3.5824142,3.386614,2.857229,2.327844,1.7966459,1.2672608,0.73787576,0.76325727,0.7868258,0.8122072,0.8375887,0.8629702,3.2035048,5.542227,7.8827615,10.223296,12.562017,10.56232,8.562622,6.5629244,4.5632267,2.561716,2.520018,2.47832,2.4348087,2.3931105,2.3495996,1.9652514,1.5790904,1.1947423,0.8103943,0.42423326,0.34083697,0.25562772,0.17041849,0.08520924,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.30276474,0.5420758,0.78319985,1.0225109,1.261822,1.0116332,0.76325727,0.51306844,0.26287958,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.94274056,1.8727903,2.8028402,3.73289,4.6629395,5.034597,5.408067,5.7797246,6.153195,6.5248523,6.8203654,7.115878,7.409578,7.705091,8.000604,8.049554,8.100317,8.149267,8.200029,8.2507925,8.0858135,7.9208336,7.755854,7.590874,7.4258947,6.3145485,5.2050157,4.0954823,2.9841363,1.8746033,1.7621996,1.649796,1.5373923,1.4249886,1.3125849,1.1530442,0.9916905,0.8321498,0.6726091,0.51306844,0.45324063,0.39159992,0.33177215,0.27194437,0.21211663,0.2030518,0.19217403,0.18310922,0.17223145,0.16316663,0.15772775,0.15228885,0.14684997,0.14322405,0.13778515,0.12690738,0.11784257,0.10696479,0.09789998,0.0870222,0.09427405,0.10333887,0.11059072,0.11784257,0.12509441,0.16497959,0.20486477,0.24474995,0.28463513,0.3245203,0.291887,0.25925365,0.22662032,0.19579996,0.16316663,0.47318324,0.78319985,1.0932164,1.403233,1.7132497,1.7567607,1.8020848,1.8474089,1.892733,1.938057,1.8165885,1.696933,1.5772774,1.4576219,1.3379664,2.2245052,3.1128569,3.9993954,4.8877473,5.774286,4.6393714,3.5044568,2.3695421,1.2346275,0.099712946,0.17767033,0.25562772,0.33177215,0.40972954,0.48768693,0.67079616,0.8520924,1.0352017,1.2183108,1.3996071,1.3724127,1.3452182,1.3180238,1.2908293,1.261822,1.0950294,0.92823684,0.75963134,0.59283876,0.42423326,0.34990177,0.2755703,0.19942589,0.12509441,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.03988518,0.07977036,0.11965553,0.15954071,0.19942589,0.19942589,0.19942589,0.19942589,0.19942589,0.19942589,0.17041849,0.13959812,0.11059072,0.07977036,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.61278135,1.1131591,1.6117238,2.1121013,2.612479,2.5399606,2.467442,2.3949237,2.322405,2.2498865,2.5943494,2.9406252,3.2850883,3.6295512,3.975827,3.299592,2.6251698,1.9507477,1.2745126,0.6000906,0.4894999,0.38072214,0.27013144,0.15954071,0.05076295,0.27013144,0.4894999,0.7106813,0.9300498,1.1494182,1.5355793,1.9199274,2.3042755,2.6904364,3.0747845,3.2633326,3.4500678,3.636803,3.825351,4.0120864,3.491766,2.9732587,2.4529383,1.9326181,1.4122978,1.1421664,0.872035,0.60190356,0.33177215,0.06164073,0.054388877,0.047137026,0.03988518,0.032633327,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.072518505,0.14503701,0.21755551,0.29007402,0.36259252,0.71430725,1.067835,1.4195497,1.7730774,2.124792,1.7368182,1.3506571,0.96268314,0.5747091,0.18673515,0.2574407,0.32814622,0.39703882,0.46774435,0.53663695,2.3133402,2.7992141,3.2869012,3.774588,4.262275,4.749962,5.125245,5.5005283,5.8758116,6.249282,6.624565,7.6380115,8.649645,9.663091,10.674724,11.6881695,12.763257,13.838344,14.91343,15.986704,17.06179,15.8743,14.68681,13.499319,12.311829,11.124338,11.836833,12.549327,13.261822,13.974316,14.68681,15.950445,17.212267,18.475903,19.737724,20.999546,22.388275,23.77519,25.162107,26.550837,27.937754,36.163166,44.386765,52.612175,60.837585,69.062996,56.56262,44.062244,31.561865,19.06149,6.5629244,5.674573,4.788034,3.8996825,3.0131438,2.124792,2.2118144,2.3006494,2.3876717,2.474694,2.561716,2.5744069,2.5870976,2.5997884,2.612479,2.6251698,3.8507326,5.0744824,6.300045,7.5256076,8.749357,7.0125394,5.275721,3.53709,1.8002719,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.3245203,0.6508536,0.97537386,1.2998942,1.6244144,2.6251698,3.6241121,4.6248674,5.6256227,6.624565,8.149267,9.675781,11.200482,12.725184,14.249886,14.525456,14.799213,15.074784,15.350354,15.624111,15.963136,16.300346,16.637558,16.97477,17.31198,15.950445,14.587097,13.225562,11.862214,10.500679,10.500679,10.500679,10.500679,10.500679,10.500679,9.137331,7.7757964,6.412449,5.049101,3.6875658,3.6005437,3.5117085,3.4246864,3.3376641,3.2506418,3.5117085,3.774588,4.0374675,4.3003473,4.5632267,5.0001507,5.4370747,5.8758116,6.3127356,6.7496595,6.3870673,6.0244746,5.661882,5.2992897,4.936697,5.6999545,6.4632115,7.224656,7.987913,8.749357,8.736667,8.725789,8.713099,8.700407,8.6877165,7.7123427,6.736969,5.7615952,4.788034,3.8126602,4.313038,4.8116026,5.3119802,5.812358,6.3127356,6.1368785,5.962834,5.7869763,5.612932,5.4370747,5.3627434,5.2865987,5.2122674,5.137936,5.0617914,6.5756154,8.087626,9.599637,11.111648,12.625471,11.088079,9.550687,8.013294,6.474089,4.936697,6.3254266,7.7123427,9.099259,10.487988,11.874905,14.349599,16.824293,19.3008,21.775494,24.250187,21.775494,19.3008,16.824293,14.349599,11.874905,12.562017,13.24913,13.938056,14.625169,15.312282,14.625169,13.938056,13.24913,12.562017,11.874905,12.699803,13.524701,14.349599,15.174497,15.999394,14.474693,12.949992,11.42529,9.900589,8.375887,7.4367723,6.4994707,5.562169,4.6248674,3.6875658,3.8869917,4.0882306,4.2876563,4.4870825,4.688321,5.6872635,6.688019,7.686961,8.6877165,9.686659,9.762803,9.837135,9.91328,9.987611,10.061942,9.211663,8.363196,7.512917,6.6626377,5.812358,7.512917,9.211663,10.912222,12.612781,14.313339,17.237648,20.161957,23.088078,26.012386,28.936695,26.66324,24.387972,22.112705,19.837437,17.562168,16.813416,16.062849,15.312282,14.561715,13.812962,11.624716,9.438283,7.250037,5.0617914,2.8753586,3.6241121,4.3746786,5.125245,5.8758116,6.624565,5.750717,4.8750563,3.9993954,3.1255474,2.2498865,1.9743162,1.7005589,1.4249886,1.1494182,0.87566096,1.5120108,2.1501737,2.7883365,3.4246864,4.062849,4.550536,5.038223,5.52591,6.011784,6.4994707,6.350808,6.200332,6.049856,5.89938,5.750717,4.599486,3.4500678,2.3006494,1.1494182,0.0,0.0,0.0,0.0,0.0,0.0,2.5744069,5.1506267,7.7250338,10.29944,12.87566,11.361836,9.849826,8.337815,6.825804,5.3119802,4.5632267,3.8126602,3.0620937,2.3133402,1.5627737,1.7132497,1.8619126,2.0123885,2.1628644,2.3133402,4.8496747,7.3878226,9.92597,12.462305,15.000452,12.513068,10.025683,7.5382986,5.049101,2.561716,2.2245052,1.887294,1.550083,1.2128719,0.87566096,1.6371052,2.4003625,3.1618068,3.925064,4.688321,4.2242026,3.7618973,3.299592,2.8372865,2.374981,1.8999848,1.4249886,0.9499924,0.4749962,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,3.049403,5.975525,8.899834,11.8241415,14.750263,12.436923,10.125396,7.8120556,5.5005283,3.1871881,2.6378605,2.08672,1.5373923,0.9880646,0.43692398,0.44961473,0.46230546,0.4749962,0.48768693,0.50037766,0.40066472,0.2991388,0.19942589,0.099712946,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.36259252,0.66173136,0.96268314,1.261822,1.5627737,1.2491312,0.93730164,0.62547207,0.31182957,0.0,0.0,0.0,0.0,0.0,0.0,0.76325727,1.5247015,2.2879589,3.049403,3.8126602,4.2876563,4.762653,5.237649,5.712645,6.187641,6.6626377,7.137634,7.61263,8.087626,8.562622,8.662335,8.762048,8.861761,8.963287,9.063,8.825501,8.588004,8.350506,8.113008,7.8755093,6.7623506,5.6491914,4.537845,3.4246864,2.3133402,2.175555,2.03777,1.8999848,1.7621996,1.6244144,1.4249886,1.2255627,1.0243238,0.824898,0.62547207,0.5493277,0.4749962,0.40066472,0.3245203,0.25018883,0.2374981,0.22480737,0.21211663,0.19942589,0.18673515,0.17585737,0.16316663,0.15047589,0.13778515,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.0870222,0.11240368,0.13778515,0.16316663,0.18673515,0.18673515,0.18673515,0.18673515,0.18673515,0.18673515,0.5747091,0.96268314,1.3506571,1.7368182,2.124792,1.7132497,1.2998942,0.8883517,0.4749962,0.06164073,0.2991388,0.53663695,0.774135,1.0116332,1.2491312,2.1501737,3.049403,3.9504454,4.8496747,5.750717,4.612177,3.4754493,2.3369088,1.2001812,0.06164073,0.16316663,0.26287958,0.36259252,0.46230546,0.5620184,0.44961473,0.33721104,0.22480737,0.11240368,0.0,0.06164073,0.12509441,0.18673515,0.25018883,0.31182957,0.25018883,0.18673515,0.12509441,0.06164073,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,0.25018883,0.25018883,0.25018883,0.25018883,0.25018883,0.21211663,0.17585737,0.13778515,0.099712946,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.37528324,0.7505665,1.1258497,1.49932,1.8746033,1.6117238,1.3506571,1.0877775,0.824898,0.5620184,0.89922947,1.2382535,1.5754645,1.9126755,2.2498865,1.9507477,1.649796,1.3506571,1.0497054,0.7505665,0.61278135,0.4749962,0.33721104,0.19942589,0.06164073,0.16316663,0.26287958,0.36259252,0.46230546,0.5620184,1.1367276,1.7132497,2.2879589,2.8626678,3.437377,3.3757362,3.3122826,3.2506418,3.1871881,3.1255474,2.8372865,2.5508385,2.2625773,1.9743162,1.6878681,1.3633479,1.0370146,0.7124943,0.387974,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06164073,0.12509441,0.18673515,0.25018883,0.31182957,0.28826106,0.26287958,0.2374981,0.21211663,0.18673515,0.16316663,0.13778515,0.11240368,0.0870222,0.06164073,0.11240368,0.16316663,0.21211663,0.26287958,0.31182957,2.2625773,2.6849976,3.1074178,3.529838,3.9522583,4.3746786,4.652062,4.9294453,5.2068286,5.484212,5.7615952,6.892884,8.02236,9.151835,10.283124,11.4126,12.467744,13.522888,14.5780325,15.633177,16.68832,15.798156,14.907991,14.017827,13.127662,12.237497,12.971747,13.70781,14.4420595,15.1781225,15.912373,16.887747,17.863121,18.836681,19.812056,20.78743,22.9231,25.056955,27.192625,29.328295,31.462152,37.18749,42.912823,48.63816,54.361683,60.087017,49.214684,38.342346,27.470009,16.597672,5.7253356,5.179634,4.6357455,4.0900435,3.5443418,3.000453,2.9279346,2.855416,2.7828975,2.7103791,2.6378605,2.5399606,2.4420607,2.3441606,2.2480736,2.1501737,3.1273603,4.1045475,5.081734,6.060734,7.037921,5.6401267,4.2423325,2.8445382,1.4467441,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.11421664,0.16679256,0.21936847,0.27194437,0.3245203,0.52032024,0.71430725,0.9101072,1.1059072,1.2998942,2.4819458,3.6658103,4.847862,6.0299134,7.211965,8.455658,9.697536,10.939416,12.183108,13.424988,13.8147745,14.204562,14.594349,14.984136,15.375735,15.616859,15.859797,16.102734,16.34567,16.586794,15.410182,14.231756,13.055143,11.876718,10.700105,10.667472,10.634838,10.602205,10.5695715,10.536939,9.267865,7.996978,6.7279043,5.4570174,4.1879435,4.1498713,4.1117992,4.07554,4.0374675,3.9993954,4.4145637,4.8297324,5.2449007,5.660069,6.0752378,6.4033837,6.7297173,7.057863,7.3841968,7.7123427,7.311678,6.9128265,6.5121617,6.11331,5.712645,6.5030966,7.2917356,8.082188,8.872639,9.663091,9.452786,9.242483,9.03218,8.821876,8.613385,7.652515,6.6916447,5.732588,4.7717175,3.8126602,4.122677,4.4326935,4.74271,5.0527267,5.3627434,5.2503395,5.137936,5.0255322,4.9131284,4.800725,4.7680917,4.7354584,4.702825,4.670192,4.6375585,6.169512,7.703278,9.235231,10.767185,12.299138,10.999244,9.699349,8.399456,7.0995617,5.7996674,7.2971745,8.794682,10.292189,11.789696,13.287203,15.384801,17.482399,19.579996,21.677593,23.77519,21.44916,19.124943,16.800724,14.474693,12.1504755,12.685299,13.220123,13.754947,14.289771,14.824595,14.097597,13.370599,12.6417885,11.91479,11.187792,12.027194,12.866595,13.70781,14.547212,15.386614,14.010575,12.632723,11.254871,9.87702,8.499168,7.5219817,6.544795,5.567608,4.590421,3.6132345,3.8525455,4.0918565,4.3329806,4.572292,4.8116026,5.65463,6.497658,7.3406854,8.1819,9.024928,9.077503,9.130079,9.182655,9.235231,9.287807,8.685904,8.082188,7.4802837,6.87838,6.2746634,7.7395372,9.2044115,10.669285,12.134158,13.600845,16.458075,19.315304,22.172533,25.029762,27.88699,25.740442,23.592083,21.445534,19.297174,17.150625,16.642996,16.135366,15.627737,15.120108,14.612478,12.264692,9.916905,7.569119,5.223145,2.8753586,3.7492065,4.6248674,5.5005283,6.3743763,7.250037,6.205771,5.1596913,4.115425,3.0693457,2.0250793,1.7730774,1.5192627,1.2672608,1.015259,0.76325727,1.4358664,2.1066625,2.7792716,3.4518807,4.12449,4.8297324,5.5349746,6.240217,6.94546,7.650702,7.0524244,6.454147,5.857682,5.2594047,4.6629395,4.572292,4.4816437,4.3928084,4.3021603,4.213325,3.6531196,3.092914,2.5327086,1.9725033,1.4122978,3.4573197,5.5023413,7.5473633,9.592385,11.637406,10.277685,8.917963,7.558241,6.1967063,4.836984,4.655688,4.4725785,4.2894692,4.1081734,3.925064,3.8597972,3.7945306,3.729264,3.6658103,3.6005437,6.472276,9.345822,12.217555,15.089288,17.962833,15.227073,12.493125,9.757364,7.021604,4.2876563,3.8869917,3.48814,3.0874753,2.6868105,2.2879589,5.565795,8.841819,12.119655,15.397491,18.675327,15.386614,12.099712,8.812811,5.524097,2.2371957,3.6676233,5.0980506,6.526665,7.957093,9.38752,7.6216946,5.857682,4.0918565,2.327844,0.5620184,2.810092,5.0581656,7.304426,9.5525,11.800573,11.352772,10.90497,10.457169,10.009366,9.563377,7.7195945,5.8776245,4.0356545,2.1918716,0.34990177,0.37165734,0.39522585,0.4169814,0.4405499,0.46230546,0.36984438,0.27738327,0.18492219,0.092461094,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.291887,0.53482395,0.7777609,1.020698,1.261822,1.0098201,0.75781834,0.5058166,0.2520018,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.81583315,1.5301404,2.2444477,2.960568,3.6748753,4.0846047,4.494334,4.9058766,5.315606,5.7253356,6.4233265,7.119504,7.817495,8.515485,9.211663,8.917963,8.62245,8.326937,8.033237,7.7377243,7.8301854,7.9226465,8.015107,8.107569,8.200029,7.2482243,6.294606,5.3428006,4.3891826,3.437377,3.1255474,2.811905,2.5000753,2.1882458,1.8746033,1.647983,1.4195497,1.1929294,0.9644961,0.73787576,0.6345369,0.533011,0.42967212,0.32814622,0.22480737,0.21574254,0.20486477,0.19579996,0.18492219,0.17585737,0.16497959,0.15410182,0.14503701,0.13415924,0.12509441,0.11059072,0.09427405,0.07977036,0.065266654,0.05076295,0.07070554,0.09064813,0.11059072,0.13053331,0.15047589,0.3825351,0.61459434,0.8466535,1.0805258,1.3125849,1.0805258,0.8466535,0.61459434,0.3825351,0.15047589,0.47318324,0.79589057,1.1167849,1.4394923,1.7621996,1.4304274,1.0968424,0.7650702,0.43329805,0.099712946,0.46955732,0.83940166,1.209246,1.5809034,1.9507477,2.617918,3.2850883,3.9522583,4.6194286,5.2865987,4.360175,3.4319382,2.5055144,1.5772774,0.6508536,0.6653573,0.67986095,0.69436467,0.7106813,0.72518504,0.5873999,0.44961473,0.31182957,0.17585737,0.038072214,0.07977036,0.12328146,0.16497959,0.20667773,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.052575916,0.04169814,0.032633327,0.02175555,0.012690738,0.058014803,0.10333887,0.14684997,0.19217403,0.2374981,0.24837588,0.2574407,0.26831847,0.27738327,0.28826106,0.25562772,0.2229944,0.19036107,0.15772775,0.12509441,0.10515183,0.08520924,0.065266654,0.045324065,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.2991388,0.6000906,0.89922947,1.2001812,1.49932,1.2926424,1.0841516,0.8774739,0.67079616,0.46230546,0.8520924,1.2418793,1.6316663,2.0232663,2.4130533,2.5907235,2.7683938,2.9442513,3.1219215,3.299592,2.8953013,2.4891977,2.084907,1.6806163,1.2745126,1.1874905,1.1004683,1.0116332,0.9246109,0.8375887,1.2291887,1.6226015,2.0142014,2.4076142,2.7992141,2.9297476,3.0602808,3.1908143,3.3195345,3.4500678,3.73289,4.0157123,4.2967215,4.5795436,4.8623657,4.0555973,3.247016,2.4402475,1.6316663,0.824898,0.66173136,0.50037766,0.33721104,0.17585737,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.052575916,0.10515183,0.15772775,0.21030366,0.26287958,0.23931105,0.21755551,0.19579996,0.17223145,0.15047589,0.16679256,0.18492219,0.2030518,0.21936847,0.2374981,0.533011,0.82671094,1.1222239,1.4177368,1.7132497,2.2118144,2.570781,2.9279346,3.2850883,3.6422417,3.9993954,4.1806917,4.360175,4.539658,4.7191415,4.900438,6.147756,7.3950744,8.642392,9.88971,11.137029,12.172231,13.207433,14.242634,15.277836,16.313038,15.720199,15.127359,14.534521,13.941682,13.3506565,14.106662,14.86448,15.622298,16.380117,17.137936,17.825048,18.512161,19.199274,19.888199,20.575312,23.457922,26.340534,29.223145,32.105755,34.988365,38.21181,41.437073,44.662334,47.887592,51.112854,41.866745,32.622448,23.376339,14.132043,4.8877473,4.6846952,4.4816437,4.2804046,4.077353,3.874301,3.6422417,3.4101827,3.1781235,2.9442513,2.712192,2.5055144,2.2970235,2.0903459,1.8818551,1.6751775,2.4058013,3.1346123,3.8652363,4.59586,5.3246713,4.267714,3.2107568,2.1519866,1.0950294,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.23024625,0.33539808,0.4405499,0.54570174,0.6508536,0.71430725,0.7795739,0.8448406,0.9101072,0.97537386,2.3405347,3.7056956,5.0708566,6.434204,7.799365,8.760235,9.719293,10.680162,11.63922,12.60009,13.104094,13.60991,14.115726,14.61973,15.125546,15.272397,15.419247,15.567909,15.71476,15.861609,14.869919,13.878228,12.884725,11.893035,10.899531,10.834265,10.770811,10.705544,10.640278,10.57501,9.398398,8.219973,7.0433598,5.864934,4.688321,4.699199,4.7118897,4.7245803,4.7372713,4.749962,5.317419,5.8848767,6.452334,7.019791,7.5872483,7.804804,8.02236,8.239915,8.457471,8.675026,8.238102,7.799365,7.362441,6.925517,6.48678,7.304426,8.122072,8.939718,9.757364,10.57501,10.167094,9.759177,9.353074,8.945157,8.537241,7.592687,6.6481338,5.7017674,4.7572136,3.8126602,3.9323158,4.0519714,4.171627,4.2930956,4.4127507,4.361988,4.313038,4.262275,4.213325,4.162562,4.171627,4.1825047,4.1933823,4.2024474,4.213325,5.765221,7.317117,8.870826,10.422722,11.974618,10.912222,9.849826,8.78743,7.7250338,6.6626377,8.270736,9.87702,11.485118,13.093216,14.699501,16.420002,18.140503,19.859192,21.579693,23.300196,21.12464,18.950897,16.775343,14.599788,12.4242325,12.806767,13.189302,13.571837,13.954373,14.336908,13.5700245,12.803142,12.034446,11.267563,10.500679,11.354585,12.210303,13.064208,13.919927,14.775645,13.544643,12.3154545,11.084454,9.855265,8.624263,7.607191,6.590119,5.573047,4.554162,3.53709,3.8180993,4.0972953,4.3783045,4.6575007,4.936697,5.621997,6.3072968,6.9925966,7.6778965,8.363196,8.392203,8.423024,8.452031,8.482852,8.511859,8.158332,7.802991,7.4476504,7.0923095,6.736969,7.9679704,9.197159,10.428161,11.65735,12.888351,15.676687,18.466837,21.256987,24.047136,26.837286,24.817644,22.798004,20.77655,18.75691,16.73727,16.472578,16.207886,15.9431925,15.676687,15.411995,12.904668,10.397341,7.890013,5.382686,2.8753586,3.874301,4.8750563,5.8758116,6.874754,7.8755093,6.6608243,5.4443264,4.229642,3.0149567,1.8002719,1.5700256,1.3397794,1.1095331,0.8792868,0.6508536,1.357909,2.0649643,2.7720199,3.4808881,4.1879435,5.1107416,6.0317264,6.9545245,7.877322,8.80012,7.755854,6.7097745,5.6655083,4.6194286,3.5751622,4.5450974,5.5150323,6.484967,7.454902,8.424837,7.304426,6.185828,5.0654173,3.9450066,2.8245957,4.3402324,5.8540564,7.369693,8.885329,10.399154,9.19172,7.9842873,6.776854,5.569421,4.361988,4.748149,5.132497,5.516845,5.903006,6.2873545,6.008158,5.727149,5.4479527,5.1669436,4.8877473,8.094878,11.302009,14.510953,17.718082,20.925215,17.94289,14.960567,11.978244,8.994107,6.011784,5.5494785,5.087173,4.6248674,4.162562,3.7002566,9.492672,15.285088,21.077503,26.869919,32.662334,26.549025,20.437527,14.324218,8.212721,2.0994108,5.4352617,8.7693,12.105151,15.441002,18.77504,15.219821,11.664601,8.109382,4.554162,1.0007553,2.570781,4.1408067,5.710832,7.2808576,8.8508835,10.266808,11.684544,13.102281,14.520018,15.937754,12.803142,9.6685295,6.532104,3.397492,0.26287958,0.2955129,0.32814622,0.36077955,0.39159992,0.42423326,0.34083697,0.25562772,0.17041849,0.08520924,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.2229944,0.40791658,0.59283876,0.7777609,0.96268314,0.7705091,0.57833505,0.38434806,0.19217403,0.0,0.03988518,0.07977036,0.11965553,0.15954071,0.19942589,0.8684091,1.5355793,2.2027495,2.8699198,3.53709,3.8833659,4.227829,4.572292,4.9167547,5.2630305,6.1822023,7.1031876,8.02236,8.943344,9.862516,9.171778,8.482852,7.7921133,7.1031876,6.412449,6.834869,7.2572894,7.6797094,8.10213,8.52455,7.7322855,6.9400206,6.147756,5.3554916,4.5632267,4.07554,3.587853,3.100166,2.612479,2.124792,1.8691645,1.6153497,1.3597219,1.1040943,0.85027945,0.7197462,0.58921283,0.4604925,0.32995918,0.19942589,0.19217403,0.18492219,0.17767033,0.17041849,0.16316663,0.15410182,0.14684997,0.13959812,0.13234627,0.12509441,0.10696479,0.09064813,0.072518505,0.054388877,0.038072214,0.07795739,0.11784257,0.15772775,0.19761293,0.2374981,0.678048,1.1167849,1.5573349,1.9978848,2.4366217,1.9725033,1.5083848,1.0424535,0.57833505,0.11240368,0.36984438,0.62728506,0.88472575,1.1421664,1.3996071,1.1476053,0.89560354,0.6417888,0.38978696,0.13778515,0.6399758,1.1421664,1.6443571,2.1483607,2.6505513,3.0856624,3.5207734,3.9558845,4.3891826,4.8242936,4.1081734,3.39024,2.6723068,1.9543737,1.2382535,1.167548,1.0968424,1.0279498,0.9572442,0.8883517,0.72518504,0.5620184,0.40066472,0.2374981,0.07433146,0.09789998,0.11965553,0.14322405,0.16497959,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.054388877,0.047137026,0.03988518,0.032633327,0.025381476,0.065266654,0.10515183,0.14503701,0.18492219,0.22480737,0.24474995,0.26469254,0.28463513,0.3045777,0.3245203,0.29732585,0.27013144,0.24293698,0.21574254,0.18673515,0.15954071,0.13234627,0.10515183,0.07795739,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.22480737,0.44961473,0.6744221,0.89922947,1.1258497,0.97174793,0.8194591,0.6671702,0.5148814,0.36259252,0.80495536,1.2473183,1.6896812,2.132044,2.5744069,3.2306993,3.8851788,4.539658,5.1941376,5.8504305,5.177821,4.505212,3.832603,3.159994,2.4873846,2.2118144,1.938057,1.6624867,1.3869164,1.1131591,1.3216497,1.5319533,1.742257,1.9525607,2.1628644,2.4855716,2.808279,3.1291735,3.4518807,3.774588,4.6266804,5.480586,6.3326783,7.1847706,8.036863,6.7478466,5.4570174,4.168001,2.8771715,1.5881553,1.2745126,0.96268314,0.6508536,0.33721104,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.04169814,0.08520924,0.12690738,0.17041849,0.21211663,0.19217403,0.17223145,0.15228885,0.13234627,0.11240368,0.17223145,0.23205921,0.291887,0.35171473,0.41335547,0.95180535,1.4920682,2.032331,2.572594,3.1128569,2.1628644,2.4547513,2.7466383,3.0403383,3.3322253,3.6241121,3.7075086,3.7909048,3.872488,3.9558845,4.0374675,5.4026284,6.7677894,8.13295,9.498111,10.863272,11.876718,12.891977,13.907236,14.922495,15.937754,15.6422415,15.346728,15.053028,14.757515,14.462003,15.241576,16.022963,16.802538,17.582111,18.361685,18.76235,19.163015,19.561867,19.96253,20.363195,23.992746,27.622297,31.251848,34.883213,38.512764,39.23795,39.963135,40.68832,41.41169,42.136875,34.520622,26.902552,19.284483,11.668227,4.0501585,4.1897564,4.329355,4.4707656,4.610364,4.749962,4.358362,3.9649491,3.5733492,3.1799364,2.7883365,2.469255,2.1519866,1.8347181,1.5174497,1.2001812,1.6824293,2.1646774,2.6469254,3.1291735,3.6132345,2.8953013,2.1773682,1.4594349,0.7433147,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.3444629,0.50219065,0.65991837,0.81764615,0.97537386,0.9101072,0.8448406,0.7795739,0.71430725,0.6508536,2.1973107,3.7455807,5.292038,6.8403077,8.386765,9.064813,9.742861,10.420909,11.097144,11.775192,12.395226,13.015259,13.635292,14.255324,14.875358,14.927934,14.98051,15.033086,15.085662,15.138238,14.329657,13.522888,12.714307,11.907538,11.10077,11.00287,10.90497,10.80707,10.70917,10.613083,9.527119,8.442966,7.3570023,6.2728505,5.186886,5.2503395,5.3119802,5.375434,5.4370747,5.5005283,6.2202744,6.9400206,7.6597667,8.379513,9.099259,9.208037,9.3150015,9.421967,9.530745,9.637709,9.162713,8.6877165,8.212721,7.7377243,7.262728,8.107569,8.952409,9.79725,10.642091,11.486931,10.883214,10.277685,9.672155,9.066626,8.46291,7.5328593,6.60281,5.67276,4.74271,3.8126602,3.7419548,3.673062,3.6023567,3.531651,3.4627585,3.4754493,3.48814,3.5008307,3.5117085,3.5243993,3.576975,3.6295512,3.682127,3.7347028,3.787279,5.3591175,6.932769,8.504607,10.078259,11.650098,10.825199,10.000301,9.175404,8.350506,7.5256076,9.242483,10.959359,12.678047,14.394923,16.1118,17.455204,18.796797,20.140202,21.481794,22.8252,20.80012,18.77504,16.749962,14.724882,12.699803,12.930049,13.1602955,13.390542,13.620788,13.849221,13.042453,12.235684,11.427103,10.620335,9.811753,10.681975,11.552197,12.42242,13.292642,14.162864,13.080525,11.998186,10.915848,9.8316965,8.749357,7.6924005,6.635443,5.576673,4.519716,3.4627585,3.7818398,4.102734,4.421816,4.74271,5.0617914,5.5893636,6.1169357,6.644508,7.17208,7.699652,7.706904,7.7141557,7.723221,7.7304726,7.7377243,7.6307597,7.5219817,7.415017,7.308052,7.1992745,8.194591,9.189907,10.185224,11.18054,12.175857,14.897114,17.620184,20.343254,23.06451,25.78758,23.894846,22.002113,20.10938,18.216648,16.325727,16.30216,16.280403,16.256836,16.23508,16.213324,13.544643,10.877775,8.209095,5.542227,2.8753586,3.9993954,5.125245,6.249282,7.3751316,8.499168,7.115878,5.730775,4.345671,2.960568,1.5754645,1.3669738,1.1602961,0.95180535,0.7451276,0.53663695,1.2799516,2.0232663,2.764768,3.5080826,4.249584,5.389938,6.530291,7.6706448,8.809185,9.949538,8.457471,6.965402,5.473334,3.9794528,2.4873846,4.517903,6.546608,8.577126,10.607644,12.638163,10.957546,9.27693,7.5981264,5.91751,4.2368937,5.223145,6.207584,7.192023,8.178274,9.162713,8.107569,7.0524244,5.99728,4.942136,3.8869917,4.84061,5.7924156,6.7442207,7.6978393,8.649645,8.154706,7.6597667,7.1648283,6.6698895,6.1749506,9.71748,13.260008,16.802538,20.345066,23.887594,20.656897,17.428009,14.19731,10.966611,7.7377243,7.211965,6.688019,6.16226,5.638314,5.1125546,13.421362,21.726543,30.03535,38.342346,46.64934,37.711433,28.775343,19.837437,10.899531,1.9616255,7.2029004,12.442362,17.681824,22.9231,28.162561,22.817947,17.473333,12.126906,6.782293,1.4376793,2.3296568,3.2216346,4.115425,5.0074024,5.89938,9.182655,12.464118,15.747393,19.030668,22.31213,17.884876,13.457622,9.030367,4.603112,0.17585737,0.21755551,0.25925365,0.30276474,0.3444629,0.387974,0.3100166,0.23205921,0.15410182,0.07795739,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.15228885,0.27919623,0.40791658,0.53482395,0.66173136,0.5293851,0.39703882,0.26469254,0.13234627,0.0,0.059827764,0.11965553,0.1794833,0.23931105,0.2991388,0.91917205,1.5392052,2.1592383,2.7792716,3.3993049,3.680314,3.9595103,4.2405195,4.519716,4.800725,5.942891,7.0850577,8.227224,9.3693905,10.51337,9.427405,8.343254,7.2572894,6.1731377,5.087173,5.8395524,6.591932,7.344311,8.096691,8.8508835,8.21816,7.5854354,6.9527116,6.319988,5.6872635,5.0255322,4.361988,3.7002566,3.0367124,2.374981,2.0921588,1.8093367,1.5283275,1.2455053,0.96268314,0.80495536,0.64722764,0.4894999,0.33177215,0.17585737,0.17041849,0.16497959,0.15954071,0.15410182,0.15047589,0.14503701,0.13959812,0.13415924,0.13053331,0.12509441,0.10515183,0.08520924,0.065266654,0.045324065,0.025381476,0.08520924,0.14503701,0.20486477,0.26469254,0.3245203,0.97174793,1.6207886,2.268016,2.9152439,3.5624714,2.864481,2.1683033,1.4703126,0.77232206,0.07433146,0.26831847,0.4604925,0.6526665,0.8448406,1.0370146,0.86478317,0.69255173,0.52032024,0.3480888,0.17585737,0.8103943,1.4449311,2.079468,2.715818,3.350355,3.5534067,3.7546456,3.9576974,4.160749,4.361988,3.8543584,3.346729,2.8390994,2.333283,1.8256533,1.6697385,1.5156367,1.3597219,1.2056202,1.0497054,0.8629702,0.6744221,0.48768693,0.2991388,0.11240368,0.11421664,0.11784257,0.11965553,0.12328146,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.058014803,0.052575916,0.047137026,0.04169814,0.038072214,0.072518505,0.10696479,0.14322405,0.17767033,0.21211663,0.24293698,0.27194437,0.30276474,0.33177215,0.36259252,0.34083697,0.31726846,0.2955129,0.27194437,0.25018883,0.21574254,0.1794833,0.14503701,0.11059072,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.15047589,0.2991388,0.44961473,0.6000906,0.7505665,0.6526665,0.55476654,0.45686656,0.36077955,0.26287958,0.75781834,1.2527572,1.7476959,2.2426348,2.7375734,3.870675,5.0019636,6.1350656,7.268167,8.399456,7.460341,6.5194135,5.580299,4.6393714,3.7002566,3.2379513,2.7756457,2.3133402,1.8492218,1.3869164,1.4141108,1.4431182,1.4703126,1.4975071,1.5247015,2.039583,2.5544643,3.0693457,3.584227,4.099108,5.522284,6.94546,8.366822,9.789998,11.213174,9.440096,7.667019,5.8957543,4.122677,2.3495996,1.887294,1.4249886,0.96268314,0.50037766,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.032633327,0.065266654,0.09789998,0.13053331,0.16316663,0.14503701,0.12690738,0.11059072,0.092461094,0.07433146,0.17767033,0.27919623,0.3825351,0.48587397,0.5873999,1.3724127,2.1574254,2.9424384,3.727451,4.512464,2.1121013,2.3405347,2.5671551,2.7955883,3.0222087,3.2506418,3.2343252,3.2198215,3.2053177,3.1908143,3.1744974,4.6575007,6.1405044,7.6216946,9.104698,10.587702,11.583018,12.578335,13.571837,14.567154,15.56247,15.564283,15.567909,15.569723,15.573349,15.575162,16.378304,17.179634,17.982777,18.78592,19.587248,19.699652,19.812056,19.92446,20.036863,20.149265,24.52757,28.904062,33.282368,37.66067,42.037163,40.26227,38.48738,36.712494,34.937603,33.162712,27.172684,21.182655,15.192626,9.202598,3.2125697,3.6948178,4.177066,4.6593137,5.143375,5.6256227,5.0726695,4.519716,3.966762,3.4156215,2.8626678,2.4348087,2.0069497,1.5790904,1.1530442,0.72518504,0.96087015,1.1947423,1.4304274,1.6642996,1.8999848,1.5228885,1.1457924,0.7668832,0.38978696,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,0.4604925,0.67079616,0.8792868,1.0895905,1.2998942,1.1059072,0.9101072,0.71430725,0.52032024,0.3245203,2.0540867,3.785466,5.5150323,7.2445984,8.974165,9.3693905,9.764616,10.1598425,10.555068,10.950294,11.684544,12.420607,13.154857,13.889107,14.625169,14.581658,14.53996,14.498261,14.454751,14.413053,13.789393,13.167547,12.545701,11.922042,11.300196,11.169662,11.039129,10.910409,10.779876,10.649343,9.657652,8.664148,7.6724577,6.680767,5.6872635,5.7996674,5.9120708,6.0244746,6.1368785,6.249282,7.12313,7.995165,8.8672,9.739235,10.613083,10.609457,10.607644,10.605831,10.602205,10.600392,10.087324,9.574255,9.063,8.549932,8.036863,8.910711,9.782746,10.654781,11.526816,12.400664,11.597522,10.794379,9.99305,9.189907,8.386765,7.473032,6.5574856,5.6419396,4.7282066,3.8126602,3.5534067,3.29234,3.0330863,2.7720199,2.5127661,2.5870976,2.663242,2.7375734,2.811905,2.8880494,2.9823234,3.0765975,3.1726844,3.2669585,3.3630457,4.954827,6.546608,8.140202,9.731983,11.325577,10.738177,10.150778,9.563377,8.974165,8.386765,10.2142315,12.0416975,13.870976,15.698443,17.52591,18.490406,19.4549,20.419397,21.385706,22.350203,20.4756,18.599184,16.72458,14.849977,12.975373,13.05333,13.129475,13.207433,13.28539,13.363347,12.514881,11.668227,10.81976,9.973107,9.12464,10.009366,10.894093,11.780631,12.665357,13.550082,12.6145935,11.680918,10.745429,9.80994,8.874452,7.7776093,6.680767,5.582112,4.4852695,3.386614,3.7473936,4.1081734,4.4671397,4.8279195,5.186886,5.5567303,5.9283876,6.298232,6.6680765,7.037921,7.021604,7.0071006,6.9925966,6.978093,6.9617763,7.1031876,7.2427855,7.382384,7.5219817,7.663393,8.423024,9.182655,9.9422865,10.701918,11.463363,14.117539,16.771717,19.427708,22.081884,24.737875,22.97205,21.208036,19.442211,17.678198,15.912373,16.13174,16.352922,16.57229,16.79166,17.01284,14.184619,11.358211,8.529989,5.7017674,2.8753586,4.12449,5.375434,6.624565,7.8755093,9.12464,7.570932,6.01541,4.459888,2.904366,1.3506571,1.1657349,0.9808127,0.79589057,0.6091554,0.42423326,1.2019942,1.9797552,2.7575161,3.5352771,4.313038,5.669134,7.027043,8.384952,9.742861,11.10077,9.1609,7.219217,5.279347,3.339477,1.3996071,4.4907084,7.5799966,10.669285,13.760386,16.849674,14.610665,12.3698435,10.130835,7.890013,5.6491914,6.104245,6.5592985,7.0143523,7.4694057,7.9244595,7.021604,6.1205616,5.217706,4.314851,3.4119956,4.933071,6.452334,7.9734097,9.492672,11.011934,10.303066,9.592385,8.881703,8.172835,7.462154,11.340081,15.218008,19.095936,22.97205,26.849976,23.372713,19.89545,16.41819,12.939114,9.461852,8.874452,8.287052,7.699652,7.112252,6.5248523,17.34824,28.169813,38.9932,49.814774,60.63816,48.873844,37.113155,25.348843,13.588155,1.8256533,8.970539,16.115425,23.26031,30.405195,37.55008,30.41426,23.280252,16.144432,9.010424,1.8746033,2.0903459,2.3042755,2.520018,2.7357605,2.94969,8.098504,13.245504,18.392506,23.539507,28.68832,22.96661,17.248526,11.526816,5.806919,0.0870222,0.13959812,0.19217403,0.24474995,0.29732585,0.34990177,0.27919623,0.21030366,0.13959812,0.07070554,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.08339628,0.15228885,0.2229944,0.291887,0.36259252,0.29007402,0.21755551,0.14503701,0.072518505,0.0,0.07977036,0.15954071,0.23931105,0.3208944,0.40066472,0.97174793,1.5446441,2.1175404,2.6904364,3.2633326,3.4772623,3.6930048,3.9069343,4.122677,4.3366065,5.7017674,7.066928,8.432089,9.79725,11.162411,9.683033,8.201842,6.722465,5.243088,3.7618973,4.844236,5.9265747,7.0107265,8.093065,9.175404,8.70222,8.23085,7.757667,7.2844834,6.813113,5.975525,5.137936,4.3003473,3.4627585,2.6251698,2.3151531,2.0051367,1.69512,1.3851035,1.0750868,0.8901646,0.70524246,0.52032024,0.33539808,0.15047589,0.14684997,0.14503701,0.14322405,0.13959812,0.13778515,0.13415924,0.13234627,0.13053331,0.12690738,0.12509441,0.10333887,0.07977036,0.058014803,0.034446288,0.012690738,0.092461094,0.17223145,0.2520018,0.33177215,0.41335547,1.2672608,2.1229792,2.9768846,3.832603,4.688321,3.7582715,2.8282216,1.8981718,0.968122,0.038072214,0.16497959,0.291887,0.42060733,0.5475147,0.6744221,0.581961,0.4894999,0.39703882,0.3045777,0.21211663,0.9808127,1.7476959,2.514579,3.2832751,4.0501585,4.019338,3.9903307,3.9595103,3.930503,3.8996825,3.6023567,3.3050308,3.007705,2.7103791,2.4130533,2.1719291,1.9326181,1.693307,1.452183,1.2128719,1.0007553,0.7868258,0.5747091,0.36259252,0.15047589,0.13234627,0.11421664,0.09789998,0.07977036,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.059827764,0.058014803,0.054388877,0.052575916,0.05076295,0.07977036,0.11059072,0.13959812,0.17041849,0.19942589,0.23931105,0.27919623,0.3208944,0.36077955,0.40066472,0.3825351,0.36440548,0.3480888,0.32995918,0.31182957,0.27013144,0.22662032,0.18492219,0.14322405,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0,0.0,0.0,0.0,0.0,0.07433146,0.15047589,0.22480737,0.2991388,0.37528324,0.33177215,0.29007402,0.24837588,0.20486477,0.16316663,0.7106813,1.258196,1.8057107,2.3532255,2.9007401,4.510651,6.1205616,7.7304726,9.340384,10.950294,9.742861,8.535428,7.327995,6.1205616,4.9131284,4.262275,3.6132345,2.962381,2.3133402,1.6624867,1.5083848,1.35247,1.1983683,1.0424535,0.8883517,1.5954071,2.3024626,3.009518,3.7165732,4.4254417,6.4178877,8.410334,10.40278,12.395226,14.387671,12.132345,9.87702,7.6216946,5.368182,3.1128569,2.5000753,1.887294,1.2745126,0.66173136,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.09789998,0.08339628,0.06707962,0.052575916,0.038072214,0.18310922,0.32814622,0.47318324,0.61822027,0.76325727,1.79302,2.8227828,3.8525455,4.882308,5.9120708,2.0631514,2.2245052,2.3876717,2.5508385,2.712192,2.8753586,2.762955,2.6505513,2.5381477,2.4257438,2.3133402,3.9123733,5.5132194,7.112252,8.713099,10.312131,11.287505,12.262879,13.238253,14.211814,15.187187,15.488139,15.787278,16.08823,16.38737,16.68832,17.513218,18.338116,19.163015,19.987913,20.81281,20.636953,20.462908,20.287052,20.113007,19.93715,25.062395,30.18764,35.312885,40.43813,45.563377,41.28841,37.013443,32.736664,28.4617,24.186733,19.824745,15.462758,11.10077,6.736969,2.374981,3.199879,4.024777,4.8496747,5.674573,6.4994707,5.7869763,5.0744824,4.361988,3.6494937,2.9369993,2.4003625,1.8619126,1.3252757,0.7868258,0.25018883,0.2374981,0.22480737,0.21211663,0.19942589,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06164073,0.12509441,0.18673515,0.25018883,0.31182957,0.5747091,0.8375887,1.1004683,1.3633479,1.6244144,1.2998942,0.97537386,0.6508536,0.3245203,0.0,1.9126755,3.825351,5.7380266,7.650702,9.563377,9.675781,9.788185,9.900589,10.012992,10.125396,10.975676,11.8241415,12.674421,13.524701,14.37498,14.237195,14.09941,13.961625,13.825653,13.687867,13.24913,12.812206,12.375282,11.938358,11.499621,11.338268,11.175101,11.011934,10.850581,10.687414,9.788185,8.887142,7.987913,7.0868707,6.187641,6.350808,6.5121617,6.6753283,6.836682,6.9998484,8.024173,9.050309,10.074633,11.10077,12.125093,12.012691,11.900287,11.787883,11.675479,11.563075,11.011934,10.462607,9.91328,9.362139,8.812811,9.712041,10.613083,11.512312,12.413355,13.312584,12.311829,11.312886,10.312131,9.313189,8.312433,7.413204,6.5121617,5.612932,4.7118897,3.8126602,3.3630457,2.911618,2.4620032,2.0123885,1.5627737,1.7005589,1.8383441,1.9743162,2.1121013,2.2498865,2.3876717,2.525457,2.663242,2.7992141,2.9369993,4.550536,6.16226,7.7757964,9.38752,10.999244,10.649343,10.29944,9.949538,9.599637,9.249735,11.187792,13.124036,15.062093,17.00015,18.938208,19.525606,20.113007,20.700407,21.287807,21.875206,20.149265,18.425138,16.699198,14.975071,13.24913,13.174799,13.100468,13.024323,12.949992,12.87566,11.9873085,11.10077,10.212419,9.325879,8.437528,9.336758,10.2378,11.137029,12.038072,12.937301,12.1504755,11.361836,10.57501,9.788185,8.999546,7.8628187,6.7242785,5.5875506,4.4508233,3.3122826,3.7129474,4.1117992,4.512464,4.9131284,5.3119802,5.524097,5.7380266,5.9501433,6.16226,6.3743763,6.338117,6.300045,6.261973,6.2257137,6.187641,6.5756154,6.9617763,7.3497505,7.7377243,8.125698,8.649645,9.175404,9.699349,10.225109,10.750868,13.337966,15.925063,18.512161,21.099258,23.68817,22.049252,20.412146,18.77504,17.137936,15.50083,15.963136,16.425442,16.887747,17.350052,17.812357,14.824595,11.836833,8.849071,5.863121,2.8753586,4.249584,5.6256227,6.9998484,8.375887,9.750113,8.024173,6.300045,4.574105,2.8499773,1.1258497,0.96268314,0.7995165,0.63816285,0.4749962,0.31182957,1.1258497,1.938057,2.7502642,3.5624714,4.3746786,5.9501433,7.5256076,9.099259,10.674724,12.250188,9.862516,7.474845,5.087173,2.6995013,0.31182957,4.461701,8.611572,12.763257,16.913128,21.063,18.261972,15.462758,12.661731,9.862516,7.063302,6.987158,6.9128265,6.836682,6.7623506,6.688019,5.9374523,5.186886,4.4381323,3.6875658,2.9369993,5.0255322,7.112252,9.200785,11.287505,13.374225,12.449615,11.525003,10.600392,9.675781,8.749357,12.962683,17.174194,21.38752,25.600845,29.812357,26.08672,22.362894,18.637255,14.911617,11.187792,10.536939,9.8878975,9.237044,8.588004,7.93715,21.275116,34.611267,47.951046,61.2872,74.62517,60.036255,45.450974,30.862062,16.274965,1.6878681,10.738177,19.786674,28.836983,37.88729,46.937603,38.012386,29.087172,20.161957,11.236742,2.3133402,1.8492218,1.3869164,0.9246109,0.46230546,0.0,7.0125394,14.025079,21.037619,28.050158,35.062695,28.050158,21.037619,14.025079,7.0125394,0.0,0.06164073,0.12509441,0.18673515,0.25018883,0.31182957,0.25018883,0.18673515,0.12509441,0.06164073,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.099712946,0.19942589,0.2991388,0.40066472,0.50037766,1.0243238,1.550083,2.0758421,2.5997884,3.1255474,3.2742105,3.4246864,3.5751622,3.7256382,3.874301,5.462456,7.0506115,8.636953,10.225109,11.813264,9.936848,8.062244,6.187641,4.313038,2.4366217,3.8507326,5.2630305,6.6753283,8.087626,9.499924,9.188094,8.874452,8.562622,8.2507925,7.93715,6.925517,5.9120708,4.900438,3.8869917,2.8753586,2.5381477,2.1991236,1.8619126,1.5247015,1.1874905,0.97537386,0.76325727,0.5493277,0.33721104,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.099712946,0.19942589,0.2991388,0.40066472,0.50037766,1.5627737,2.6251698,3.6875658,4.749962,5.812358,4.650249,3.48814,2.324218,1.162109,0.0,0.06164073,0.12509441,0.18673515,0.25018883,0.31182957,0.2991388,0.28826106,0.2755703,0.26287958,0.25018883,1.1494182,2.0504606,2.94969,3.8507326,4.749962,4.4870825,4.2242026,3.9631362,3.7002566,3.437377,3.350355,3.2633326,3.1744974,3.0874753,3.000453,2.6741197,2.3495996,2.0250793,1.7005589,1.3742256,1.1367276,0.89922947,0.66173136,0.42423326,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.0870222,0.11240368,0.13778515,0.16316663,0.18673515,0.2374981,0.28826106,0.33721104,0.387974,0.43692398,0.42423326,0.41335547,0.40066472,0.387974,0.37528324,0.3245203,0.2755703,0.22480737,0.17585737,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.66173136,1.261822,1.8619126,2.4620032,3.0620937,5.1506267,7.2373466,9.325879,11.4126,13.499319,12.025381,10.549629,9.07569,7.5999393,6.1241875,5.2865987,4.4508233,3.6132345,2.7756457,1.938057,1.6008459,1.261822,0.9246109,0.5873999,0.25018883,1.1494182,2.0504606,2.94969,3.8507326,4.749962,7.313491,9.875207,12.436923,15.000452,17.562168,14.824595,12.087022,9.349448,6.6118746,3.874301,3.1128569,2.3495996,1.5881553,0.824898,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.18673515,0.37528324,0.5620184,0.7505665,0.93730164,2.2118144,3.48814,4.762653,6.037165,7.311678,2.2498865,2.427557,2.6052272,2.7828975,2.960568,3.1382382,3.2053177,3.2723975,3.339477,3.4083695,3.4754493,5.2032027,6.929143,8.656897,10.384649,12.112403,13.100468,14.0867195,15.074784,16.062849,17.050913,17.027344,17.005589,16.982021,16.960264,16.936697,17.50778,18.07705,18.648132,19.217403,19.786674,20.015106,20.241728,20.470161,20.696781,20.925215,25.852846,30.78048,35.70811,40.635742,45.563377,40.57773,35.592083,30.608248,25.6226,20.636953,17.052727,13.468499,9.882459,6.298232,2.712192,3.2850883,3.8579843,4.4308805,5.0019636,5.57486,5.1941376,4.8152285,4.4345064,4.0555973,3.6748753,3.5008307,3.3249733,3.149116,2.9750717,2.7992141,2.2970235,1.794833,1.2926424,0.7904517,0.28826106,0.23024625,0.17223145,0.11421664,0.058014803,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.11784257,0.23568514,0.35171473,0.46955732,0.5873999,0.78319985,0.97718686,1.1729867,1.3669738,1.5627737,1.2491312,0.93730164,0.62547207,0.31182957,0.0,1.8999848,3.7999697,5.6999545,7.5999393,9.499924,9.670342,9.840761,10.009366,10.179785,10.3502035,11.030065,11.709926,12.389787,13.069647,13.749508,13.6244135,13.499319,13.374225,13.24913,13.125849,12.658105,12.19036,11.722616,11.254871,10.7871275,10.674724,10.56232,10.449916,10.337513,10.225109,9.52168,8.820063,8.116633,7.415017,6.7134004,6.8602505,7.0071006,7.155763,7.3026133,7.4494634,8.497355,9.545248,10.593141,11.63922,12.687112,12.737875,12.786825,12.837588,12.888351,12.937301,12.351714,11.7679405,11.182353,10.596766,10.012992,10.6783495,11.341894,12.007251,12.672608,13.337966,12.389787,11.443419,10.49524,9.547061,8.600695,7.552802,6.5049095,5.4570174,4.409125,3.3630457,3.0167696,2.6723068,2.327844,1.983381,1.6371052,1.7205015,1.8020848,1.8854811,1.9670644,2.0504606,2.3405347,2.6306088,2.9206827,3.2107568,3.5008307,4.695573,5.8903155,7.0850577,8.2798,9.474543,9.32044,9.164526,9.010424,8.854509,8.700407,11.4126,14.124791,16.836983,19.549175,22.26318,22.179785,22.098202,22.014805,21.933222,21.849825,20.252605,18.655384,17.058165,15.459132,13.861912,13.845595,13.827466,13.809336,13.793019,13.77489,12.645414,11.515939,10.384649,9.255174,8.125698,8.807372,9.490859,10.172533,10.854207,11.537694,10.957546,10.377398,9.79725,9.217102,8.636953,7.6398244,6.642695,5.6455655,4.646623,3.6494937,4.0519714,4.454449,4.856927,5.2594047,5.661882,5.6655083,5.667321,5.669134,5.67276,5.674573,5.661882,5.6491914,5.638314,5.6256227,5.612932,6.0244746,6.43783,6.849373,7.262728,7.6742706,8.330563,8.985043,9.639522,10.2958145,10.950294,13.000754,15.049402,17.099863,19.150324,21.200785,19.797552,18.394318,16.992899,15.589665,14.188245,14.512766,14.837286,15.161806,15.488139,15.812659,13.207433,10.602205,7.996978,5.391751,2.7883365,3.7890918,4.7916603,5.7942286,6.796797,7.799365,6.4632115,5.125245,3.787279,2.4493124,1.1131591,1.0497054,0.9880646,0.9246109,0.8629702,0.7995165,1.3470312,1.8945459,2.4420607,2.9895754,3.53709,5.1071157,6.677141,8.247167,9.817192,11.3872175,9.255174,7.12313,4.989273,2.857229,0.72518504,4.2477713,7.7703576,11.292944,14.81553,18.338116,16.115425,13.892733,11.67004,9.447348,7.224656,7.083245,6.9400206,6.796797,6.6553855,6.5121617,5.6800117,4.847862,4.0157123,3.1817493,2.3495996,4.022964,5.6945157,7.36788,9.039432,10.712796,9.987611,9.262425,8.537241,7.8120556,7.0868707,10.792566,14.498261,18.202145,21.90784,25.611723,22.355642,19.097748,15.839854,12.581961,9.325879,10.125396,10.924912,11.724429,12.525759,13.325275,22.640276,31.955278,41.27028,50.58528,59.900284,49.116783,38.335094,27.551592,16.769903,5.9882154,12.300951,18.611874,24.92461,31.237345,37.55008,30.630003,23.709925,16.789846,9.869768,2.94969,3.6132345,4.274966,4.936697,5.600241,6.261973,10.620335,14.976884,19.335245,23.691795,28.050158,22.439037,16.829731,11.220426,5.6093063,0.0,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.13778515,0.22480737,0.31182957,0.40066472,0.48768693,0.72337204,0.9572442,1.1929294,1.4268016,1.6624867,1.8818551,2.1030366,2.322405,2.5417736,2.762955,3.2397642,3.7183862,4.195195,4.6720047,5.1506267,6.3072968,7.46578,8.62245,9.77912,10.937603,9.24067,7.5419245,5.844991,4.1480584,2.4493124,3.5624714,4.6756306,5.7869763,6.9001355,8.013294,7.746789,7.4820967,7.217404,6.9527116,6.688019,6.0679855,5.4479527,4.8279195,4.207886,3.587853,3.2651455,2.9424384,2.619731,2.2970235,1.9743162,1.6026589,1.2291887,0.8575313,0.48587397,0.11240368,0.11784257,0.12328146,0.12690738,0.13234627,0.13778515,0.13234627,0.12690738,0.12328146,0.11784257,0.11240368,0.12690738,0.14322405,0.15772775,0.17223145,0.18673515,0.23205921,0.27738327,0.32270733,0.3680314,0.41335547,1.35247,2.2915847,3.2325122,4.171627,5.1125546,4.0918565,3.0729716,2.0522738,1.0333886,0.012690738,0.06164073,0.11240368,0.16316663,0.21211663,0.26287958,0.2755703,0.28826106,0.2991388,0.31182957,0.3245203,1.0841516,1.845596,2.6052272,3.3648586,4.12449,4.0102735,3.8942437,3.780027,3.6658103,3.5497808,3.3793623,3.2107568,3.0403383,2.8699198,2.6995013,2.4058013,2.1102884,1.8147756,1.5192627,1.2255627,1.015259,0.80495536,0.5946517,0.38434806,0.17585737,0.13959812,0.10515183,0.07070554,0.034446288,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.07433146,0.07433146,0.07433146,0.07433146,0.07433146,0.07433146,0.10333887,0.13053331,0.15772775,0.18492219,0.21211663,0.25925365,0.30820364,0.35534066,0.40247768,0.44961473,0.43329805,0.41516843,0.39703882,0.38072214,0.36259252,0.3245203,0.28826106,0.25018883,0.21211663,0.17585737,0.15410182,0.13415924,0.11421664,0.09427405,0.07433146,0.387974,0.69980353,1.0116332,1.3252757,1.6371052,1.5972201,1.5573349,1.5174497,1.4775645,1.4376793,1.1602961,0.88291276,0.6055295,0.32814622,0.05076295,0.6345369,1.2201238,1.8057107,2.3894846,2.9750717,5.4932766,8.009668,10.527874,13.044266,15.56247,14.0323305,12.50219,10.97205,9.441909,7.911769,6.7152133,5.516845,4.3202896,3.1219215,1.9253663,1.649796,1.3742256,1.1004683,0.824898,0.5493277,1.3071461,2.0649643,2.8227828,3.5806012,4.3366065,6.8203654,9.302311,11.784257,14.268016,16.749962,14.190058,11.630155,9.070251,6.510349,3.9504454,3.1744974,2.4003625,1.6244144,0.85027945,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.15954071,0.2574407,0.35534066,0.45324063,0.5493277,0.7469406,0.9445535,1.1421664,1.3397794,1.5373923,2.6505513,3.7618973,4.8750563,5.9882154,7.0995617,2.4366217,2.6306088,2.8227828,3.0149567,3.207131,3.3993049,3.6476808,3.8942437,4.1426196,4.3891826,4.6375585,6.492219,8.34688,10.203354,12.058014,13.912675,14.911617,15.912373,16.913128,17.912071,18.912827,18.568363,18.222088,17.877625,17.533161,17.186886,17.50234,17.817797,18.133251,18.446894,18.76235,19.393261,20.022358,20.653269,21.282368,21.913279,26.643297,31.371504,36.103336,40.833355,45.563377,39.867046,34.17253,28.478016,22.781689,17.087172,14.280706,11.472427,8.664148,5.857682,3.049403,3.3702974,3.6893787,4.0102735,4.329355,4.650249,4.603112,4.554162,4.507025,4.459888,4.4127507,4.599486,4.788034,4.974769,5.163317,5.3500524,4.358362,3.3648586,2.373168,1.3796645,0.387974,0.3100166,0.23205921,0.15410182,0.07795739,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.17223145,0.3444629,0.5166943,0.69073874,0.8629702,0.9898776,1.1167849,1.2455053,1.3724127,1.49932,1.2001812,0.89922947,0.6000906,0.2991388,0.0,1.887294,3.774588,5.661882,7.549176,9.438283,9.664904,9.893337,10.119957,10.348391,10.57501,11.084454,11.595709,12.105151,12.6145935,13.125849,13.011633,12.899229,12.786825,12.674421,12.562017,12.065266,11.566701,11.069949,10.573197,10.074633,10.012992,9.949538,9.8878975,9.824444,9.762803,9.256987,8.752983,8.247167,7.743163,7.2373466,7.369693,7.502039,7.6343856,7.7667317,7.900891,8.970539,10.040187,11.109835,12.179482,13.24913,13.46306,13.675177,13.887294,14.09941,14.313339,13.693306,13.073273,12.45324,11.833207,11.213174,11.642846,12.072517,12.50219,12.931862,13.363347,12.467744,11.57214,10.6783495,9.782746,8.887142,7.6924005,6.497658,5.3029156,4.1081734,2.911618,2.6723068,2.4329958,2.1918716,1.9525607,1.7132497,1.7404441,1.7676386,1.794833,1.8220274,1.8492218,2.2933977,2.7357605,3.1781235,3.6204863,4.062849,4.84061,5.618371,6.394319,7.17208,7.949841,7.989726,8.029612,8.069496,8.109382,8.149267,11.637406,15.125546,18.611874,22.100014,25.588154,24.835773,24.083395,23.329203,22.576822,21.824444,20.354132,18.885632,17.41532,15.945006,14.474693,14.514579,14.554463,14.594349,14.634234,14.674119,13.301706,11.929294,10.556881,9.184468,7.8120556,8.2779875,8.7421055,9.208037,9.672155,10.138086,9.764616,9.39296,9.019489,8.647832,8.274362,7.41683,6.5592985,5.7017674,4.844236,3.9867048,4.3928084,4.797099,5.2032027,5.6074934,6.011784,5.805106,5.5966153,5.389938,5.18326,4.974769,4.98746,5.0001507,5.0128417,5.0255322,5.038223,5.475147,5.9120708,6.350808,6.787732,7.224656,8.009668,8.794682,9.579695,10.364707,11.14972,12.661731,14.175554,15.687565,17.199575,18.711586,17.545853,16.378304,15.210756,14.043208,12.87566,13.062395,13.24913,13.437678,13.6244135,13.812962,11.59027,9.367578,7.1448855,4.9221935,2.6995013,3.3304121,3.9595103,4.590421,5.219519,5.8504305,4.900438,3.9504454,3.000453,2.0504606,1.1004683,1.1367276,1.1747998,1.2128719,1.2491312,1.2872034,1.5700256,1.8528478,2.13567,2.4166791,2.6995013,4.264088,5.8304877,7.3950744,8.9596615,10.524248,8.647832,6.7696023,4.893186,3.0149567,1.1367276,4.0320287,6.92733,9.822631,12.717933,15.613234,13.967064,12.322706,10.676537,9.03218,7.3878226,7.177519,6.967215,6.7569118,6.546608,6.338117,5.422571,4.507025,3.5932918,2.6777458,1.7621996,3.0203958,4.2767787,5.5349746,6.793171,8.049554,7.5256076,6.9998484,6.474089,5.9501433,5.424384,8.62245,11.820516,15.016769,18.214834,21.4129,18.622751,15.8326025,13.042453,10.252303,7.462154,9.712041,11.961927,14.211814,16.4617,18.7134,24.005438,29.297476,34.58951,39.883366,45.1754,38.197308,31.22103,24.242935,17.264843,10.28675,13.861912,17.437075,21.012236,24.587399,28.162561,23.24762,18.332678,13.417736,8.502794,3.587853,5.375434,7.1630154,8.950596,10.738177,12.525759,14.22813,15.930502,17.632874,19.335245,21.037619,16.829731,12.621845,8.4139595,4.207886,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.22480737,0.41335547,0.6000906,0.7868258,0.97537386,1.3452182,1.7150626,2.084907,2.4547513,2.8245957,2.7393866,2.6541772,2.570781,2.4855716,2.4003625,3.2053177,4.0102735,4.8152285,5.620184,6.4251394,7.1521373,7.8791356,8.607946,9.334945,10.061942,8.54268,7.023417,5.5023413,3.9830787,2.4620032,3.2742105,4.0882306,4.900438,5.712645,6.5248523,6.3072968,6.089741,5.8721857,5.65463,5.4370747,5.2104545,4.9820213,4.7554007,4.5269675,4.3003473,3.9921436,3.6857529,3.3775494,3.0693457,2.762955,2.229944,1.696933,1.1657349,0.6327239,0.099712946,0.11059072,0.11965553,0.13053331,0.13959812,0.15047589,0.13959812,0.13053331,0.11965553,0.11059072,0.099712946,0.15410182,0.21030366,0.26469254,0.3208944,0.37528324,0.36440548,0.35534066,0.3444629,0.33539808,0.3245203,1.1421664,1.9598125,2.7774587,3.5951047,4.4127507,3.5352771,2.657803,1.7803292,0.90285534,0.025381476,0.06164073,0.099712946,0.13778515,0.17585737,0.21211663,0.25018883,0.28826106,0.3245203,0.36259252,0.40066472,1.020698,1.6407311,2.2607644,2.8807976,3.5008307,3.531651,3.5642843,3.5969179,3.6295512,3.6621845,3.4101827,3.1581807,2.904366,2.6523643,2.4003625,2.13567,1.8691645,1.6044719,1.3397794,1.0750868,0.8919776,0.7106813,0.5275721,0.3444629,0.16316663,0.13053331,0.09789998,0.065266654,0.032633327,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.038072214,0.05076295,0.06164073,0.07433146,0.0870222,0.0870222,0.0870222,0.0870222,0.0870222,0.0870222,0.11784257,0.14684997,0.17767033,0.20667773,0.2374981,0.28282216,0.32814622,0.37165734,0.4169814,0.46230546,0.4405499,0.4169814,0.39522585,0.37165734,0.34990177,0.3245203,0.2991388,0.2755703,0.25018883,0.22480737,0.21030366,0.19579996,0.1794833,0.16497959,0.15047589,0.774135,1.3996071,2.0250793,2.6505513,3.2742105,3.1944401,3.1146698,3.0348995,2.955129,2.8753586,2.3079014,1.7404441,1.1729867,0.6055295,0.038072214,0.6073425,1.1766127,1.7476959,2.3169663,2.8880494,5.8359265,8.781991,11.729868,14.677745,17.625622,16.03928,14.454751,12.870221,11.285692,9.699349,8.1420145,6.58468,5.027345,3.4700103,1.9126755,1.7005589,1.4866294,1.2745126,1.062396,0.85027945,1.4648738,2.079468,2.6958754,3.3104696,3.925064,6.3272395,8.729415,11.133403,13.535579,15.937754,13.555521,11.171475,8.789243,6.4070096,4.024777,3.2379513,2.4493124,1.6624867,0.87566096,0.0870222,0.07070554,0.052575916,0.034446288,0.018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.27013144,0.47680917,0.6852999,0.8919776,1.1004683,1.3071461,1.5156367,1.7223145,1.9308052,2.137483,3.0874753,4.0374675,4.98746,5.9374523,6.887445,2.6251698,2.8318477,3.0403383,3.247016,3.4555066,3.6621845,4.0900435,4.517903,4.945762,5.371808,5.7996674,7.783048,9.764616,11.747997,13.729566,15.712947,16.72458,17.738026,18.749659,19.763105,20.774738,20.107569,19.440397,18.773228,18.104244,17.437075,17.496902,17.55673,17.61837,17.678198,17.738026,18.769602,19.80299,20.834566,21.867954,22.89953,27.431936,31.964344,36.49675,41.030968,45.563377,39.15818,32.752983,26.347786,19.942589,13.537392,11.506873,9.4781685,7.4476504,5.4171324,3.386614,3.4555066,3.5225863,3.589666,3.6567454,3.7256382,4.0102735,4.2949085,4.5795436,4.8641787,5.1506267,5.6999545,6.249282,6.8004227,7.3497505,7.899078,6.4178877,4.934884,3.4518807,1.9706904,0.48768693,0.38978696,0.291887,0.19579996,0.09789998,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.22662032,0.4550536,0.68167394,0.9101072,1.1367276,1.1983683,1.258196,1.3180238,1.3778516,1.4376793,1.1494182,0.8629702,0.5747091,0.28826106,0.0,1.8746033,3.7492065,5.6256227,7.500226,9.374829,9.659465,9.944099,10.230548,10.515183,10.799818,11.1406555,11.479679,11.820516,12.15954,12.500377,12.400664,12.299138,12.199425,12.099712,11.999999,11.472427,10.944855,10.417283,9.88971,9.362139,9.349448,9.336758,9.325879,9.313189,9.300498,8.992294,8.685904,8.3777,8.069496,7.763106,7.8791356,7.996978,8.1148205,8.232663,8.350506,9.441909,10.535126,11.628342,12.719746,13.812962,14.188245,14.561715,14.936998,15.312282,15.687565,15.033086,14.376793,13.722314,13.067834,12.413355,12.607342,12.803142,12.9971285,13.192928,13.386916,12.545701,11.702674,10.859646,10.016619,9.175404,7.8319983,6.490406,5.147001,3.8054085,2.4620032,2.327844,2.1918716,2.0577126,1.9217403,1.7875811,1.7603867,1.7331922,1.7041848,1.6769904,1.649796,2.2444477,2.8390994,3.435564,4.0302157,4.6248674,4.985647,5.3446136,5.7053933,6.0643597,6.4251394,6.6608243,6.8946967,7.130382,7.364254,7.5999393,11.862214,16.124489,20.386765,24.650852,28.913128,27.489952,26.066776,24.645412,23.222239,21.800875,20.45747,19.115877,17.772472,16.43088,15.087475,15.185374,15.283275,15.379361,15.477262,15.575162,13.959812,12.344462,10.729113,9.115576,7.500226,7.746789,7.995165,8.241728,8.490104,8.736667,8.571687,8.406708,8.241728,8.076748,7.911769,7.1956487,6.4777155,5.7597823,5.041849,4.325729,4.7318325,5.139749,5.5476656,5.955582,6.3616858,5.9447045,5.527723,5.1107416,4.691947,4.274966,4.313038,4.349297,4.3873696,4.4254417,4.461701,4.9258194,5.388125,5.8504305,6.3127356,6.775041,7.690587,8.604321,9.519867,10.435412,11.349146,12.32452,13.299893,14.275268,15.250641,16.224201,15.292339,14.3604765,13.426801,12.494938,11.563075,11.612025,11.662788,11.711739,11.762501,11.813264,9.973107,8.13295,6.2927933,4.4526362,2.612479,2.8699198,3.1273603,3.3848011,3.6422417,3.8996825,3.3376641,2.7756457,2.2118144,1.649796,1.0877775,1.2255627,1.3633479,1.49932,1.6371052,1.7748904,1.79302,1.8093367,1.8274662,1.845596,1.8619126,3.4228733,4.9820213,6.542982,8.10213,9.663091,8.040489,6.4178877,4.795286,3.1726844,1.550083,3.8180993,6.0843024,8.352319,10.620335,12.888351,11.820516,10.752681,9.684846,8.617011,7.549176,7.271793,6.9944096,6.717026,6.439643,6.16226,5.1651306,4.168001,3.1708715,2.1719291,1.1747998,2.0178273,2.8608549,3.7020695,4.5450974,5.388125,5.0617914,4.7372713,4.4127507,4.0882306,3.7618973,6.452334,9.142771,11.833207,14.521831,17.212267,14.889862,12.567456,10.245051,7.9226465,5.600241,9.300498,13.000754,16.699198,20.399454,24.099712,25.370598,26.639671,27.910559,29.179632,30.45052,27.277836,24.10515,20.932467,17.75978,14.587097,15.4246855,16.262274,17.099863,17.937452,18.77504,15.865235,12.955431,10.045626,7.135821,4.2242026,7.137634,10.049252,12.962683,15.8743,18.787731,17.834112,16.882307,15.930502,14.976884,14.025079,11.220426,8.415772,5.6093063,2.8046532,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.31182957,0.6000906,0.8883517,1.1747998,1.4630609,1.9670644,2.472881,2.9768846,3.482701,3.9867048,3.5969179,3.207131,2.817344,2.427557,2.03777,3.1708715,4.3021603,5.4352617,6.5683637,7.699652,7.996978,8.294304,8.59163,8.890768,9.188094,7.844689,6.5030966,5.1596913,3.8180993,2.474694,2.9877625,3.5008307,4.0120864,4.5251546,5.038223,4.8678045,4.6973863,4.5269675,4.358362,4.1879435,4.3529234,4.517903,4.6828823,4.847862,5.0128417,4.7191415,4.4272547,4.135368,3.8416677,3.5497808,2.857229,2.1646774,1.4721256,0.7795739,0.0870222,0.10333887,0.11784257,0.13234627,0.14684997,0.16316663,0.14684997,0.13234627,0.11784257,0.10333887,0.0870222,0.18310922,0.27738327,0.37165734,0.46774435,0.5620184,0.49675176,0.43329805,0.3680314,0.30276474,0.2374981,0.9318628,1.6280404,2.322405,3.0167696,3.7129474,2.9768846,2.2426348,1.5083848,0.77232206,0.038072214,0.06164073,0.0870222,0.11240368,0.13778515,0.16316663,0.22480737,0.28826106,0.34990177,0.41335547,0.4749962,0.9554313,1.4358664,1.9144884,2.3949237,2.8753586,3.054842,3.2343252,3.4156215,3.5951047,3.774588,3.43919,3.105605,2.770207,2.4348087,2.0994108,1.8655385,1.6298534,1.3941683,1.1602961,0.9246109,0.7705091,0.61459434,0.4604925,0.3045777,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.05076295,0.06164073,0.07433146,0.0870222,0.099712946,0.099712946,0.099712946,0.099712946,0.099712946,0.099712946,0.13234627,0.16497959,0.19761293,0.23024625,0.26287958,0.3045777,0.3480888,0.38978696,0.43329805,0.4749962,0.44780177,0.42060733,0.39159992,0.36440548,0.33721104,0.3245203,0.31182957,0.2991388,0.28826106,0.2755703,0.26469254,0.25562772,0.24474995,0.23568514,0.22480737,1.162109,2.0994108,3.0367124,3.975827,4.9131284,4.7916603,4.6720047,4.552349,4.4326935,4.313038,3.4555066,2.5979755,1.7404441,0.88291276,0.025381476,0.58014804,1.1349145,1.6896812,2.2444477,2.7992141,6.1785765,9.554313,12.931862,16.309412,19.68696,18.048042,16.40731,14.766581,13.127662,11.486931,9.570629,7.652515,5.7344007,3.8180993,1.8999848,1.7495089,1.6008459,1.4503701,1.2998942,1.1494182,1.6226015,2.0957847,2.5671551,3.0403383,3.5117085,5.8359265,8.158332,10.480737,12.803142,15.125546,12.919171,10.714609,8.510046,6.305484,4.099108,3.299592,2.5000753,1.7005589,0.89922947,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.38072214,0.6979906,1.015259,1.3325275,1.649796,1.8673514,2.084907,2.3024626,2.520018,2.7375734,3.5243993,4.313038,5.0998635,5.8866897,6.6753283,2.811905,3.0348995,3.2578938,3.4808881,3.7020695,3.925064,4.5324063,5.139749,5.7470913,6.354434,6.9617763,9.072064,11.182353,13.292642,15.40293,17.513218,18.537542,19.561867,20.588003,21.612328,22.63665,21.646772,20.656897,19.667019,18.677141,17.687263,17.493277,17.297476,17.101677,16.907688,16.71189,18.147755,19.581808,21.017675,22.451729,23.887594,28.22239,32.557182,36.891975,41.22677,45.563377,38.4475,31.333433,24.217554,17.101677,9.987611,8.734854,7.4820967,6.2293396,4.976582,3.7256382,3.540716,3.3557937,3.1708715,2.9841363,2.7992141,3.4174345,4.0356545,4.652062,5.2702823,5.8866897,6.8004227,7.7123427,8.624263,9.537996,10.449916,8.477413,6.5049095,4.5324063,2.5599031,0.5873999,0.46955732,0.35171473,0.23568514,0.11784257,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.28282216,0.5656443,0.8466535,1.1294757,1.4122978,1.405046,1.3977941,1.3905423,1.3832904,1.3742256,1.1004683,0.824898,0.5493277,0.2755703,0.0,1.8619126,3.7256382,5.5875506,7.4494634,9.313189,9.655839,9.9966755,10.339326,10.681975,11.024626,11.195044,11.365462,11.535881,11.704487,11.874905,11.787883,11.700861,11.612025,11.525003,11.437981,10.879588,10.323009,9.764616,9.208037,8.649645,8.6877165,8.725789,8.762048,8.80012,8.838193,8.727602,8.617011,8.508233,8.397643,8.287052,8.39039,8.491917,8.595256,8.696781,8.80012,9.915092,11.030065,12.145037,13.260008,14.37498,14.911617,15.4500675,15.986704,16.525154,17.06179,16.372866,15.682126,14.9932,14.302462,13.611723,13.571837,13.531953,13.492067,13.452183,13.412297,12.621845,11.833207,11.042755,10.252303,9.461852,7.9734097,6.4831543,4.992899,3.5026438,2.0123885,1.983381,1.9525607,1.9217403,1.892733,1.8619126,1.7803292,1.696933,1.6153497,1.5319533,1.4503701,2.1973107,2.9442513,3.6930048,4.439945,5.186886,5.130684,5.0726695,5.0146546,4.95664,4.900438,5.33011,5.7597823,6.189454,6.6191263,7.0506115,12.087022,17.125244,22.163467,27.199877,32.238102,30.145943,28.05197,25.959812,23.867653,21.775494,20.560808,19.34431,18.129625,16.914942,15.700256,15.854358,16.010273,16.164375,16.32029,16.474392,14.617917,12.75963,10.903157,9.04487,7.1883965,7.217404,7.2482243,7.2772317,7.308052,7.3370595,7.380571,7.422269,7.46578,7.507478,7.549176,6.972654,6.394319,5.8177967,5.239462,4.6629395,5.0726695,5.482399,5.8921285,6.301858,6.7134004,6.0843024,5.4570174,4.8297324,4.2024474,3.5751622,3.636803,3.7002566,3.7618973,3.825351,3.8869917,4.3746786,4.8623657,5.3500524,5.8377395,6.3254266,7.369693,8.415772,9.460039,10.504305,11.5503845,11.9873085,12.4242325,12.862969,13.299893,13.736817,13.04064,12.342649,11.644659,10.946668,10.25049,10.161655,10.074633,9.987611,9.900589,9.811753,8.354132,6.8983226,5.4407005,3.9830787,2.525457,2.4094272,2.2952106,2.179181,2.0649643,1.9507477,1.7748904,1.6008459,1.4249886,1.2491312,1.0750868,1.3125849,1.550083,1.7875811,2.0250793,2.2625773,2.0142014,1.7676386,1.5192627,1.2726997,1.0243238,2.5798457,4.135368,5.6908894,7.2445984,8.80012,7.4331465,6.0643597,4.6973863,3.3304121,1.9616255,3.6023567,5.243088,6.882006,8.5227375,10.161655,9.672155,9.182655,8.693155,8.201842,7.7123427,7.36788,7.023417,6.677141,6.3326783,5.9882154,4.9076896,3.827164,2.7466383,1.6679256,0.5873999,1.015259,1.4431182,1.8691645,2.2970235,2.7248828,2.5997884,2.474694,2.3495996,2.2245052,2.0994108,4.2822175,6.4650245,8.647832,10.830639,13.011633,11.156972,9.302311,7.4476504,5.5929894,3.738329,8.887142,14.037769,19.188396,24.33721,29.487837,26.73576,23.981869,21.229792,18.477715,15.725637,16.356548,16.989273,17.621996,18.25472,18.887444,16.98746,15.087475,13.1874895,11.287505,9.38752,8.482852,7.5781837,6.6717024,5.767034,4.8623657,8.899834,12.937301,16.97477,21.012236,25.049704,21.441908,17.835926,14.22813,10.620335,7.0125394,5.6093063,4.207886,2.8046532,1.403233,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.40066472,0.7868258,1.1747998,1.5627737,1.9507477,2.5907235,3.2306993,3.870675,4.510651,5.1506267,4.454449,3.7600844,3.0657198,2.3695421,1.6751775,3.1346123,4.59586,6.055295,7.51473,8.974165,8.841819,8.709473,8.577126,8.444779,8.312433,7.1466985,5.9827766,4.8170414,3.6531196,2.4873846,2.6995013,2.911618,3.1255474,3.3376641,3.5497808,3.4283123,3.3050308,3.1817493,3.0602808,2.9369993,3.4953918,4.0519714,4.610364,5.1669436,5.7253356,5.4479527,5.1705694,4.893186,4.615803,4.3366065,3.484514,2.6324217,1.7803292,0.92823684,0.07433146,0.09427405,0.11421664,0.13415924,0.15410182,0.17585737,0.15410182,0.13415924,0.11421664,0.09427405,0.07433146,0.21030366,0.3444629,0.48043507,0.61459434,0.7505665,0.629098,0.5094425,0.38978696,0.27013144,0.15047589,0.72337204,1.2944553,1.8673514,2.4402475,3.0131438,2.420305,1.8274662,1.2346275,0.6417888,0.05076295,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.19942589,0.28826106,0.37528324,0.46230546,0.5493277,0.8901646,1.2291887,1.5700256,1.9108626,2.2498865,2.5780327,2.904366,3.2325122,3.5606585,3.8869917,3.4700103,3.053029,2.6342347,2.2172532,1.8002719,1.5954071,1.3905423,1.1856775,0.9808127,0.774135,0.64722764,0.52032024,0.39159992,0.26469254,0.13778515,0.11059072,0.08339628,0.054388877,0.027194439,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.11240368,0.11240368,0.11240368,0.11240368,0.11240368,0.14684997,0.18310922,0.21755551,0.2520018,0.28826106,0.32814622,0.3680314,0.40791658,0.44780177,0.48768693,0.4550536,0.4224203,0.38978696,0.35715362,0.3245203,0.3245203,0.3245203,0.3245203,0.3245203,0.3245203,0.3208944,0.3154555,0.3100166,0.3045777,0.2991388,1.550083,2.7992141,4.0501585,5.2992897,6.550234,6.390693,6.2293396,6.069799,5.910258,5.750717,4.603112,3.4555066,2.3079014,1.1602961,0.012690738,0.5529536,1.0932164,1.6316663,2.1719291,2.712192,6.5194135,10.326634,14.13567,17.94289,21.750113,20.054993,18.359873,16.664753,14.969632,13.274512,10.997431,8.72035,6.4432693,4.164375,1.887294,1.8002719,1.7132497,1.6244144,1.5373923,1.4503701,1.7803292,2.1102884,2.4402475,2.770207,3.100166,5.3428006,7.5854354,9.82807,12.070704,14.313339,12.284635,10.257742,8.229037,6.202145,4.175253,3.3630457,2.5490253,1.7368182,0.9246109,0.11240368,0.09064813,0.06707962,0.045324065,0.02175555,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.4894999,0.91735905,1.3452182,1.7730774,2.1991236,2.427557,2.6541772,2.8826106,3.1092308,3.3376641,3.9631362,4.5867953,5.2122674,5.8377395,6.4632115,3.000453,3.2379513,3.4754493,3.7129474,3.9504454,4.1879435,4.974769,5.7615952,6.550234,7.3370595,8.125698,10.362894,12.60009,14.837286,17.074482,19.311678,20.350506,21.38752,22.424534,23.463362,24.500376,23.187792,21.875206,20.562622,19.250036,17.937452,17.487837,17.038223,16.586794,16.13718,15.687565,17.524096,19.36244,21.200785,23.037315,24.87566,29.01284,33.15002,37.2872,41.42438,45.563377,37.736816,29.91207,22.087322,14.262577,6.43783,5.962834,5.487838,5.0128417,4.537845,4.062849,3.6241121,3.1871881,2.7502642,2.3133402,1.8746033,2.8245957,3.774588,4.7245803,5.674573,6.624565,7.899078,9.175404,10.449916,11.724429,13.000754,10.536939,8.074935,5.612932,3.149116,0.6871128,0.5493277,0.41335547,0.2755703,0.13778515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.33721104,0.6744221,1.0116332,1.3506571,1.6878681,1.6117238,1.5373923,1.4630609,1.3869164,1.3125849,1.0497054,0.7868258,0.52575916,0.26287958,0.0,1.8492218,3.7002566,5.5494785,7.400513,9.249735,9.6504,10.049252,10.449916,10.850581,11.249433,11.249433,11.249433,11.249433,11.249433,11.249433,11.175101,11.10077,11.024626,10.950294,10.874149,10.28675,9.699349,9.11195,8.52455,7.93715,8.024173,8.113008,8.200029,8.287052,8.375887,8.46291,8.549932,8.636953,8.725789,8.812811,8.899834,8.9868555,9.07569,9.162713,9.249735,10.388275,11.525003,12.661731,13.800271,14.936998,15.636803,16.336605,17.038223,17.738026,18.43783,17.712645,16.98746,16.262274,15.537089,14.811904,14.538147,14.262577,13.987006,13.713249,13.437678,12.699803,11.961927,11.225864,10.487988,9.750113,8.113008,6.4759026,4.836984,3.199879,1.5627737,1.6371052,1.7132497,1.7875811,1.8619126,1.938057,1.8002719,1.6624867,1.5247015,1.3869164,1.2491312,2.1501737,3.049403,3.9504454,4.8496747,5.750717,5.275721,4.800725,4.325729,3.8507326,3.3757362,3.9993954,4.6248674,5.2503395,5.8758116,6.4994707,12.311829,18.124187,23.938358,29.750715,35.563072,32.800117,30.037165,27.27421,24.513067,21.750113,20.662334,19.574556,18.48678,17.400814,16.313038,16.525154,16.73727,16.949387,17.163317,17.375433,15.27421,13.174799,11.075388,8.974165,6.874754,6.688019,6.4994707,6.3127356,6.1241875,5.9374523,6.187641,6.43783,6.688019,6.9382076,7.1883965,6.7496595,6.3127356,5.8758116,5.4370747,5.0001507,5.411693,5.825049,6.2384043,6.6499467,7.063302,6.2257137,5.388125,4.550536,3.7129474,2.8753586,2.962381,3.049403,3.1382382,3.2252605,3.3122826,3.825351,4.3366065,4.8496747,5.3627434,5.8758116,7.0506115,8.225411,9.400211,10.57501,11.74981,11.650098,11.5503845,11.450671,11.349146,11.249433,10.7871275,10.324821,9.862516,9.400211,8.937905,8.713099,8.488291,8.26167,8.036863,7.8120556,6.736969,5.661882,4.5867953,3.5117085,2.4366217,1.9507477,1.4630609,0.97537386,0.48768693,0.0,0.21211663,0.42423326,0.63816285,0.85027945,1.062396,1.3996071,1.7368182,2.0758421,2.4130533,2.7502642,2.2371957,1.7241274,1.2128719,0.69980353,0.18673515,1.7368182,3.2869012,4.836984,6.3870673,7.93715,6.825804,5.712645,4.599486,3.48814,2.374981,3.386614,4.40006,5.411693,6.4251394,7.4367723,7.5256076,7.61263,7.699652,7.7866745,7.8755093,7.462154,7.0506115,6.637256,6.2257137,5.812358,4.650249,3.48814,2.324218,1.162109,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.13778515,0.21211663,0.28826106,0.36259252,0.43692398,2.1121013,3.787279,5.462456,7.137634,8.812811,7.424082,6.037165,4.650249,3.2633326,1.8746033,8.4756,15.074784,21.675781,28.274965,34.87415,28.099108,21.325878,14.549025,7.7757964,1.0007553,5.4370747,9.875207,14.313339,18.749659,23.187792,18.550234,13.912675,9.275117,4.6375585,0.0,1.1004683,2.1991236,3.299592,4.40006,5.5005283,10.662033,15.825351,20.986855,26.150173,31.311676,25.049704,18.787731,12.523946,6.261973,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.48768693,0.97537386,1.4630609,1.9507477,2.4366217,3.2125697,3.9867048,4.762653,5.5367875,6.3127356,5.3119802,4.313038,3.3122826,2.3133402,1.3125849,3.100166,4.8877473,6.6753283,8.46291,10.25049,9.686659,9.12464,8.562622,8.000604,7.4367723,6.450521,5.462456,4.4743915,3.48814,2.5000753,2.4130533,2.324218,2.2371957,2.1501737,2.0631514,1.987007,1.9126755,1.8383441,1.7621996,1.6878681,2.6378605,3.587853,4.537845,5.487838,6.43783,6.1749506,5.9120708,5.6491914,5.388125,5.125245,4.1117992,3.100166,2.08672,1.0750868,0.06164073,0.0870222,0.11240368,0.13778515,0.16316663,0.18673515,0.16316663,0.13778515,0.11240368,0.0870222,0.06164073,0.2374981,0.41335547,0.5873999,0.76325727,0.93730164,0.76325727,0.5873999,0.41335547,0.2374981,0.06164073,0.51306844,0.96268314,1.4122978,1.8619126,2.3133402,1.8619126,1.4122978,0.96268314,0.51306844,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.17585737,0.28826106,0.40066472,0.51306844,0.62547207,0.824898,1.0243238,1.2255627,1.4249886,1.6244144,2.0994108,2.5744069,3.049403,3.5243993,3.9993954,3.5008307,3.000453,2.5000753,1.9996977,1.49932,1.3252757,1.1494182,0.97537386,0.7995165,0.62547207,0.52575916,0.42423326,0.3245203,0.22480737,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.16316663,0.19942589,0.2374981,0.2755703,0.31182957,0.34990177,0.387974,0.42423326,0.46230546,0.50037766,0.46230546,0.42423326,0.387974,0.34990177,0.31182957,0.3245203,0.33721104,0.34990177,0.36259252,0.37528324,0.37528324,0.37528324,0.37528324,0.37528324,0.37528324,1.938057,3.5008307,5.0617914,6.624565,8.187339,7.987913,7.7866745,7.5872483,7.3878226,7.1883965,5.750717,4.313038,2.8753586,1.4376793,0.0,0.52575916,1.0497054,1.5754645,2.0994108,2.6251698,6.8620634,11.10077,15.337664,19.574556,23.813263,22.061941,20.312433,18.562923,16.813416,15.062093,12.4242325,9.788185,7.1503243,4.512464,1.8746033,1.8492218,1.8256533,1.8002719,1.7748904,1.7495089,1.938057,2.124792,2.3133402,2.5000753,2.6868105,4.8496747,7.0125394,9.175404,11.338268,13.499319,11.650098,9.799063,7.949841,6.1006193,4.249584,3.4246864,2.5997884,1.7748904,0.9499924,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.6000906,1.1367276,1.6751775,2.2118144,2.7502642,2.9877625,3.2252605,3.4627585,3.7002566,3.9377546,4.40006,4.8623657,5.3246713,5.7869763,6.249282,3.000453,3.245203,3.489953,3.7347028,3.9794528,4.2242026,5.032784,5.8395524,6.6481338,7.454902,8.26167,10.440851,12.618219,14.795588,16.972956,19.150324,20.209093,21.269676,22.33026,23.390842,24.449614,23.160597,21.869768,20.580751,19.289923,18.000906,17.185072,16.36924,15.555219,14.739386,13.925365,16.965704,20.004229,23.044567,26.084906,29.125244,31.759478,34.395527,37.029762,39.66581,42.30004,34.982925,27.66581,20.34688,13.029762,5.712645,5.424384,5.137936,4.8496747,4.5632267,4.274966,3.787279,3.299592,2.811905,2.324218,1.8383441,2.904366,3.972201,5.040036,6.107871,7.175706,8.01692,8.859948,9.702975,10.54419,11.3872175,9.275117,7.1630154,5.049101,2.9369993,0.824898,0.65991837,0.4949388,0.32995918,0.16497959,0.0,0.058014803,0.11421664,0.17223145,0.23024625,0.28826106,0.23024625,0.17223145,0.11421664,0.058014803,0.0,0.3100166,0.6200332,0.9300498,1.2400664,1.550083,1.5627737,1.5754645,1.5881553,1.6008459,1.6117238,1.2926424,0.97174793,0.6526665,0.33177215,0.012690738,1.8582866,3.7020695,5.5476656,7.3932614,9.237044,9.699349,10.161655,10.625773,11.088079,11.5503845,11.6881695,11.8241415,11.961927,12.099712,12.237497,12.337211,12.436923,12.536636,12.638163,12.737875,12.125093,11.512312,10.899531,10.28675,9.675781,9.550687,9.425592,9.300498,9.175404,9.050309,8.927028,8.805559,8.682278,8.560809,8.437528,8.609759,8.781991,8.954222,9.128266,9.300498,10.339326,11.379966,12.420607,13.4594345,14.500074,15.23795,15.975826,16.71189,17.449764,18.187641,17.741652,17.297476,16.8533,16.40731,15.963136,15.584227,15.20713,14.830034,14.452938,14.075842,13.254569,12.43511,11.615651,10.794379,9.97492,8.306994,6.640882,4.972956,3.3050308,1.6371052,1.7331922,1.8274662,1.9217403,2.0178273,2.1121013,2.0142014,1.9181144,1.8202144,1.7223145,1.6244144,2.3296568,3.0348995,3.7401419,4.445384,5.1506267,4.8170414,4.4852695,4.1516843,3.8199122,3.48814,4.1444325,4.802538,5.4606433,6.1169357,6.775041,12.522133,18.269224,24.018127,29.765219,35.51231,32.560806,29.607492,26.654177,23.702673,20.749357,19.822933,18.894695,17.968271,17.040035,16.1118,16.15531,16.197008,16.240519,16.282217,16.325727,14.313339,12.300951,10.28675,8.274362,6.261973,6.249282,6.2384043,6.2257137,6.2130227,6.200332,6.58468,6.970841,7.3551893,7.7395372,8.125698,7.6416373,7.159389,6.677141,6.1948934,5.712645,6.0643597,6.4178877,6.7696023,7.12313,7.474845,6.4831543,5.4896507,4.49796,3.5044568,2.5127661,2.5744069,2.6378605,2.6995013,2.762955,2.8245957,3.5044568,4.1843176,4.8641787,5.5458527,6.2257137,7.1448855,8.06587,8.985043,9.904215,10.825199,10.680162,10.535126,10.390089,10.245051,10.100015,10.165281,10.230548,10.2958145,10.359268,10.424535,9.8878975,9.349448,8.812811,8.274362,7.7377243,6.736969,5.7380266,4.7372713,3.738329,2.7375734,2.2843328,1.8329052,1.3796645,0.92823684,0.4749962,1.0478923,1.6207886,2.1918716,2.764768,3.3376641,3.1128569,2.8880494,2.663242,2.4366217,2.2118144,1.840157,1.4666867,1.0950294,0.72337204,0.34990177,1.6298534,2.909805,4.1897564,5.469708,6.7496595,5.823236,4.894999,3.966762,3.0403383,2.1121013,3.105605,4.0972953,5.090799,6.0824895,7.07418,7.0850577,7.0941224,7.1050005,7.115878,7.124943,6.697084,6.2692246,5.8431783,5.4153194,4.98746,3.9903307,2.9932013,1.9942589,0.99712944,0.0,0.045324065,0.09064813,0.13415924,0.1794833,0.22480737,0.2755703,0.3245203,0.37528324,0.42423326,0.4749962,2.1084754,3.7401419,5.371808,7.0052876,8.636953,7.5292335,6.4233265,5.315606,4.207886,3.100166,8.669587,14.239008,19.810242,25.379663,30.949083,24.939114,18.930956,12.919171,6.9092,0.89922947,4.6629395,8.424837,12.186734,15.950445,19.712341,15.939567,12.166792,8.394017,4.6230545,0.85027945,1.5627737,2.275268,2.9877625,3.7002566,4.4127507,8.540867,12.66717,16.795286,20.9234,25.049704,20.042301,15.034899,10.027496,5.0200934,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.027194439,0.04169814,0.058014803,0.072518505,0.0870222,0.5058166,0.922798,1.3397794,1.7567607,2.175555,2.7502642,3.3249733,3.8996825,4.4743915,5.049101,4.459888,3.870675,3.2796493,2.6904364,2.0994108,3.7981565,5.4950895,7.192023,8.890768,10.587702,9.795437,9.003172,8.209095,7.41683,6.624565,5.772473,4.9203806,4.068288,3.2143826,2.3622901,2.2408218,2.1175404,1.9942589,1.8727903,1.7495089,1.9978848,2.2444477,2.4928236,2.7393866,2.9877625,3.6930048,4.3982472,5.101677,5.806919,6.5121617,6.281915,6.051669,5.823236,5.5929894,5.3627434,4.7300196,4.0972953,3.4645715,2.8318477,2.1991236,1.794833,1.3905423,0.98443866,0.58014804,0.17585737,0.15228885,0.13053331,0.10696479,0.08520924,0.06164073,0.5166943,0.97174793,1.4268016,1.8818551,2.3369088,1.8818551,1.4268016,0.97174793,0.5166943,0.06164073,0.65810543,1.2527572,1.8474089,2.4420607,3.0367124,2.4801328,1.9217403,1.3651608,0.80676836,0.25018883,0.6200332,0.9898776,1.3597219,1.7295663,2.0994108,2.228131,2.3550384,2.4819458,2.610666,2.7375734,2.8155308,2.8916752,2.9696326,3.04759,3.1255474,3.6857529,4.2441454,4.804351,5.3645563,5.924762,5.424384,4.9258194,4.4254417,3.925064,3.4246864,2.8499773,2.275268,1.7005589,1.1258497,0.5493277,0.4604925,0.36984438,0.27919623,0.19036107,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.065266654,0.07977036,0.09427405,0.11059072,0.12509441,0.13415924,0.14503701,0.15410182,0.16497959,0.17585737,0.21574254,0.25562772,0.2955129,0.33539808,0.37528324,0.41335547,0.44961473,0.48768693,0.52575916,0.5620184,0.5275721,0.49312583,0.45686656,0.4224203,0.387974,0.40066472,0.41335547,0.42423326,0.43692398,0.44961473,1.1729867,1.8945459,2.617918,3.339477,4.062849,5.382686,6.7025228,8.02236,9.342196,10.662033,10.477111,10.292189,10.107266,9.922344,9.737422,8.254418,6.773228,5.290225,3.8072214,2.324218,2.762955,3.199879,3.636803,4.07554,4.512464,7.8247466,11.137029,14.449312,17.761595,21.07569,19.797552,18.519413,17.243088,15.964949,14.68681,12.618219,10.547816,8.477413,6.4070096,4.3366065,3.9903307,3.6422417,3.294153,2.9478772,2.5997884,3.0729716,3.5443418,4.017525,4.4907084,4.9620786,6.5973706,8.232663,9.867955,11.503247,13.136727,11.193231,9.247922,7.3026133,5.3573046,3.4119956,2.7502642,2.08672,1.4249886,0.76325727,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.13053331,0.19761293,0.26469254,0.33177215,0.40066472,1.0279498,1.6552348,2.2825198,2.909805,3.53709,3.7492065,3.9631362,4.175253,4.3873696,4.599486,4.764466,4.9294453,5.0944247,5.2594047,5.424384,3.000453,3.2524548,3.5044568,3.7582715,4.0102735,4.262275,5.090799,5.91751,6.7442207,7.572745,8.399456,10.516996,12.634536,14.752076,16.869617,18.987158,20.069496,21.151834,22.234173,23.318325,24.400663,23.133402,21.864328,20.597069,19.329807,18.062546,16.882307,15.702069,14.521831,13.341592,12.163166,16.405499,20.647831,24.890163,29.132496,33.37483,34.50793,35.639217,36.77232,37.905422,39.03671,32.227222,25.417736,18.606436,11.7969475,4.98746,4.8877473,4.788034,4.688321,4.5867953,4.4870825,3.9504454,3.4119956,2.8753586,2.3369088,1.8002719,2.9841363,4.169814,5.3554916,6.539356,7.7250338,8.134763,8.544493,8.954222,9.365765,9.775495,8.013294,6.249282,4.4870825,2.7248828,0.96268314,0.7705091,0.57833505,0.38434806,0.19217403,0.0,0.11421664,0.23024625,0.3444629,0.4604925,0.5747091,0.4604925,0.3444629,0.23024625,0.11421664,0.0,0.28282216,0.5656443,0.8466535,1.1294757,1.4122978,1.5120108,1.6117238,1.7132497,1.8129625,1.9126755,1.5355793,1.1566701,0.7795739,0.40247768,0.025381476,1.8655385,3.7056956,5.5458527,7.3841968,9.224354,9.750113,10.275872,10.799818,11.325577,11.849524,12.125093,12.400664,12.674421,12.949992,13.225562,13.499319,13.77489,14.05046,14.324218,14.599788,13.961625,13.325275,12.687112,12.050762,11.4126,11.075388,10.738177,10.399154,10.061942,9.724731,9.39296,9.059374,8.727602,8.39583,8.062244,8.319685,8.577126,8.834567,9.092008,9.349448,10.292189,11.234929,12.17767,13.12041,14.06315,14.837286,15.613234,16.38737,17.163317,17.937452,17.772472,17.607492,17.442513,17.277533,17.112555,16.632118,16.151684,15.673061,15.192626,14.712192,13.809336,12.908294,12.005438,11.102583,10.199727,8.502794,6.8058615,5.1071157,3.4101827,1.7132497,1.8274662,1.9416829,2.0577126,2.1719291,2.2879589,2.229944,2.1719291,2.1157274,2.0577126,1.9996977,2.5091403,3.0203958,3.529838,4.0392804,4.550536,4.360175,4.169814,3.9794528,3.7890918,3.6005437,4.2894692,4.9802084,5.669134,6.359873,7.0506115,12.732436,18.41426,24.097898,29.779724,35.46336,32.319683,29.17782,26.034143,22.892279,19.750414,18.981718,18.214834,17.447952,16.679256,15.912373,15.785465,15.656745,15.529838,15.40293,15.27421,13.3506565,11.42529,9.499924,7.574558,5.6491914,5.812358,5.975525,6.1368785,6.300045,6.4632115,6.981719,7.502039,8.02236,8.54268,9.063,8.535428,8.007855,7.4802837,6.9527116,6.4251394,6.717026,7.0107265,7.3026133,7.5945,7.8882003,6.740595,5.5929894,4.445384,3.2977788,2.1501737,2.1882458,2.2245052,2.2625773,2.3006494,2.3369088,3.1853752,4.0320287,4.880495,5.727149,6.5756154,7.2391596,7.9045167,8.569874,9.235231,9.900589,9.710228,9.519867,9.329506,9.139144,8.950596,9.541622,10.13446,10.7273,11.320138,11.912977,11.062697,10.212419,9.362139,8.511859,7.663393,6.736969,5.812358,4.8877473,3.9631362,3.0367124,2.619731,2.2027495,1.7857682,1.3669738,0.9499924,1.8818551,2.8155308,3.7473936,4.6792564,5.612932,4.8242936,4.0374675,3.2506418,2.4620032,1.6751775,1.4431182,1.209246,0.97718686,0.7451276,0.51306844,1.5228885,2.5327086,3.5425289,4.552349,5.562169,4.8206677,4.077353,3.3358512,2.5925364,1.8492218,2.8227828,3.7945306,4.7680917,5.7398396,6.7134004,6.644508,6.5774283,6.510349,6.4432693,6.3743763,5.9320135,5.4896507,5.047288,4.604925,4.162562,3.3304121,2.4982624,1.6642996,0.8321498,0.0,0.07795739,0.15410182,0.23205921,0.3100166,0.387974,0.41335547,0.43692398,0.46230546,0.48768693,0.51306844,2.1030366,3.6930048,5.282973,6.872941,8.46291,7.6343856,6.8076744,5.979151,5.1524396,4.325729,8.865387,13.4050455,17.944704,22.484362,27.025833,21.77912,16.536032,11.289318,6.0444174,0.7995165,3.8869917,6.9744673,10.061942,13.149418,16.236893,13.328901,10.422722,7.51473,4.606738,1.7005589,2.0250793,2.3495996,2.6741197,3.000453,3.3249733,6.4178877,9.508988,12.601903,15.694818,18.787731,15.034899,11.282066,7.5292335,3.778214,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.054388877,0.08520924,0.11421664,0.14503701,0.17585737,0.52213323,0.87022203,1.2183108,1.5645868,1.9126755,2.2879589,2.663242,3.0367124,3.4119956,3.787279,3.6077955,3.4283123,3.247016,3.0675328,2.8880494,4.494334,6.1024323,7.71053,9.316814,10.924912,9.902402,8.87989,7.85738,6.834869,5.812358,5.0944247,4.3783045,3.6603715,2.9424384,2.2245052,2.0667772,1.9108626,1.7531348,1.5954071,1.4376793,2.0069497,2.5780327,3.147303,3.7183862,4.2876563,4.748149,5.2068286,5.667321,6.1278133,6.588306,6.390693,6.19308,5.995467,5.7978544,5.600241,5.3482394,5.0944247,4.842423,4.590421,4.3384194,3.5026438,2.666868,1.8329052,0.99712944,0.16316663,0.14322405,0.12328146,0.10333887,0.08339628,0.06164073,0.79770356,1.5319533,2.268016,3.002266,3.738329,3.002266,2.268016,1.5319533,0.79770356,0.06164073,0.8031424,1.5428312,2.2825198,3.0222087,3.7618973,3.0983531,2.4329958,1.7676386,1.1022812,0.43692398,1.1784257,1.9181144,2.657803,3.397492,4.137181,4.2804046,4.421816,4.5650396,4.708264,4.8496747,4.804351,4.76084,4.7155156,4.670192,4.6248674,5.2702823,5.915697,6.5592985,7.2047133,7.850128,7.3497505,6.849373,6.350808,5.8504305,5.3500524,4.3746786,3.3993049,2.4257438,1.4503701,0.4749962,0.39522585,0.3154555,0.23568514,0.15410182,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.054388877,0.072518505,0.09064813,0.10696479,0.12509441,0.14503701,0.16497959,0.18492219,0.20486477,0.22480737,0.26831847,0.3100166,0.35171473,0.39522585,0.43692398,0.4749962,0.51306844,0.5493277,0.5873999,0.62547207,0.59283876,0.56020546,0.5275721,0.4949388,0.46230546,0.4749962,0.48768693,0.50037766,0.51306844,0.52575916,1.9706904,3.4156215,4.860553,6.305484,7.750415,8.827314,9.904215,10.982927,12.059827,13.136727,12.968122,12.797703,12.627284,12.456866,12.28826,10.7599325,9.233418,7.705091,6.1767635,4.650249,5.0001507,5.3500524,5.6999545,6.049856,6.399758,8.78743,11.175101,13.562773,15.950445,18.338116,17.533161,16.728207,15.92325,15.118295,14.313339,12.810393,11.307447,9.804502,8.303369,6.8004227,6.1296263,5.4606433,4.7898474,4.120864,3.4500678,4.207886,4.9657044,5.7217097,6.4795284,7.2373466,8.345067,9.452786,10.560507,11.668227,12.774135,10.734551,8.694968,6.6553855,4.615803,2.5744069,2.0758421,1.5754645,1.0750868,0.5747091,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.24837588,0.36984438,0.49312583,0.61459434,0.73787576,1.455809,2.1719291,2.8898623,3.6077955,4.325729,4.512464,4.699199,4.8877473,5.0744824,5.2630305,5.130684,4.9983377,4.8641787,4.7318325,4.599486,3.000453,3.2597067,3.5207734,3.780027,4.0392804,4.3003473,5.147001,5.995467,6.8421206,7.690587,8.537241,10.594954,12.652666,14.710379,16.768091,18.825804,19.929897,21.035805,22.139898,23.245806,24.349901,23.104395,21.860703,20.615198,19.369692,18.124187,16.579542,15.034899,13.490254,11.94561,10.399154,15.845293,21.28962,26.73576,32.180084,37.624413,37.25457,36.884724,36.51488,36.145035,35.775192,29.473333,23.169662,16.867804,10.564133,4.262275,4.349297,4.4381323,4.5251546,4.612177,4.699199,4.1117992,3.5243993,2.9369993,2.3495996,1.7621996,3.0657198,4.367427,5.669134,6.972654,8.274362,8.252605,8.23085,8.207282,8.185526,8.161958,6.7496595,5.337362,3.925064,2.5127661,1.1004683,0.8792868,0.65991837,0.4405499,0.21936847,0.0,0.17223145,0.3444629,0.5166943,0.69073874,0.8629702,0.69073874,0.5166943,0.3444629,0.17223145,0.0,0.25562772,0.5094425,0.7650702,1.020698,1.2745126,1.4630609,1.649796,1.8383441,2.0250793,2.2118144,1.7767034,1.3434052,0.90829426,0.47318324,0.038072214,1.8727903,3.7075086,5.542227,7.3769445,9.211663,9.800876,10.388275,10.975676,11.563075,12.1504755,12.562017,12.975373,13.386916,13.800271,14.211814,14.663241,15.112856,15.56247,16.012085,16.4617,15.799969,15.138238,14.474693,13.812962,13.149418,12.60009,12.050762,11.499621,10.950294,10.399154,9.857078,9.3150015,8.772926,8.23085,7.686961,8.029612,8.372261,8.714911,9.057561,9.400211,10.245051,11.089892,11.934732,12.779573,13.6244135,14.436621,15.250641,16.062849,16.875055,17.687263,17.803293,17.91751,18.031725,18.147755,18.261972,17.680012,17.09805,16.514277,15.932315,15.350354,14.365915,13.379663,12.395226,11.410787,10.424535,8.696781,6.970841,5.243088,3.5153344,1.7875811,1.9217403,2.0577126,2.1918716,2.327844,2.4620032,2.4456866,2.427557,2.4094272,2.3931105,2.374981,2.6904364,3.005892,3.3195345,3.63499,3.9504454,3.9033084,3.8543584,3.8072214,3.7600844,3.7129474,4.4345064,5.1578784,5.8794374,6.60281,7.324369,12.9427395,18.559298,24.17767,29.794228,35.412598,32.08037,28.748148,25.41411,22.081884,18.749659,18.142317,17.534973,16.927631,16.32029,15.712947,15.415621,15.118295,14.819156,14.521831,14.224504,12.387974,10.549629,8.713099,6.874754,5.038223,5.375434,5.712645,6.049856,6.3870673,6.7242785,7.380571,8.03505,8.689529,9.345822,10.000301,9.427405,8.854509,8.281613,7.71053,7.137634,7.369693,7.6017523,7.835624,8.067683,8.299743,6.9980354,5.6945157,4.3928084,3.0892882,1.7875811,1.8002719,1.8129625,1.8256533,1.8383441,1.8492218,2.864481,3.87974,4.894999,5.910258,6.925517,7.3352466,7.744976,8.154706,8.564435,8.974165,8.740293,8.504607,8.270736,8.03505,7.799365,8.919776,10.040187,11.160598,12.279196,13.399607,12.237497,11.075388,9.91328,8.749357,7.5872483,6.736969,5.8866897,5.038223,4.1879435,3.3376641,2.955129,2.572594,2.1900587,1.8075237,1.4249886,2.7176309,4.0102735,5.3029156,6.5955577,7.8882003,6.5375433,5.186886,3.8380418,2.4873846,1.1367276,1.0442665,0.95180535,0.85934424,0.7668832,0.6744221,1.4141108,2.1556125,2.8953013,3.63499,4.3746786,3.8180993,3.2597067,2.7031271,2.1447346,1.5881553,2.5399606,3.491766,4.445384,5.3971896,6.350808,6.205771,6.060734,5.915697,5.77066,5.6256227,5.1669436,4.710077,4.25321,3.7945306,3.3376641,2.6704938,2.0033236,1.3343405,0.6671702,0.0,0.11059072,0.21936847,0.32995918,0.4405499,0.5493277,0.5493277,0.5493277,0.5493277,0.5493277,0.5493277,2.0975976,3.644055,5.1923246,6.740595,8.287052,7.7395372,7.192023,6.644508,6.096993,5.5494785,9.059374,12.569269,16.080978,19.590874,23.100769,18.619125,14.139296,9.659465,5.179634,0.69980353,3.1128569,5.524097,7.93715,10.3502035,12.763257,10.720048,8.676839,6.635443,4.592234,2.5508385,2.4873846,2.4257438,2.3622901,2.3006494,2.2371957,4.2949085,6.352621,8.410334,10.468046,12.525759,10.027496,7.5292335,5.032784,2.5345216,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.08339628,0.12690738,0.17223145,0.21755551,0.26287958,0.5402629,0.81764615,1.0950294,1.3724127,1.649796,1.8256533,1.9996977,2.175555,2.3495996,2.525457,2.7557032,2.9841363,3.2143826,3.444629,3.6748753,5.1923246,6.7097745,8.227224,9.744674,11.262123,10.009366,8.758422,7.5056653,6.2529078,5.0001507,4.41819,3.834416,3.2524548,2.6704938,2.08672,1.8945459,1.7023718,1.5101979,1.3180238,1.1258497,2.0178273,2.909805,3.8017826,4.695573,5.5875506,5.803293,6.017223,6.2329655,6.446895,6.6626377,6.497658,6.3326783,6.167699,6.002719,5.8377395,5.964647,6.093367,6.2202744,6.347182,6.474089,5.2104545,3.9450066,2.6795588,1.4141108,0.15047589,0.13234627,0.11421664,0.09789998,0.07977036,0.06164073,1.0768998,2.0921588,3.1074178,4.122677,5.137936,4.122677,3.1074178,2.0921588,1.0768998,0.06164073,0.9481794,1.8329052,2.7176309,3.6023567,4.4870825,3.7147603,2.9424384,2.1701162,1.3977941,0.62547207,1.7350051,2.8445382,3.9558845,5.0654173,6.1749506,6.3326783,6.490406,6.6481338,6.8058615,6.9617763,6.794984,6.628191,6.4595857,6.2927933,6.1241875,6.8548117,7.5854354,8.314246,9.04487,9.775495,9.275117,8.774739,8.274362,7.7757964,7.2754188,5.89938,4.5251546,3.149116,1.7748904,0.40066472,0.32995918,0.25925365,0.19036107,0.11965553,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.045324065,0.065266654,0.08520924,0.10515183,0.12509441,0.15410182,0.18492219,0.21574254,0.24474995,0.2755703,0.3208944,0.36440548,0.40972954,0.4550536,0.50037766,0.53663695,0.5747091,0.61278135,0.6508536,0.6871128,0.65810543,0.62728506,0.5982776,0.56745726,0.53663695,0.5493277,0.5620184,0.5747091,0.5873999,0.6000906,2.7683938,4.934884,7.1031876,9.269678,11.437981,12.271944,13.107719,13.941682,14.777458,15.613234,15.457319,15.303217,15.147303,14.9932,14.837286,13.265448,11.691795,10.119957,8.548119,6.9744673,7.2373466,7.500226,7.763106,8.024173,8.287052,9.750113,11.213174,12.674421,14.137483,15.600543,15.266958,14.935185,14.601601,14.269829,13.938056,13.002567,12.067079,11.13159,10.197914,9.262425,8.270736,7.2772317,6.285541,5.292038,4.3003473,5.3428006,6.3852544,7.4277077,8.470161,9.512614,10.092763,10.672911,11.253058,11.833207,12.413355,10.277685,8.1420145,6.008158,3.872488,1.7368182,1.3996071,1.062396,0.72518504,0.387974,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.36440548,0.5420758,0.7197462,0.8974165,1.0750868,1.8818551,2.6904364,3.4972048,4.305786,5.1125546,5.275721,5.4370747,5.600241,5.7615952,5.924762,5.4950895,5.0654173,4.6357455,4.2042603,3.774588,3.000453,3.2669585,3.5352771,3.8017826,4.070101,4.3366065,5.2050157,6.071612,6.9400206,7.806617,8.675026,10.672911,12.670795,14.666867,16.664753,18.662638,19.7903,20.917963,22.045626,23.173288,24.299137,23.0772,21.855265,20.633327,19.409578,18.187641,16.276777,14.367728,12.456866,10.547816,8.636953,15.285088,21.931408,28.579542,35.227676,41.87581,40.00302,38.13023,36.25744,34.384647,32.51186,26.71763,20.9234,15.127359,9.333132,3.53709,3.8126602,4.0882306,4.361988,4.6375585,4.9131284,4.274966,3.636803,3.000453,2.3622901,1.7241274,3.1454902,4.5650396,5.9845896,7.404139,8.825501,8.370448,7.915395,7.460341,7.0052876,6.550234,5.487838,4.4254417,3.3630457,2.3006494,1.2382535,0.9898776,0.7433147,0.4949388,0.24837588,0.0,0.23024625,0.4604925,0.69073874,0.91917205,1.1494182,0.91917205,0.69073874,0.4604925,0.23024625,0.0,0.22662032,0.4550536,0.68167394,0.9101072,1.1367276,1.4122978,1.6878681,1.9616255,2.2371957,2.5127661,2.0196402,1.5283275,1.0352017,0.5420758,0.05076295,1.8800422,3.7093215,5.540414,7.369693,9.200785,9.849826,10.500679,11.14972,11.800573,12.449615,13.000754,13.550082,14.09941,14.650551,15.199879,15.825351,16.450823,17.074482,17.699953,18.325426,17.638313,16.949387,16.262274,15.575162,14.888049,14.124791,13.363347,12.60009,11.836833,11.075388,10.323009,9.570629,8.81825,8.06587,7.311678,7.7395372,8.167397,8.595256,9.023115,9.449161,10.197914,10.944855,11.691795,12.440549,13.1874895,14.037769,14.888049,15.738328,16.586794,17.437075,17.8323,18.227526,18.622751,19.017977,19.413204,18.727903,18.042604,17.357304,16.672005,15.986704,14.920682,13.852847,12.785012,11.717177,10.649343,8.892582,7.135821,5.377247,3.6204863,1.8619126,2.0178273,2.1719291,2.327844,2.4819458,2.6378605,2.659616,2.6831846,2.70494,2.7266958,2.7502642,2.8699198,2.9895754,3.1092308,3.2306993,3.350355,3.444629,3.540716,3.63499,3.729264,3.825351,4.5795436,5.335549,6.089741,6.8457465,7.5999393,13.153044,18.704334,24.257439,29.810543,35.361835,31.839249,28.318476,24.794077,21.273302,17.750717,17.302916,16.855114,16.40731,15.95951,15.511708,15.045776,14.5780325,14.110288,13.642544,13.174799,11.42529,9.675781,7.9244595,6.1749506,4.4254417,4.936697,5.4497657,5.962834,6.4759026,6.987158,7.7776093,8.568061,9.3567,10.147152,10.937603,10.319383,9.702975,9.084756,8.4683485,7.850128,8.02236,8.194591,8.366822,8.540867,8.713099,7.2554765,5.7978544,4.3402324,2.8826106,1.4249886,1.4122978,1.3996071,1.3869164,1.3742256,1.3633479,2.5453994,3.727451,4.9095025,6.093367,7.2754188,7.4295206,7.5854354,7.7395372,7.895452,8.049554,7.7703576,7.4893484,7.210152,6.929143,6.6499467,8.29793,9.944099,11.592083,13.240066,14.888049,13.412297,11.938358,10.462607,8.9868555,7.512917,6.736969,5.962834,5.186886,4.4127507,3.636803,3.290527,2.9424384,2.5943494,2.2480736,1.8999848,3.5515938,5.2050157,6.8584375,8.510046,10.161655,8.2507925,6.338117,4.4254417,2.5127661,0.6000906,0.64722764,0.69436467,0.7433147,0.7904517,0.8375887,1.3071461,1.7767034,2.2480736,2.7176309,3.1871881,2.8155308,2.4420607,2.0704033,1.696933,1.3252757,2.2571385,3.1908143,4.122677,5.0545397,5.9882154,5.765221,5.542227,5.319232,5.0980506,4.8750563,4.401873,3.930503,3.4573197,2.9841363,2.5127661,2.0105755,1.5083848,1.0043813,0.50219065,0.0,0.14322405,0.28463513,0.42785916,0.56927025,0.7124943,0.6871128,0.66173136,0.63816285,0.61278135,0.5873999,2.0921588,3.5969179,5.101677,6.6082487,8.113008,7.844689,7.5781837,7.309865,7.0433598,6.775041,9.255174,11.735307,14.21544,16.695572,19.175705,15.459132,11.744371,8.029612,4.314851,0.6000906,2.3369088,4.07554,5.812358,7.549176,9.287807,8.109382,6.932769,5.754343,4.5777307,3.3993049,2.94969,2.5000753,2.0504606,1.6008459,1.1494182,2.1719291,3.1944401,4.216951,5.239462,6.261973,5.0200934,3.778214,2.5345216,1.2926424,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.11059072,0.17041849,0.23024625,0.29007402,0.34990177,0.55839247,0.7650702,0.97174793,1.1802386,1.3869164,1.3633479,1.3379664,1.3125849,1.2872034,1.261822,1.9017978,2.5417736,3.1817493,3.8217251,4.461701,5.8903155,7.317117,8.745731,10.172533,11.599335,10.118144,8.63514,7.1521373,5.669134,4.1879435,3.7401419,3.29234,2.8445382,2.3967366,1.9507477,1.7223145,1.4956942,1.2672608,1.0406405,0.8122072,2.0268922,3.2415771,4.458075,5.67276,6.887445,6.8566246,6.827617,6.796797,6.7677894,6.736969,6.604623,6.472276,6.33993,6.207584,6.0752378,6.582867,7.0904965,7.5981264,8.105756,8.613385,6.9182653,5.223145,3.5280252,1.8329052,0.13778515,0.12328146,0.10696479,0.092461094,0.07795739,0.06164073,1.357909,2.6523643,3.9468195,5.243088,6.5375433,5.243088,3.9468195,2.6523643,1.357909,0.06164073,1.0932164,2.1229792,3.152742,4.1825047,5.2122674,4.3329806,3.4518807,2.572594,1.693307,0.8122072,2.2933977,3.7727752,5.2521524,6.733343,8.212721,8.384952,8.557183,8.729415,8.901647,9.07569,8.785617,8.495543,8.205468,7.915395,7.6253204,8.439341,9.255174,10.069194,10.885027,11.700861,11.200482,10.700105,10.199727,9.699349,9.200785,7.424082,5.6491914,3.874301,2.0994108,0.3245203,0.26469254,0.20486477,0.14503701,0.08520924,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.034446288,0.058014803,0.07977036,0.10333887,0.12509441,0.16497959,0.20486477,0.24474995,0.28463513,0.3245203,0.37165734,0.42060733,0.46774435,0.5148814,0.5620184,0.6000906,0.63816285,0.6744221,0.7124943,0.7505665,0.72337204,0.69436467,0.6671702,0.6399758,0.61278135,0.62547207,0.63816285,0.6508536,0.66173136,0.6744221,3.5642843,6.454147,9.345822,12.235684,15.125546,15.718386,16.309412,16.90225,17.495089,18.087927,17.94833,17.80692,17.66732,17.527721,17.388124,15.769149,14.151986,12.534823,10.917661,9.300498,9.474543,9.6504,9.824444,10.000301,10.174346,10.712796,11.249433,11.787883,12.32452,12.862969,13.002567,13.142166,13.281764,13.423175,13.562773,13.194741,12.826711,12.460492,12.092461,11.724429,10.410031,9.0956335,7.7794223,6.4650245,5.1506267,6.4777155,7.804804,9.131892,10.460794,11.787883,11.840459,11.893035,11.94561,11.998186,12.050762,9.819005,7.5890613,5.3591175,3.1309865,0.89922947,0.72518504,0.5493277,0.37528324,0.19942589,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,0.48224804,0.71430725,0.9481794,1.1802386,1.4122978,2.3097143,3.207131,4.1045475,5.0019636,5.89938,6.037165,6.1749506,6.3127356,6.450521,6.588306,5.859495,5.132497,4.405499,3.6766882,2.94969,3.000453,3.2742105,3.5497808,3.825351,4.099108,4.3746786,5.2630305,6.149569,7.037921,7.9244595,8.812811,10.750868,12.687112,14.625169,16.563227,18.49947,19.650702,20.80012,21.949537,23.100769,24.250187,23.050007,21.849825,20.649643,19.449463,18.24928,15.975826,13.700559,11.42529,9.1500225,6.874754,14.724882,22.57501,30.425138,38.275265,46.125393,42.749657,39.375732,35.999996,32.62426,29.250338,23.961926,18.675327,13.386916,8.100317,2.811905,3.2742105,3.738329,4.2006345,4.6629395,5.125245,4.4381323,3.7492065,3.0620937,2.374981,1.6878681,3.2252605,4.762653,6.300045,7.837437,9.374829,8.488291,7.5999393,6.7115874,5.825049,4.936697,4.2242026,3.5117085,2.7992141,2.08672,1.3742256,1.1004683,0.824898,0.5493277,0.2755703,0.0,0.28826106,0.5747091,0.8629702,1.1494182,1.4376793,1.1494182,0.8629702,0.5747091,0.28826106,0.0,0.19942589,0.40066472,0.6000906,0.7995165,1.0007553,1.3633479,1.7241274,2.08672,2.4493124,2.811905,2.2625773,1.7132497,1.162109,0.61278135,0.06164073,1.887294,3.7129474,5.5367875,7.362441,9.188094,9.900589,10.613083,11.325577,12.038072,12.750566,13.437678,14.124791,14.811904,15.50083,16.187943,16.98746,17.786976,18.588305,19.387821,20.187338,19.474844,18.76235,18.049856,17.33736,16.624866,15.649493,14.675932,13.700559,12.725184,11.74981,10.7871275,9.824444,8.861761,7.900891,6.9382076,7.4494634,7.9625316,8.4756,8.9868555,9.499924,10.150778,10.799818,11.450671,12.099712,12.750566,13.637105,14.525456,15.411995,16.300346,17.186886,17.863121,18.537542,19.211964,19.888199,20.562622,19.775795,18.987158,18.20033,17.411694,16.624866,15.475449,14.324218,13.174799,12.025381,10.874149,9.088382,7.3008003,5.5132194,3.7256382,1.938057,2.1121013,2.2879589,2.4620032,2.6378605,2.811905,2.8753586,2.9369993,3.000453,3.0620937,3.1255474,3.049403,2.9750717,2.9007401,2.8245957,2.7502642,2.9877625,3.2252605,3.4627585,3.7002566,3.9377546,4.7245803,5.5132194,6.300045,7.0868707,7.8755093,13.361534,18.849373,24.33721,29.825047,35.312885,31.599937,27.88699,24.174044,20.462908,16.749962,16.4617,16.175253,15.8869915,15.600543,15.312282,14.674119,14.037769,13.399607,12.763257,12.125093,10.462607,8.80012,7.137634,5.475147,3.8126602,4.499773,5.186886,5.8758116,6.5629244,7.250037,8.174648,9.099259,10.025683,10.950294,11.874905,11.213174,10.549629,9.8878975,9.224354,8.562622,8.675026,8.78743,8.899834,9.012237,9.12464,7.512917,5.89938,4.2876563,2.6741197,1.062396,1.0243238,0.9880646,0.9499924,0.9119202,0.87566096,2.2245052,3.5751622,4.9258194,6.2746634,7.6253204,7.5256076,7.4258947,7.324369,7.224656,7.124943,6.8004227,6.4759026,6.149569,5.825049,5.5005283,7.6742706,9.849826,12.025381,14.200936,16.374678,14.587097,12.799516,11.011934,9.224354,7.4367723,6.736969,6.037165,5.337362,4.6375585,3.9377546,3.6241121,3.3122826,3.000453,2.6868105,2.374981,4.3873696,6.399758,8.412147,10.424535,12.436923,9.96223,7.4875355,5.0128417,2.5381477,0.06164073,0.25018883,0.43692398,0.62547207,0.8122072,1.0007553,1.2001812,1.3996071,1.6008459,1.8002719,1.9996977,1.8129625,1.6244144,1.4376793,1.2491312,1.062396,1.9743162,2.8880494,3.7999697,4.7118897,5.6256227,5.3246713,5.0255322,4.7245803,4.4254417,4.12449,3.636803,3.149116,2.663242,2.175555,1.6878681,1.3506571,1.0116332,0.6744221,0.33721104,0.0,0.17585737,0.34990177,0.52575916,0.69980353,0.87566096,0.824898,0.774135,0.72518504,0.6744221,0.62547207,2.08672,3.5497808,5.0128417,6.4759026,7.93715,7.949841,7.9625316,7.9752226,7.987913,8.000604,9.4509735,10.899531,12.349901,13.800271,15.250641,12.299138,9.349448,6.399758,3.4500678,0.50037766,1.5627737,2.6251698,3.6875658,4.749962,5.812358,5.5005283,5.186886,4.8750563,4.5632267,4.249584,3.4119956,2.5744069,1.7368182,0.89922947,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.13778515,0.21211663,0.28826106,0.36259252,0.43692398,0.5747091,0.7124943,0.85027945,0.9880646,1.1258497,0.89922947,0.6744221,0.44961473,0.22480737,0.0,1.0497054,2.0994108,3.150929,4.2006345,5.2503395,6.588306,7.9244595,9.262425,10.600392,11.938358,10.225109,8.511859,6.8004227,5.087173,3.3757362,3.0620937,2.7502642,2.4366217,2.124792,1.8129625,1.550083,1.2872034,1.0243238,0.76325727,0.50037766,2.03777,3.5751622,5.1125546,6.6499467,8.187339,7.911769,7.6380115,7.362441,7.0868707,6.813113,6.7134004,6.6118746,6.5121617,6.412449,6.3127356,7.1992745,8.087626,8.974165,9.862516,10.750868,8.624263,6.4994707,4.3746786,2.2498865,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,1.6371052,3.2125697,4.788034,6.3616858,7.93715,6.3616858,4.788034,3.2125697,1.6371052,0.06164073,1.2382535,2.4130533,3.587853,4.762653,5.9374523,4.949388,3.9631362,2.9750717,1.987007,1.0007553,2.8499773,4.699199,6.550234,8.399456,10.25049,10.437225,10.625773,10.812509,10.999244,11.187792,10.774437,10.362894,9.949538,9.537996,9.12464,10.025683,10.924912,11.8241415,12.725184,13.6244135,13.125849,12.625471,12.125093,11.624716,11.124338,8.950596,6.775041,4.599486,2.4257438,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.17585737,0.22480737,0.2755703,0.3245203,0.37528324,0.42423326,0.4749962,0.52575916,0.5747091,0.62547207,0.66173136,0.69980353,0.73787576,0.774135,0.8122072,0.7868258,0.76325727,0.73787576,0.7124943,0.6871128,0.69980353,0.7124943,0.72518504,0.73787576,0.7505665,4.361988,7.9752226,11.588457,15.199879,18.813112,19.163015,19.512917,19.862818,20.212719,20.562622,20.437527,20.312433,20.187338,20.062244,19.93715,18.274662,16.612177,14.94969,13.287203,11.624716,11.711739,11.800573,11.887595,11.974618,12.06164,11.675479,11.287505,10.899531,10.51337,10.125396,10.738177,11.349146,11.961927,12.574709,13.1874895,13.386916,13.588155,13.7875805,13.987006,14.188245,12.549327,10.912222,9.275117,7.6380115,6.000906,7.61263,9.224354,10.837891,12.449615,14.06315,13.588155,13.113158,12.638163,12.163166,11.6881695,9.362139,7.037921,4.7118897,2.3876717,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06164073,0.12509441,0.18673515,0.25018883,0.31182957,0.6000906,0.8883517,1.1747998,1.4630609,1.7495089,2.7375734,3.7256382,4.7118897,5.6999545,6.688019,6.8004227,6.9128265,7.02523,7.137634,7.250037,6.2257137,5.199577,4.175253,3.150929,2.124792,3.0131438,3.245203,3.4772623,3.7093215,3.9431937,4.175253,5.009216,5.844991,6.680767,7.51473,8.350506,10.80707,13.265448,15.722012,18.18039,20.636953,21.217102,21.797249,22.377398,22.957544,23.537693,22.533312,21.527117,20.522736,19.518354,18.512161,16.517902,14.521831,12.527572,10.533313,8.537241,16.67563,24.812206,32.950596,41.08717,49.22556,44.569874,39.915997,35.26031,30.604622,25.950747,21.325878,16.701012,12.07433,7.4494634,2.8245957,3.303218,3.780027,4.256836,4.7354584,5.2122674,4.860553,4.507025,4.15531,3.8017826,3.4500678,4.7118897,5.975525,7.2373466,8.499168,9.762803,9.177217,8.59163,8.007855,7.422269,6.836682,5.6981416,4.557788,3.4174345,2.277081,1.1367276,0.9499924,0.76325727,0.5747091,0.387974,0.19942589,0.38978696,0.58014804,0.7705091,0.96087015,1.1494182,1.0243238,0.89922947,0.774135,0.6508536,0.52575916,0.6852999,0.8448406,1.0043813,1.1657349,1.3252757,1.6153497,1.9054236,2.1954978,2.4855716,2.7756457,2.2516994,1.7295663,1.2074331,0.6852999,0.16316663,1.6733645,3.1817493,4.691947,6.202145,7.7123427,8.406708,9.102885,9.79725,10.491614,11.187792,11.999999,12.812206,13.6244135,14.436621,15.250641,15.870674,16.490707,17.11074,17.730774,18.350807,17.638313,16.92582,16.213324,15.50083,14.788336,14.0323305,13.278138,12.522133,11.7679405,11.011934,10.179785,9.347635,8.515485,7.6833353,6.849373,7.315304,7.7794223,8.245354,8.709473,9.175404,9.77912,10.384649,10.990179,11.595709,12.199425,13.002567,13.80571,14.607039,15.410182,16.213324,16.800724,17.388124,17.975525,18.562923,19.150324,18.53573,17.919323,17.304728,16.690134,16.075539,15.219821,14.365915,13.510198,12.654479,11.800573,10.032935,8.265296,6.497658,4.7300196,2.962381,3.0167696,3.0729716,3.1273603,3.1817493,3.2379513,3.2306993,3.2216346,3.2143826,3.207131,3.199879,3.1273603,3.054842,2.9823234,2.909805,2.8372865,3.101979,3.3666716,3.633177,3.8978696,4.162562,4.795286,5.42801,6.060734,6.6916447,7.324369,12.469557,17.614744,22.759932,27.90512,33.05031,29.814169,26.579844,23.34552,20.10938,16.875055,16.717327,16.5596,16.401873,16.244144,16.08823,15.190813,14.293397,13.394168,12.496751,11.599335,10.020245,8.439341,6.8602505,5.279347,3.7002566,4.4272547,5.1542525,5.883064,6.6100616,7.3370595,7.902704,8.4683485,9.03218,9.597824,10.161655,9.655839,9.14821,8.640579,8.13295,7.6253204,7.9045167,8.185526,8.464723,8.745731,9.024928,7.520169,6.01541,4.510651,3.004079,1.49932,1.4666867,1.4358664,1.403233,1.3705997,1.3379664,2.3894846,3.442816,4.494334,5.5476656,6.599184,6.695271,6.789545,6.885632,6.979906,7.07418,7.0071006,6.9400206,6.872941,6.8058615,6.736969,8.709473,10.681975,12.654479,14.626982,16.599485,14.755702,12.910107,11.06451,9.220728,7.3751316,6.7097745,6.0444174,5.3808727,4.7155156,4.0501585,3.7256382,3.3993049,3.0747845,2.7502642,2.4257438,4.1825047,5.9392653,7.6978393,9.4546,11.213174,9.017676,6.8221784,4.6266804,2.4329958,0.2374981,0.36259252,0.48768693,0.61278135,0.73787576,0.8629702,1.0116332,1.162109,1.3125849,1.4630609,1.6117238,1.5319533,1.452183,1.3724127,1.2926424,1.2128719,1.8727903,2.5327086,3.1926272,3.8525455,4.512464,4.612177,4.7118897,4.8116026,4.9131284,5.0128417,4.2822175,3.5534067,2.8227828,2.0921588,1.3633479,1.2998942,1.2382535,1.1747998,1.1131591,1.0497054,1.3434052,1.6352923,1.9271792,2.220879,2.5127661,2.1121013,1.7132497,1.3125849,0.9119202,0.51306844,1.6824293,2.8517902,4.022964,5.1923246,6.3616858,6.882006,7.402326,7.9226465,8.442966,8.963287,10.429974,11.896661,13.36516,14.831847,16.300346,15.431937,14.565341,13.696932,12.830337,11.961927,10.924912,9.8878975,8.8508835,7.8120556,6.775041,6.2746634,5.774286,5.275721,4.7753434,4.274966,3.5932918,2.909805,2.228131,1.5446441,0.8629702,0.9354887,1.0080072,1.0805258,1.1530442,1.2255627,0.9898776,0.7541924,0.52032024,0.28463513,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.11240368,0.17585737,0.2374981,0.2991388,0.36259252,0.47318324,0.581961,0.69255173,0.8031424,0.9119202,0.7324369,0.5529536,0.37165734,0.19217403,0.012690738,1.1403534,2.268016,3.395679,4.5233417,5.6491914,6.7134004,7.7757964,8.838193,9.900589,10.962985,9.860703,8.758422,7.654328,6.552047,5.4497657,5.045475,4.6393714,4.2350807,3.83079,3.4246864,3.0620937,2.6995013,2.3369088,1.9743162,1.6117238,3.2198215,4.8279195,6.434204,8.042302,9.6504,9.004985,8.3595705,7.7141557,7.0705543,6.4251394,6.446895,6.4704633,6.492219,6.5157876,6.5375433,7.3370595,8.136576,8.937905,9.737422,10.536939,8.662335,6.787732,4.9131284,3.0367124,1.162109,0.94274056,0.72337204,0.50219065,0.28282216,0.06164073,1.8057107,3.5479677,5.290225,7.0324817,8.774739,7.2899227,5.805106,4.3202896,2.8354735,1.3506571,2.2933977,3.2343252,4.177066,5.1198063,6.0625467,5.0146546,3.966762,2.9206827,1.8727903,0.824898,2.5417736,4.2604623,5.977338,7.6942134,9.412902,9.402024,9.39296,9.382081,9.373016,9.362139,9.48542,9.606889,9.73017,9.851639,9.97492,10.420909,10.865085,11.30926,11.755249,12.199425,11.896661,11.595709,11.292944,10.990179,10.687414,8.649645,6.6118746,4.574105,2.5381477,0.50037766,0.40066472,0.2991388,0.19942589,0.099712946,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.034446288,0.058014803,0.07977036,0.10333887,0.12509441,0.16679256,0.21030366,0.2520018,0.2955129,0.33721104,0.37528324,0.41335547,0.44961473,0.48768693,0.52575916,0.55476654,0.5855869,0.61459434,0.64541465,0.6744221,0.68167394,0.69073874,0.6979906,0.70524246,0.7124943,0.7433147,0.77232206,0.8031424,0.8321498,0.8629702,4.307599,7.752228,11.1968565,14.641486,18.087927,18.278288,18.466837,18.657198,18.847559,19.03792,19.244598,19.453089,19.659767,19.868258,20.074934,18.684393,17.295664,15.905121,14.514579,13.125849,13.240066,13.354282,13.470312,13.584529,13.700559,13.029762,12.360779,11.689982,11.019187,10.3502035,10.801631,11.254871,11.708113,12.15954,12.612781,12.743314,12.872034,13.002567,13.1331005,13.261822,11.925668,10.587702,9.249735,7.911769,6.5756154,8.317872,10.060129,11.802386,13.544643,15.2869005,14.364102,13.443117,12.52032,11.597522,10.674724,8.549932,6.4251394,4.3003473,2.175555,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.027194439,0.054388877,0.08339628,0.11059072,0.13778515,0.48043507,0.823085,1.1657349,1.5083848,1.8492218,1.789394,1.7295663,1.6697385,1.6099107,1.550083,2.5399606,3.529838,4.519716,5.5095935,6.4994707,6.588306,6.6753283,6.7623506,6.849373,6.9382076,5.922949,4.9076896,3.8924308,2.8771715,1.8619126,3.0258346,3.2143826,3.4047437,3.5951047,3.785466,3.975827,4.7572136,5.540414,6.3218007,7.1050005,7.8882003,10.865085,13.8419695,16.820667,19.797552,22.774435,22.785315,22.794378,22.805256,22.814322,22.8252,22.014805,21.20441,20.395828,19.585434,18.77504,17.059978,15.344915,13.629852,11.91479,10.199727,18.624565,27.049402,35.47605,43.90089,52.325726,46.390087,40.45445,34.520622,28.584982,22.649342,18.688019,14.724882,10.761745,6.8004227,2.8372865,3.3304121,3.8217251,4.314851,4.8079767,5.2992897,5.282973,5.2648435,5.2467136,5.230397,5.2122674,6.200332,7.1865835,8.174648,9.162713,10.150778,9.867955,9.585134,9.302311,9.019489,8.736667,7.170267,5.6020546,4.0356545,2.467442,0.89922947,0.7995165,0.69980353,0.6000906,0.50037766,0.40066472,0.49312583,0.5855869,0.678048,0.7705091,0.8629702,0.89922947,0.93730164,0.97537386,1.0116332,1.0497054,1.1693609,1.2908293,1.4104849,1.5301404,1.649796,1.8673514,2.084907,2.3024626,2.520018,2.7375734,2.2426348,1.7476959,1.2527572,0.75781834,0.26287958,1.4576219,2.6523643,3.8471067,5.041849,6.2365913,6.9146395,7.592687,8.270736,8.94697,9.625018,10.56232,11.499621,12.436923,13.374225,14.313339,14.752076,15.192626,15.633177,16.071913,16.512463,15.799969,15.087475,14.37498,13.662486,12.949992,12.415168,11.880343,11.34552,10.810696,10.275872,9.572442,8.870826,8.167397,7.46578,6.7623506,7.179332,7.5981264,8.015107,8.432089,8.8508835,9.409276,9.969481,10.529687,11.089892,11.650098,12.368031,13.084151,13.802084,14.520018,15.23795,15.738328,16.236893,16.73727,17.237648,17.738026,17.295664,16.8533,16.409124,15.966762,15.524399,14.964193,14.405801,13.845595,13.28539,12.725184,10.9774885,9.229793,7.4820967,5.7344007,3.9867048,3.923251,3.8579843,3.7927177,3.727451,3.6621845,3.584227,3.5080826,3.4301252,3.3521678,3.2742105,3.2053177,3.1346123,3.0657198,2.9950142,2.9243085,3.2180085,3.5098956,3.8017826,4.0954823,4.3873696,4.8641787,5.3428006,5.81961,6.298232,6.775041,11.5775795,16.380117,21.182655,25.985193,30.787731,28.030214,25.272697,22.515182,19.757666,17.00015,16.972956,16.94576,16.916754,16.889559,16.862366,15.705695,14.547212,13.390542,12.232059,11.075388,9.577881,8.080374,6.582867,5.08536,3.587853,4.3547363,5.121619,5.8903155,6.6571984,7.4258947,7.6307597,7.835624,8.040489,8.245354,8.450218,8.096691,7.744976,7.3932614,7.039734,6.688019,7.135821,7.5818095,8.029612,8.477413,8.925215,7.5274205,6.1296263,4.7318325,3.3358512,1.938057,1.9108626,1.8818551,1.8546607,1.8274662,1.8002719,2.5544643,3.3104696,4.064662,4.8206677,5.57486,5.864934,6.155008,6.445082,6.735156,7.02523,7.215591,7.404139,7.5945,7.7848616,7.9752226,9.744674,11.514126,13.28539,15.054841,16.824293,14.922495,13.020698,11.117086,9.215289,7.311678,6.68258,6.051669,5.422571,4.7916603,4.162562,3.825351,3.48814,3.149116,2.811905,2.474694,3.97764,5.480586,6.981719,8.484665,9.987611,8.073122,6.156821,4.2423325,2.327844,0.41335547,0.4749962,0.53663695,0.6000906,0.66173136,0.72518504,0.824898,0.9246109,1.0243238,1.1258497,1.2255627,1.2527572,1.2799516,1.3071461,1.3343405,1.3633479,1.7694515,2.1773682,2.5852847,2.9932013,3.3993049,3.8996825,4.40006,4.900438,5.4008155,5.89938,4.9276323,3.9558845,2.9823234,2.0105755,1.0370146,1.2491312,1.4630609,1.6751775,1.887294,2.0994108,2.5091403,2.9206827,3.3304121,3.7401419,4.1498713,3.3993049,2.6505513,1.8999848,1.1494182,0.40066472,1.2781386,2.1556125,3.0330863,3.9105604,4.788034,5.814171,6.8421206,7.8700705,8.898021,9.924157,11.410787,12.895603,14.380419,15.865235,17.350052,18.564737,19.77942,20.99592,22.210604,23.42529,20.287052,17.150625,14.012388,10.874149,7.7377243,7.0506115,6.3616858,5.674573,4.98746,4.3003473,3.7727752,3.245203,2.7176309,2.1900587,1.6624867,1.8202144,1.9779422,2.13567,2.2933977,2.4493124,1.9670644,1.4848163,1.0025684,0.52032024,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.0870222,0.13778515,0.18673515,0.2374981,0.28826106,0.36984438,0.45324063,0.53482395,0.61822027,0.69980353,0.5656443,0.42967212,0.2955129,0.15954071,0.025381476,1.2291887,2.4348087,3.6404288,4.844236,6.049856,6.836682,7.6253204,8.412147,9.200785,9.987611,9.494485,9.003172,8.510046,8.01692,7.5256076,7.027043,6.530291,6.0317264,5.5349746,5.038223,4.574105,4.1117992,3.6494937,3.1871881,2.7248828,4.401873,6.0806766,7.757667,9.434657,11.111648,10.098202,9.082943,8.067683,7.0524244,6.037165,6.1822023,6.3272395,6.472276,6.6173134,6.7623506,7.474845,8.187339,8.899834,9.612328,10.324821,8.700407,7.07418,5.4497657,3.825351,2.1991236,1.7730774,1.3452182,0.91735905,0.4894999,0.06164073,1.9725033,3.881553,5.7924156,7.703278,9.612328,8.21816,6.8221784,5.42801,4.0320287,2.6378605,3.346729,4.0574102,4.7680917,5.47696,6.187641,5.0799212,3.972201,2.864481,1.7567607,0.6508536,2.2353828,3.8199122,5.4044414,6.9907837,8.575313,8.366822,8.160145,7.951654,7.744976,7.5382986,8.194591,8.852696,9.510801,10.167094,10.825199,10.8143215,10.805257,10.794379,10.785315,10.774437,10.669285,10.564133,10.460794,10.355642,10.25049,8.350506,6.450521,4.550536,2.6505513,0.7505665,0.6000906,0.44961473,0.2991388,0.15047589,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.045324065,0.065266654,0.08520924,0.10515183,0.12509441,0.15954071,0.19579996,0.23024625,0.26469254,0.2991388,0.3245203,0.34990177,0.37528324,0.40066472,0.42423326,0.44780177,0.46955732,0.49312583,0.5148814,0.53663695,0.57833505,0.61822027,0.65810543,0.6979906,0.73787576,0.7850128,0.8321498,0.8792868,0.92823684,0.97537386,4.25321,7.5292335,10.80707,14.084907,17.362743,17.39175,17.422571,17.45339,17.482399,17.513218,18.051668,18.59193,19.132195,19.672457,20.212719,19.094122,17.977337,16.860552,15.741954,14.625169,14.7683935,14.909804,15.053028,15.194439,15.337664,14.385859,13.43224,12.480434,11.526816,10.57501,10.866898,11.160598,11.452485,11.744371,12.038072,12.097899,12.157727,12.217555,12.277383,12.337211,11.300196,10.263181,9.224354,8.187339,7.1503243,9.023115,10.894093,12.766883,14.639673,16.512463,15.141864,13.773077,12.402477,11.0318775,9.663091,7.7377243,5.812358,3.8869917,1.9634385,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.054388877,0.11059072,0.16497959,0.21936847,0.2755703,0.8974165,1.5192627,2.1429217,2.764768,3.386614,2.9805105,2.572594,2.1646774,1.7567607,1.3506571,2.3423476,3.3358512,4.327542,5.319232,6.3127356,6.3743763,6.43783,6.4994707,6.5629244,6.624565,5.620184,4.61399,3.6096084,2.6052272,1.6008459,3.0367124,3.1853752,3.3322253,3.4808881,3.6277382,3.774588,4.505212,5.235836,5.964647,6.695271,7.4258947,10.9230995,14.420304,17.91751,21.414715,24.911919,24.351713,23.793322,23.233116,22.67291,22.112705,21.49811,20.881702,20.267109,19.652514,19.03792,17.602055,16.168001,14.732134,13.29808,11.862214,20.575312,29.286598,37.999695,46.712795,55.42408,48.2103,40.99471,33.779118,26.56534,19.34975,16.050158,12.750566,9.449161,6.149569,2.8499773,3.3576066,3.8652363,4.3728657,4.880495,5.388125,5.7053933,6.0226617,6.33993,6.6571984,6.9744673,7.686961,8.399456,9.11195,9.824444,10.536939,10.556881,10.576823,10.596766,10.616709,10.636651,8.642392,6.6481338,4.652062,2.657803,0.66173136,0.6508536,0.63816285,0.62547207,0.61278135,0.6000906,0.5946517,0.58921283,0.5855869,0.58014804,0.5747091,0.774135,0.97537386,1.1747998,1.3742256,1.5754645,1.6552348,1.7350051,1.8147756,1.8945459,1.9743162,2.1193533,2.2643902,2.4094272,2.5544643,2.6995013,2.231757,1.7658255,1.2980812,0.83033687,0.36259252,1.2418793,2.1229792,3.002266,3.8833659,4.762653,5.422571,6.0824895,6.742408,7.402326,8.062244,9.12464,10.1870365,11.249433,12.311829,13.374225,13.635292,13.894546,14.155612,14.4148655,14.674119,13.961625,13.24913,12.536636,11.8241415,11.111648,10.798005,10.48255,10.167094,9.851639,9.537996,8.9651,8.392203,7.819308,7.2482243,6.6753283,7.0451727,7.415017,7.7848616,8.154706,8.52455,9.039432,9.554313,10.069194,10.585889,11.10077,11.731681,12.364405,12.9971285,13.629852,14.262577,14.674119,15.087475,15.50083,15.912373,16.325727,16.055597,15.785465,15.515334,15.245202,14.975071,14.710379,14.445685,14.17918,13.914488,13.649796,11.922042,10.194288,8.466536,6.740595,5.0128417,4.8279195,4.6429973,4.458075,4.273153,4.0882306,3.9395678,3.7927177,3.6458678,3.4972048,3.350355,3.2832751,3.2143826,3.147303,3.0802233,3.0131438,3.3322253,3.6531196,3.972201,4.2930956,4.612177,4.934884,5.2575917,5.580299,5.903006,6.2257137,10.685601,15.14549,19.605377,24.065266,28.525154,26.244446,23.965553,21.684845,19.404139,17.125244,17.22677,17.330109,17.431635,17.534973,17.638313,16.220575,14.802839,13.385102,11.967366,10.549629,9.135518,7.7195945,6.305484,4.88956,3.4754493,4.2822175,5.090799,5.8975673,6.7043357,7.512917,7.3570023,7.2029004,7.0469856,6.892884,6.736969,6.539356,6.341743,6.14413,5.9483304,5.750717,6.3653116,6.979906,7.5945,8.210908,8.825501,7.5346723,6.245656,4.954827,3.6658103,2.374981,2.3532255,2.3296568,2.3079014,2.2843328,2.2625773,2.7194438,3.1781235,3.63499,4.0918565,4.550536,5.034597,5.520471,6.004532,6.490406,6.9744673,7.422269,7.8700705,8.317872,8.765674,9.211663,10.779876,12.348088,13.914488,15.4827,17.0491,15.089288,13.129475,11.169662,9.20985,7.250037,6.6553855,6.060734,5.464269,4.8696175,4.274966,3.925064,3.5751622,3.2252605,2.8753586,2.525457,3.7727752,5.0200934,6.2674117,7.51473,8.762048,7.1267557,5.4932766,3.8579843,2.222692,0.5873999,0.5873999,0.5873999,0.5873999,0.5873999,0.5873999,0.63816285,0.6871128,0.73787576,0.7868258,0.8375887,0.97174793,1.1077201,1.2418793,1.3778516,1.5120108,1.6679256,1.8220274,1.9779422,2.132044,2.2879589,3.1871881,4.0882306,4.98746,5.8866897,6.787732,5.573047,4.358362,3.141864,1.9271792,0.7124943,1.2001812,1.6878681,2.175555,2.663242,3.149116,3.6766882,4.2042603,4.7318325,5.2594047,5.7869763,4.688321,3.587853,2.4873846,1.3869164,0.28826106,0.872035,1.4576219,2.0432088,2.6269827,3.2125697,4.748149,6.281915,7.817495,9.353074,10.88684,12.389787,13.892733,15.3956785,16.89681,18.399757,21.697536,24.995316,28.293095,31.590874,34.88684,29.64919,24.413355,19.175705,13.938056,8.700407,7.8247466,6.9508986,6.0752378,5.199577,4.325729,3.9522583,3.5806012,3.207131,2.8354735,2.4620032,2.70494,2.9478772,3.1908143,3.4319382,3.6748753,2.9442513,2.2154403,1.4848163,0.7541924,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.06164073,0.099712946,0.13778515,0.17585737,0.21211663,0.26831847,0.32270733,0.3770962,0.43329805,0.48768693,0.39703882,0.30820364,0.21755551,0.12690738,0.038072214,1.3198367,2.6016014,3.8851788,5.1669436,6.450521,6.9617763,7.474845,7.987913,8.499168,9.012237,9.130079,9.247922,9.365765,9.481794,9.599637,9.010424,8.419398,7.8301854,7.2391596,6.6499467,6.0879283,5.52591,4.9620786,4.40006,3.8380418,5.5857377,7.3316207,9.079316,10.827013,12.574709,11.189605,9.804502,8.419398,7.0342946,5.6491914,5.91751,6.185828,6.452334,6.720652,6.987158,7.61263,8.238102,8.861761,9.487233,10.112705,8.736667,7.362441,5.9882154,4.612177,3.2379513,2.6016014,1.9670644,1.3325275,0.6979906,0.06164073,2.1392958,4.216951,6.294606,8.372261,10.449916,9.144584,7.83925,6.53573,5.230397,3.925064,4.401873,4.880495,5.3573046,5.8341136,6.3127356,5.145188,3.97764,2.810092,1.6425442,0.4749962,1.9271792,3.3793623,4.8333583,6.285541,7.7377243,7.3316207,6.92733,6.5230393,6.1169357,5.712645,6.9055743,8.096691,9.28962,10.48255,11.675479,11.209548,10.745429,10.279498,9.815379,9.349448,9.441909,9.53437,9.626831,9.719293,9.811753,8.049554,6.2873545,4.5251546,2.762955,1.0007553,0.7995165,0.6000906,0.40066472,0.19942589,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.054388877,0.072518505,0.09064813,0.10696479,0.12509441,0.15228885,0.1794833,0.20667773,0.23568514,0.26287958,0.2755703,0.28826106,0.2991388,0.31182957,0.3245203,0.34083697,0.35534066,0.36984438,0.38434806,0.40066472,0.47318324,0.54570174,0.61822027,0.69073874,0.76325727,0.82671094,0.8919776,0.9572442,1.0225109,1.0877775,4.1970086,7.308052,10.417283,13.526514,16.637558,16.507025,16.378304,16.24777,16.117237,15.986704,16.860552,17.732588,18.604622,19.476658,20.350506,19.505665,18.660824,17.81417,16.96933,16.124489,16.294909,16.465326,16.635744,16.80435,16.97477,15.740141,14.505513,13.2690735,12.034446,10.799818,10.932164,11.06451,11.1968565,11.329204,11.463363,11.452485,11.4416065,11.432542,11.421664,11.4126,10.674724,9.936848,9.200785,8.46291,7.7250338,9.728357,11.729868,13.7331915,15.734702,17.738026,15.919624,14.103036,12.284635,10.468046,8.649645,6.925517,5.199577,3.4754493,1.7495089,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08339628,0.16497959,0.24837588,0.32995918,0.41335547,1.3143979,2.2172532,3.1201086,4.022964,4.9258194,4.169814,3.4156215,2.659616,1.9054236,1.1494182,2.1447346,3.1400511,4.135368,5.130684,6.1241875,6.16226,6.200332,6.2384043,6.2746634,6.3127356,5.317419,4.322103,3.3267863,2.333283,1.3379664,3.049403,3.1545548,3.2597067,3.3648586,3.4700103,3.5751622,4.25321,4.9294453,5.6074934,6.285541,6.9617763,10.979301,14.996826,19.01435,23.031878,27.049402,25.919926,24.790451,23.659163,22.529686,21.40021,20.979603,20.560808,20.140202,19.719595,19.3008,18.144129,16.989273,15.834415,14.679558,13.524701,22.524246,31.525606,40.525154,49.5247,58.524246,50.030514,41.534973,33.03943,24.5457,16.050158,13.412297,10.774437,8.136576,5.5005283,2.8626678,3.3848011,3.9069343,4.4308805,4.953014,5.475147,6.1278133,6.78048,7.4331465,8.0858135,8.736667,9.175404,9.612328,10.049252,10.487988,10.924912,11.24762,11.570327,11.893035,12.215742,12.536636,10.114518,7.6924005,5.2702823,2.8481643,0.42423326,0.50037766,0.5747091,0.6508536,0.72518504,0.7995165,0.6979906,0.5946517,0.49312583,0.38978696,0.28826106,0.6508536,1.0116332,1.3742256,1.7368182,2.0994108,2.1392958,2.179181,2.220879,2.2607644,2.3006494,2.373168,2.4456866,2.518205,2.5907235,2.663242,2.222692,1.7821422,1.3415923,0.90285534,0.46230546,1.0279498,1.5917811,2.1574254,2.72307,3.2869012,3.930503,4.572292,5.2158933,5.857682,6.4994707,7.686961,8.874452,10.061942,11.249433,12.436923,12.516694,12.598277,12.678047,12.757817,12.837588,12.125093,11.4126,10.700105,9.987611,9.275117,9.180842,9.084756,8.990481,8.894395,8.80012,8.357758,7.915395,7.473032,7.0306687,6.588306,6.9092,7.231908,7.554615,7.877322,8.200029,8.669587,9.139144,9.610515,10.080072,10.549629,11.097144,11.644659,12.192173,12.739688,13.287203,13.611723,13.938056,14.262577,14.587097,14.911617,14.81553,14.71763,14.61973,14.521831,14.425743,14.454751,14.485571,14.514579,14.545399,14.574407,12.868408,11.160598,9.452786,7.744976,6.037165,5.732588,5.42801,5.121619,4.8170414,4.512464,4.2949085,4.077353,3.8597972,3.6422417,3.4246864,3.3594196,3.294153,3.2306993,3.1654327,3.100166,3.4482548,3.7945306,4.1426196,4.4907084,4.836984,5.0055895,5.1723824,5.3391747,5.5077806,5.674573,9.791811,13.909049,18.0281,22.145338,26.262575,24.460491,22.658407,20.85451,19.052423,17.25034,17.482399,17.714457,17.94833,18.18039,18.412449,16.735458,15.056654,13.379663,11.702674,10.025683,8.693155,7.360628,6.0281005,4.695573,3.3630457,4.209699,5.0581656,5.904819,6.7532854,7.5999393,7.0850577,6.5701766,6.055295,5.540414,5.0255322,4.9820213,4.940323,4.896812,4.855114,4.8116026,5.5948024,6.378002,7.159389,7.9425893,8.725789,7.5419245,6.359873,5.177821,3.9957695,2.811905,2.7955883,2.7774587,2.759329,2.7430124,2.7248828,2.8844235,3.045777,3.2053177,3.3648586,3.5243993,4.2042603,4.8841214,5.565795,6.245656,6.925517,7.6307597,8.334189,9.039432,9.744674,10.449916,11.815077,13.180238,14.545399,15.91056,17.27572,15.257894,13.240066,11.222239,9.2044115,7.1883965,6.628191,6.0679855,5.5077806,4.947575,4.3873696,4.024777,3.6621845,3.299592,2.9369993,2.5744069,3.5679104,4.559601,5.5531044,6.544795,7.5382986,6.1822023,4.8279195,3.4718235,2.1175404,0.76325727,0.69980353,0.63816285,0.5747091,0.51306844,0.44961473,0.44961473,0.44961473,0.44961473,0.44961473,0.44961473,0.69255173,0.9354887,1.1766127,1.4195497,1.6624867,1.5645868,1.4666867,1.3705997,1.2726997,1.1747998,2.474694,3.774588,5.0744824,6.3743763,7.6742706,6.2166486,4.76084,3.303218,1.845596,0.387974,1.1494182,1.9126755,2.675933,3.437377,4.2006345,4.844236,5.4896507,6.1350656,6.78048,7.4258947,5.975525,4.5251546,3.0747845,1.6244144,0.17585737,0.46774435,0.75963134,1.0533313,1.3452182,1.6371052,3.680314,5.7217097,7.764919,9.808127,11.849524,13.370599,14.889862,16.410936,17.9302,19.449463,24.830336,30.209396,35.590267,40.96933,46.3502,39.01133,31.676083,24.33721,17.00015,9.663091,8.600695,7.5382986,6.474089,5.411693,4.349297,4.1317415,3.9141862,3.6966307,3.4808881,3.2633326,3.589666,3.917812,4.2441454,4.572292,4.900438,3.923251,2.9442513,1.9670644,0.9898776,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.038072214,0.06164073,0.0870222,0.11240368,0.13778515,0.16497959,0.19217403,0.21936847,0.24837588,0.2755703,0.23024625,0.18492219,0.13959812,0.09427405,0.05076295,1.4104849,2.770207,4.1299286,5.4896507,6.849373,7.0868707,7.324369,7.5618668,7.799365,8.036863,8.765674,9.492672,10.21967,10.946668,11.675479,10.991992,10.310318,9.626831,8.945157,8.26167,7.5999393,6.9382076,6.2746634,5.612932,4.949388,6.7677894,8.584378,10.40278,12.219368,14.037769,12.282822,10.527874,8.772926,7.017978,5.2630305,5.6528172,6.0426044,6.432391,6.8221784,7.211965,7.750415,8.287052,8.825501,9.362139,9.900589,8.774739,7.650702,6.5248523,5.4008155,4.274966,3.4319382,2.5907235,1.7476959,0.90466833,0.06164073,2.3079014,4.552349,6.796797,9.043057,11.287505,10.07282,8.858135,7.6416373,6.4269524,5.2122674,5.4570174,5.7017674,5.9483304,6.19308,6.43783,5.2104545,3.9830787,2.7557032,1.5283275,0.2991388,1.6207886,2.9406252,4.2604623,5.580299,6.9001355,6.298232,5.6945157,5.092612,4.4907084,3.8869917,5.614745,7.3424983,9.070251,10.798005,12.525759,11.6047735,10.685601,9.764616,8.845445,7.9244595,8.214534,8.504607,8.794682,9.084756,9.374829,7.750415,6.1241875,4.499773,2.8753586,1.2491312,1.0007553,0.7505665,0.50037766,0.25018883,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.065266654,0.07977036,0.09427405,0.11059072,0.12509441,0.14503701,0.16497959,0.18492219,0.20486477,0.22480737,0.22480737,0.22480737,0.22480737,0.22480737,0.22480737,0.23205921,0.23931105,0.24837588,0.25562772,0.26287958,0.3680314,0.47318324,0.57833505,0.68167394,0.7868258,0.87022203,0.95180535,1.0352017,1.1167849,1.2001812,4.1426196,7.0850577,10.027496,12.969934,15.912373,15.622298,15.332225,15.0421505,14.752076,14.462003,15.667623,16.873243,18.07705,19.282671,20.48829,19.915394,19.342497,18.769602,18.196705,17.625622,17.823235,18.020847,18.216648,18.41426,18.611874,17.094423,15.576975,14.059525,12.542075,11.024626,10.997431,10.970237,10.943042,10.915848,10.88684,10.80707,10.7273,10.64753,10.567759,10.487988,10.049252,9.612328,9.175404,8.736667,8.299743,10.431787,12.565643,14.697688,16.829731,18.961775,16.697386,14.432995,12.166792,9.902402,7.6380115,6.111497,4.5867953,3.0620937,1.5373923,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.11059072,0.21936847,0.32995918,0.4405499,0.5493277,1.7331922,2.9152439,4.0972953,5.279347,6.4632115,5.3591175,4.256836,3.1545548,2.0522738,0.9499924,1.9471219,2.9442513,3.9431937,4.940323,5.9374523,5.9501433,5.962834,5.975525,5.9882154,5.999093,5.0146546,4.0302157,3.045777,2.0595255,1.0750868,3.0620937,3.1255474,3.1871881,3.2506418,3.3122826,3.3757362,3.9993954,4.6248674,5.2503395,5.8758116,6.4994707,11.037316,15.575162,20.113007,24.650852,29.186884,27.488138,25.78758,24.08702,22.388275,20.687716,20.462908,20.238102,20.013294,19.786674,19.561867,18.688019,17.812357,16.936697,16.062849,15.187187,24.474995,33.762802,43.05061,52.338417,61.624413,51.85073,42.075237,32.29974,22.524246,12.750566,10.774437,8.80012,6.825804,4.8496747,2.8753586,3.4119956,3.9504454,4.4870825,5.0255322,5.562169,6.550234,7.5382986,8.52455,9.512614,10.500679,10.662033,10.825199,10.988366,11.14972,11.312886,11.938358,12.562017,13.1874895,13.812962,14.436621,11.586644,8.73848,5.8866897,3.0367124,0.18673515,0.34990177,0.51306844,0.6744221,0.8375887,1.0007553,0.7995165,0.6000906,0.40066472,0.19942589,0.0,0.52575916,1.0497054,1.5754645,2.0994108,2.6251698,2.6251698,2.6251698,2.6251698,2.6251698,2.6251698,2.6251698,2.6251698,2.6251698,2.6251698,2.6251698,2.2118144,1.8002719,1.3869164,0.97537386,0.5620184,0.8122072,1.062396,1.3125849,1.5627737,1.8129625,2.4366217,3.0620937,3.6875658,4.313038,4.936697,6.249282,7.5618668,8.874452,10.1870365,11.499621,11.399909,11.300196,11.200482,11.10077,10.999244,10.28675,9.574255,8.861761,8.149267,7.4367723,7.5618668,7.686961,7.8120556,7.93715,8.062244,7.750415,7.4367723,7.124943,6.813113,6.4994707,6.775041,7.0506115,7.324369,7.5999393,7.8755093,8.299743,8.725789,9.1500225,9.574255,10.000301,10.462607,10.924912,11.3872175,11.849524,12.311829,12.549327,12.786825,13.024323,13.261822,13.499319,13.575464,13.649796,13.724127,13.800271,13.874602,14.199123,14.525456,14.849977,15.174497,15.50083,13.812962,12.125093,10.437225,8.749357,7.063302,6.637256,6.2130227,5.7869763,5.3627434,4.936697,4.650249,4.361988,4.07554,3.787279,3.5008307,3.437377,3.3757362,3.3122826,3.2506418,3.1871881,3.5624714,3.9377546,4.313038,4.688321,5.0617914,5.0744824,5.087173,5.0998635,5.1125546,5.125245,8.899834,12.674421,16.450823,20.22541,23.999998,22.674723,21.349447,20.024172,18.700708,17.375433,17.738026,18.100618,18.463211,18.825804,19.188396,17.25034,15.312282,13.374225,11.437981,9.499924,8.2507925,6.9998484,5.750717,4.499773,3.2506418,4.137181,5.0255322,5.9120708,6.8004227,7.686961,6.813113,5.9374523,5.0617914,4.1879435,3.3122826,3.4246864,3.53709,3.6494937,3.7618973,3.874301,4.8242936,5.774286,6.7242785,7.6742706,8.624263,7.549176,6.4759026,5.4008155,4.325729,3.2506418,3.2379513,3.2252605,3.2125697,3.199879,3.1871881,3.049403,2.911618,2.7756457,2.6378605,2.5000753,3.3757362,4.249584,5.125245,6.000906,6.874754,7.837437,8.80012,9.762803,10.725487,11.6881695,12.850279,14.012388,15.174497,16.338419,17.500528,15.4246855,13.3506565,11.274815,9.200785,7.124943,6.599184,6.0752378,5.5494785,5.0255322,4.499773,4.12449,3.7492065,3.3757362,3.000453,2.6251698,3.3630457,4.099108,4.836984,5.57486,6.3127356,5.237649,4.162562,3.0874753,2.0123885,0.93730164,0.8122072,0.6871128,0.5620184,0.43692398,0.31182957,0.26287958,0.21211663,0.16316663,0.11240368,0.06164073,0.41335547,0.76325727,1.1131591,1.4630609,1.8129625,1.4630609,1.1131591,0.76325727,0.41335547,0.06164073,1.7621996,3.4627585,5.163317,6.8620634,8.562622,6.8620634,5.163317,3.4627585,1.7621996,0.06164073,1.1004683,2.137483,3.1744974,4.213325,5.2503395,6.011784,6.775041,7.5382986,8.299743,9.063,7.262728,5.462456,3.6621845,1.8619126,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,2.612479,5.163317,7.7123427,10.263181,12.812206,14.349599,15.8869915,17.424383,18.961775,20.499168,27.963135,35.42529,42.887444,50.349598,57.811752,48.375282,38.936996,29.500526,20.062244,10.625773,9.374829,8.125698,6.874754,5.6256227,4.3746786,4.313038,4.249584,4.1879435,4.12449,4.062849,4.4743915,4.8877473,5.2992897,5.712645,6.1241875,4.900438,3.6748753,2.4493124,1.2255627,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,1.49932,2.9369993,4.3746786,5.812358,7.250037,7.211965,7.175706,7.137634,7.0995617,7.063302,8.399456,9.737422,11.075388,12.413355,13.749508,12.975373,12.199425,11.42529,10.649343,9.875207,9.11195,8.350506,7.5872483,6.825804,6.0625467,7.949841,9.837135,11.724429,13.611723,15.50083,13.374225,11.249433,9.12464,6.9998484,4.8750563,5.388125,5.89938,6.412449,6.925517,7.4367723,7.8882003,8.337815,8.78743,9.237044,9.686659,8.812811,7.93715,7.063302,6.187641,5.3119802,4.262275,3.2125697,2.1628644,1.1131591,0.06164073,2.474694,4.8877473,7.3008003,9.712041,12.125093,10.999244,9.875207,8.749357,7.6253204,6.4994707,6.5121617,6.5248523,6.5375433,6.550234,6.5629244,5.275721,3.9867048,2.6995013,1.4122978,0.12509441,1.3125849,2.5000753,3.6875658,4.8750563,6.0625467,5.2630305,4.461701,3.6621845,2.8626678,2.0631514,4.325729,6.588306,8.8508835,11.111648,13.374225,11.999999,10.625773,9.249735,7.8755093,6.4994707,6.987158,7.474845,7.9625316,8.450218,8.937905,7.4494634,5.962834,4.4743915,2.9877625,1.49932,1.2001812,0.89922947,0.6000906,0.2991388,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.13778515,0.15047589,0.16316663,0.17585737,0.18673515,0.17585737,0.16316663,0.15047589,0.13778515,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.26287958,0.40066472,0.53663695,0.6744221,0.8122072,0.9119202,1.0116332,1.1131591,1.2128719,1.3125849,4.0882306,6.8620634,9.637709,12.411542,15.187187,14.737573,14.287958,13.838344,13.386916,12.937301,14.474693,16.012085,17.549479,19.08687,20.624262,20.325123,20.024172,19.725033,19.425894,19.124943,19.34975,19.574556,19.799364,20.024172,20.250792,18.45052,16.650248,14.849977,13.049705,11.249433,11.062697,10.874149,10.687414,10.500679,10.312131,10.161655,10.012992,9.862516,9.712041,9.563377,9.425592,9.287807,9.1500225,9.012237,8.874452,11.137029,13.399607,15.662184,17.92476,20.187338,17.475147,14.762955,12.050762,9.338571,6.624565,5.2992897,3.974014,2.6505513,1.3252757,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13778515,0.2755703,0.41335547,0.5493277,0.6871128,2.1501737,3.6132345,5.0744824,6.5375433,8.000604,6.550234,5.0998635,3.6494937,2.2009366,0.7505665,1.7495089,2.7502642,3.7492065,4.749962,5.750717,5.7380266,5.7253356,5.712645,5.6999545,5.6872635,4.7118897,3.736516,2.762955,1.7875811,0.8122072,3.1744974,3.2343252,3.294153,3.3557937,3.4156215,3.4754493,4.2006345,4.9258194,5.6491914,6.3743763,7.0995617,11.724429,16.349297,20.975977,25.600845,30.225712,28.369238,26.514578,24.659918,22.805256,20.950596,20.907085,20.865387,20.821875,20.780178,20.736666,19.77942,18.822178,17.864933,16.907688,15.950445,24.224806,32.49917,40.77534,49.0497,57.32588,48.110588,38.895298,29.68001,20.464722,11.249433,9.712041,8.174648,6.637256,5.0998635,3.5624714,4.0102735,4.458075,4.9058766,5.351866,5.7996674,6.492219,7.1847706,7.877322,8.569874,9.262425,9.354887,9.447348,9.539809,9.63227,9.724731,10.205167,10.685601,11.164224,11.644659,12.125093,9.936848,7.750415,5.562169,3.3757362,1.1874905,1.1802386,1.1729867,1.1657349,1.1566701,1.1494182,1.017072,0.88472575,0.7523795,0.6200332,0.48768693,0.823085,1.1566701,1.4920682,1.8274662,2.1628644,2.1556125,2.1483607,2.1392958,2.132044,2.124792,2.1229792,2.1193533,2.1175404,2.1157274,2.1121013,2.077655,2.0432088,2.0069497,1.9725033,1.938057,2.0196402,2.1030366,2.18462,2.268016,2.3495996,2.6976883,3.045777,3.392053,3.7401419,4.0882306,5.3591175,6.6318173,7.9045167,9.177217,10.449916,10.203354,9.954978,9.706602,9.460039,9.211663,8.72035,8.227224,7.7340984,7.2427855,6.7496595,6.787732,6.825804,6.8620634,6.9001355,6.9382076,6.7134004,6.48678,6.261973,6.037165,5.812358,6.115123,6.4178877,6.720652,7.021604,7.324369,7.6724577,8.020547,8.366822,8.714911,9.063,9.644961,10.226922,10.810696,11.392657,11.974618,12.106964,12.23931,12.371656,12.5058155,12.638163,12.830337,13.022511,13.2146845,13.406858,13.600845,13.715062,13.829279,13.945308,14.059525,14.175554,12.754191,11.334642,9.915092,8.495543,7.07418,6.7025228,6.3308654,5.957395,5.5857377,5.2122674,4.7717175,4.3329806,3.8924308,3.4518807,3.0131438,3.005892,2.9968271,2.9895754,2.9823234,2.9750717,3.3267863,3.680314,4.0320287,4.3855567,4.7372713,4.797099,4.856927,4.9167547,4.9783955,5.038223,8.372261,11.708113,15.0421505,18.378002,21.71204,21.097446,20.482851,19.868258,19.25185,18.637255,18.622751,18.608248,18.59193,18.577427,18.562923,16.840609,15.118295,13.394168,11.671853,9.949538,8.624263,7.3008003,5.975525,4.650249,3.3249733,4.322103,5.319232,6.3181744,7.315304,8.312433,7.2047133,6.096993,4.989273,3.8833659,2.7756457,2.9224956,3.0693457,3.2180085,3.3648586,3.5117085,4.554162,5.5966153,6.640882,7.6833353,8.725789,7.8120556,6.9001355,5.9882154,5.0744824,4.162562,4.1099863,4.0574102,4.004834,3.9522583,3.8996825,4.2441454,4.590421,4.934884,5.279347,5.6256227,6.089741,6.5556726,7.019791,7.4857225,7.949841,8.497355,9.04487,9.592385,10.139899,10.687414,12.134158,13.582716,15.02946,16.478018,17.92476,15.693004,13.4594345,11.227677,8.994107,6.7623506,6.3091097,5.857682,5.4044414,4.953014,4.499773,4.3166637,4.135368,3.9522583,3.7691493,3.587853,4.3547363,5.121619,5.8903155,6.6571984,7.4258947,6.1278133,4.8297324,3.531651,2.2353828,0.93730164,0.87566096,0.8122072,0.7505665,0.6871128,0.62547207,0.5094425,0.39522585,0.27919623,0.16497959,0.05076295,1.1004683,2.1501737,3.199879,4.249584,5.2992897,4.853301,4.405499,3.9576974,3.5098956,3.0620937,3.8199122,4.5777307,5.335549,6.093367,6.849373,5.6655083,4.4798307,3.294153,2.1102884,0.9246109,1.79302,2.659616,3.5280252,4.3946214,5.2630305,5.812358,6.3616858,6.9128265,7.462154,8.013294,6.4197006,4.8279195,3.2343252,1.6425442,0.05076295,0.20486477,0.36077955,0.5148814,0.67079616,0.824898,2.864481,4.9040637,6.94546,8.985043,11.024626,12.329959,13.635292,14.940624,16.244144,17.549479,23.354584,29.15969,34.964798,40.7699,46.57501,38.95875,31.34431,23.729868,16.115425,8.499168,7.567306,6.635443,5.7017674,4.7699046,3.8380418,3.720199,3.6023567,3.484514,3.3666716,3.2506418,3.5806012,3.9105604,4.2405195,4.5704784,4.900438,3.9431937,2.9841363,2.0268922,1.0696479,0.11240368,0.15228885,0.19217403,0.23205921,0.27194437,0.31182957,0.2955129,0.27738327,0.25925365,0.24293698,0.22480737,0.1794833,0.13415924,0.09064813,0.045324065,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.02175555,0.032633327,0.04169814,0.052575916,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.14503701,0.22662032,0.3100166,0.39159992,0.4749962,1.551896,2.6306088,3.7075086,4.784408,5.863121,5.89938,5.9374523,5.975525,6.011784,6.049856,7.170267,8.290678,9.409276,10.529687,11.650098,11.18054,10.70917,10.239613,9.770056,9.300498,8.94697,8.595256,8.241728,7.890013,7.5382986,9.052122,10.567759,12.083396,13.597219,15.112856,12.9427395,10.772624,8.602508,6.432391,4.262275,4.974769,5.6872635,6.399758,7.112252,7.8247466,7.9081426,7.989726,8.073122,8.154706,8.238102,7.647076,7.057863,6.4668374,5.8776245,5.2865987,4.3366065,3.388427,2.4366217,1.4866294,0.53663695,2.4474995,4.3565493,6.2674117,8.178274,10.087324,10.2142315,10.342952,10.469859,10.596766,10.725487,9.9422865,9.1609,8.3777,7.5945,6.813113,5.9392653,5.06723,4.195195,3.3231604,2.4493124,2.9805105,3.5098956,4.0392804,4.5704784,5.0998635,8.365009,11.630155,14.895301,18.160446,21.425592,19.585434,17.745277,15.905121,14.064963,12.224807,11.338268,10.449916,9.563377,8.675026,7.7866745,7.6742706,7.5618668,7.4494634,7.3370595,7.224656,6.0299134,4.835171,3.6404288,2.4456866,1.2491312,1.0007553,0.7505665,0.50037766,0.25018883,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.08520924,0.09427405,0.10515183,0.11421664,0.12509441,0.13234627,0.13959812,0.14684997,0.15410182,0.16316663,0.15228885,0.14322405,0.13234627,0.12328146,0.11240368,0.11059072,0.10696479,0.10515183,0.10333887,0.099712946,0.21755551,0.33539808,0.45324063,0.56927025,0.6871128,1.2527572,1.8165885,2.382233,2.9478772,3.5117085,5.9447045,8.3777,10.810696,13.2418785,15.674874,15.877926,16.079165,16.282217,16.48527,16.68832,17.67276,18.657198,19.641636,20.627888,21.612328,21.02674,20.442966,19.85738,19.271791,18.688019,18.677141,18.668076,18.657198,18.648132,18.637255,17.170568,15.702069,14.235382,12.766883,11.300196,11.334642,11.370901,11.405348,11.439794,11.47424,11.011934,10.549629,10.087324,9.625018,9.162713,9.354887,9.547061,9.739235,9.933222,10.125396,11.827768,13.53014,15.2325115,16.934883,18.637255,16.207886,13.776703,11.347333,8.917963,6.48678,5.1905117,3.8924308,2.5943494,1.2980812,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.42423326,0.73787576,1.0497054,1.3633479,1.6751775,2.956942,4.2405195,5.522284,6.8040485,8.087626,6.9382076,5.7869763,4.6375585,3.48814,2.3369088,3.1781235,4.017525,4.856927,5.6981416,6.5375433,6.412449,6.2873545,6.16226,6.037165,5.9120708,4.896812,3.881553,2.8681068,1.8528478,0.8375887,3.2869012,3.3449159,3.4029307,3.4591327,3.5171473,3.5751622,4.40006,5.224958,6.049856,6.874754,7.699652,12.411542,17.125244,21.837133,26.550837,31.262726,29.252151,27.24339,25.232813,23.222239,21.211662,21.353073,21.492672,21.632269,21.771868,21.913279,20.872639,19.831997,18.79317,17.75253,16.71189,23.974617,31.237345,38.500072,45.762802,53.025528,44.370445,35.715363,27.06028,18.405195,9.750113,8.649645,7.549176,6.450521,5.3500524,4.249584,4.606738,4.9657044,5.3228583,5.6800117,6.037165,6.434204,6.833056,7.230095,7.6271334,8.024173,8.047741,8.069496,8.093065,8.1148205,8.138389,8.471974,8.807372,9.142771,9.4781685,9.811753,8.287052,6.7623506,5.237649,3.7129474,2.1882458,2.0105755,1.8329052,1.6552348,1.4775645,1.2998942,1.2346275,1.1693609,1.1059072,1.0406405,0.97537386,1.1204109,1.2654479,1.4104849,1.5555218,1.7005589,1.6842422,1.6697385,1.6552348,1.6407311,1.6244144,1.6207886,1.6153497,1.6099107,1.6044719,1.6008459,1.9416829,2.2843328,2.6269827,2.9696326,3.3122826,3.2270734,3.141864,3.056655,2.9732587,2.8880494,2.956942,3.0276475,3.0983531,3.1672456,3.2379513,4.4707656,5.7017674,6.9345818,8.167397,9.400211,9.004985,8.609759,8.214534,7.819308,7.424082,7.1521373,6.880193,6.6082487,6.3344913,6.0625467,6.011784,5.962834,5.9120708,5.863121,5.812358,5.674573,5.5367875,5.4008155,5.2630305,5.125245,5.4552045,5.7851634,6.115123,6.445082,6.775041,7.0451727,7.315304,7.5854354,7.855567,8.125698,8.827314,9.530745,10.232361,10.93579,11.637406,11.664601,11.691795,11.720803,11.747997,11.775192,12.085209,12.395226,12.705242,13.015259,13.325275,13.229188,13.134913,13.04064,12.944552,12.850279,11.697234,10.54419,9.39296,8.239915,7.0868707,6.7677894,6.446895,6.1278133,5.806919,5.487838,4.894999,4.3021603,3.7093215,3.1182957,2.525457,2.572594,2.619731,2.666868,2.715818,2.762955,3.092914,3.4228733,3.7528327,4.082792,4.4127507,4.519716,4.6266804,4.7354584,4.842423,4.949388,7.844689,10.73999,13.635292,16.530592,19.424082,19.520168,19.614443,19.71053,19.804804,19.90089,19.507477,19.115877,18.722466,18.330864,17.937452,16.43088,14.922495,13.41411,11.907538,10.399154,8.999546,7.5999393,6.200332,4.800725,3.3993049,4.507025,5.614745,6.722465,7.8301854,8.937905,7.5981264,6.258347,4.9167547,3.576975,2.2371957,2.420305,2.6016014,2.7847104,2.9678197,3.149116,4.2858434,5.4207582,6.5556726,7.690587,8.825501,8.074935,7.324369,6.5756154,5.825049,5.0744824,4.9820213,4.88956,4.797099,4.704638,4.612177,5.4407005,6.2674117,7.0959353,7.9226465,8.749357,8.805559,8.859948,8.914337,8.970539,9.024928,9.157274,9.28962,9.421967,9.554313,9.686659,11.419851,13.153044,14.884423,16.617615,18.350807,15.95951,13.5700245,11.18054,8.789243,6.399758,6.0208488,5.6401267,5.2594047,4.880495,4.499773,4.510651,4.519716,4.5305934,4.539658,4.550536,5.3482394,6.14413,6.9418335,7.7395372,8.537241,7.017978,5.4969025,3.97764,2.4583774,0.93730164,0.93730164,0.93730164,0.93730164,0.93730164,0.93730164,0.75781834,0.57833505,0.39703882,0.21755551,0.038072214,1.7875811,3.53709,5.2884116,7.037921,8.78743,8.241728,7.6978393,7.1521373,6.6082487,6.0625467,5.8776245,5.6927023,5.5077806,5.3228583,5.137936,4.4671397,3.7981565,3.1273603,2.4583774,1.7875811,2.4855716,3.1817493,3.87974,4.5777307,5.275721,5.612932,5.9501433,6.2873545,6.624565,6.9617763,5.576673,4.1933823,2.808279,1.4231756,0.038072214,0.3480888,0.65810543,0.968122,1.2781386,1.5881553,3.1182957,4.646623,6.1767635,7.706904,9.237044,10.310318,11.381779,12.455053,13.528327,14.599788,18.747847,22.89409,27.04215,31.190208,35.33827,29.544039,23.753435,17.959208,12.166792,6.3743763,5.7597823,5.145188,4.5305934,3.9141862,3.299592,3.1273603,2.955129,2.7828975,2.610666,2.4366217,2.6849976,2.9333735,3.1799364,3.4283123,3.6748753,2.9841363,2.2952106,1.6044719,0.9155461,0.22480737,0.3045777,0.38434806,0.46411842,0.54570174,0.62547207,0.58921283,0.55476654,0.52032024,0.48587397,0.44961473,0.36077955,0.27013144,0.1794833,0.09064813,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.032633327,0.03988518,0.047137026,0.054388877,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.22662032,0.39159992,0.55839247,0.72337204,0.8883517,1.6044719,2.322405,3.0403383,3.7582715,4.4743915,4.5867953,4.699199,4.8116026,4.9258194,5.038223,5.9392653,6.8421206,7.744976,8.647832,9.550687,9.385707,9.220728,9.055748,8.890768,8.725789,8.781991,8.840006,8.898021,8.954222,9.012237,10.154404,11.29657,12.440549,13.582716,14.724882,12.509441,10.2958145,8.080374,5.864934,3.6494937,4.5632267,5.475147,6.3870673,7.3008003,8.212721,7.9280853,7.6416373,7.3570023,7.072367,6.787732,6.4831543,6.1767635,5.8721857,5.567608,5.2630305,4.4127507,3.5624714,2.712192,1.8619126,1.0116332,2.420305,3.827164,5.235836,6.642695,8.049554,9.429218,10.810696,12.19036,13.5700245,14.94969,13.372412,11.795135,10.217857,8.640579,7.063302,6.604623,6.147756,5.6908894,5.23221,4.7753434,4.646623,4.519716,4.3928084,4.265901,4.137181,11.4688015,18.796797,26.128416,33.458225,40.788033,34.845142,28.90225,22.959358,17.01828,11.075388,10.674724,10.275872,9.875207,9.474543,9.07569,8.363196,7.650702,6.9382076,6.2257137,5.5132194,4.610364,3.7075086,2.8046532,1.9017978,1.0007553,0.7995165,0.6000906,0.40066472,0.19942589,0.0,0.0,0.0,0.0,0.0,0.0,0.018129626,0.034446288,0.052575916,0.07070554,0.0870222,0.09427405,0.10333887,0.11059072,0.11784257,0.12509441,0.12690738,0.13053331,0.13234627,0.13415924,0.13778515,0.13053331,0.12328146,0.11421664,0.10696479,0.099712946,0.09427405,0.09064813,0.08520924,0.07977036,0.07433146,0.17223145,0.27013144,0.3680314,0.46411842,0.5620184,1.5917811,2.6233568,3.6531196,4.6828823,5.712645,7.802991,9.893337,11.98187,14.072216,16.162561,17.01828,17.872185,18.727903,19.581808,20.437527,20.870825,21.30231,21.73561,22.167093,22.600391,21.73017,20.859947,19.989725,19.119503,18.24928,18.004532,17.75978,17.515032,17.27028,17.025532,15.890617,14.755702,13.620788,12.485873,11.349146,11.608399,11.86584,12.123281,12.380721,12.638163,11.862214,11.088079,10.312131,9.537996,8.762048,9.284182,9.808127,10.330261,10.852394,11.374527,12.516694,13.660673,14.802839,15.945006,17.087172,14.940624,12.792264,10.645717,8.497355,6.350808,5.0799212,3.8090343,2.5399606,1.2708868,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.045324065,0.09064813,0.13415924,0.1794833,0.22480737,0.7124943,1.2001812,1.6878681,2.175555,2.663242,3.7655232,4.8678045,5.9700856,7.072367,8.174648,7.324369,6.474089,5.6256227,4.7753434,3.925064,4.604925,5.2847857,5.964647,6.644508,7.324369,7.0868707,6.849373,6.6118746,6.3743763,6.1368785,5.081734,4.02659,2.9732587,1.9181144,0.8629702,3.3993049,3.4555066,3.5098956,3.5642843,3.6204863,3.6748753,4.599486,5.524097,6.450521,7.3751316,8.299743,13.100468,17.89938,22.700104,27.50083,32.29974,30.135063,27.970387,25.80571,23.63922,21.474543,21.797249,22.119957,22.442663,22.765371,23.088078,21.965855,20.841818,19.719595,10258.0,17.475147,23.724428,29.975523,36.224804,42.4759,48.72518,40.630306,32.535427,24.440548,16.34567,8.2507925,7.5872483,6.925517,6.261973,5.600241,4.936697,5.2050157,5.473334,5.7398396,6.008158,6.2746634,6.378002,6.4795284,6.582867,6.684393,6.787732,6.740595,6.6916447,6.644508,6.5973706,6.550234,6.740595,6.929143,7.119504,7.309865,7.500226,6.637256,5.774286,4.9131284,4.0501585,3.1871881,2.8409123,2.4928236,2.1447346,1.7966459,1.4503701,1.452183,1.455809,1.4576219,1.4594349,1.4630609,1.4177368,1.3724127,1.3270886,1.2817645,1.2382535,1.214685,1.1929294,1.1693609,1.1476053,1.1258497,1.1167849,1.1095331,1.1022812,1.0950294,1.0877775,1.8075237,2.5272698,3.247016,3.966762,4.688321,4.4345064,4.1825047,3.930503,3.6766882,3.4246864,3.2180085,3.009518,2.8028402,2.5943494,2.3876717,3.5806012,4.7717175,5.964647,7.157576,8.350506,7.806617,7.264541,6.722465,6.1803894,5.638314,5.5857377,5.5331616,5.480586,5.42801,5.375434,5.237649,5.0998635,4.9620786,4.8242936,4.688321,4.6375585,4.5867953,4.537845,4.4870825,4.4381323,4.795286,5.1524396,5.5095935,5.866747,6.2257137,6.4178877,6.6100616,6.8022356,6.9944096,7.1865835,8.009668,8.832754,9.655839,10.477111,11.300196,11.222239,11.144281,11.068136,10.990179,10.912222,11.340081,11.7679405,12.195799,12.621845,13.049705,12.745127,12.440549,12.134158,11.829581,11.525003,10.640278,9.755551,8.870826,7.9842873,7.0995617,6.833056,6.5647373,6.298232,6.0299134,5.763408,5.0182805,4.273153,3.5280252,2.7828975,2.03777,2.1392958,2.2426348,2.3441606,2.4474995,2.5508385,2.857229,3.1654327,3.4718235,3.780027,4.0882306,4.2423325,4.3982472,4.552349,4.708264,4.8623657,7.317117,9.771869,12.228433,14.683184,17.137936,17.94289,18.747847,19.552801,20.357758,21.162712,20.392202,19.621695,18.852999,18.082489,17.31198,16.019337,14.726695,13.435865,12.143224,10.850581,9.374829,7.900891,6.4251394,4.949388,3.4754493,4.691947,5.910258,7.1267557,8.345067,9.563377,7.989726,6.4178877,4.844236,3.2723975,1.7005589,1.9181144,2.13567,2.3532255,2.570781,2.7883365,4.0157123,5.243088,6.4704633,7.6978393,8.925215,8.337815,7.750415,7.1630154,6.5756154,5.9882154,5.8558693,5.7217097,5.5893636,5.4570174,5.3246713,6.635443,7.944402,9.255174,10.565946,11.874905,11.519565,11.164224,10.810696,10.455356,10.100015,9.817192,9.53437,9.253361,8.970539,8.6877165,10.705544,12.721559,14.739386,16.757214,18.77504,16.227829,13.680615,11.13159,8.584378,6.037165,5.730775,5.422571,5.1143675,4.8079767,4.499773,4.702825,4.9058766,5.1071157,5.3101673,5.5132194,6.33993,7.166641,7.995165,8.821876,9.6504,7.9081426,6.165886,4.421816,2.6795588,0.93730164,1.0007553,1.062396,1.1258497,1.1874905,1.2491312,1.0043813,0.75963134,0.5148814,0.27013144,0.025381476,2.474694,4.9258194,7.3751316,9.824444,12.27557,11.631968,10.990179,10.348391,9.704789,9.063,7.935337,6.8076744,5.6800117,4.552349,3.4246864,3.2705846,3.1146698,2.960568,2.8046532,2.6505513,3.1781235,3.7056956,4.233268,4.76084,5.2865987,5.411693,5.5367875,5.661882,5.7869763,5.9120708,4.7354584,3.5570326,2.38042,1.2019942,0.025381476,0.4894999,0.9554313,1.4195497,1.8854811,2.3495996,3.3702974,4.3891826,5.40988,6.430578,7.4494634,8.290678,9.130079,9.969481,10.810696,11.650098,14.139296,16.630306,19.119503,21.610514,24.099712,20.129324,16.160748,12.19036,8.219973,4.249584,3.9522583,3.6549325,3.3576066,3.0602808,2.762955,2.5345216,2.3079014,2.079468,1.8528478,1.6244144,1.789394,1.9543737,2.1193533,2.2843328,2.4493124,2.0268922,1.6044719,1.1820517,0.75963134,0.33721104,0.45686656,0.57833505,0.6979906,0.81764615,0.93730164,0.88472575,0.8321498,0.7795739,0.726998,0.6744221,0.5402629,0.40429065,0.27013144,0.13415924,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.04169814,0.047137026,0.052575916,0.058014803,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.3100166,0.55839247,0.80495536,1.0533313,1.2998942,1.6570477,2.0142014,2.373168,2.7303216,3.0874753,3.2742105,3.4627585,3.6494937,3.8380418,4.024777,4.710077,5.3953767,6.0806766,6.7641635,7.4494634,7.590874,7.7304726,7.8700705,8.009668,8.149267,8.617011,9.084756,9.5525,10.020245,10.487988,11.256684,12.027194,12.797703,13.568212,14.336908,12.077957,9.817192,7.558241,5.297477,3.0367124,4.1498713,5.2630305,6.3743763,7.4875355,8.600695,7.948028,7.2953615,6.642695,5.9900284,5.337362,5.317419,5.297477,5.277534,5.2575917,5.237649,4.4870825,3.738329,2.9877625,2.2371957,1.4866294,2.3931105,3.2977788,4.2024474,5.1071157,6.011784,8.646019,11.276628,13.910862,16.543283,19.175705,16.802538,14.429369,12.058014,9.684846,7.311678,7.26998,7.228282,7.1847706,7.1430726,7.0995617,6.3145485,5.529536,4.744523,3.9595103,3.1744974,14.57078,25.96525,37.35972,48.756004,60.15047,50.104847,40.061035,30.015408,19.969784,9.924157,10.012992,10.100015,10.1870365,10.275872,10.362894,9.050309,7.7377243,6.4251394,5.1125546,3.7999697,3.1908143,2.5798457,1.9706904,1.3597219,0.7505665,0.6000906,0.44961473,0.2991388,0.15047589,0.0,0.0,0.0,0.0,0.0,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.10515183,0.11059072,0.11421664,0.11965553,0.12509441,0.12328146,0.11965553,0.11784257,0.11421664,0.11240368,0.10696479,0.10333887,0.09789998,0.092461094,0.0870222,0.07977036,0.072518505,0.065266654,0.058014803,0.05076295,0.12690738,0.20486477,0.28282216,0.36077955,0.43692398,1.9326181,3.4283123,4.9221935,6.4178877,7.911769,9.659465,11.407161,13.154857,14.902553,16.650248,18.15682,19.665205,21.171778,22.680162,24.186733,24.067078,23.947422,23.827766,23.70811,23.586643,22.431786,21.276928,20.122072,18.967215,17.812357,17.331923,16.8533,16.372866,15.89243,15.411995,14.610665,13.807523,13.00438,12.203052,11.399909,11.880343,12.360779,12.839401,13.319836,13.800271,12.712494,11.624716,10.536939,9.449161,8.363196,9.215289,10.067381,10.919474,11.771566,12.625471,13.207433,13.789393,14.373167,14.955129,15.537089,13.671551,11.807825,9.9422865,8.076748,6.2130227,4.9693303,3.727451,2.4855716,1.2418793,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.06707962,0.13415924,0.2030518,0.27013144,0.33721104,1.0007553,1.6624867,2.324218,2.9877625,3.6494937,4.572292,5.4950895,6.4178877,7.3406854,8.26167,7.7123427,7.1630154,6.6118746,6.0625467,5.5132194,6.0317264,6.552047,7.072367,7.592687,8.113008,7.763106,7.413204,7.063302,6.7134004,6.3616858,5.2666564,4.171627,3.0765975,1.983381,0.8883517,3.5117085,3.5642843,3.6168604,3.6694362,3.7220123,3.774588,4.800725,5.825049,6.849373,7.8755093,8.899834,13.7875805,18.675327,23.563074,28.45082,33.336758,31.017977,28.697384,26.376793,24.058014,21.737421,22.243238,22.747242,23.253057,23.757061,24.262878,23.057259,21.851639,20.647831,19.442211,18.238403,23.47424,28.71189,33.94954,39.187187,44.424835,36.890163,29.35549,21.819004,14.284332,6.7496595,6.5248523,6.300045,6.0752378,5.8504305,5.6256227,5.803293,5.979151,6.156821,6.3344913,6.5121617,6.319988,6.1278133,5.9356394,5.7416525,5.5494785,5.431636,5.315606,5.197764,5.0799212,4.9620786,5.0074024,5.0527267,5.0980506,5.143375,5.186886,4.98746,4.788034,4.5867953,4.3873696,4.1879435,3.6694362,3.152742,2.6342347,2.1175404,1.6008459,1.6697385,1.7404441,1.8093367,1.8800422,1.9507477,1.7150626,1.4793775,1.2455053,1.0098201,0.774135,0.7451276,0.71430725,0.6852999,0.6544795,0.62547207,0.61459434,0.6055295,0.5946517,0.5855869,0.5747091,1.6733645,2.770207,3.8670492,4.9657044,6.0625467,5.6419396,5.223145,4.802538,4.3819304,3.9631362,3.4772623,2.9932013,2.5073273,2.0232663,1.5373923,2.6904364,3.8416677,4.994712,6.147756,7.3008003,6.6100616,5.919323,5.230397,4.539658,3.8507326,4.017525,4.1843176,4.3529234,4.519716,4.688321,4.461701,4.2368937,4.0120864,3.787279,3.5624714,3.6005437,3.636803,3.6748753,3.7129474,3.7492065,4.135368,4.519716,4.9058766,5.290225,5.674573,5.7906027,5.904819,6.0208488,6.1350656,6.249282,7.192023,8.134763,9.077503,10.020245,10.962985,10.779876,10.596766,10.41547,10.232361,10.049252,10.594954,11.1406555,11.684544,12.230246,12.774135,12.259253,11.744371,11.22949,10.714609,10.199727,9.583321,8.9651,8.34688,7.7304726,7.112252,6.8983226,6.68258,6.4668374,6.2529078,6.037165,5.139749,4.2423325,3.3449159,2.4474995,1.550083,1.7078108,1.8655385,2.0232663,2.179181,2.3369088,2.6233568,2.907992,3.1926272,3.4772623,3.7618973,3.9649491,4.168001,4.36924,4.572292,4.7753434,6.789545,8.805559,10.81976,12.835775,14.849977,16.365614,17.879436,19.395073,20.910711,22.424534,21.276928,20.129324,18.981718,17.834112,16.68832,15.609608,14.532708,13.455809,12.377095,11.300196,9.750113,8.200029,6.6499467,5.0998635,3.5497808,4.876869,6.205771,7.5328593,8.859948,10.1870365,8.383139,6.5774283,4.7717175,2.9678197,1.162109,1.4141108,1.6679256,1.9199274,2.1719291,2.4257438,3.7455807,5.0654173,6.3852544,7.705091,9.024928,8.600695,8.174648,7.750415,7.324369,6.9001355,6.7279043,6.5556726,6.3816285,6.209397,6.037165,7.8301854,9.623205,11.4144125,13.207433,15.000452,14.235382,13.470312,12.705242,11.940171,11.175101,10.477111,9.77912,9.082943,8.384952,7.686961,9.989424,12.291886,14.594349,16.89681,19.199274,16.494333,13.789393,11.084454,8.379513,5.674573,5.4407005,5.2050157,4.9693303,4.7354584,4.499773,4.894999,5.290225,5.6854506,6.0806766,6.4759026,7.3316207,8.189152,9.046683,9.904215,10.761745,8.798307,6.833056,4.8678045,2.902553,0.93730164,1.062396,1.1874905,1.3125849,1.4376793,1.5627737,1.2527572,0.94274056,0.6327239,0.32270733,0.012690738,3.1618068,6.3127356,9.461852,12.612781,15.761897,15.022208,14.282519,13.54283,12.803142,12.06164,9.99305,7.9226465,5.8522434,3.7818398,1.7132497,2.0722163,2.4329958,2.7919624,3.152742,3.5117085,3.870675,4.227829,4.5849824,4.942136,5.2992897,5.2122674,5.125245,5.038223,4.949388,4.8623657,3.8924308,2.9224956,1.9525607,0.9826257,0.012690738,0.6327239,1.2527572,1.8727903,2.4928236,3.1128569,3.6222992,4.1317415,4.6429973,5.1524396,5.661882,6.2692246,6.87838,7.4857225,8.093065,8.700407,9.5325575,10.364707,11.1968565,12.03082,12.862969,10.714609,8.568061,6.4197006,4.273153,2.124792,2.1447346,2.1646774,2.18462,2.2045624,2.2245052,1.9416829,1.6606737,1.3778516,1.0950294,0.8122072,0.89560354,0.97718686,1.0605831,1.1421664,1.2255627,1.0696479,0.9155461,0.75963134,0.6055295,0.44961473,0.6091554,0.7705091,0.9300498,1.0895905,1.2491312,1.1802386,1.1095331,1.0406405,0.969935,0.89922947,0.7197462,0.5402629,0.36077955,0.1794833,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.052575916,0.054388877,0.058014803,0.059827764,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.3934129,0.72337204,1.0533313,1.3832904,1.7132497,1.7096237,1.7078108,1.7041848,1.7023718,1.7005589,1.9616255,2.2245052,2.4873846,2.7502642,3.0131438,3.4808881,3.9468195,4.4145637,4.882308,5.3500524,5.7942286,6.240217,6.684393,7.130382,7.574558,8.452031,9.329506,10.20698,11.084454,11.961927,12.360779,12.757817,13.154857,13.551895,13.9507475,11.644659,9.340384,7.0342946,4.7300196,2.4257438,3.738329,5.049101,6.3616858,7.6742706,8.9868555,7.9679704,6.947273,5.9265747,4.9076896,3.8869917,4.1516843,4.41819,4.6828823,4.947575,5.2122674,4.5632267,3.9123733,3.2633326,2.612479,1.9616255,2.3659163,2.7683938,3.1708715,3.5733492,3.975827,7.861006,11.744371,15.62955,19.514729,23.399908,20.232662,17.065416,13.898171,10.729113,7.5618668,7.935337,8.306994,8.680465,9.052122,9.425592,7.9824743,6.539356,5.0980506,3.6549325,2.2118144,17.67276,33.13189,48.592834,64.05197,79.51292,65.364555,51.218006,37.069645,22.9231,8.774739,9.349448,9.924157,10.500679,11.075388,11.650098,9.737422,7.8247466,5.9120708,3.9993954,2.08672,1.7694515,1.452183,1.1349145,0.81764615,0.50037766,0.40066472,0.2991388,0.19942589,0.099712946,0.0,0.0,0.0,0.0,0.0,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.11421664,0.11784257,0.11965553,0.12328146,0.12509441,0.11784257,0.11059072,0.10333887,0.09427405,0.0870222,0.08520924,0.08339628,0.07977036,0.07795739,0.07433146,0.065266654,0.054388877,0.045324065,0.034446288,0.025381476,0.08339628,0.13959812,0.19761293,0.25562772,0.31182957,2.2734551,4.233268,6.19308,8.152893,10.112705,11.517752,12.922797,14.327844,15.732889,17.137936,19.297174,21.458225,23.617464,25.776703,27.937754,27.265144,26.592535,25.919926,25.247316,24.574707,23.135216,21.695723,20.254417,18.814926,17.375433,16.659313,15.945006,15.230699,14.514579,13.800271,13.330714,12.859344,12.389787,11.920229,11.450671,12.152288,12.855718,13.557334,14.260764,14.96238,13.562773,12.163166,10.761745,9.362139,7.9625316,9.144584,10.326634,11.510499,12.692551,13.874602,13.898171,13.919927,13.941682,13.965251,13.987006,12.40429,10.823386,9.24067,7.6579537,6.0752378,4.860553,3.644055,2.42937,1.214685,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.09064813,0.1794833,0.27013144,0.36077955,0.44961473,1.2872034,2.124792,2.962381,3.7999697,4.6375585,5.3808727,6.1223745,6.8656893,7.607191,8.350506,8.100317,7.850128,7.5999393,7.3497505,7.0995617,7.460341,7.819308,8.180087,8.540867,8.899834,8.437528,7.9752226,7.512917,7.0506115,6.588306,5.4515786,4.3166637,3.1817493,2.0468347,0.9119202,3.6241121,3.6748753,3.7256382,3.774588,3.825351,3.874301,5.0001507,6.1241875,7.250037,8.375887,9.499924,14.474693,19.449463,24.426044,29.400814,34.375584,31.90089,29.424383,26.949688,24.474995,22.000301,22.687414,23.374527,24.06164,24.750565,25.437677,24.150475,22.863272,21.574255,20.287052,18.999847,23.22405,27.450066,31.674269,35.900284,40.12449,33.15002,26.175554,19.199274,12.224807,5.2503395,5.462456,5.674573,5.8866897,6.1006193,6.3127356,6.399758,6.48678,6.5756154,6.6626377,6.7496595,6.261973,5.774286,5.2865987,4.800725,4.313038,4.12449,3.9377546,3.7492065,3.5624714,3.3757362,3.2742105,3.1744974,3.0747845,2.9750717,2.8753586,3.3376641,3.7999697,4.262275,4.7245803,5.186886,4.499773,3.8126602,3.1255474,2.4366217,1.7495089,1.887294,2.0250793,2.1628644,2.3006494,2.4366217,2.0123885,1.5881553,1.162109,0.73787576,0.31182957,0.2755703,0.2374981,0.19942589,0.16316663,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,1.5373923,3.0131438,4.4870825,5.962834,7.4367723,6.849373,6.261973,5.674573,5.087173,4.499773,3.738329,2.9750717,2.2118144,1.4503701,0.6871128,1.8002719,2.911618,4.024777,5.137936,6.249282,5.411693,4.5759177,3.738329,2.9007401,2.0631514,2.4493124,2.8372865,3.2252605,3.6132345,3.9993954,3.6875658,3.3757362,3.0620937,2.7502642,2.4366217,2.561716,2.6868105,2.811905,2.9369993,3.0620937,3.4754493,3.8869917,4.3003473,4.7118897,5.125245,5.163317,5.199577,5.237649,5.275721,5.3119802,6.3743763,7.4367723,8.499168,9.563377,10.625773,10.337513,10.049252,9.762803,9.474543,9.188094,9.849826,10.51337,11.175101,11.836833,12.500377,11.775192,11.050007,10.324821,9.599637,8.874452,8.52455,8.174648,7.8247466,7.474845,7.124943,6.9617763,6.8004227,6.637256,6.4759026,6.3127356,5.2630305,4.213325,3.1618068,2.1121013,1.062396,1.2745126,1.4866294,1.7005589,1.9126755,2.124792,2.3876717,2.6505513,2.911618,3.1744974,3.437377,3.6875658,3.9377546,4.1879435,4.4381323,4.688321,6.261973,7.837437,9.412902,10.988366,12.562017,14.788336,17.01284,19.237347,21.461851,23.68817,22.161655,20.636953,19.112251,17.58755,16.062849,15.199879,14.336908,13.475751,12.612781,11.74981,10.125396,8.499168,6.874754,5.2503395,3.6241121,5.0617914,6.4994707,7.93715,9.374829,10.812509,8.774739,6.736969,4.699199,2.663242,0.62547207,0.9119202,1.2001812,1.4866294,1.7748904,2.0631514,3.4754493,4.8877473,6.300045,7.7123427,9.12464,8.861761,8.600695,8.337815,8.074935,7.8120556,7.5999393,7.3878226,7.175706,6.9617763,6.7496595,9.024928,11.300196,13.575464,15.850732,18.124187,16.949387,15.774588,14.599788,13.424988,12.250188,11.137029,10.025683,8.912524,7.799365,6.688019,9.275117,11.862214,14.449312,17.038223,19.62532,16.762651,13.899984,11.037316,8.174648,5.3119802,5.1506267,4.98746,4.8242936,4.6629395,4.499773,5.087173,5.674573,6.261973,6.849373,7.4367723,8.325124,9.211663,10.100015,10.988366,11.874905,9.686659,7.500226,5.3119802,3.1255474,0.93730164,1.1258497,1.3125849,1.49932,1.6878681,1.8746033,1.49932,1.1258497,0.7505665,0.37528324,0.0,3.8507326,7.699652,11.5503845,15.399304,19.250036,18.412449,17.57486,16.73727,15.899682,15.062093,12.050762,9.037619,6.0244746,3.0131438,0.0,0.87566096,1.7495089,2.6251698,3.5008307,4.3746786,4.5632267,4.749962,4.936697,5.125245,5.3119802,5.0128417,4.7118897,4.4127507,4.1117992,3.8126602,3.049403,2.2879589,1.5247015,0.76325727,0.0,0.775948,1.550083,2.324218,3.100166,3.874301,3.874301,3.874301,3.874301,3.874301,3.874301,4.249584,4.6248674,5.0001507,5.375434,5.750717,4.9258194,4.100921,3.2742105,2.4493124,1.6244144,1.2998942,0.97537386,0.6508536,0.3245203,0.0,0.33721104,0.6744221,1.0116332,1.3506571,1.6878681,1.3506571,1.0116332,0.6744221,0.33721104,0.0,0.0,0.0,0.0,0.0,0.0,0.11240368,0.22480737,0.33721104,0.44961473,0.5620184,0.76325727,0.96268314,1.162109,1.3633479,1.5627737,1.4757515,1.3869164,1.2998942,1.2128719,1.1258497,0.89922947,0.6744221,0.44961473,0.22480737,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.4749962,0.8883517,1.2998942,1.7132497,2.124792,1.7621996,1.3996071,1.0370146,0.6744221,0.31182957,0.6508536,0.9880646,1.3252757,1.6624867,1.9996977,2.2498865,2.5000753,2.7502642,3.000453,3.2506418,3.9993954,4.749962,5.5005283,6.249282,6.9998484,8.287052,9.574255,10.863272,12.1504755,13.437678,13.46306,13.486629,13.512011,13.537392,13.562773,11.213174,8.861761,6.5121617,4.162562,1.8129625,3.3249733,4.836984,6.350808,7.8628187,9.374829,7.987913,6.599184,5.2122674,3.825351,2.4366217,2.9877625,3.53709,4.0882306,4.6375585,5.186886,4.6375585,4.0882306,3.53709,2.9877625,2.4366217,2.3369088,2.2371957,2.137483,2.03777,1.938057,7.075993,12.212116,17.350052,22.487988,27.624111,23.662788,19.699652,15.736515,11.775192,7.8120556,8.600695,9.38752,10.174346,10.962985,11.74981,9.6504,7.549176,5.4497657,3.350355,1.2491312,20.77655,40.29853,59.82595,79.34975,98.87535,80.62426,62.374977,44.123882,25.874601,7.6253204,8.6877165,9.750113,10.812509,11.874905,12.937301,10.424535,7.911769,5.4008155,2.8880494,0.37528324,0.34990177,0.3245203,0.2991388,0.2755703,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,2.612479,5.038223,7.462154,9.8878975,12.311829,13.374225,14.436621,15.50083,16.563227,17.625622,20.437527,23.249432,26.06315,28.875055,31.68696,30.463211,29.237648,28.012085,26.788336,25.562773,23.836832,22.112705,20.386765,18.662638,16.936697,15.986704,15.036712,14.0867195,13.136727,12.186734,12.050762,11.912977,11.775192,11.637406,11.499621,12.4242325,13.3506565,14.275268,15.199879,16.124489,14.413053,12.699803,10.986553,9.275117,7.5618668,9.07569,10.587702,12.099712,13.611723,15.125546,14.587097,14.05046,13.512011,12.975373,12.436923,11.137029,9.837135,8.537241,7.2373466,5.9374523,4.749962,3.5624714,2.374981,1.1874905,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.11240368,0.22480737,0.33721104,0.44961473,0.5620184,1.5754645,2.5870976,3.6005437,4.612177,5.6256227,6.187641,6.7496595,7.311678,7.8755093,8.437528,8.488291,8.537241,8.588004,8.636953,8.6877165,8.887142,9.088382,9.287807,9.487233,9.686659,9.11195,8.537241,7.9625316,7.3878226,6.813113,5.638314,4.461701,3.2869012,2.1121013,0.93730164,3.48814,3.5806012,3.673062,3.7655232,3.8579843,3.9504454,5.08536,6.2202744,7.3551893,8.490104,9.625018,14.462003,19.298986,24.137783,28.974768,33.811752,31.376944,28.942135,26.507326,24.072517,21.637709,22.087322,22.536938,22.988365,23.43798,23.887594,23.445232,23.002869,22.560507,22.118143,21.675781,24.629097,27.584227,30.539354,33.494484,36.44961,30.115122,23.78063,17.444326,11.109835,4.7753434,5.0998635,5.424384,5.750717,6.0752378,6.399758,6.2220874,6.0444174,5.866747,5.6908894,5.5132194,5.1179934,4.7227674,4.327542,3.9323158,3.53709,3.587853,3.636803,3.6875658,3.738329,3.787279,4.1444325,4.503399,4.860553,5.217706,5.57486,5.7978544,6.0208488,6.24203,6.4650245,6.688019,6.0770507,5.467895,4.856927,4.2477713,3.636803,3.4228733,3.207131,2.9932013,2.7774587,2.561716,2.1483607,1.7331922,1.3180238,0.90285534,0.48768693,0.40972954,0.33177215,0.25562772,0.17767033,0.099712946,0.10333887,0.10515183,0.10696479,0.11059072,0.11240368,1.49932,2.8880494,4.274966,5.661882,7.0506115,6.359873,5.669134,4.9802084,4.2894692,3.6005437,2.9950142,2.3894846,1.7857682,1.1802386,0.5747091,1.5174497,2.4601903,3.4029307,4.345671,5.2865987,4.5632267,3.8380418,3.1128569,2.3876717,1.6624867,2.0123885,2.3622901,2.712192,3.0620937,3.4119956,3.3068438,3.2016919,3.0983531,2.9932013,2.8880494,2.9224956,2.956942,2.9932013,3.0276475,3.0620937,3.3702974,3.6766882,3.9848917,4.2930956,4.599486,4.7191415,4.84061,4.9602656,5.0799212,5.199577,6.1006193,6.9998484,7.900891,8.80012,9.699349,9.512614,9.325879,9.137331,8.950596,8.762048,9.20985,9.657652,10.1054535,10.553255,10.999244,10.352016,9.704789,9.057561,8.410334,7.763106,7.5328593,7.3026133,7.072367,6.8421206,6.6118746,6.492219,6.3725634,6.2529078,6.1332526,6.011784,5.041849,4.071914,3.101979,2.132044,1.162109,1.5120108,1.8619126,2.2118144,2.561716,2.911618,2.9968271,3.0820365,3.1672456,3.2524548,3.3376641,3.5697234,3.8017826,4.0356545,4.267714,4.499773,5.844991,7.1902094,8.535428,9.880646,11.225864,13.41411,15.604169,17.794228,19.984287,22.174345,20.73304,19.289923,17.846804,16.405499,14.96238,14.380419,13.796645,13.2146845,12.632723,12.050762,10.7273,9.40565,8.082188,6.7605376,5.4370747,7.0506115,8.662335,10.275872,11.887595,13.499319,11.1968565,8.894395,6.591932,4.2894692,1.987007,2.132044,2.277081,2.422118,2.5671551,2.712192,4.0882306,5.462456,6.836682,8.212721,9.5869465,9.135518,8.682278,8.23085,7.7776093,7.324369,7.231908,7.1394467,7.0469856,6.9545245,6.8620634,9.108324,11.352772,13.597219,15.841667,18.087927,16.79166,15.497204,14.202749,12.908294,11.612025,10.8143215,10.018432,9.220728,8.423024,7.6253204,9.980359,12.335398,14.690435,17.045475,19.400513,16.820667,14.240821,11.6591625,9.079316,6.4994707,6.149569,5.7996674,5.4497657,5.0998635,4.749962,5.009216,5.2702823,5.529536,5.7906027,6.049856,6.825804,7.5999393,8.375887,9.1500225,9.924157,8.178274,6.430578,4.6828823,2.9351864,1.1874905,1.3017071,1.4177368,1.5319533,1.647983,1.7621996,1.4141108,1.067835,0.7197462,0.37165734,0.025381476,3.7147603,7.404139,11.095331,14.78471,18.475903,17.190512,15.905121,14.61973,13.33434,12.050762,9.657652,7.264541,4.8732433,2.4801328,0.0870222,0.7904517,1.4920682,2.1954978,2.8971143,3.6005437,3.8217251,4.0447197,4.267714,4.4907084,4.7118897,4.8206677,4.9276323,5.034597,5.143375,5.2503395,4.5324063,3.8144734,3.0983531,2.38042,1.6624867,2.2571385,2.8517902,3.4482548,4.0429068,4.6375585,4.407312,4.177066,3.9468195,3.7183862,3.48814,3.7582715,4.02659,4.2967215,4.5668526,4.836984,4.1317415,3.4283123,2.72307,2.0178273,1.3125849,1.0497054,0.7868258,0.52575916,0.26287958,0.0,0.27013144,0.5402629,0.8103943,1.0805258,1.3506571,1.0841516,0.8194591,0.55476654,0.29007402,0.025381476,0.10696479,0.19036107,0.27194437,0.35534066,0.43692398,0.64541465,0.8520924,1.0605831,1.2672608,1.4757515,1.5283275,1.5809034,1.6316663,1.6842422,1.7368182,1.5954071,1.452183,1.310772,1.167548,1.0243238,0.8194591,0.61459434,0.40972954,0.20486477,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.07433146,0.072518505,0.07070554,0.06707962,0.065266654,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.0870222,0.11240368,0.13778515,0.16316663,0.18673515,0.38978696,0.59283876,0.79589057,0.99712944,1.2001812,1.4177368,1.6352923,1.8528478,2.0704033,2.2879589,1.9217403,1.5573349,1.1929294,0.82671094,0.46230546,0.9155461,1.3669738,1.8202144,2.2716422,2.7248828,2.9641938,3.2053177,3.444629,3.6857529,3.925064,4.327542,4.7300196,5.132497,5.5349746,5.9374523,7.065115,8.192778,9.32044,10.448103,11.575767,12.070704,12.565643,13.060582,13.555521,14.05046,11.5503845,9.050309,6.550234,4.0501585,1.550083,2.8753586,4.2006345,5.52591,6.849373,8.174648,7.07418,5.975525,4.8750563,3.774588,2.6741197,3.0675328,3.4591327,3.8525455,4.2441454,4.6375585,4.2042603,3.7727752,3.339477,2.907992,2.474694,2.3205922,2.1646774,2.0105755,1.8546607,1.7005589,7.5382986,13.374225,19.211964,25.049704,30.887444,26.05771,21.22798,16.398247,11.566701,6.736969,9.026741,11.318325,13.608097,15.897869,18.187641,14.891675,11.597522,8.301556,5.0074024,1.7132497,17.190512,32.667774,48.145035,63.622295,79.099556,64.57591,50.055897,35.532253,21.010424,6.48678,7.752228,9.017676,10.283124,11.546759,12.812206,10.342952,7.8718834,5.4026284,2.9315605,0.46230546,0.40972954,0.35715362,0.3045777,0.2520018,0.19942589,0.15954071,0.11965553,0.07977036,0.03988518,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.034446288,0.058014803,0.07977036,0.10333887,0.12509441,0.12328146,0.11965553,0.11784257,0.11421664,0.11240368,0.10333887,0.092461094,0.08339628,0.072518505,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.09064813,0.1794833,0.27013144,0.36077955,0.44961473,3.6077955,6.7641635,9.922344,13.080525,16.236893,16.885933,17.533161,18.18039,18.827616,19.474844,21.452785,23.430729,25.406858,27.3848,29.362741,28.157122,26.953314,25.747694,24.542074,23.338266,22.402779,21.46729,20.531801,19.598125,18.662638,17.48965,16.316664,15.14549,13.972503,12.799516,12.547514,12.295512,12.0416975,11.789696,11.537694,12.707055,13.878228,15.047589,16.21695,17.388124,15.792717,14.19731,12.601903,11.008308,9.412902,10.323009,11.233116,12.143224,13.05333,13.961625,13.397794,12.8321495,12.268318,11.702674,11.137029,9.869768,8.602508,7.3352466,6.0679855,4.800725,3.8398547,2.8789847,1.9199274,0.96087015,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.38072214,0.6852999,0.9898776,1.2944553,1.6008459,2.666868,3.7347028,4.802538,5.870373,6.9382076,7.1466985,7.3570023,7.567306,7.7776093,7.987913,8.161958,8.337815,8.511859,8.6877165,8.861761,9.200785,9.537996,9.875207,10.212419,10.549629,10.025683,9.499924,8.974165,8.450218,7.9244595,6.6571984,5.389938,4.122677,2.855416,1.5881553,3.350355,3.484514,3.6204863,3.7546456,3.8906176,4.024777,5.1705694,6.3145485,7.460341,8.604321,9.750113,14.449312,19.150324,23.849524,28.550535,33.249733,30.85481,28.459887,26.064962,23.67004,21.275116,21.487232,21.699348,21.913279,22.125395,22.337511,22.73999,23.142467,23.544945,23.947422,24.349901,26.034143,27.720198,29.40444,31.090496,32.77474,27.080221,21.385706,15.689378,9.994863,4.3003473,4.7372713,5.1741953,5.612932,6.049856,6.48678,6.0444174,5.6020546,5.1596913,4.7173285,4.274966,3.972201,3.6694362,3.3666716,3.0657198,2.762955,3.049403,3.3376641,3.6241121,3.9123733,4.2006345,5.0146546,5.8304877,6.644508,7.460341,8.274362,8.258044,8.239915,8.221786,8.205468,8.187339,7.654328,7.12313,6.590119,6.057108,5.52591,4.95664,4.3891826,3.8217251,3.254268,2.6868105,2.2825198,1.8782293,1.4721256,1.067835,0.66173136,0.54570174,0.42785916,0.3100166,0.19217403,0.07433146,0.092461094,0.11059072,0.12690738,0.14503701,0.16316663,1.4630609,2.762955,4.062849,5.3627434,6.6626377,5.870373,5.0781083,4.2858434,3.491766,2.6995013,2.2516994,1.8057107,1.357909,0.9101072,0.46230546,1.2346275,2.0069497,2.7792716,3.5534067,4.325729,3.7129474,3.100166,2.4873846,1.8746033,1.261822,1.5754645,1.887294,2.1991236,2.5127661,2.8245957,2.9279346,3.0294604,3.1327994,3.2343252,3.3376641,3.2832751,3.2270734,3.1726844,3.1182957,3.0620937,3.2651455,3.4681973,3.6694362,3.872488,4.07554,4.2767787,4.4798307,4.6828823,4.8841214,5.087173,5.825049,6.5629244,7.3008003,8.036863,8.774739,8.6877165,8.600695,8.511859,8.424837,8.337815,8.569874,8.801933,9.035806,9.267865,9.499924,8.930654,8.3595705,7.7903004,7.219217,6.6499467,6.539356,6.430578,6.319988,6.209397,6.1006193,6.0226617,5.9447045,5.866747,5.7906027,5.712645,4.8224807,3.9323158,3.0421512,2.1519866,1.261822,1.7495089,2.2371957,2.7248828,3.2125697,3.7002566,3.6077955,3.5153344,3.4228733,3.3304121,3.2379513,3.4518807,3.6676233,3.8833659,4.0972953,4.313038,5.42801,6.542982,7.6579537,8.772926,9.8878975,12.0416975,14.19731,16.352922,18.506721,20.662334,19.302612,17.94289,16.583168,15.221634,13.861912,13.559147,13.258195,12.955431,12.652666,12.349901,11.329204,10.310318,9.28962,8.270736,7.250037,9.037619,10.825199,12.612781,14.400362,16.187943,13.620788,11.05182,8.484665,5.91751,3.350355,3.3521678,3.3557937,3.3576066,3.3594196,3.3630457,4.699199,6.037165,7.3751316,8.713099,10.049252,9.407463,8.765674,8.122072,7.4802837,6.836682,6.8656893,6.892884,6.9200783,6.947273,6.9744673,9.189907,11.405348,13.620788,15.834415,18.049856,16.635744,15.219821,13.80571,12.389787,10.975676,10.491614,10.009366,9.527119,9.04487,8.562622,10.685601,12.806767,14.929747,17.052727,19.175705,16.87687,14.579845,12.282822,9.985798,7.686961,7.1503243,6.6118746,6.0752378,5.5367875,5.0001507,4.933071,4.8641787,4.797099,4.7300196,4.6629395,5.3246713,5.9882154,6.6499467,7.311678,7.9752226,6.6680765,5.3609304,4.0519714,2.7448254,1.4376793,1.4793775,1.5228885,1.5645868,1.6080978,1.649796,1.3307146,1.0098201,0.69073874,0.36984438,0.05076295,3.5806012,7.1104393,10.640278,14.170115,17.699953,15.966762,14.235382,12.50219,10.770811,9.037619,7.264541,5.4932766,3.720199,1.9471219,0.17585737,0.70524246,1.2346275,1.7658255,2.2952106,2.8245957,3.0820365,3.339477,3.5969179,3.8543584,4.1117992,4.6266804,5.143375,5.658256,6.1731377,6.688019,6.01541,5.3428006,4.670192,3.9975824,3.3249733,3.7401419,4.15531,4.5704784,4.985647,5.4008155,4.940323,4.4798307,4.019338,3.5606585,3.100166,3.2651455,3.4301252,3.5951047,3.7600844,3.925064,3.339477,2.7557032,2.1701162,1.5845293,1.0007553,0.7995165,0.6000906,0.40066472,0.19942589,0.0,0.2030518,0.40429065,0.6073425,0.8103943,1.0116332,0.8194591,0.62728506,0.43511102,0.24293698,0.05076295,0.21574254,0.38072214,0.54570174,0.7106813,0.87566096,1.1784257,1.4793775,1.7821422,2.084907,2.3876717,2.2933977,2.1973107,2.1030366,2.0069497,1.9126755,1.7150626,1.5174497,1.3198367,1.1222239,0.9246109,0.73968875,0.55476654,0.36984438,0.18492219,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.038072214,0.05076295,0.06164073,0.07433146,0.0870222,0.08339628,0.07795739,0.072518505,0.06707962,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.11240368,0.16316663,0.21211663,0.26287958,0.31182957,0.7179332,1.1222239,1.5283275,1.9326181,2.3369088,2.3604772,2.382233,2.4058013,2.427557,2.4493124,2.0830941,1.7150626,1.3470312,0.9808127,0.61278135,1.1802386,1.7476959,2.3151531,2.8826106,3.4500678,3.680314,3.9105604,4.1408067,4.36924,4.599486,4.655688,4.710077,4.764466,4.8206677,4.8750563,5.8431783,6.8094873,7.7776093,8.745731,9.712041,10.6783495,11.642846,12.607342,13.571837,14.538147,11.887595,9.237044,6.588306,3.9377546,1.2872034,2.4257438,3.5624714,4.699199,5.8377395,6.9744673,6.16226,5.3500524,4.537845,3.7256382,2.911618,3.147303,3.3829882,3.6168604,3.8525455,4.0882306,3.7727752,3.4573197,3.141864,2.8282216,2.5127661,2.3024626,2.0921588,1.8818551,1.6733645,1.4630609,8.000604,14.538147,21.07569,27.613234,34.150776,28.452635,22.754494,17.058165,11.3600235,5.661882,9.4546,13.247317,17.040035,20.832752,24.625471,20.134762,15.645867,11.155159,6.6644506,2.175555,13.606284,25.0352,36.46593,47.894844,59.325573,48.52938,37.735004,26.93881,16.144432,5.3500524,6.816739,8.285239,9.751925,11.220426,12.687112,10.259555,7.8319983,5.4044414,2.9768846,0.5493277,0.46955732,0.38978696,0.3100166,0.23024625,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.045324065,0.065266654,0.08520924,0.10515183,0.12509441,0.11965553,0.11421664,0.11059072,0.10515183,0.099712946,0.092461094,0.08520924,0.07795739,0.07070554,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.14322405,0.28463513,0.42785916,0.56927025,0.7124943,4.603112,8.491917,12.382534,16.273151,20.161957,20.395828,20.627888,20.859947,21.092007,21.325878,22.468046,23.610212,24.752378,25.894545,27.03671,25.852846,24.66717,23.483305,22.297626,21.11195,20.966911,20.821875,20.676838,20.531801,20.386765,18.992596,17.598429,16.202446,14.808278,13.412297,13.044266,12.678047,12.310016,11.941984,11.575767,12.989877,14.405801,15.819912,17.234022,18.649946,17.172382,15.694818,14.217253,12.739688,11.262123,11.570327,11.876718,12.184921,12.493125,12.799516,12.206677,11.615651,11.022813,10.429974,9.837135,8.602508,7.36788,6.1332526,4.896812,3.6621845,2.9297476,2.1973107,1.4648738,0.7324369,0.0,0.0,0.0,0.0,0.0,0.0,0.018129626,0.034446288,0.052575916,0.07070554,0.0870222,0.07070554,0.052575916,0.034446288,0.018129626,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.64722764,1.1457924,1.6425442,2.1392958,2.6378605,3.7600844,4.882308,6.004532,7.1267557,8.2507925,8.107569,7.9643445,7.8229337,7.6797094,7.5382986,7.837437,8.138389,8.437528,8.736667,9.037619,9.512614,9.987611,10.462607,10.937603,11.4126,10.937603,10.462607,9.987611,9.512614,9.037619,7.6778965,6.3181744,4.95664,3.5969179,2.2371957,3.2125697,3.39024,3.5679104,3.7455807,3.923251,4.099108,5.2557783,6.4106355,7.5654926,8.72035,9.875207,14.436621,18.999847,23.563074,28.124489,32.687714,30.332678,27.977638,25.6226,23.267561,20.912523,20.887142,20.861761,20.838192,20.81281,20.78743,22.034748,23.282066,24.529385,25.776703,27.025833,27.439188,27.854357,28.269526,28.684694,29.099863,24.045322,18.990784,13.93443,8.87989,3.825351,4.3746786,4.9258194,5.475147,6.0244746,6.5756154,5.866747,5.1596913,4.4526362,3.7455807,3.0367124,2.8282216,2.617918,2.4076142,2.1973107,1.987007,2.5127661,3.0367124,3.5624714,4.0882306,4.612177,5.8848767,7.157576,8.430276,9.702975,10.975676,10.718235,10.460794,10.203354,9.945912,9.686659,9.233418,8.778365,8.323311,7.8682575,7.413204,6.492219,5.573047,4.652062,3.73289,2.811905,2.4166791,2.0232663,1.6280404,1.2328146,0.8375887,0.67986095,0.52213323,0.36440548,0.20667773,0.05076295,0.08339628,0.11421664,0.14684997,0.1794833,0.21211663,1.4249886,2.6378605,3.8507326,5.0617914,6.2746634,5.3808727,4.4852695,3.589666,2.6958754,1.8002719,1.5101979,1.2201238,0.9300498,0.6399758,0.34990177,0.95180535,1.5555218,2.1574254,2.759329,3.3630457,2.8626678,2.3622901,1.8619126,1.3633479,0.8629702,1.1367276,1.4122978,1.6878681,1.9616255,2.2371957,2.5472124,2.857229,3.1672456,3.4772623,3.787279,3.6422417,3.4972048,3.3521678,3.207131,3.0620937,3.159994,3.2578938,3.3557937,3.4518807,3.5497808,3.834416,4.120864,4.405499,4.690134,4.974769,5.5494785,6.1241875,6.70071,7.2754188,7.850128,7.8628187,7.8755093,7.8882003,7.900891,7.911769,7.9298983,7.948028,7.9643445,7.9824743,8.000604,7.507478,7.0143523,6.5230393,6.0299134,5.5367875,5.5476656,5.5567303,5.567608,5.576673,5.5875506,5.5531044,5.516845,5.482399,5.4479527,5.411693,4.603112,3.7927177,2.9823234,2.1719291,1.3633479,1.987007,2.612479,3.2379513,3.8634233,4.4870825,4.216951,3.9468195,3.6766882,3.4083695,3.1382382,3.3358512,3.531651,3.729264,3.926877,4.12449,5.009216,5.8957543,6.78048,7.665206,8.549932,10.669285,12.790451,14.909804,17.029158,19.150324,17.872185,16.59586,15.31772,14.039582,12.763257,12.739688,12.717933,12.694364,12.672608,12.650853,11.9329195,11.214987,10.497053,9.77912,9.063,11.024626,12.988064,14.94969,16.913128,18.874754,16.042906,13.209246,10.377398,7.5455503,4.7118897,4.572292,4.4326935,4.2930956,4.1516843,4.0120864,5.3119802,6.6118746,7.911769,9.211663,10.51337,9.679407,8.847258,8.015107,7.1829576,6.350808,6.497658,6.644508,6.793171,6.9400206,7.0868707,9.273304,11.457924,13.642544,15.827164,18.011784,16.478018,14.942437,13.406858,11.873092,10.337513,10.17072,10.002114,9.835322,9.666717,9.499924,11.390844,13.279951,15.170871,17.059978,18.950897,16.934883,14.920682,12.904668,10.890467,8.874452,8.149267,7.4258947,6.70071,5.975525,5.2503395,4.855114,4.459888,4.064662,3.6694362,3.2742105,3.825351,4.3746786,4.9258194,5.475147,6.0244746,5.1578784,4.2894692,3.4228733,2.5544643,1.6878681,1.6570477,1.6280404,1.5972201,1.5682126,1.5373923,1.2455053,0.95180535,0.65991837,0.3680314,0.07433146,3.444629,6.814926,10.185224,13.555521,16.92582,14.744824,12.565643,10.384649,8.205468,6.0244746,4.8732433,3.720199,2.5671551,1.4141108,0.26287958,0.6200332,0.97718686,1.3343405,1.693307,2.0504606,2.3423476,2.6342347,2.9279346,3.2198215,3.5117085,4.4345064,5.3573046,6.2801023,7.2029004,8.125698,7.4966,6.869315,6.24203,5.614745,4.98746,5.223145,5.4570174,5.6927023,5.9283876,6.16226,5.473334,4.782595,4.0918565,3.4029307,2.712192,2.7720199,2.8318477,2.8916752,2.953316,3.0131438,2.5472124,2.0830941,1.6171626,1.1530442,0.6871128,0.5493277,0.41335547,0.2755703,0.13778515,0.0,0.13415924,0.27013144,0.40429065,0.5402629,0.6744221,0.55476654,0.43511102,0.3154555,0.19579996,0.07433146,0.32270733,0.56927025,0.81764615,1.064209,1.3125849,1.7096237,2.1066625,2.5055144,2.902553,3.299592,3.056655,2.8155308,2.572594,2.3296568,2.08672,1.8347181,1.5827163,1.3307146,1.0768998,0.824898,0.65991837,0.4949388,0.32995918,0.16497959,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.05076295,0.06164073,0.07433146,0.0870222,0.099712946,0.092461094,0.08520924,0.07795739,0.07070554,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.13778515,0.21211663,0.28826106,0.36259252,0.43692398,1.0442665,1.651609,2.2607644,2.8681068,3.4754493,3.303218,3.1291735,2.956942,2.7847104,2.612479,2.2426348,1.8727903,1.502946,1.1331016,0.76325727,1.4449311,2.126605,2.810092,3.491766,4.175253,4.3946214,4.615803,4.835171,5.0545397,5.275721,4.9820213,4.690134,4.3982472,4.1045475,3.8126602,4.6194286,5.42801,6.2347784,7.0433598,7.850128,9.284182,10.720048,12.155914,13.589968,15.025834,12.224807,9.425592,6.624565,3.825351,1.0243238,1.9743162,2.9243085,3.874301,4.8242936,5.774286,5.2503395,4.7245803,4.2006345,3.6748753,3.149116,3.2270734,3.3050308,3.3829882,3.4591327,3.53709,3.339477,3.141864,2.9442513,2.7466383,2.5508385,2.2843328,2.0196402,1.7549478,1.4902552,1.2255627,8.46291,15.700256,22.937603,30.17495,37.412296,30.847559,24.282822,17.718082,11.151533,4.5867953,9.882459,15.1781225,20.471973,25.767637,31.063301,25.37785,19.6924,14.006948,8.323311,2.6378605,10.020245,17.402628,24.785011,32.167397,39.549778,32.481037,25.415922,18.347181,11.280253,4.213325,5.883064,7.552802,9.222541,10.89228,12.562017,10.177972,7.7921133,5.408067,3.0222087,0.63816285,0.5293851,0.4224203,0.3154555,0.20667773,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.054388877,0.072518505,0.09064813,0.10696479,0.12509441,0.11784257,0.11059072,0.10333887,0.09427405,0.0870222,0.08339628,0.07795739,0.072518505,0.06707962,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.19579996,0.38978696,0.5855869,0.7795739,0.97537386,5.5984282,10.21967,14.842725,19.463966,24.08702,23.905725,23.722616,23.539507,23.35821,23.1751,23.483305,23.789696,24.097898,24.40429,24.712494,23.546759,22.382835,21.217102,20.053179,18.887444,19.53286,20.178274,20.821875,21.46729,22.112705,20.495543,18.87838,17.259403,15.6422415,14.025079,13.54283,13.060582,12.578335,12.094274,11.612025,13.272699,14.93156,16.592234,18.252907,19.911768,18.552046,17.192324,15.8326025,14.47288,13.113158,12.817645,12.522133,12.22662,11.9329195,11.637406,11.017374,10.397341,9.7773075,9.157274,8.537241,7.3352466,6.1332526,4.9294453,3.727451,2.525457,2.0196402,1.5156367,1.0098201,0.5058166,0.0,0.0,0.0,0.0,0.0,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.045324065,0.09064813,0.13415924,0.1794833,0.22480737,0.9155461,1.6044719,2.2952106,2.9841363,3.6748753,4.853301,6.0299134,7.208339,8.384952,9.563377,9.066626,8.571687,8.076748,7.5818095,7.0868707,7.512917,7.93715,8.363196,8.78743,9.211663,9.824444,10.437225,11.050007,11.662788,12.27557,11.849524,11.42529,10.999244,10.57501,10.150778,8.696781,7.2445984,5.7924156,4.3402324,2.8880494,3.0747845,3.294153,3.5153344,3.7347028,3.9558845,4.175253,5.3391747,6.5049095,7.6706448,8.834567,10.000301,14.425743,18.849373,23.274813,27.700254,32.125698,29.810543,27.49539,25.180237,22.865084,20.54993,20.287052,20.024172,19.763105,19.500225,19.237347,21.329504,23.421663,25.515635,27.607794,29.699953,28.844234,27.99033,27.134611,26.280706,25.424988,21.010424,16.59586,12.179482,7.764919,3.350355,4.0120864,4.6756306,5.337362,6.000906,6.6626377,5.6908894,4.7173285,3.7455807,2.7720199,1.8002719,1.6824293,1.5645868,1.4467441,1.3307146,1.2128719,1.9743162,2.7375734,3.5008307,4.262275,5.0255322,6.755099,8.484665,10.2142315,11.94561,13.675177,13.176612,12.67986,12.183108,11.684544,11.187792,10.810696,10.431787,10.05469,9.677594,9.300498,8.027799,6.755099,5.482399,4.209699,2.9369993,2.5526514,2.1683033,1.7821422,1.3977941,1.0116332,0.81583315,0.61822027,0.42060733,0.2229944,0.025381476,0.072518505,0.11965553,0.16679256,0.21574254,0.26287958,1.3869164,2.5127661,3.636803,4.762653,5.8866897,4.88956,3.8924308,2.8953013,1.8981718,0.89922947,0.7668832,0.6345369,0.50219065,0.36984438,0.2374981,0.67079616,1.1022812,1.5355793,1.9670644,2.4003625,2.0123885,1.6244144,1.2382535,0.85027945,0.46230546,0.69980353,0.93730164,1.1747998,1.4122978,1.649796,2.1683033,2.6849976,3.2016919,3.720199,4.2368937,4.0030212,3.7673361,3.531651,3.2977788,3.0620937,3.054842,3.04759,3.0403383,3.0330863,3.0258346,3.392053,3.7600844,4.1281157,4.494334,4.8623657,5.275721,5.6872635,6.1006193,6.5121617,6.925517,7.037921,7.1503243,7.262728,7.3751316,7.4875355,7.2899227,7.0923095,6.8946967,6.697084,6.4994707,6.0843024,5.669134,5.2557783,4.84061,4.4254417,4.554162,4.6846952,4.8152285,4.945762,5.0744824,5.081734,5.090799,5.0980506,5.105303,5.1125546,4.3819304,3.6531196,2.9224956,2.1918716,1.4630609,2.2245052,2.9877625,3.7492065,4.512464,5.275721,4.8279195,4.3801174,3.9323158,3.484514,3.0367124,3.2180085,3.397492,3.576975,3.7582715,3.9377546,4.592234,5.2467136,5.903006,6.5574856,7.211965,9.296872,11.381779,13.466686,15.553406,17.638313,16.441757,15.247015,14.052273,12.857531,11.662788,11.920229,12.17767,12.43511,12.692551,12.949992,12.534823,12.119655,11.704487,11.289318,10.874149,13.011633,15.149116,17.288412,19.425894,21.563377,18.465023,15.368484,12.270131,9.171778,6.0752378,5.7924156,5.5095935,5.2267714,4.945762,4.6629395,5.924762,7.1865835,8.450218,9.712041,10.975676,9.953164,8.930654,7.9081426,6.885632,5.863121,6.1296263,6.397945,6.6644506,6.932769,7.1992745,9.354887,11.510499,13.664299,15.819912,17.975525,16.32029,14.665054,13.009819,11.354585,9.699349,9.848013,9.994863,10.141713,10.290376,10.437225,12.094274,13.753134,15.410182,17.06723,18.724277,16.992899,15.2597065,13.528327,11.795135,10.061942,9.1500225,8.238102,7.324369,6.412449,5.5005283,4.7771564,4.0555973,3.3322253,2.610666,1.887294,2.324218,2.762955,3.199879,3.636803,4.07554,3.6476808,3.2198215,2.7919624,2.3641033,1.938057,1.8347181,1.7331922,1.6298534,1.5283275,1.4249886,1.1602961,0.89560354,0.629098,0.36440548,0.099712946,3.3104696,6.5194135,9.73017,12.940927,16.14987,13.522888,10.8959055,8.267109,5.6401267,3.0131438,2.4801328,1.9471219,1.4141108,0.88291276,0.34990177,0.53482395,0.7197462,0.90466833,1.0895905,1.2745126,1.6026589,1.9308052,2.2571385,2.5852847,2.911618,4.2423325,5.573047,6.9019485,8.232663,9.563377,8.979604,8.397643,7.8156815,7.231908,6.6499467,6.7043357,6.7605376,6.814926,6.869315,6.925517,6.004532,5.08536,4.164375,3.245203,2.324218,2.280707,2.2353828,2.1900587,2.1447346,2.0994108,1.7549478,1.4104849,1.064209,0.7197462,0.37528324,0.2991388,0.22480737,0.15047589,0.07433146,0.0,0.06707962,0.13415924,0.2030518,0.27013144,0.33721104,0.29007402,0.24293698,0.19579996,0.14684997,0.099712946,0.42967212,0.75963134,1.0895905,1.4195497,1.7495089,2.2426348,2.7357605,3.2270734,3.720199,4.213325,3.8217251,3.4319382,3.0421512,2.6523643,2.2625773,1.9543737,1.647983,1.3397794,1.0333886,0.72518504,0.58014804,0.43511102,0.29007402,0.14503701,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.10333887,0.092461094,0.08339628,0.072518505,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.16316663,0.26287958,0.36259252,0.46230546,0.5620184,1.3724127,2.182807,2.9932013,3.8017826,4.612177,4.2441454,3.877927,3.5098956,3.141864,2.7756457,2.4021754,2.030518,1.6570477,1.2853905,0.9119202,1.7096237,2.5073273,3.3050308,4.102734,4.900438,5.1107416,5.319232,5.529536,5.7398396,5.9501433,5.3101673,4.670192,4.0302157,3.39024,2.7502642,3.397492,4.0447197,4.691947,5.3391747,5.9882154,7.891826,9.79725,11.702674,13.608097,15.511708,12.562017,9.612328,6.6626377,3.7129474,0.76325727,1.5247015,2.2879589,3.049403,3.8126602,4.574105,4.3366065,4.099108,3.8616104,3.6241121,3.386614,3.3068438,3.2270734,3.147303,3.0675328,2.9877625,2.907992,2.8282216,2.7466383,2.666868,2.5870976,2.268016,1.9471219,1.6280404,1.3071461,0.9880646,8.925215,16.862366,24.799515,32.73848,40.67563,33.24248,25.809336,18.378002,10.944855,3.5117085,10.310318,17.107115,23.905725,30.702522,37.499317,30.619125,23.740746,16.860552,9.980359,3.100166,6.436017,9.770056,13.1059065,16.439945,19.775795,16.434505,13.095029,9.755551,6.414262,3.0747845,4.947575,6.8203654,8.693155,10.564133,12.436923,10.094576,7.752228,5.40988,3.0675328,0.72518504,0.58921283,0.4550536,0.3208944,0.18492219,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.065266654,0.07977036,0.09427405,0.11059072,0.12509441,0.11421664,0.10515183,0.09427405,0.08520924,0.07433146,0.072518505,0.07070554,0.06707962,0.065266654,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.24837588,0.4949388,0.7433147,0.9898776,1.2382535,6.591932,11.947423,17.302916,22.656593,28.012085,27.41562,26.817343,26.220879,25.6226,25.024323,24.49675,23.96918,23.441607,22.915848,22.388275,21.242483,20.096691,18.952711,17.80692,16.66294,18.096992,19.53286,20.966911,22.402779,23.836832,21.996675,20.15833,18.318174,16.478018,14.63786,14.039582,13.443117,12.84484,12.248375,11.650098,13.555521,15.459132,17.364555,19.26998,21.175404,19.931711,18.68983,17.447952,16.20426,14.96238,14.064963,13.167547,12.270131,11.372714,10.475298,9.82807,9.180842,8.531802,7.8845744,7.2373466,6.0679855,4.896812,3.727451,2.5580902,1.3869164,1.1095331,0.8321498,0.55476654,0.27738327,0.0,0.0,0.0,0.0,0.0,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.09064813,0.06707962,0.045324065,0.02175555,0.0,0.059827764,0.11965553,0.1794833,0.23931105,0.2991388,1.1820517,2.0649643,2.9478772,3.83079,4.7118897,5.9447045,7.177519,8.410334,9.643148,10.874149,10.027496,9.179029,8.3323765,7.4857225,6.637256,7.1883965,7.7377243,8.287052,8.838193,9.38752,10.138086,10.88684,11.637406,12.387974,13.136727,12.763257,12.387974,12.012691,11.637406,11.262123,9.71748,8.172835,6.628191,5.081734,3.53709,2.9369993,3.199879,3.4627585,3.7256382,3.9867048,4.249584,5.424384,6.599184,7.7757964,8.950596,10.125396,14.413053,18.700708,22.988365,27.27421,31.561865,29.28841,27.013142,24.737875,22.462606,20.187338,19.68696,19.188396,18.688019,18.187641,17.687263,20.624262,23.563074,26.500074,29.437073,32.375885,30.24928,28.124489,25.999697,23.874905,21.750113,17.975525,14.200936,10.424535,6.6499467,2.8753586,3.6494937,4.4254417,5.199577,5.975525,6.7496595,5.5132194,4.274966,3.0367124,1.8002719,0.5620184,0.53663695,0.51306844,0.48768693,0.46230546,0.43692398,1.4376793,2.4366217,3.437377,4.4381323,5.4370747,7.6253204,9.811753,11.999999,14.188245,16.374678,15.636803,14.90074,14.162864,13.424988,12.687112,12.387974,12.087022,11.787883,11.486931,11.187792,9.563377,7.93715,6.3127356,4.688321,3.0620937,2.6868105,2.3133402,1.938057,1.5627737,1.1874905,0.9499924,0.7124943,0.4749962,0.2374981,0.0,0.06164073,0.12509441,0.18673515,0.25018883,0.31182957,1.3506571,2.3876717,3.4246864,4.461701,5.5005283,4.40006,3.299592,2.1991236,1.1004683,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.387974,0.6508536,0.9119202,1.1747998,1.4376793,1.162109,0.8883517,0.61278135,0.33721104,0.06164073,0.26287958,0.46230546,0.66173136,0.8629702,1.062396,1.7875811,2.5127661,3.2379513,3.9631362,4.688321,4.361988,4.0374675,3.7129474,3.386614,3.0620937,2.94969,2.8372865,2.7248828,2.612479,2.5000753,2.94969,3.3993049,3.8507326,4.3003473,4.749962,5.0001507,5.2503395,5.5005283,5.750717,6.000906,6.2130227,6.4251394,6.637256,6.849373,7.063302,6.6499467,6.2384043,5.825049,5.411693,5.0001507,4.6629395,4.325729,3.9867048,3.6494937,3.3122826,3.5624714,3.8126602,4.062849,4.313038,4.5632267,4.612177,4.6629395,4.7118897,4.762653,4.8116026,4.162562,3.5117085,2.8626678,2.2118144,1.5627737,2.4620032,3.3630457,4.262275,5.163317,6.0625467,5.4370747,4.8134155,4.1879435,3.5624714,2.9369993,3.100166,3.2633326,3.4246864,3.587853,3.7492065,4.175253,4.599486,5.0255322,5.4497657,5.8758116,7.9244595,9.97492,12.025381,14.075842,16.124489,15.013144,13.899984,12.786825,11.675479,10.56232,11.10077,11.637406,12.175857,12.712494,13.24913,13.136727,13.024323,12.91192,12.799516,12.687112,15.000452,17.31198,19.62532,21.936848,24.250187,20.887142,17.52591,14.162864,10.799818,7.4367723,7.0125394,6.588306,6.16226,5.7380266,5.3119802,6.5375433,7.763106,8.9868555,10.212419,11.437981,10.225109,9.012237,7.799365,6.588306,5.375434,5.7615952,6.149569,6.5375433,6.925517,7.311678,9.438283,11.563075,13.687867,15.812659,17.937452,16.162561,14.387671,12.612781,10.837891,9.063,9.525306,9.987611,10.449916,10.912222,11.374527,12.799516,14.224504,15.649493,17.074482,18.49947,17.050913,15.600543,14.150173,12.699803,11.249433,10.150778,9.050309,7.949841,6.849373,5.750717,4.699199,3.6494937,2.5997884,1.550083,0.50037766,0.824898,1.1494182,1.4757515,1.8002719,2.124792,2.137483,2.1501737,2.1628644,2.175555,2.1882458,2.0123885,1.8383441,1.6624867,1.4866294,1.3125849,1.0750868,0.8375887,0.6000906,0.36259252,0.12509441,3.1744974,6.2257137,9.275117,12.32452,15.375735,12.300951,9.224354,6.149569,3.0747845,0.0,0.0870222,0.17585737,0.26287958,0.34990177,0.43692398,0.44961473,0.46230546,0.4749962,0.48768693,0.50037766,0.8629702,1.2255627,1.5881553,1.9507477,2.3133402,4.0501585,5.7869763,7.5256076,9.262425,10.999244,10.462607,9.924157,9.38752,8.8508835,8.312433,8.187339,8.062244,7.93715,7.8120556,7.686961,6.5375433,5.388125,4.2368937,3.0874753,1.938057,1.7875811,1.6371052,1.4866294,1.3379664,1.1874905,0.96268314,0.73787576,0.51306844,0.28826106,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.53663695,0.9499924,1.3633479,1.7748904,2.1882458,2.7756457,3.3630457,3.9504454,4.537845,5.125245,4.5867953,4.0501585,3.5117085,2.9750717,2.4366217,2.0758421,1.7132497,1.3506571,0.9880646,0.62547207,0.50037766,0.37528324,0.25018883,0.12509441,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.18673515,0.31182957,0.43692398,0.5620184,0.6871128,1.7005589,2.712192,3.7256382,4.7372713,5.750717,5.186886,4.6248674,4.062849,3.5008307,2.9369993,2.561716,2.1882458,1.8129625,1.4376793,1.062396,1.9743162,2.8880494,3.7999697,4.7118897,5.6256227,5.825049,6.0244746,6.2257137,6.4251394,6.624565,5.638314,4.650249,3.6621845,2.6741197,1.6878681,2.175555,2.663242,3.149116,3.636803,4.12449,6.4994707,8.874452,11.249433,13.6244135,15.999394,12.899229,9.800876,6.70071,3.6005437,0.50037766,1.0750868,1.649796,2.2245052,2.7992141,3.3757362,3.4246864,3.4754493,3.5243993,3.5751622,3.6241121,3.386614,3.149116,2.911618,2.6741197,2.4366217,2.474694,2.5127661,2.5508385,2.5870976,2.6251698,2.2498865,1.8746033,1.49932,1.1258497,0.7505665,9.38752,18.024473,26.66324,35.300194,43.93715,35.637405,27.337664,19.03792,10.738177,2.4366217,10.738177,19.03792,27.337664,35.637405,43.93715,35.862213,27.787277,19.712341,11.637406,3.5624714,2.8499773,2.137483,1.4249886,0.7124943,0.0,0.387974,0.774135,1.162109,1.550083,1.938057,4.0120864,6.0879283,8.161958,10.2378,12.311829,10.012992,7.7123427,5.411693,3.1128569,0.8122072,0.6508536,0.48768693,0.3245203,0.16316663,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.2991388,0.6000906,0.89922947,1.2001812,1.49932,7.5872483,13.675177,19.763105,25.84922,31.93715,30.925516,29.91207,28.900436,27.88699,26.875357,25.512009,24.150475,22.787127,21.425592,20.062244,18.938208,17.812357,16.68832,15.56247,14.436621,16.66294,18.887444,21.11195,23.338266,25.562773,23.49962,21.438282,19.375132,17.31198,15.250641,14.538147,13.825653,13.113158,12.400664,11.6881695,13.838344,15.986704,18.136877,20.287052,22.437225,21.313189,20.187338,19.063301,17.937452,16.811602,15.312282,13.812962,12.311829,10.812509,9.313189,8.636953,7.9625316,7.28811,6.6118746,5.9374523,4.800725,3.6621845,2.525457,1.3869164,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.07433146,0.15047589,0.22480737,0.2991388,0.37528324,1.4503701,2.525457,3.6005437,4.6756306,5.750717,7.037921,8.325124,9.612328,10.899531,12.186734,10.986553,9.788185,8.588004,7.3878226,6.187641,6.8620634,7.5382986,8.212721,8.887142,9.563377,10.449916,11.338268,12.224807,13.113158,13.999697,13.675177,13.3506565,13.024323,12.699803,12.375282,10.738177,9.099259,7.462154,5.825049,4.1879435,2.7883365,3.0276475,3.2669585,3.5080826,3.7473936,3.9867048,4.9276323,5.866747,6.8076744,7.746789,8.6877165,13.232814,17.77791,22.323008,26.868105,31.413202,29.302914,27.192625,25.082336,22.97205,20.861761,20.676838,20.491917,20.306993,20.122072,19.93715,22.727299,25.517448,28.307598,31.097748,33.887897,31.09956,28.313036,25.5247,22.738176,19.94984,16.51065,13.069647,9.630457,6.189454,2.7502642,3.4953918,4.2405195,4.985647,5.730775,6.4759026,5.331923,4.1897564,3.04759,1.9054236,0.76325727,1.0007553,1.2382535,1.4757515,1.7132497,1.9507477,2.8771715,3.8054085,4.7318325,5.660069,6.588306,7.949841,9.313189,10.674724,12.038072,13.399607,13.049705,12.699803,12.349901,11.999999,11.650098,11.292944,10.93579,10.576823,10.21967,9.862516,8.508233,7.1521373,5.7978544,4.441758,3.0874753,2.659616,2.231757,1.8057107,1.3778516,0.9499924,0.75963134,0.56927025,0.38072214,0.19036107,0.0,0.08339628,0.16497959,0.24837588,0.32995918,0.41335547,1.2853905,2.1574254,3.0294604,3.9033084,4.7753434,4.1879435,3.6005437,3.0131438,2.4257438,1.8383441,2.1628644,2.4873846,2.811905,3.1382382,3.4627585,3.1853752,2.907992,2.6306088,2.3532255,2.0758421,1.6697385,1.2654479,0.85934424,0.4550536,0.05076295,0.21030366,0.36984438,0.5293851,0.69073874,0.85027945,1.4304274,2.0105755,2.5907235,3.1708715,3.7492065,3.7347028,3.720199,3.7056956,3.6893787,3.6748753,3.5824142,3.489953,3.397492,3.3050308,3.2125697,3.5515938,3.8924308,4.233268,4.572292,4.9131284,5.185073,5.4570174,5.730775,6.002719,6.2746634,6.347182,6.4197006,6.492219,6.5647373,6.637256,6.2220874,5.806919,5.391751,4.9783955,4.5632267,4.441758,4.322103,4.2024474,4.082792,3.9631362,4.004834,4.0483456,4.0900435,4.1317415,4.175253,4.25321,4.329355,4.407312,4.4852695,4.5632267,3.9504454,3.3376641,2.7248828,2.1121013,1.49932,2.275268,3.049403,3.825351,4.599486,5.375434,4.8732433,4.36924,3.8670492,3.3648586,2.8626678,3.005892,3.147303,3.290527,3.4319382,3.5751622,3.919625,4.264088,4.610364,4.954827,5.2992897,7.2373466,9.175404,11.113461,13.049705,14.9877615,13.974316,12.962683,11.949236,10.937603,9.924157,10.257742,10.589515,10.9230995,11.254871,11.586644,12.230246,12.872034,13.515636,14.157425,14.799213,16.358362,17.915697,19.473032,21.030367,22.5877,19.565493,16.543283,13.519262,10.497053,7.474845,7.137634,6.8004227,6.4632115,6.1241875,5.7869763,6.965402,8.1420145,9.32044,10.497053,11.675479,10.5695715,9.465478,8.3595705,7.2554765,6.149569,6.7677894,7.3841968,8.002417,8.620637,9.237044,11.095331,12.951805,14.810091,16.668379,18.52485,16.472578,14.420304,12.368031,10.315757,8.26167,8.696781,9.131892,9.567003,10.002114,10.437225,11.889409,13.341592,14.795588,16.24777,17.699953,16.104548,14.50914,12.915545,11.320138,9.724731,8.999546,8.274362,7.549176,6.825804,6.1006193,5.4570174,4.8152285,4.171627,3.529838,2.8880494,2.7847104,2.6831846,2.5798457,2.47832,2.374981,2.4166791,2.4601903,2.5018883,2.5453994,2.5870976,2.3042755,2.0232663,1.7404441,1.4576219,1.1747998,0.9880646,0.7995165,0.61278135,0.42423326,0.2374981,2.8517902,5.467895,8.082188,10.698292,13.312584,10.6783495,8.042302,5.408067,2.7720199,0.13778515,0.18310922,0.22662032,0.27194437,0.31726846,0.36259252,0.52575916,0.6871128,0.85027945,1.0116332,1.1747998,1.3832904,1.5899682,1.7966459,2.0051367,2.2118144,3.529838,4.847862,6.165886,7.4820967,8.80012,8.450218,8.100317,7.750415,7.400513,7.0506115,6.925517,6.8004227,6.6753283,6.550234,6.4251394,5.560356,4.695573,3.83079,2.9641938,2.0994108,1.8691645,1.6407311,1.4104849,1.1802386,0.9499924,0.7777609,0.6055295,0.43329805,0.25925365,0.0870222,0.07070554,0.052575916,0.034446288,0.018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.09789998,0.19579996,0.291887,0.38978696,0.48768693,0.8321498,1.1766127,1.5228885,1.8673514,2.2118144,2.8499773,3.48814,4.12449,4.762653,5.4008155,4.8279195,4.255023,3.682127,3.1092308,2.5381477,2.1574254,1.7767034,1.3977941,1.017072,0.63816285,0.51306844,0.387974,0.26287958,0.13778515,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.07433146,0.08520924,0.09427405,0.10515183,0.11421664,0.12509441,0.11421664,0.10515183,0.09427405,0.08520924,0.07433146,0.072518505,0.07070554,0.06707962,0.065266654,0.06164073,0.16316663,0.26287958,0.36259252,0.46230546,0.5620184,1.452183,2.3423476,3.2325122,4.122677,5.0128417,4.4816437,3.9522583,3.4228733,2.8916752,2.3622901,2.0631514,1.7621996,1.4630609,1.162109,0.8629702,1.5917811,2.322405,3.053029,3.7818398,4.512464,4.9076896,5.3029156,5.6981416,6.093367,6.48678,6.0824895,5.678199,5.272095,4.8678045,4.461701,4.358362,4.25321,4.1480584,4.0429068,3.9377546,6.053482,8.167397,10.283124,12.397038,14.512766,11.704487,8.898021,6.089741,3.2832751,0.4749962,1.0768998,1.6806163,2.2825198,2.8844235,3.48814,3.6948178,3.9033084,4.1099863,4.3166637,4.5251546,4.267714,4.0102735,3.7528327,3.4953918,3.2379513,3.2796493,3.3231604,3.3648586,3.4083695,3.4500678,2.9877625,2.525457,2.0631514,1.6008459,1.1367276,9.246109,17.351866,25.459433,33.567,41.674572,33.85889,26.045021,18.22934,10.41547,2.5997884,10.315757,18.029913,25.745882,33.460037,41.174194,33.52893,25.885479,18.240217,10.594954,2.94969,5.2449007,7.5401115,9.835322,12.130532,14.425743,11.98187,9.539809,7.0977483,4.655688,2.2118144,3.9975824,5.7833505,7.567306,9.353074,11.137029,9.063,6.987158,4.9131284,2.8372865,0.76325727,0.6091554,0.45686656,0.3045777,0.15228885,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.13778515,0.13053331,0.12328146,0.11421664,0.10696479,0.099712946,0.09427405,0.09064813,0.08520924,0.07977036,0.07433146,0.072518505,0.07070554,0.06707962,0.065266654,0.06164073,0.059827764,0.058014803,0.054388877,0.052575916,0.05076295,0.6544795,1.260009,1.8655385,2.469255,3.0747845,8.528176,13.979754,19.433146,24.884724,30.338116,29.081734,27.827162,26.572592,25.318022,24.06164,22.584074,21.108324,19.630758,18.153194,16.67563,16.095482,15.515334,14.935185,14.355038,13.77489,16.140806,18.50491,20.870825,23.234928,25.600845,24.487686,23.374527,22.26318,21.15002,20.036863,19.204712,18.372562,17.540413,16.708263,15.8743,17.567608,19.259102,20.952408,22.645716,24.33721,22.810696,21.282368,19.755854,18.227526,16.699198,15.3956785,14.090345,12.785012,11.479679,10.174346,9.460039,8.745731,8.029612,7.315304,6.599184,5.335549,4.070101,2.8046532,1.5392052,0.2755703,0.21936847,0.16497959,0.11059072,0.054388877,0.0,0.0,0.0,0.0,0.0,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.09427405,0.07795739,0.059827764,0.04169814,0.025381476,0.30276474,0.58014804,0.8575313,1.1349145,1.4122978,2.333283,3.2524548,4.171627,5.092612,6.011784,7.1031876,8.192778,9.282369,10.371959,11.463363,10.700105,9.936848,9.175404,8.412147,7.650702,8.885329,10.119957,11.354585,12.589212,13.825653,15.147303,16.470764,17.792416,19.114065,20.437527,18.465023,16.492521,14.520018,12.547514,10.57501,9.282369,7.989726,6.697084,5.4044414,4.1117992,2.6378605,2.855416,3.0729716,3.290527,3.5080826,3.7256382,4.4308805,5.1343102,5.8395524,6.544795,7.250037,12.052575,16.855114,21.657652,26.46019,31.262726,29.317417,27.372108,25.4268,23.483305,21.537996,21.666716,21.797249,21.927782,22.058315,22.187037,24.830336,27.471823,30.115122,32.75842,35.399906,31.949839,28.499771,25.049704,21.599636,18.149569,15.045776,11.940171,8.834567,5.730775,2.6251698,3.339477,4.0555973,4.7699046,5.484212,6.200332,5.1524396,4.1045475,3.056655,2.0105755,0.96268314,1.4630609,1.9616255,2.4620032,2.962381,3.4627585,4.3166637,5.1723824,6.0281005,6.882006,7.7377243,8.274362,8.812811,9.349448,9.8878975,10.424535,10.462607,10.500679,10.536939,10.57501,10.613083,10.197914,9.782746,9.367578,8.952409,8.537241,7.453089,6.3671246,5.282973,4.1970086,3.1128569,2.6324217,2.1519866,1.6733645,1.1929294,0.7124943,0.56927025,0.42785916,0.28463513,0.14322405,0.0,0.10333887,0.20486477,0.30820364,0.40972954,0.51306844,1.2201238,1.9271792,2.6342347,3.343103,4.0501585,3.975827,3.8996825,3.825351,3.7492065,3.6748753,4.3003473,4.9258194,5.5494785,6.1749506,6.8004227,5.9827766,5.1651306,4.347484,3.529838,2.712192,2.1773682,1.6425442,1.1077201,0.5728962,0.038072214,0.15772775,0.27738327,0.39703882,0.5166943,0.63816285,1.0732739,1.5083848,1.9416829,2.3767939,2.811905,3.1074178,3.4029307,3.6966307,3.9921436,4.2876563,4.215138,4.1426196,4.070101,3.9975824,3.925064,4.15531,4.3855567,4.615803,4.844236,5.0744824,5.369995,5.6655083,5.959208,6.2547207,6.550234,6.4831543,6.414262,6.347182,6.2801023,6.2130227,5.7942286,5.377247,4.9602656,4.5432844,4.12449,4.2223897,4.3202896,4.41819,4.514277,4.612177,4.4471974,4.2822175,4.117238,3.9522583,3.787279,3.8924308,3.9975824,4.102734,4.207886,4.313038,3.738329,3.1618068,2.5870976,2.0123885,1.4376793,2.08672,2.7375734,3.386614,4.0374675,4.688321,4.307599,3.926877,3.5479677,3.1672456,2.7883365,2.909805,3.0330863,3.1545548,3.2778363,3.3993049,3.6658103,3.930503,4.195195,4.459888,4.7245803,6.550234,8.374074,10.199727,12.025381,13.849221,12.937301,12.025381,11.111648,10.199727,9.287807,9.414715,9.541622,9.670342,9.79725,9.924157,11.321951,12.719746,14.117539,15.515334,16.913128,17.714457,18.5176,19.320742,20.122072,20.925215,18.24203,15.5606575,12.877473,10.194288,7.512917,7.262728,7.0125394,6.7623506,6.5121617,6.261973,7.3932614,8.5227375,9.652213,10.781689,11.912977,10.915848,9.916905,8.919776,7.9226465,6.925517,7.7721705,8.620637,9.467291,10.315757,11.162411,12.752378,14.342347,15.932315,17.522284,19.112251,16.782595,14.452938,12.123281,9.791811,7.462154,7.8700705,8.2779875,8.685904,9.092008,9.499924,10.979301,12.460492,13.939869,15.419247,16.900436,15.159993,13.419549,11.679105,9.940474,8.200029,7.850128,7.500226,7.1503243,6.8004227,6.450521,6.2148356,5.979151,5.7452784,5.5095935,5.275721,4.744523,4.215138,3.6857529,3.1545548,2.6251698,2.6976883,2.770207,2.8427253,2.9152439,2.9877625,2.5979755,2.2081885,1.8165885,1.4268016,1.0370146,0.89922947,0.76325727,0.62547207,0.48768693,0.34990177,2.5290828,4.710077,6.889258,9.070251,11.249433,9.055748,6.8602505,4.664753,2.469255,0.2755703,0.27738327,0.27919623,0.28282216,0.28463513,0.28826106,0.6000906,0.9119202,1.2255627,1.5373923,1.8492218,1.9017978,1.9543737,2.0069497,2.0595255,2.1121013,3.009518,3.9069343,4.804351,5.7017674,6.599184,6.43783,6.2746634,6.11331,5.9501433,5.7869763,5.661882,5.5367875,5.411693,5.2865987,5.163317,4.5831695,4.0030212,3.4228733,2.8427253,2.2625773,1.9525607,1.6425442,1.3325275,1.0225109,0.7124943,0.59283876,0.47318324,0.35171473,0.23205921,0.11240368,0.09064813,0.06707962,0.045324065,0.02175555,0.0,0.0,0.0,0.0,0.0,0.0,0.17041849,0.34083697,0.5094425,0.67986095,0.85027945,1.1276628,1.405046,1.6824293,1.9598125,2.2371957,2.9243085,3.6132345,4.3003473,4.98746,5.674573,5.06723,4.459888,3.8525455,3.245203,2.6378605,2.2408218,1.84197,1.4449311,1.0478923,0.6508536,0.52575916,0.40066472,0.2755703,0.15047589,0.025381476,0.038072214,0.05076295,0.06164073,0.07433146,0.0870222,0.09427405,0.10333887,0.11059072,0.11784257,0.12509441,0.11784257,0.11059072,0.10333887,0.09427405,0.0870222,0.08339628,0.07795739,0.072518505,0.06707962,0.06164073,0.13778515,0.21211663,0.28826106,0.36259252,0.43692398,1.2056202,1.9725033,2.7393866,3.5080826,4.274966,3.778214,3.2796493,2.7828975,2.2843328,1.7875811,1.5627737,1.3379664,1.1131591,0.8883517,0.66173136,1.209246,1.7567607,2.3042755,2.8517902,3.3993049,3.9903307,4.5795436,5.1705694,5.7597823,6.350808,6.526665,6.7043357,6.882006,7.059676,7.2373466,6.539356,5.8431783,5.145188,4.4471974,3.7492065,5.6056805,7.460341,9.3150015,11.169662,13.024323,10.509744,7.995165,5.480586,2.9641938,0.44961473,1.0805258,1.7096237,2.3405347,2.9696326,3.6005437,3.9649491,4.329355,4.695573,5.0599785,5.424384,5.147001,4.8696175,4.592234,4.314851,4.0374675,4.0846047,4.1317415,4.1806917,4.227829,4.274966,3.7256382,3.1744974,2.6251698,2.0758421,1.5247015,9.102885,16.679256,24.257439,31.835623,39.411995,32.082188,24.752378,17.422571,10.092763,2.762955,9.893337,17.021906,24.152288,31.28267,38.41305,31.19746,23.981869,16.768091,9.5525,2.3369088,7.6398244,12.9427395,18.245655,23.54857,28.849674,23.577578,18.305483,13.031575,7.75948,2.4873846,3.9830787,5.47696,6.972654,8.4683485,9.96223,8.113008,6.261973,4.4127507,2.561716,0.7124943,0.56927025,0.42785916,0.28463513,0.14322405,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.038072214,0.05076295,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.13778515,0.15047589,0.14684997,0.14503701,0.14322405,0.13959812,0.13778515,0.12690738,0.11784257,0.10696479,0.09789998,0.0870222,0.08339628,0.07795739,0.072518505,0.06707962,0.06164073,0.07070554,0.07795739,0.08520924,0.092461094,0.099712946,1.0098201,1.9199274,2.8300345,3.7401419,4.650249,9.467291,14.284332,19.103188,23.920229,28.73727,27.239763,25.742256,24.24475,22.747242,21.249735,19.657953,18.06436,16.472578,14.880796,13.287203,13.252756,13.21831,13.182051,13.147605,13.113158,15.616859,18.122374,20.627888,23.13159,25.637104,25.47575,25.312584,25.149418,24.988064,24.824896,23.87309,22.919474,21.967669,21.015862,20.062244,21.296871,22.533312,23.767939,25.002567,26.237194,24.308203,22.377398,20.446592,18.5176,16.586794,15.477262,14.367728,13.258195,12.14685,11.037316,10.283124,9.527119,8.772926,8.01692,7.262728,5.870373,4.478018,3.0856624,1.693307,0.2991388,0.23931105,0.1794833,0.11965553,0.059827764,0.0,0.0,0.0,0.0,0.0,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.09064813,0.07977036,0.07070554,0.059827764,0.05076295,0.5293851,1.0098201,1.4902552,1.9706904,2.4493124,3.2143826,3.9794528,4.744523,5.5095935,6.2746634,7.168454,8.0604315,8.952409,9.844387,10.738177,10.411844,10.087324,9.762803,9.438283,9.11195,10.906783,12.703429,14.498261,16.293095,18.087927,19.844688,21.603262,23.360023,25.116783,26.875357,23.254871,19.634384,16.01571,12.395226,8.774739,7.8265595,6.880193,5.9320135,4.985647,4.0374675,2.4873846,2.6831846,2.8771715,3.0729716,3.2669585,3.4627585,3.9323158,4.401873,4.8732433,5.3428006,5.812358,10.872336,15.932315,20.992294,26.052273,31.112251,29.331923,27.553406,25.773077,23.992746,22.212418,22.658407,23.102583,23.546759,23.992746,24.436922,26.933372,29.428009,31.922646,34.417282,36.91192,32.800117,28.68832,24.574707,20.462908,16.349297,13.580903,10.810696,8.040489,5.2702823,2.5000753,3.1853752,3.870675,4.554162,5.239462,5.924762,4.972956,4.019338,3.0675328,2.1157274,1.162109,1.9253663,2.6868105,3.4500678,4.213325,4.974769,5.7579694,6.539356,7.322556,8.105756,8.887142,8.600695,8.312433,8.024173,7.7377243,7.4494634,7.8755093,8.299743,8.725789,9.1500225,9.574255,9.102885,8.629702,8.158332,7.6851482,7.211965,6.397945,5.582112,4.7680917,3.9522583,3.1382382,2.6052272,2.0722163,1.5392052,1.0080072,0.4749962,0.38072214,0.28463513,0.19036107,0.09427405,0.0,0.12328146,0.24474995,0.3680314,0.4894999,0.61278135,1.1548572,1.696933,2.2408218,2.7828975,3.3249733,3.7618973,4.2006345,4.6375585,5.0744824,5.5132194,6.43783,7.362441,8.287052,9.211663,10.138086,8.780178,7.422269,6.0643597,4.708264,3.350355,2.6849976,2.0196402,1.3542831,0.69073874,0.025381476,0.10515183,0.18492219,0.26469254,0.3444629,0.42423326,0.71430725,1.0043813,1.2944553,1.5845293,1.8746033,2.4801328,3.0856624,3.6893787,4.2949085,4.900438,4.847862,4.795286,4.74271,4.690134,4.6375585,4.7572136,4.876869,4.9983377,5.1179934,5.237649,5.5549173,5.8721857,6.189454,6.506723,6.825804,6.6173134,6.4106355,6.202145,5.995467,5.7869763,5.368182,4.947575,4.5269675,4.1081734,3.6875658,4.0030212,4.3166637,4.632119,4.947575,5.2630305,4.88956,4.517903,4.1444325,3.7727752,3.3993049,3.531651,3.6658103,3.7981565,3.930503,4.062849,3.5243993,2.9877625,2.4493124,1.9126755,1.3742256,1.8999848,2.4257438,2.94969,3.4754493,3.9993954,3.7419548,3.484514,3.2270734,2.9696326,2.712192,2.8155308,2.9170568,3.0203958,3.1219215,3.2252605,3.4101827,3.5951047,3.780027,3.9649491,4.1498713,5.863121,7.574558,9.287807,10.999244,12.712494,11.900287,11.088079,10.275872,9.461852,8.649645,8.571687,8.495543,8.417585,8.339628,8.26167,10.41547,12.567456,14.719443,16.873243,19.025229,19.072367,19.119503,19.166641,19.21559,19.262728,16.92038,14.5780325,12.235684,9.893337,7.549176,7.3878226,7.224656,7.063302,6.9001355,6.736969,7.819308,8.901647,9.985798,11.068136,12.1504755,11.26031,10.370146,9.479981,8.589817,7.699652,8.778365,9.855265,10.932164,12.010877,13.087777,14.409427,15.732889,17.054539,18.378002,19.699652,17.092611,14.485571,11.876718,9.269678,6.6626377,7.0433598,7.422269,7.802991,8.1819,8.562622,10.069194,11.5775795,13.084151,14.592536,16.099108,14.21544,12.329959,10.444477,8.560809,6.6753283,6.70071,6.7242785,6.7496595,6.775041,6.8004227,6.972654,7.1448855,7.317117,7.4893484,7.663393,6.7043357,5.7470913,4.7898474,3.832603,2.8753586,2.9768846,3.0802233,3.1817493,3.2850883,3.386614,2.8898623,2.3931105,1.8945459,1.3977941,0.89922947,0.8122072,0.72518504,0.63816285,0.5493277,0.46230546,2.2081885,3.9522583,5.6981416,7.4422116,9.188094,7.4331465,5.678199,3.923251,2.1683033,0.41335547,0.37165734,0.33177215,0.291887,0.2520018,0.21211663,0.6744221,1.1367276,1.6008459,2.0631514,2.525457,2.422118,2.3205922,2.2172532,2.1157274,2.0123885,2.4891977,2.9678197,3.444629,3.923251,4.40006,4.4254417,4.4508233,4.4743915,4.499773,4.5251546,4.40006,4.274966,4.1498713,4.024777,3.8996825,3.6041696,3.3104696,3.0149567,2.7194438,2.4257438,2.034144,1.6443571,1.2545701,0.86478317,0.4749962,0.40791658,0.34083697,0.27194437,0.20486477,0.13778515,0.11059072,0.08339628,0.054388877,0.027194439,0.0,0.0,0.0,0.0,0.0,0.0,0.24293698,0.48587397,0.726998,0.969935,1.2128719,1.4231756,1.6316663,1.84197,2.0522738,2.2625773,3.000453,3.738329,4.4743915,5.2122674,5.9501433,5.3083544,4.664753,4.022964,3.3793623,2.7375734,2.322405,1.9072367,1.4920682,1.0768998,0.66173136,0.53663695,0.41335547,0.28826106,0.16316663,0.038072214,0.05076295,0.06164073,0.07433146,0.0870222,0.099712946,0.10515183,0.11059072,0.11421664,0.11965553,0.12509441,0.11965553,0.11421664,0.11059072,0.10515183,0.099712946,0.092461094,0.08520924,0.07795739,0.07070554,0.06164073,0.11240368,0.16316663,0.21211663,0.26287958,0.31182957,0.9572442,1.6026589,2.2480736,2.8916752,3.53709,3.0729716,2.6070402,2.1429217,1.6769904,1.2128719,1.062396,0.9119202,0.76325727,0.61278135,0.46230546,0.82671094,1.1929294,1.5573349,1.9217403,2.2879589,3.0729716,3.8579843,4.6429973,5.42801,6.2130227,6.972654,7.7322855,8.491917,9.253361,10.012992,8.722163,7.4331465,6.1423173,4.853301,3.5624714,5.1578784,6.7532854,8.34688,9.9422865,11.537694,9.3150015,7.0923095,4.8696175,2.6469254,0.42423326,1.0823387,1.7404441,2.3967366,3.054842,3.7129474,4.2350807,4.7572136,5.279347,5.803293,6.3254266,6.0281005,5.730775,5.431636,5.1343102,4.836984,4.88956,4.942136,4.994712,5.047288,5.0998635,4.461701,3.825351,3.1871881,2.5508385,1.9126755,8.9596615,16.006647,23.055445,30.10243,37.149418,30.303669,23.459736,16.613989,9.770056,2.9243085,9.470917,16.013899,22.560507,29.1053,35.650097,28.864178,22.08007,15.294152,8.510046,1.7241274,10.034748,18.345367,26.655989,34.964798,43.275417,35.171474,27.071157,18.967215,10.865085,2.762955,3.966762,5.1723824,6.378002,7.5818095,8.78743,7.1630154,5.5367875,3.9123733,2.2879589,0.66173136,0.5293851,0.39703882,0.26469254,0.13234627,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.05076295,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.13778515,0.15047589,0.16316663,0.16497959,0.16679256,0.17041849,0.17223145,0.17585737,0.15954071,0.14503701,0.13053331,0.11421664,0.099712946,0.092461094,0.08520924,0.07795739,0.07070554,0.06164073,0.07977036,0.09789998,0.11421664,0.13234627,0.15047589,1.3651608,2.5798457,3.7945306,5.009216,6.2257137,10.408218,14.590723,18.773228,22.953918,27.138237,25.397793,23.657349,21.916904,20.178274,18.43783,16.730019,15.022208,13.314397,11.608399,9.900589,10.410031,10.919474,11.430729,11.940171,12.449615,15.094727,17.73984,20.38495,23.030064,25.675177,26.462002,27.25064,28.037466,28.824291,29.61293,28.539658,27.468197,26.394922,25.323462,24.250187,25.027948,25.80571,26.581657,27.359419,28.137178,25.80571,23.472427,21.139143,18.807674,16.474392,15.5606575,14.645112,13.729566,12.815832,11.900287,11.104396,10.310318,9.514427,8.72035,7.9244595,6.4051967,4.8859344,3.3648586,1.845596,0.3245203,0.25925365,0.19579996,0.13053331,0.065266654,0.0,0.0,0.0,0.0,0.0,0.0,0.018129626,0.034446288,0.052575916,0.07070554,0.0870222,0.08520924,0.08339628,0.07977036,0.07795739,0.07433146,0.75781834,1.4394923,2.1229792,2.8046532,3.48814,4.0972953,4.708264,5.317419,5.9265747,6.5375433,7.231908,7.9280853,8.62245,9.316814,10.012992,10.125396,10.2378,10.3502035,10.462607,10.57501,12.930049,15.285088,17.640125,19.995165,22.350203,24.542074,26.73576,28.927631,31.119503,33.313187,28.044718,22.776249,17.509592,12.242936,6.9744673,6.3725634,5.77066,5.1669436,4.5650396,3.9631362,2.3369088,2.5091403,2.6831846,2.855416,3.0276475,3.199879,3.435564,3.6694362,3.9051213,4.1408067,4.3746786,9.692098,15.009518,20.326937,25.644356,30.961775,29.348238,27.73289,26.117538,24.50219,22.886839,23.648283,24.407915,25.167547,25.927177,26.68681,29.034595,31.382381,33.730167,36.077957,38.425743,33.6504,28.875055,24.099712,19.324368,14.5508375,12.114216,9.679407,7.2445984,4.8097897,2.374981,3.0294604,3.6857529,4.3402324,4.994712,5.6491914,4.7916603,3.9341288,3.0765975,2.220879,1.3633479,2.3876717,3.4119956,4.4381323,5.462456,6.48678,7.1974616,7.9081426,8.617011,9.327692,10.038374,8.925215,7.8120556,6.70071,5.5875506,4.4743915,5.2865987,6.1006193,6.9128265,7.7250338,8.537241,8.007855,7.476658,6.947273,6.4178877,5.8866897,5.3428006,4.797099,4.25321,3.7075086,3.1618068,2.5780327,1.9924458,1.4068589,0.823085,0.2374981,0.19036107,0.14322405,0.09427405,0.047137026,0.0,0.14322405,0.28463513,0.42785916,0.56927025,0.7124943,1.0895905,1.4666867,1.845596,2.222692,2.5997884,3.5497808,4.499773,5.4497657,6.399758,7.3497505,8.575313,9.799063,11.024626,12.250188,13.475751,11.5775795,9.679407,7.783048,5.8848767,3.9867048,3.1926272,2.3967366,1.6026589,0.80676836,0.012690738,0.052575916,0.092461094,0.13234627,0.17223145,0.21211663,0.35715362,0.50219065,0.64722764,0.79226464,0.93730164,1.8528478,2.7665808,3.682127,4.597673,5.5132194,5.480586,5.4479527,5.4153194,5.382686,5.3500524,5.3591175,5.369995,5.3808727,5.389938,5.4008155,5.7398396,6.0806766,6.4197006,6.7605376,7.0995617,6.7532854,6.4051967,6.057108,5.710832,5.3627434,4.940323,4.517903,4.0954823,3.673062,3.2506418,3.7818398,4.314851,4.847862,5.3808727,5.9120708,5.331923,4.751775,4.171627,3.5932918,3.0131438,3.1726844,3.3322253,3.491766,3.6531196,3.8126602,3.3122826,2.811905,2.3133402,1.8129625,1.3125849,1.7132497,2.1121013,2.5127661,2.911618,3.3122826,3.1781235,3.0421512,2.907992,2.7720199,2.6378605,2.7194438,2.8028402,2.8844235,2.9678197,3.049403,3.1545548,3.2597067,3.3648586,3.4700103,3.5751622,5.1741953,6.775041,8.375887,9.97492,11.575767,10.863272,10.150778,9.438283,8.725789,8.013294,7.7304726,7.4476504,7.1648283,6.882006,6.599184,9.507175,12.415168,15.32316,18.22934,21.137331,20.430275,19.72322,19.01435,18.307297,17.60024,15.596917,13.595407,11.592083,9.590572,7.5872483,7.512917,7.4367723,7.362441,7.28811,7.211965,8.247167,9.282369,10.31757,11.352772,12.387974,11.6047735,10.823386,10.040187,9.256987,8.4756,9.782746,11.089892,12.397038,13.704185,15.013144,16.068287,17.121618,18.176764,19.231907,20.287052,17.402628,14.518205,11.631968,8.747544,5.863121,6.2148356,6.5683637,6.9200783,7.271793,7.6253204,9.159087,10.694666,12.230246,13.765825,15.299591,13.270886,11.240368,9.20985,7.179332,5.1506267,5.5494785,5.9501433,6.350808,6.7496595,7.1503243,7.7304726,8.31062,8.890768,9.469104,10.049252,8.664148,7.2808576,5.8957543,4.510651,3.1255474,3.2578938,3.39024,3.5225863,3.6549325,3.787279,3.1817493,2.5780327,1.9725033,1.3669738,0.76325727,0.72518504,0.6871128,0.6508536,0.61278135,0.5747091,1.8854811,3.1944401,4.505212,5.814171,7.124943,5.810545,4.494334,3.1799364,1.8655385,0.5493277,0.46774435,0.38434806,0.30276474,0.21936847,0.13778515,0.7505665,1.3633479,1.9743162,2.5870976,3.199879,2.9424384,2.6849976,2.427557,2.1701162,1.9126755,1.9706904,2.0268922,2.084907,2.1429217,2.1991236,2.4130533,2.6251698,2.8372865,3.049403,3.2633326,3.1382382,3.0131438,2.8880494,2.762955,2.6378605,2.6269827,2.617918,2.6070402,2.5979755,2.5870976,2.1175404,1.647983,1.1766127,0.7070554,0.2374981,0.2229944,0.20667773,0.19217403,0.17767033,0.16316663,0.13053331,0.09789998,0.065266654,0.032633327,0.0,0.0,0.0,0.0,0.0,0.0,0.3154555,0.629098,0.9445535,1.260009,1.5754645,1.7168756,1.8600996,2.0033236,2.1447346,2.2879589,3.0747845,3.8616104,4.650249,5.4370747,6.2257137,5.5476656,4.8696175,4.1933823,3.5153344,2.8372865,2.4058013,1.9725033,1.5392052,1.1077201,0.6744221,0.5493277,0.42423326,0.2991388,0.17585737,0.05076295,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.11421664,0.11784257,0.11965553,0.12328146,0.12509441,0.12328146,0.11965553,0.11784257,0.11421664,0.11240368,0.10333887,0.092461094,0.08339628,0.072518505,0.06164073,0.0870222,0.11240368,0.13778515,0.16316663,0.18673515,0.7106813,1.2328146,1.7549478,2.277081,2.7992141,2.3677292,1.9344311,1.502946,1.0696479,0.63816285,0.5620184,0.48768693,0.41335547,0.33721104,0.26287958,0.44417584,0.62728506,0.8103943,0.9916905,1.1747998,2.1556125,3.1346123,4.115425,5.0944247,6.0752378,7.41683,8.760235,10.101828,11.445232,12.786825,10.90497,9.023115,7.1394467,5.2575917,3.3757362,4.710077,6.0444174,7.380571,8.714911,10.049252,8.120259,6.189454,4.2604623,2.3296568,0.40066472,1.0841516,1.7694515,2.4547513,3.1400511,3.825351,4.505212,5.185073,5.864934,6.544795,7.224656,6.9073873,6.590119,6.2728505,5.955582,5.638314,5.6945157,5.75253,5.810545,5.866747,5.924762,5.199577,4.4743915,3.7492065,3.0258346,2.3006494,8.81825,15.334038,21.85345,28.369238,34.88684,28.526966,22.167093,15.80722,9.447348,3.0874753,9.048496,15.007704,20.966911,26.927933,32.887142,26.532707,20.178274,13.822026,7.4675927,1.1131591,12.431484,23.747997,35.06451,46.382835,57.69935,46.76718,35.83502,24.902855,13.97069,3.0367124,3.9522583,4.8678045,5.7833505,6.697084,7.61263,6.2130227,4.8134155,3.4119956,2.0123885,0.61278135,0.4894999,0.3680314,0.24474995,0.12328146,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.13778515,0.15047589,0.16316663,0.17585737,0.18310922,0.19036107,0.19761293,0.20486477,0.21211663,0.19217403,0.17223145,0.15228885,0.13234627,0.11240368,0.10333887,0.092461094,0.08339628,0.072518505,0.06164073,0.09064813,0.11784257,0.14503701,0.17223145,0.19942589,1.7205015,3.2397642,4.76084,6.2801023,7.799365,11.347333,14.895301,18.443268,21.989424,25.537392,23.55401,21.572441,19.58906,17.607492,15.624111,13.802084,11.980057,10.15803,8.336002,6.5121617,7.567306,8.62245,9.677594,10.7327385,11.787883,14.572594,17.357304,20.142014,22.926725,25.71325,27.450066,29.186884,30.925516,32.662334,34.39915,33.208035,32.015106,30.822176,29.629248,28.438131,28.757212,29.078106,29.397188,29.718082,30.037165,27.303217,24.567455,21.831696,19.097748,16.361988,15.6422415,14.922495,14.202749,13.483003,12.763257,11.927481,11.091705,10.257742,9.421967,8.588004,6.9400206,5.292038,3.644055,1.9978848,0.34990177,0.27919623,0.21030366,0.13959812,0.07070554,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.07977036,0.08520924,0.09064813,0.09427405,0.099712946,0.98443866,1.8709774,2.7557032,3.6404288,4.5251546,4.9802084,5.4352617,5.8903155,6.345369,6.8004227,7.2971745,7.795739,8.292491,8.789243,9.287807,9.837135,10.388275,10.937603,11.486931,12.038072,14.953316,17.868559,20.78199,23.697233,26.612478,29.23946,31.868256,34.49524,37.122223,39.749203,32.834564,25.919926,19.005287,12.090648,5.1741953,4.9167547,4.6593137,4.401873,4.1444325,3.8869917,2.1882458,2.3369088,2.4873846,2.6378605,2.7883365,2.9369993,2.9369993,2.9369993,2.9369993,2.9369993,2.9369993,8.511859,14.0867195,19.663393,25.238253,30.813112,29.362741,27.912373,26.462002,25.011631,23.563074,24.63816,25.71325,26.788336,27.863422,28.936695,31.137632,33.336758,35.537693,37.736816,39.93775,34.50068,29.06179,23.624716,18.187641,12.750566,10.649343,8.549932,6.450521,4.349297,2.2498865,2.8753586,3.5008307,4.12449,4.749962,5.375434,4.612177,3.8507326,3.0874753,2.324218,1.5627737,2.8499773,4.137181,5.424384,6.7134004,8.000604,8.636953,9.275117,9.91328,10.549629,11.187792,9.249735,7.311678,5.375434,3.437377,1.49932,2.6995013,3.8996825,5.0998635,6.300045,7.500226,6.9128265,6.3254266,5.7380266,5.1506267,4.5632267,4.2876563,4.0120864,3.738329,3.4627585,3.1871881,2.5508385,1.9126755,1.2745126,0.63816285,0.0,0.0,0.0,0.0,0.0,0.0,0.16316663,0.3245203,0.48768693,0.6508536,0.8122072,1.0243238,1.2382535,1.4503701,1.6624867,1.8746033,3.3376641,4.800725,6.261973,7.7250338,9.188094,10.712796,12.237497,13.762199,15.2869005,16.811602,14.37498,11.938358,9.499924,7.063302,4.6248674,3.7002566,2.7756457,1.8492218,0.9246109,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.2255627,2.4493124,3.6748753,4.900438,6.1241875,6.11331,6.1006193,6.0879283,6.0752378,6.0625467,5.962834,5.863121,5.7615952,5.661882,5.562169,5.924762,6.2873545,6.6499467,7.0125394,7.3751316,6.887445,6.399758,5.9120708,5.424384,4.936697,4.512464,4.0882306,3.6621845,3.2379513,2.811905,3.5624714,4.313038,5.0617914,5.812358,6.5629244,5.774286,4.98746,4.2006345,3.4119956,2.6251698,2.811905,3.000453,3.1871881,3.3757362,3.5624714,3.100166,2.6378605,2.175555,1.7132497,1.2491312,1.5247015,1.8002719,2.0758421,2.3495996,2.6251698,2.612479,2.5997884,2.5870976,2.5744069,2.561716,2.6251698,2.6868105,2.7502642,2.811905,2.8753586,2.9007401,2.9243085,2.94969,2.9750717,3.000453,4.4870825,5.975525,7.462154,8.950596,10.437225,9.824444,9.211663,8.600695,7.987913,7.3751316,6.887445,6.399758,5.9120708,5.424384,4.936697,8.600695,12.262879,15.925063,19.587248,23.249432,21.788185,20.325123,18.862062,17.400814,15.937754,14.275268,12.612781,10.950294,9.287807,7.6253204,7.6380115,7.650702,7.663393,7.6742706,7.686961,8.675026,9.663091,10.649343,11.637406,12.625471,11.949236,11.274815,10.600392,9.924157,9.249735,10.7871275,12.32452,13.861912,15.399304,16.936697,17.725336,18.512161,19.3008,20.087626,20.87445,17.712645,14.5508375,11.3872175,8.225411,5.0617914,5.388125,5.712645,6.037165,6.3616858,6.688019,8.2507925,9.811753,11.374527,12.937301,14.500074,12.32452,10.150778,7.9752226,5.7996674,3.6241121,4.40006,5.1741953,5.9501433,6.7242785,7.500226,8.488291,9.474543,10.462607,11.450671,12.436923,10.625773,8.812811,6.9998484,5.186886,3.3757362,3.53709,3.7002566,3.8616104,4.024777,4.1879435,3.4754493,2.762955,2.0504606,1.3379664,0.62547207,0.63816285,0.6508536,0.66173136,0.6744221,0.6871128,1.5627737,2.4366217,3.3122826,4.1879435,5.0617914,4.1879435,3.3122826,2.4366217,1.5627737,0.6871128,0.5620184,0.43692398,0.31182957,0.18673515,0.06164073,0.824898,1.5881553,2.3495996,3.1128569,3.874301,3.4627585,3.049403,2.6378605,2.2245052,1.8129625,1.4503701,1.0877775,0.72518504,0.36259252,0.0,0.40066472,0.7995165,1.2001812,1.6008459,1.9996977,1.8746033,1.7495089,1.6244144,1.49932,1.3742256,1.649796,1.9253663,2.1991236,2.474694,2.7502642,2.1991236,1.649796,1.1004683,0.5493277,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.0,0.0,0.0,0.0,0.0,0.387974,0.774135,1.162109,1.550083,1.938057,2.0123885,2.08672,2.1628644,2.2371957,2.3133402,3.150929,3.9867048,4.8242936,5.661882,6.4994707,5.7869763,5.0744824,4.361988,3.6494937,2.9369993,2.4873846,2.03777,1.5881553,1.1367276,0.6871128,0.5620184,0.43692398,0.31182957,0.18673515,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.46230546,0.8629702,1.261822,1.6624867,2.0631514,1.6624867,1.261822,0.8629702,0.46230546,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,1.2382535,2.4130533,3.587853,4.762653,5.9374523,7.8628187,9.788185,11.711739,13.637105,15.56247,13.087777,10.613083,8.136576,5.661882,3.1871881,4.262275,5.337362,6.412449,7.4875355,8.562622,6.925517,5.2884116,3.6494937,2.0123885,0.37528324,1.0877775,1.8002719,2.5127661,3.2252605,3.9377546,4.7753434,5.612932,6.450521,7.28811,8.125698,7.7866745,7.4494634,7.112252,6.775041,6.43783,6.4994707,6.5629244,6.624565,6.688019,6.7496595,5.9374523,5.125245,4.313038,3.5008307,2.6868105,8.675026,14.661428,20.649643,26.63786,32.62426,26.750263,20.87445,15.000452,9.12464,3.2506418,8.626076,13.999697,19.375132,24.750565,30.124186,24.199425,18.274662,12.349901,6.4251394,0.50037766,14.826408,29.148813,43.474842,57.800873,72.12509,58.36108,44.600693,30.836681,17.074482,3.3122826,3.9377546,4.5632267,5.186886,5.812358,6.43783,5.2630305,4.0882306,2.911618,1.7368182,0.5620184,0.44961473,0.33721104,0.22480737,0.11240368,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.13778515,0.15047589,0.16316663,0.17585737,0.18673515,0.19942589,0.21211663,0.22480737,0.2374981,0.25018883,0.22480737,0.19942589,0.17585737,0.15047589,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.099712946,0.13778515,0.17585737,0.21211663,0.25018883,2.0758421,3.8996825,5.7253356,7.549176,9.374829,12.28826,15.199879,18.11331,21.024927,23.938358,21.71204,19.487535,17.26303,15.038525,12.812206,10.874149,8.937905,6.9998484,5.0617914,3.1255474,4.7245803,6.3254266,7.9244595,9.525306,11.124338,14.05046,16.97477,19.90089,22.8252,25.749508,28.438131,31.12494,33.811752,36.500374,39.187187,37.8746,36.562016,35.24943,33.936848,32.62426,32.48829,32.350506,32.21272,32.074936,31.93715,28.79891,25.662485,22.524246,19.387821,16.249584,15.725637,15.199879,14.674119,14.150173,13.6244135,12.750566,11.874905,10.999244,10.125396,9.249735,7.474845,5.6999545,3.925064,2.1501737,0.37528324,0.2991388,0.22480737,0.15047589,0.07433146,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,1.2128719,2.3006494,3.388427,4.4743915,5.562169,5.863121,6.16226,6.4632115,6.7623506,7.063302,7.362441,7.663393,7.9625316,8.26167,8.562622,9.550687,10.536939,11.525003,12.513068,13.499319,16.97477,20.450218,23.925667,27.399303,30.874752,33.936848,37.00075,40.062847,43.124943,46.187035,37.624413,29.06179,20.499168,11.938358,3.3757362,3.4627585,3.5497808,3.636803,3.7256382,3.8126602,2.4366217,2.565342,2.6922495,2.819157,2.9478772,3.0747845,3.0856624,3.094727,3.105605,3.1146698,3.1255474,8.760235,14.394923,20.02961,25.664299,31.300798,30.247467,29.194136,28.142618,27.089287,26.03777,26.597975,27.15818,27.718386,28.276777,28.836983,31.445835,34.052876,36.659916,39.266956,41.87581,36.065266,30.254719,24.444174,18.635443,12.824898,10.805257,8.785617,6.7641635,4.744523,2.7248828,3.1871881,3.6494937,4.1117992,4.574105,5.038223,4.3946214,3.7528327,3.1092308,2.467442,1.8256533,2.9696326,4.115425,5.2594047,6.4051967,7.549176,7.9715962,8.39583,8.81825,9.24067,9.663091,8.113008,6.5629244,5.0128417,3.4627585,1.9126755,3.1726844,4.4326935,5.6927023,6.9527116,8.212721,7.415017,6.6173134,5.81961,5.0219064,4.2242026,3.9522583,3.680314,3.4083695,3.1346123,2.8626678,2.3405347,1.8184015,1.2944553,0.77232206,0.25018883,0.26469254,0.27919623,0.2955129,0.3100166,0.3245203,0.4169814,0.5094425,0.60190356,0.69436467,0.7868258,1.0750868,1.3633479,1.649796,1.938057,2.2245052,3.4573197,4.690134,5.922949,7.155763,8.386765,9.594198,10.801631,12.010877,13.21831,14.425743,12.449615,10.475298,8.499168,6.5248523,4.550536,3.9450066,3.339477,2.7357605,2.1302311,1.5247015,1.452183,1.3796645,1.3071461,1.2346275,1.162109,0.9318628,0.7016165,0.47318324,0.24293698,0.012690738,0.9898776,1.9670644,2.9442513,3.923251,4.900438,5.027345,5.1542525,5.282973,5.40988,5.5367875,5.922949,6.3072968,6.6916447,7.077806,7.462154,7.554615,7.647076,7.7395372,7.8319983,7.9244595,7.2826705,6.640882,5.99728,5.3554916,4.7118897,4.249584,3.787279,3.3249733,2.8626678,2.4003625,3.105605,3.8108473,4.514277,5.219519,5.924762,5.23221,4.539658,3.8471067,3.1545548,2.4620032,2.6378605,2.811905,2.9877625,3.1618068,3.3376641,2.9641938,2.5925364,2.220879,1.8474089,1.4757515,1.7404441,2.0051367,2.269829,2.5345216,2.7992141,2.770207,2.7393866,2.7103791,2.6795588,2.6505513,2.6505513,2.6505513,2.6505513,2.6505513,2.6505513,2.6995013,2.7502642,2.7992141,2.8499773,2.9007401,4.169814,5.4407005,6.7097745,7.9806614,9.249735,8.841819,8.435715,8.027799,7.6198816,7.211965,6.8403077,6.4668374,6.09518,5.7217097,5.3500524,8.636953,11.925668,15.212569,18.49947,21.788185,20.430275,19.072367,17.714457,16.358362,15.000452,13.366973,11.735307,10.101828,8.470161,6.836682,7.17208,7.507478,7.842876,8.178274,8.511859,9.24067,9.967669,10.694666,11.421664,12.1504755,11.327391,10.504305,9.683033,8.859948,8.036863,9.499924,10.962985,12.4242325,13.887294,15.350354,16.342045,17.335548,18.327238,19.320742,20.312433,17.292038,14.273455,11.253058,8.232663,5.2122674,5.337362,5.462456,5.5875506,5.712645,5.8377395,7.2029004,8.568061,9.933222,11.298383,12.661731,11.300196,9.936848,8.575313,7.211965,5.8504305,6.4994707,7.1503243,7.799365,8.450218,9.099259,9.768243,10.435412,11.102583,11.769753,12.436923,10.81976,9.202598,7.5854354,5.9682727,4.349297,4.329355,4.309412,4.2894692,4.269527,4.249584,3.5624714,2.8753586,2.1882458,1.49932,0.8122072,0.7904517,0.7668832,0.7451276,0.72337204,0.69980353,1.4503701,2.1991236,2.94969,3.7002566,4.4508233,3.6948178,2.9406252,2.18462,1.4304274,0.6744221,0.581961,0.4894999,0.39703882,0.3045777,0.21211663,0.8321498,1.452183,2.0722163,2.6922495,3.3122826,3.045777,2.7774587,2.5091403,2.2426348,1.9743162,1.5790904,1.1856775,0.7904517,0.39522585,0.0,0.44417584,0.8901646,1.3343405,1.7803292,2.2245052,2.0033236,1.7803292,1.5573349,1.3343405,1.1131591,1.3307146,1.54827,1.7658255,1.983381,2.1991236,1.8945459,1.5899682,1.2853905,0.9808127,0.6744221,0.56927025,0.46411842,0.36077955,0.25562772,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.0,0.0,0.0,0.0,0.0,0.3100166,0.6200332,0.9300498,1.2400664,1.550083,1.6896812,1.8292793,1.9706904,2.1102884,2.2498865,3.000453,3.7492065,4.499773,5.2503395,5.999093,5.6093063,5.219519,4.8297324,4.439945,4.0501585,3.3557937,2.659616,1.9652514,1.2708868,0.5747091,0.47680917,0.38072214,0.28282216,0.18492219,0.0870222,0.092461094,0.09789998,0.10333887,0.10696479,0.11240368,0.11240368,0.11240368,0.11240368,0.11240368,0.11240368,0.11421664,0.11784257,0.11965553,0.12328146,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.6345369,1.2074331,1.7803292,2.3532255,2.9243085,2.3532255,1.7803292,1.2074331,0.6345369,0.06164073,0.059827764,0.058014803,0.054388877,0.052575916,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.99712944,1.9453088,2.8916752,3.8398547,4.788034,6.755099,8.722163,10.689227,12.658105,14.625169,12.978999,11.334642,9.690285,8.044115,6.399758,6.7859187,7.170267,7.554615,7.9407763,8.325124,6.932769,5.540414,4.1480584,2.7557032,1.3633479,2.3604772,3.3576066,4.3547363,5.351866,6.350808,6.967215,7.5854354,8.201842,8.820063,9.438283,8.937905,8.437528,7.93715,7.4367723,6.9382076,6.9617763,6.987158,7.0125394,7.037921,7.063302,6.261973,5.462456,4.6629395,3.8616104,3.0620937,8.930654,14.7974,20.66596,26.532707,32.399456,26.440247,20.48104,14.520018,8.560809,2.5997884,7.5219817,12.444175,17.368181,22.290375,27.212568,22.194288,17.17782,12.15954,7.1430726,2.124792,13.976129,25.82384,37.675175,49.5247,61.37422,50.151985,38.929745,27.707508,16.48527,5.2630305,5.522284,5.7833505,6.0426044,6.301858,6.5629244,5.3391747,4.117238,2.8953013,1.6733645,0.44961473,0.36077955,0.27013144,0.1794833,0.09064813,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.13959812,0.15410182,0.17041849,0.18492219,0.19942589,0.21030366,0.21936847,0.23024625,0.23931105,0.25018883,0.2229944,0.19579996,0.16679256,0.13959812,0.11240368,0.15772775,0.2030518,0.24837588,0.291887,0.33721104,0.65810543,0.97718686,1.2980812,1.6171626,1.938057,3.0620937,4.1879435,5.3119802,6.43783,7.5618668,9.994863,12.427858,14.860854,17.292038,19.725033,18.289167,16.855114,15.419247,13.985193,12.549327,11.432542,10.315757,9.197159,8.080374,6.9617763,8.424837,9.8878975,11.350959,12.812206,14.275268,16.862366,19.449463,22.038374,24.625471,27.212568,29.112553,31.012537,32.91252,34.812508,36.712494,35.069946,33.427402,31.78486,30.142317,28.499771,28.659313,28.820665,28.980207,29.139748,29.299288,26.976883,24.654478,22.332073,20.009668,17.687263,16.80979,15.932315,15.054841,14.177367,13.299893,12.429671,11.559449,10.689227,9.820818,8.950596,7.304426,5.660069,4.0157123,2.3695421,0.72518504,0.58014804,0.43511102,0.29007402,0.14503701,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.20667773,0.3154555,0.4224203,0.5293851,0.63816285,0.53482395,0.43329805,0.32995918,0.22662032,0.12509441,1.2328146,2.3405347,3.4482548,4.554162,5.661882,5.995467,6.3272395,6.6608243,6.9925966,7.324369,7.7123427,8.100317,8.488291,8.874452,9.262425,9.935035,10.607644,11.280253,11.952863,12.625471,15.790904,18.954523,22.119957,25.285389,28.45082,30.990782,33.530743,36.070705,38.610664,41.150623,33.9024,26.654177,19.407764,12.15954,4.9131284,4.7554007,4.597673,4.439945,4.2822175,4.12449,2.6868105,2.7919624,2.8971143,3.002266,3.1074178,3.2125697,3.2325122,3.2524548,3.2723975,3.29234,3.3122826,9.006798,14.703127,20.397642,26.092157,31.786673,31.132193,30.477715,29.823235,29.166943,28.512463,28.557787,28.603111,28.646622,28.691946,28.73727,31.752226,34.767185,37.78214,40.797096,43.812054,37.629852,31.447649,25.265446,19.083244,12.899229,10.959359,9.019489,7.079619,5.139749,3.199879,3.5008307,3.7999697,4.099108,4.40006,4.699199,4.177066,3.6549325,3.1327994,2.610666,2.08672,3.0892882,4.0918565,5.0944247,6.096993,7.0995617,7.308052,7.51473,7.723221,7.9298983,8.138389,6.9744673,5.812358,4.650249,3.48814,2.324218,3.6458678,4.9657044,6.285541,7.605378,8.925215,7.9172077,6.9092,5.903006,4.894999,3.8869917,3.6168604,3.346729,3.0765975,2.808279,2.5381477,2.1302311,1.7223145,1.3143979,0.90829426,0.50037766,0.5293851,0.56020546,0.58921283,0.6200332,0.6508536,0.6726091,0.69436467,0.7179332,0.73968875,0.76325727,1.1258497,1.4866294,1.8492218,2.2118144,2.5744069,3.576975,4.5795436,5.582112,6.58468,7.5872483,8.477413,9.367578,10.257742,11.147907,12.038072,10.524248,9.012237,7.500226,5.9882154,4.4743915,4.1897564,3.9051213,3.6204863,3.3358512,3.049403,2.904366,2.759329,2.6142921,2.469255,2.324218,1.8655385,1.405046,0.9445535,0.48587397,0.025381476,0.7541924,1.4848163,2.2154403,2.9442513,3.6748753,3.9431937,4.209699,4.478018,4.744523,5.0128417,5.883064,6.7532854,7.6216946,8.491917,9.362139,9.184468,9.006798,8.829127,8.653271,8.4756,7.6778965,6.880193,6.0824895,5.2847857,4.4870825,3.9867048,3.48814,2.9877625,2.4873846,1.987007,2.6469254,3.3068438,3.966762,4.6266804,5.2865987,4.690134,4.0918565,3.4953918,2.8971143,2.3006494,2.4620032,2.6251698,2.7883365,2.94969,3.1128569,2.8300345,2.5472124,2.2643902,1.983381,1.7005589,1.9543737,2.2100015,2.465629,2.7194438,2.9750717,2.9279346,2.8807976,2.8318477,2.7847104,2.7375734,2.6741197,2.612479,2.5508385,2.4873846,2.4257438,2.5000753,2.5744069,2.6505513,2.7248828,2.7992141,3.8525455,4.9040637,5.957395,7.0107265,8.062244,7.859193,7.6579537,7.454902,7.25185,7.0506115,6.793171,6.53573,6.2782893,6.0208488,5.763408,8.675026,11.586644,14.500074,17.411694,20.325123,19.072367,17.819609,16.566853,15.314095,14.06315,12.460492,10.857833,9.255174,7.652515,6.049856,6.7079616,7.364254,8.02236,8.680465,9.336758,9.804502,10.272246,10.73999,11.207735,11.675479,10.705544,9.735609,8.765674,7.795739,6.825804,8.212721,9.599637,10.988366,12.375282,13.762199,14.960567,16.157122,17.355492,18.552046,19.750414,16.873243,13.994258,11.117086,8.239915,5.3627434,5.2865987,5.2122674,5.137936,5.0617914,4.98746,6.155008,7.322556,8.490104,9.657652,10.825199,10.275872,9.724731,9.175404,8.624263,8.074935,8.600695,9.12464,9.6504,10.174346,10.700105,11.048194,11.39447,11.7425585,12.090648,12.436923,11.015561,9.592385,8.1692095,6.7478466,5.3246713,5.121619,4.9203806,4.7173285,4.514277,4.313038,3.6494937,2.9877625,2.324218,1.6624867,1.0007553,0.94274056,0.88472575,0.82671094,0.7705091,0.7124943,1.3379664,1.9616255,2.5870976,3.2125697,3.8380418,3.2016919,2.5671551,1.9326181,1.2980812,0.66173136,0.60190356,0.5420758,0.48224804,0.4224203,0.36259252,0.83940166,1.3180238,1.794833,2.2716422,2.7502642,2.6269827,2.5055144,2.382233,2.2607644,2.137483,1.7096237,1.2817645,0.8557183,0.42785916,0.0,0.4894999,0.9808127,1.4703126,1.9598125,2.4493124,2.1302311,1.8093367,1.4902552,1.1693609,0.85027945,1.0098201,1.1693609,1.3307146,1.4902552,1.649796,1.5899682,1.5301404,1.4703126,1.4104849,1.3506571,1.1022812,0.8557183,0.6073425,0.36077955,0.11240368,0.09064813,0.06707962,0.045324065,0.02175555,0.0,0.0,0.0,0.0,0.0,0.0,0.23205921,0.46411842,0.6979906,0.9300498,1.162109,1.3669738,1.5718386,1.7767034,1.983381,2.1882458,2.8499773,3.5117085,4.175253,4.836984,5.5005283,5.431636,5.3645563,5.297477,5.230397,5.163317,4.2223897,3.2832751,2.3423476,1.403233,0.46230546,0.39159992,0.32270733,0.2520018,0.18310922,0.11240368,0.11059072,0.10696479,0.10515183,0.10333887,0.099712946,0.099712946,0.099712946,0.099712946,0.099712946,0.099712946,0.10515183,0.11059072,0.11421664,0.11965553,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.80676836,1.551896,2.2970235,3.0421512,3.787279,3.0421512,2.2970235,1.551896,0.80676836,0.06164073,0.058014803,0.052575916,0.047137026,0.04169814,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.75781834,1.4775645,2.1973107,2.9170568,3.636803,5.6473784,7.6579537,9.666717,11.677292,13.687867,12.872034,12.058014,11.242181,10.428161,9.612328,9.30775,9.003172,8.696781,8.392203,8.087626,6.9400206,5.7924156,4.64481,3.4972048,2.3495996,3.633177,4.914942,6.1967063,7.4802837,8.762048,9.1609,9.557939,9.954978,10.352016,10.750868,10.087324,9.425592,8.762048,8.100317,7.4367723,7.4258947,7.413204,7.400513,7.3878226,7.3751316,6.588306,5.7996674,5.0128417,4.2242026,3.437377,9.184468,14.93156,20.680464,26.427555,32.17465,26.13023,20.085812,14.039582,7.995165,1.9507477,6.4197006,10.890467,15.359419,19.830185,24.299137,20.189152,16.080978,11.969179,7.859193,3.7492065,13.125849,22.498865,31.875507,41.25034,50.625168,41.94108,33.260612,24.57652,15.894243,7.211965,7.1068134,7.0016613,6.8983226,6.793171,6.688019,5.4171324,4.1480584,2.8771715,1.6080978,0.33721104,0.27013144,0.2030518,0.13415924,0.06707962,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.14322405,0.15954071,0.17767033,0.19579996,0.21211663,0.21936847,0.22662032,0.23568514,0.24293698,0.25018883,0.21936847,0.19036107,0.15954071,0.13053331,0.099712946,0.2030518,0.3045777,0.40791658,0.5094425,0.61278135,1.214685,1.8165885,2.420305,3.0222087,3.6241121,4.0501585,4.4743915,4.900438,5.3246713,5.750717,7.703278,9.654026,11.608399,13.559147,15.511708,14.868106,14.222692,13.577277,12.931862,12.28826,11.989121,11.691795,11.39447,11.097144,10.799818,12.125093,13.45037,14.775645,16.099108,17.424383,19.67427,21.924156,24.175856,26.425743,28.675629,29.786976,30.900135,32.013294,33.124638,34.237797,32.265297,30.292791,28.320288,26.347786,24.375282,24.832148,25.290829,25.747694,26.204561,26.66324,25.154856,23.648283,22.139898,20.633327,19.124943,17.895754,16.664753,15.435563,14.204562,12.975373,12.11059,11.245807,10.37921,9.514427,8.649645,7.134008,5.620184,4.1045475,2.5907235,1.0750868,0.85934424,0.64541465,0.42967212,0.21574254,0.0,0.03988518,0.07977036,0.11965553,0.15954071,0.19942589,0.40247768,0.6055295,0.80676836,1.0098201,1.2128719,0.99531645,0.7777609,0.56020546,0.34264994,0.12509441,1.2527572,2.38042,3.5080826,4.6357455,5.7615952,6.1278133,6.492219,6.8566246,7.2228427,7.5872483,8.062244,8.537241,9.012237,9.487233,9.96223,10.319383,10.6783495,11.035503,11.392657,11.74981,14.6052265,17.460642,20.314245,23.169662,26.025078,28.042906,30.060732,32.076748,34.094574,36.1124,30.180387,24.246561,18.314548,12.382534,6.450521,6.0480433,5.6455655,5.243088,4.84061,4.4381323,2.9369993,3.0203958,3.101979,3.1853752,3.2669585,3.350355,3.3793623,3.4101827,3.43919,3.4700103,3.5008307,9.255174,15.009518,20.765673,26.520016,32.27436,32.01692,31.759478,31.502037,31.244596,30.987156,30.5176,30.048042,29.576672,29.107115,28.637556,32.06043,35.483303,38.904366,42.327236,45.75011,39.19444,32.64058,26.084906,19.529232,12.975373,11.115273,9.255174,7.3950744,5.5349746,3.6748753,3.8126602,3.9504454,4.0882306,4.2242026,4.361988,3.9595103,3.5570326,3.1545548,2.752077,2.3495996,3.2107568,4.070101,4.9294453,5.7906027,6.6499467,6.642695,6.635443,6.628191,6.6191263,6.6118746,5.8377395,5.0617914,4.2876563,3.5117085,2.7375734,4.117238,5.4969025,6.87838,8.258044,9.637709,8.419398,7.2029004,5.9845896,4.7680917,3.5497808,3.2832751,3.0149567,2.7466383,2.4801328,2.2118144,1.9199274,1.6280404,1.3343405,1.0424535,0.7505665,0.79589057,0.83940166,0.88472575,0.9300498,0.97537386,0.92823684,0.8792868,0.8321498,0.7850128,0.73787576,1.1747998,1.6117238,2.0504606,2.4873846,2.9243085,3.6966307,4.4707656,5.243088,6.01541,6.787732,7.360628,7.931711,8.504607,9.077503,9.6504,8.600695,7.549176,6.4994707,5.4497657,4.40006,4.4345064,4.4707656,4.505212,4.539658,4.5759177,4.358362,4.1408067,3.923251,3.7056956,3.48814,2.7974012,2.1066625,1.4177368,0.726998,0.038072214,0.52032024,1.0025684,1.4848163,1.9670644,2.4493124,2.857229,3.2651455,3.673062,4.079166,4.4870825,5.8431783,7.1974616,8.551744,9.907841,11.262123,10.8143215,10.368333,9.920531,9.47273,9.024928,8.073122,7.119504,6.167699,5.2140803,4.262275,3.7256382,3.1871881,2.6505513,2.1121013,1.5754645,2.1900587,2.8046532,3.4192474,4.0356545,4.650249,4.1480584,3.6458678,3.141864,2.6396735,2.137483,2.2879589,2.4366217,2.5870976,2.7375734,2.8880494,2.6958754,2.5018883,2.3097143,2.1175404,1.9253663,2.1701162,2.4148662,2.659616,2.904366,3.149116,3.0856624,3.0203958,2.955129,2.8898623,2.8245957,2.6995013,2.5744069,2.4493124,2.324218,2.1991236,2.3006494,2.4003625,2.5000753,2.5997884,2.6995013,3.5352771,4.36924,5.2050157,6.0407915,6.874754,6.87838,6.880193,6.882006,6.885632,6.887445,6.7442207,6.60281,6.4595857,6.3181744,6.1749506,8.713099,11.249433,13.7875805,16.325727,18.862062,17.714457,16.566853,15.419247,14.271642,13.125849,11.552197,9.980359,8.406708,6.834869,5.2630305,6.24203,7.2228427,8.201842,9.182655,10.161655,10.370146,10.576823,10.785315,10.991992,11.200482,10.081885,8.9651,7.8483152,6.7297173,5.612932,6.925517,8.238102,9.550687,10.863272,12.175857,13.577277,14.98051,16.38193,17.785164,19.188396,16.452635,13.716875,10.982927,8.247167,5.5132194,5.237649,4.9620786,4.688321,4.4127507,4.137181,5.1071157,6.0770507,7.0469856,8.01692,8.9868555,9.249735,9.512614,9.775495,10.038374,10.29944,10.700105,11.10077,11.499621,11.900287,12.299138,12.328146,12.35534,12.382534,12.409729,12.436923,11.209548,9.982172,8.754796,7.5274205,6.300045,5.915697,5.529536,5.145188,4.76084,4.3746786,3.738329,3.100166,2.4620032,1.8256533,1.1874905,1.0950294,1.0025684,0.9101072,0.81764615,0.72518504,1.2255627,1.7241274,2.2245052,2.7248828,3.2252605,2.7103791,2.1954978,1.6806163,1.1657349,0.6508536,0.62184614,0.5946517,0.56745726,0.5402629,0.51306844,0.8466535,1.1820517,1.5174497,1.8528478,2.1882458,2.2100015,2.231757,2.2553256,2.277081,2.3006494,1.840157,1.3796645,0.91917205,0.4604925,0.0,0.53482395,1.0696479,1.6044719,2.1392958,2.6741197,2.2571385,1.840157,1.4231756,1.0043813,0.5873999,0.69073874,0.79226464,0.89560354,0.99712944,1.1004683,1.2853905,1.4703126,1.6552348,1.840157,2.0250793,1.6352923,1.2455053,0.8557183,0.46411842,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.15591478,0.3100166,0.46411842,0.6200332,0.774135,1.0442665,1.3143979,1.5845293,1.8546607,2.124792,2.6995013,3.2742105,3.8507326,4.4254417,5.0001507,5.2557783,5.5095935,5.765221,6.0208488,6.2746634,5.090799,3.9051213,2.7194438,1.5355793,0.34990177,0.30820364,0.26469254,0.2229944,0.1794833,0.13778515,0.12690738,0.11784257,0.10696479,0.09789998,0.0870222,0.0870222,0.0870222,0.0870222,0.0870222,0.0870222,0.09427405,0.10333887,0.11059072,0.11784257,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.9808127,1.8981718,2.8155308,3.73289,4.650249,3.73289,2.8155308,1.8981718,0.9808127,0.06164073,0.054388877,0.047137026,0.03988518,0.032633327,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.5166943,1.0098201,1.502946,1.9942589,2.4873846,4.539658,6.591932,8.644206,10.698292,12.750566,12.76507,12.779573,12.79589,12.810393,12.824898,11.829581,10.834265,9.840761,8.845445,7.850128,6.947273,6.0444174,5.143375,4.2405195,3.3376641,4.9058766,6.472276,8.040489,9.606889,11.175101,11.352772,11.530442,11.708113,11.885782,12.06164,11.236742,10.411844,9.5869465,8.762048,7.93715,7.8882003,7.837437,7.7866745,7.7377243,7.686961,6.9128265,6.1368785,5.3627434,4.5867953,3.8126602,9.440096,15.067532,20.694967,26.322403,31.949839,25.820213,19.690586,13.559147,7.4295206,1.2998942,5.317419,9.334945,13.352469,17.369995,21.38752,18.184015,14.982323,11.780631,8.577126,5.375434,12.27557,19.173893,26.07584,32.974163,39.8743,33.731983,27.589664,21.447348,15.30503,9.162713,8.693155,8.221786,7.752228,7.2826705,6.813113,5.4950895,4.177066,2.8608549,1.5428312,0.22480737,0.1794833,0.13415924,0.09064813,0.045324065,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.14503701,0.16497959,0.18492219,0.20486477,0.22480737,0.23024625,0.23568514,0.23931105,0.24474995,0.25018883,0.21755551,0.18492219,0.15228885,0.11965553,0.0870222,0.24837588,0.40791658,0.56745726,0.726998,0.8883517,1.7730774,2.657803,3.5425289,4.4272547,5.3119802,5.038223,4.762653,4.4870825,4.213325,3.9377546,5.40988,6.882006,8.354132,9.82807,11.300196,11.445232,11.59027,11.735307,11.880343,12.025381,12.547514,13.069647,13.591781,14.115726,14.63786,15.825351,17.01284,18.20033,19.387821,20.575312,22.487988,24.400663,26.31334,28.224201,30.136877,30.463211,30.787731,31.112251,31.436771,31.763105,29.460642,27.15818,24.855717,22.553255,20.250792,21.004984,21.759176,22.515182,23.269375,24.025381,23.332829,22.640276,21.947725,21.255173,20.562622,18.979906,17.397188,15.814472,14.231756,12.650853,11.789696,10.930351,10.069194,9.20985,8.350506,6.965402,5.580299,4.195195,2.810092,1.4249886,1.1403534,0.8557183,0.56927025,0.28463513,0.0,0.059827764,0.11965553,0.1794833,0.23931105,0.2991388,0.5982776,0.89560354,1.1929294,1.4902552,1.7875811,1.455809,1.1222239,0.7904517,0.45686656,0.12509441,1.2726997,2.420305,3.5679104,4.7155156,5.863121,6.26016,6.6571984,7.0542374,7.453089,7.850128,8.412147,8.975978,9.537996,10.100015,10.662033,10.705544,10.747242,10.790753,10.832452,10.874149,13.419549,15.964949,18.510347,21.053934,23.599335,25.095028,26.590723,28.084604,29.580297,31.074179,26.456562,21.838947,17.223145,12.605529,7.987913,7.3406854,6.6916447,6.0444174,5.3971896,4.749962,3.1871881,3.247016,3.3068438,3.3666716,3.4283123,3.48814,3.5280252,3.5679104,3.6077955,3.6476808,3.6875658,9.501737,15.31772,21.131891,26.947876,32.762047,32.901646,33.043056,33.182655,33.32225,33.46185,32.477413,31.492973,30.506721,29.522284,28.537844,32.36682,36.197613,40.0284,43.857376,47.688168,40.760838,33.833508,26.904366,19.977036,13.049705,11.269376,9.490859,7.71053,5.9302006,4.1498713,4.12449,4.099108,4.07554,4.0501585,4.024777,3.7419548,3.4591327,3.1781235,2.8953013,2.612479,3.3304121,4.0483456,4.764466,5.482399,6.200332,5.977338,5.754343,5.5331616,5.3101673,5.087173,4.699199,4.313038,3.925064,3.53709,3.149116,4.590421,6.0299134,7.4694057,8.910711,10.3502035,8.923402,7.494787,6.0679855,4.6393714,3.2125697,2.9478772,2.6831846,2.4166791,2.1519866,1.887294,1.7096237,1.5319533,1.3542831,1.1766127,1.0007553,1.0605831,1.1204109,1.1802386,1.2400664,1.2998942,1.1820517,1.064209,0.9481794,0.83033687,0.7124943,1.2255627,1.7368182,2.2498865,2.762955,3.2742105,3.8180993,4.360175,4.902251,5.4443264,5.9882154,6.24203,6.497658,6.7532854,7.0071006,7.262728,6.6753283,6.0879283,5.5005283,4.9131284,4.325729,4.6792564,5.034597,5.389938,5.7452784,6.1006193,5.810545,5.520471,5.230397,4.940323,4.650249,3.729264,2.810092,1.889107,0.969935,0.05076295,0.28463513,0.52032024,0.7541924,0.9898776,1.2255627,1.7730774,2.3205922,2.8681068,3.4156215,3.9631362,5.803293,7.6416373,9.481794,11.321951,13.162108,12.444175,11.728055,11.010121,10.292189,9.574255,8.4683485,7.360628,6.2529078,5.145188,4.0374675,3.4627585,2.8880494,2.3133402,1.7368182,1.162109,1.7331922,2.3024626,2.8717327,3.442816,4.0120864,3.6041696,3.198066,2.7901495,2.382233,1.9743162,2.1121013,2.2498865,2.3876717,2.525457,2.663242,2.5599031,2.4583774,2.3550384,2.2516994,2.1501737,2.3858588,2.619731,2.855416,3.0892882,3.3249733,3.24339,3.159994,3.0765975,2.9950142,2.911618,2.7248828,2.5381477,2.3495996,2.1628644,1.9743162,2.0994108,2.2245052,2.3495996,2.474694,2.5997884,3.2180085,3.834416,4.4526362,5.0708566,5.6872635,5.8957543,6.1024323,6.3091097,6.5176005,6.7242785,6.697084,6.6698895,6.642695,6.6155005,6.588306,8.749357,10.912222,13.075087,15.23795,17.400814,16.358362,15.3159075,14.271642,13.229188,12.186734,10.645717,9.102885,7.560054,6.017223,4.4743915,5.7779117,7.079619,8.383139,9.684846,10.988366,10.93579,10.883214,10.830639,10.778063,10.725487,9.460039,8.194591,6.929143,5.6655083,4.40006,5.638314,6.874754,8.113008,9.349448,10.587702,12.195799,13.802084,15.410182,17.01828,18.624565,16.032028,13.439491,10.846955,8.254418,5.661882,5.186886,4.7118897,4.2368937,3.7618973,3.2869012,4.059223,4.8333583,5.6056805,6.378002,7.1503243,8.225411,9.300498,10.375585,11.450671,12.525759,12.799516,13.075087,13.3506565,13.6244135,13.899984,13.608097,13.314397,13.022511,12.730623,12.436923,11.405348,10.371959,9.340384,8.306994,7.2754188,6.7079616,6.1405044,5.573047,5.0055895,4.4381323,3.825351,3.2125697,2.5997884,1.987007,1.3742256,1.2473183,1.1204109,0.9916905,0.86478317,0.73787576,1.1131591,1.4866294,1.8619126,2.2371957,2.612479,2.2172532,1.8220274,1.4268016,1.0333886,0.63816285,0.6417888,0.64722764,0.6526665,0.65810543,0.66173136,0.8557183,1.0478923,1.2400664,1.4322405,1.6244144,1.79302,1.9598125,2.126605,2.2952106,2.4620032,1.9706904,1.4775645,0.98443866,0.49312583,0.0,0.58014804,1.1602961,1.7404441,2.3205922,2.9007401,2.3858588,1.8691645,1.3542831,0.83940166,0.3245203,0.36984438,0.41516843,0.4604925,0.5058166,0.5493277,0.9808127,1.4104849,1.840157,2.269829,2.6995013,2.1683033,1.6352923,1.1022812,0.56927025,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.07795739,0.15410182,0.23205921,0.3100166,0.387974,0.72337204,1.0569572,1.3923552,1.7277533,2.0631514,2.5508385,3.0367124,3.5243993,4.0120864,4.499773,5.0781083,5.65463,6.2329655,6.8094873,7.3878226,5.957395,4.5269675,3.0983531,1.6679256,0.2374981,0.2229944,0.20667773,0.19217403,0.17767033,0.16316663,0.14503701,0.12690738,0.11059072,0.092461094,0.07433146,0.07433146,0.07433146,0.07433146,0.07433146,0.07433146,0.08520924,0.09427405,0.10515183,0.11421664,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,1.1530442,2.2426348,3.3322253,4.421816,5.5132194,4.421816,3.3322253,2.2426348,1.1530442,0.06164073,0.052575916,0.04169814,0.032633327,0.02175555,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.27738327,0.5420758,0.80676836,1.0732739,1.3379664,3.4319382,5.527723,7.6216946,9.71748,11.813264,12.658105,13.502945,14.347786,15.192626,16.037468,14.353225,12.66717,10.982927,9.296872,7.61263,6.9545245,6.298232,5.6401267,4.9820213,4.325729,6.1767635,8.029612,9.882459,11.735307,13.588155,13.544643,13.502945,13.4594345,13.417736,13.374225,12.387974,11.399909,10.411844,9.425592,8.437528,8.350506,8.26167,8.174648,8.087626,8.000604,7.2373466,6.4759026,5.712645,4.949388,4.1879435,9.695724,15.201692,20.70947,26.217253,31.725033,25.510197,19.29536,13.080525,6.8656893,0.6508536,4.215138,7.7794223,11.34552,14.909804,18.475903,16.18069,13.885481,11.59027,9.295059,6.9998484,11.42529,15.850732,20.27436,24.699802,29.125244,25.522888,21.92053,18.318174,14.715817,11.111648,10.277685,9.441909,8.607946,7.7721705,6.9382076,5.573047,4.207886,2.8427253,1.4775645,0.11240368,0.09064813,0.06707962,0.045324065,0.02175555,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.14684997,0.17041849,0.19217403,0.21574254,0.2374981,0.23931105,0.24293698,0.24474995,0.24837588,0.25018883,0.21574254,0.1794833,0.14503701,0.11059072,0.07433146,0.291887,0.5094425,0.726998,0.9445535,1.162109,2.3296568,3.4972048,4.664753,5.8323007,6.9998484,6.0244746,5.050914,4.07554,3.100166,2.124792,3.1182957,4.1099863,5.101677,6.09518,7.0868707,8.02236,8.957849,9.893337,10.827013,11.762501,13.1059065,14.447499,15.790904,17.132496,18.474089,19.525606,20.575312,21.625017,22.674723,23.724428,25.299892,26.875357,28.45082,30.024473,31.599937,31.137632,30.675327,30.213022,29.750715,29.28841,26.654177,24.021753,21.389332,18.75691,16.124489,17.17782,18.22934,19.282671,20.334188,21.38752,21.510801,21.632269,21.75555,21.87702,22.000301,20.064056,18.129625,16.195194,14.260764,12.32452,11.470614,10.614896,9.759177,8.9052725,8.049554,6.794984,5.540414,4.2858434,3.0294604,1.7748904,1.4195497,1.064209,0.7106813,0.35534066,0.0,0.07977036,0.15954071,0.23931105,0.3208944,0.40066472,0.79226464,1.1856775,1.5772774,1.9706904,2.3622901,1.9144884,1.4666867,1.020698,0.5728962,0.12509441,1.2926424,2.4601903,3.6277382,4.795286,5.962834,6.392506,6.8221784,7.25185,7.6833353,8.113008,8.762048,9.412902,10.061942,10.712796,11.361836,11.089892,10.817947,10.54419,10.272246,10.000301,12.235684,14.471067,16.704638,18.94002,21.175404,22.14715,23.120712,24.09246,25.064207,26.03777,22.73455,19.431334,16.129929,12.828524,9.525306,8.6333275,7.7395372,6.8475595,5.955582,5.0617914,3.437377,3.4754493,3.5117085,3.5497808,3.587853,3.6241121,3.6748753,3.7256382,3.774588,3.825351,3.874301,9.750113,15.624111,21.499924,27.375734,33.249733,33.788185,34.32482,34.86327,35.399906,35.93836,34.437225,32.937904,31.436771,29.93745,28.438131,32.675026,36.91192,41.150623,45.38752,49.624413,42.325424,35.024624,27.725637,20.424837,13.125849,11.42529,9.724731,8.024173,6.3254266,4.6248674,4.4381323,4.249584,4.062849,3.874301,3.6875658,3.5243993,3.3630457,3.199879,3.0367124,2.8753586,3.4500678,4.024777,4.599486,5.1741953,5.750717,5.3119802,4.8750563,4.4381323,3.9993954,3.5624714,3.5624714,3.5624714,3.5624714,3.5624714,3.5624714,5.0617914,6.5629244,8.062244,9.563377,11.062697,9.425592,7.7866745,6.149569,4.512464,2.8753586,2.612479,2.3495996,2.08672,1.8256533,1.5627737,1.49932,1.4376793,1.3742256,1.3125849,1.2491312,1.3252757,1.3996071,1.4757515,1.550083,1.6244144,1.4376793,1.2491312,1.062396,0.87566096,0.6871128,1.2745126,1.8619126,2.4493124,3.0367124,3.6241121,3.9377546,4.249584,4.5632267,4.8750563,5.186886,5.125245,5.0617914,5.0001507,4.936697,4.8750563,4.749962,4.6248674,4.499773,4.3746786,4.249584,4.9258194,5.600241,6.2746634,6.9508986,7.6253204,7.262728,6.9001355,6.5375433,6.1749506,5.812358,4.6629395,3.5117085,2.3622901,1.2128719,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.6871128,1.3742256,2.0631514,2.7502642,3.437377,5.7615952,8.087626,10.411844,12.737875,15.062093,14.075842,13.087777,12.099712,11.111648,10.125396,8.861761,7.5999393,6.338117,5.0744824,3.8126602,3.199879,2.5870976,1.9743162,1.3633479,0.7505665,1.2745126,1.8002719,2.324218,2.8499773,3.3757362,3.0620937,2.7502642,2.4366217,2.124792,1.8129625,1.938057,2.0631514,2.1882458,2.3133402,2.4366217,2.4257438,2.4130533,2.4003625,2.3876717,2.374981,2.5997884,2.8245957,3.049403,3.2742105,3.5008307,3.3993049,3.299592,3.199879,3.100166,3.000453,2.7502642,2.5000753,2.2498865,1.9996977,1.7495089,1.8999848,2.0504606,2.1991236,2.3495996,2.5000753,2.9007401,3.299592,3.7002566,4.099108,4.499773,4.9131284,5.3246713,5.7380266,6.149569,6.5629244,6.6499467,6.736969,6.825804,6.9128265,6.9998484,8.78743,10.57501,12.362592,14.150173,15.937754,15.000452,14.06315,13.125849,12.186734,11.249433,9.737422,8.225411,6.7115874,5.199577,3.6875658,5.3119802,6.9382076,8.562622,10.1870365,11.813264,11.499621,11.187792,10.874149,10.56232,10.25049,8.838193,7.4258947,6.011784,4.599486,3.1871881,4.349297,5.5132194,6.6753283,7.837437,8.999546,10.812509,12.625471,14.438434,16.249584,18.062546,15.613234,13.162108,10.712796,8.26167,5.812358,5.137936,4.461701,3.787279,3.1128569,2.4366217,3.0131438,3.587853,4.162562,4.7372713,5.3119802,7.1992745,9.086569,10.975676,12.862969,14.750263,14.90074,15.049402,15.199879,15.350354,15.50083,14.888049,14.275268,13.662486,13.049705,12.436923,11.599335,10.761745,9.924157,9.088382,8.2507925,7.500226,6.7496595,5.999093,5.2503395,4.499773,3.9123733,3.3249733,2.7375734,2.1501737,1.5627737,1.3996071,1.2382535,1.0750868,0.9119202,0.7505665,1.0007553,1.2491312,1.49932,1.7495089,1.9996977,1.7241274,1.4503701,1.1747998,0.89922947,0.62547207,0.66173136,0.69980353,0.73787576,0.774135,0.8122072,0.8629702,0.9119202,0.96268314,1.0116332,1.062396,1.3742256,1.6878681,1.9996977,2.3133402,2.6251698,2.0994108,1.5754645,1.0497054,0.52575916,0.0,0.62547207,1.2491312,1.8746033,2.5000753,3.1255474,2.5127661,1.8999848,1.2872034,0.6744221,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.6744221,1.3506571,2.0250793,2.6995013,3.3757362,2.6995013,2.0250793,1.3506571,0.6744221,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.40066472,0.7995165,1.2001812,1.6008459,1.9996977,2.4003625,2.7992141,3.199879,3.6005437,3.9993954,4.900438,5.7996674,6.70071,7.5999393,8.499168,6.825804,5.1506267,3.4754493,1.8002719,0.12509441,0.13778515,0.15047589,0.16316663,0.17585737,0.18673515,0.16316663,0.13778515,0.11240368,0.0870222,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,1.3252757,2.5870976,3.8507326,5.1125546,6.3743763,5.1125546,3.8507326,2.5870976,1.3252757,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,2.326031,4.461701,6.599184,8.736667,10.874149,12.549327,14.224504,15.899682,17.57486,19.250036,16.875055,14.500074,12.125093,9.750113,7.3751316,6.9617763,6.550234,6.1368785,5.7253356,5.3119802,7.4494634,9.5869465,11.724429,13.861912,15.999394,15.738328,15.475449,15.212569,14.94969,14.68681,13.537392,12.387974,11.236742,10.087324,8.937905,8.812811,8.6877165,8.562622,8.437528,8.312433,7.5618668,6.813113,6.0625467,5.3119802,4.5632267,9.949538,15.337664,20.725788,26.1121,31.500225,25.20018,18.900135,12.60009,6.300045,0.0,3.1128569,6.2257137,9.336758,12.449615,15.56247,14.175554,12.786825,11.399909,10.012992,8.624263,10.57501,12.525759,14.474693,16.425442,18.374376,17.31198,16.249584,15.187187,14.124791,13.062395,11.862214,10.662033,9.461852,8.26167,7.063302,5.6491914,4.2368937,2.8245957,1.4122978,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.15047589,0.17585737,0.19942589,0.22480737,0.25018883,0.25018883,0.25018883,0.25018883,0.25018883,0.25018883,0.21211663,0.17585737,0.13778515,0.099712946,0.06164073,0.33721104,0.61278135,0.8883517,1.162109,1.4376793,2.8880494,4.3366065,5.7869763,7.2373466,8.6877165,7.0125394,5.337362,3.6621845,1.987007,0.31182957,0.824898,1.3379664,1.8492218,2.3622901,2.8753586,4.599486,6.3254266,8.049554,9.775495,11.499621,13.662486,15.825351,17.988214,20.149265,22.31213,23.225864,24.137783,25.049704,25.961624,26.875357,28.111797,29.350052,30.588305,31.824745,33.063,31.812054,30.562923,29.31198,28.062847,26.811903,23.849524,20.887142,17.92476,14.96238,11.999999,13.3506565,14.699501,16.050158,17.400814,18.749659,19.68696,20.624262,21.563377,22.500679,23.43798,21.15002,18.862062,16.574104,14.287958,11.999999,11.14972,10.29944,9.449161,8.600695,7.750415,6.624565,5.5005283,4.3746786,3.2506418,2.124792,1.7005589,1.2745126,0.85027945,0.42423326,0.0,0.099712946,0.19942589,0.2991388,0.40066472,0.50037766,0.9880646,1.4757515,1.9616255,2.4493124,2.9369993,2.374981,1.8129625,1.2491312,0.6871128,0.12509441,1.3125849,2.5000753,3.6875658,4.8750563,6.0625467,6.5248523,6.987158,7.4494634,7.911769,8.375887,9.11195,9.849826,10.587702,11.325577,12.06164,11.47424,10.88684,10.29944,9.712041,9.12464,11.050007,12.975373,14.90074,16.824293,18.749659,19.199274,19.650702,20.100317,20.54993,20.999546,19.012539,17.025532,15.036712,13.049705,11.062697,9.924157,8.78743,7.650702,6.5121617,5.375434,3.299592,3.3449159,3.39024,3.435564,3.4808881,3.5243993,3.6531196,3.780027,3.9069343,4.0356545,4.162562,9.3150015,14.467442,19.61988,24.77232,29.92476,30.958149,31.989725,33.023113,34.054688,35.088078,33.98942,32.892582,31.795738,30.697083,29.60024,32.87989,36.15954,39.441,42.72065,46.0003,39.395676,32.791054,26.184618,19.579996,12.975373,11.289318,9.605076,7.9208336,6.2347784,4.550536,4.690134,4.8297324,4.9693303,5.1107416,5.2503395,5.2594047,5.2702823,5.279347,5.290225,5.2992897,5.67276,6.0444174,6.4178877,6.789545,7.1630154,6.495845,5.826862,5.1596913,4.4925213,3.825351,4.1317415,4.439945,4.748149,5.0545397,5.3627434,6.526665,7.6924005,8.858135,10.022058,11.187792,9.597824,8.007855,6.4178877,4.8279195,3.2379513,3.4083695,3.576975,3.7473936,3.917812,4.0882306,3.8942437,3.7020695,3.5098956,3.3177216,3.1255474,2.8445382,2.565342,2.2843328,2.0051367,1.7241274,1.5192627,1.3143979,1.1095331,0.90466833,0.69980353,1.2726997,1.845596,2.4166791,2.9895754,3.5624714,3.870675,4.177066,4.4852695,4.7916603,5.0998635,5.0219064,4.945762,4.8678045,4.7898474,4.7118897,4.5831695,4.4526362,4.322103,4.1933823,4.062849,4.572292,5.081734,5.5929894,6.1024323,6.6118746,6.2782893,5.942891,5.6074934,5.272095,4.936697,4.022964,3.1074178,2.1918716,1.2781386,0.36259252,0.31182957,0.26287958,0.21211663,0.16316663,0.11240368,0.6399758,1.167548,1.69512,2.222692,2.7502642,4.6375585,6.5248523,8.412147,10.29944,12.186734,11.612025,11.037316,10.462607,9.8878975,9.313189,8.232663,7.1521373,6.071612,4.992899,3.9123733,3.4283123,2.9424384,2.4583774,1.9725033,1.4866294,1.8746033,2.2625773,2.6505513,3.0367124,3.4246864,3.1255474,2.8245957,2.525457,2.2245052,1.9253663,2.0450218,2.1646774,2.2843328,2.4058013,2.525457,2.565342,2.6052272,2.6451125,2.6849976,2.7248828,2.9895754,3.254268,3.5207734,3.785466,4.0501585,3.8054085,3.5606585,3.3140955,3.0693457,2.8245957,2.6396735,2.4547513,2.269829,2.084907,1.8999848,2.0975976,2.2952106,2.4928236,2.6904364,2.8880494,3.198066,3.5080826,3.8180993,4.1281157,4.4381323,4.896812,5.3573046,5.8177967,6.2782893,6.736969,6.697084,6.6571984,6.6173134,6.5774283,6.5375433,8.073122,9.606889,11.142468,12.678047,14.211814,14.112101,14.012388,13.912675,13.812962,13.713249,12.179482,10.64753,9.115576,7.5818095,6.049856,7.3551893,8.660522,9.965856,11.269376,12.574709,12.344462,12.114216,11.885782,11.655537,11.42529,9.91328,8.399456,6.887445,5.375434,3.8616104,4.550536,5.237649,5.924762,6.6118746,7.3008003,9.296872,11.294757,13.292642,15.290526,17.286598,15.107417,12.928236,10.747242,8.568061,6.3870673,5.5349746,4.6828823,3.83079,2.9768846,2.124792,3.4700103,4.8152285,6.1604466,7.5056653,8.8508835,9.7229185,10.594954,11.466989,12.340837,13.212872,13.867351,14.521831,15.1781225,15.8326025,16.487082,16.526966,16.566853,16.606737,16.646622,16.68832,14.732134,12.7777605,10.821573,8.8672,6.9128265,6.2674117,5.621997,4.976582,4.3329806,3.6875658,3.2578938,2.8282216,2.3967366,1.9670644,1.5373923,1.3996071,1.261822,1.1258497,0.9880646,0.85027945,1.0297627,1.209246,1.3905423,1.5700256,1.7495089,1.504759,1.260009,1.015259,0.7705091,0.52575916,0.56745726,0.6091554,0.6526665,0.69436467,0.73787576,0.75963134,0.78319985,0.80495536,0.82671094,0.85027945,1.1095331,1.3705997,1.6298534,1.889107,2.1501737,2.030518,1.9108626,1.789394,1.6697385,1.550083,1.7857682,2.0196402,2.2553256,2.4891977,2.7248828,2.2045624,1.6842422,1.1657349,0.64541465,0.12509441,0.10696479,0.09064813,0.072518505,0.054388877,0.038072214,0.56927025,1.1022812,1.6352923,2.1683033,2.6995013,2.1592383,1.6207886,1.0805258,0.5402629,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.4169814,0.83577573,1.2527572,1.6697385,2.08672,2.3097143,2.5327086,2.7557032,2.9768846,3.199879,3.923251,4.64481,5.368182,6.089741,6.813113,5.5494785,4.2876563,3.0258346,1.7621996,0.50037766,0.44236287,0.38434806,0.32814622,0.27013144,0.21211663,0.19217403,0.17223145,0.15228885,0.13234627,0.11240368,0.10333887,0.092461094,0.08339628,0.072518505,0.06164073,0.072518505,0.08339628,0.092461094,0.10333887,0.11240368,0.10333887,0.092461094,0.08339628,0.072518505,0.06164073,0.072518505,0.08339628,0.092461094,0.10333887,0.11240368,1.4630609,2.811905,4.162562,5.5132194,6.8620634,5.5005283,4.137181,2.7756457,1.4122978,0.05076295,0.04169814,0.034446288,0.027194439,0.01994259,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.16679256,0.33539808,0.50219065,0.67079616,0.8375887,2.8282216,4.8170414,6.8076744,8.798307,10.7871275,12.32452,13.861912,15.399304,16.936697,18.475903,16.545097,14.614291,12.685299,10.754494,8.825501,8.1819,7.5401115,6.8983226,6.2547207,5.612932,7.36788,9.122828,10.877775,12.632723,14.387671,14.217253,14.046834,13.878228,13.70781,13.537392,12.32452,11.111648,9.900589,8.6877165,7.474845,7.4893484,7.5056653,7.520169,7.5346723,7.549176,6.8221784,6.09518,5.368182,4.6393714,3.9123733,9.130079,14.347786,19.565493,24.7832,29.999092,24.00725,18.01541,12.021755,6.0299134,0.038072214,2.8372865,5.638314,8.437528,11.236742,14.037769,12.804955,11.57214,10.339326,9.108324,7.8755093,9.244296,10.614896,11.985496,13.354282,14.724882,14.0323305,13.339779,12.647227,11.954676,11.262123,10.352016,9.441909,8.531802,7.6216946,6.7134004,5.369995,4.028403,2.6849976,1.3415923,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.02175555,0.032633327,0.04169814,0.052575916,0.06164073,0.08339628,0.10333887,0.12328146,0.14322405,0.16316663,0.18673515,0.21211663,0.2374981,0.26287958,0.28826106,0.2755703,0.26287958,0.25018883,0.2374981,0.22480737,0.24474995,0.26469254,0.28463513,0.3045777,0.3245203,0.59283876,0.85934424,1.1276628,1.3941683,1.6624867,2.7248828,3.787279,4.8496747,5.9120708,6.9744673,5.6292486,4.2858434,2.9406252,1.5954071,0.25018883,1.4703126,2.6904364,3.9105604,5.130684,6.350808,8.080374,9.80994,11.539507,13.2690735,15.000452,16.189756,17.380873,18.570175,19.75948,20.950596,21.759176,22.56957,23.379965,24.19036,25.000753,26.309713,27.620485,28.929443,30.240215,31.549175,30.457771,29.364555,28.273151,27.179935,26.08672,23.285692,20.482851,17.680012,14.877171,12.07433,13.702372,15.330412,16.958452,18.584679,20.212719,21.450974,22.687414,23.925667,25.162107,26.400362,24.279196,22.159842,20.04049,17.919323,15.799969,14.29521,12.790451,11.285692,9.780933,8.274362,7.0705543,5.864934,4.6593137,3.4555066,2.2498865,2.322405,2.3949237,2.467442,2.5399606,2.612479,2.665055,2.7176309,2.770207,2.8227828,2.8753586,3.303218,3.729264,4.157123,4.5849824,5.0128417,5.0074024,5.0019636,4.9983377,4.992899,4.98746,5.6818247,6.378002,7.072367,7.7667317,8.46291,8.471974,8.482852,8.491917,8.502794,8.511859,9.104698,9.697536,10.290376,10.883214,11.47424,10.9230995,10.370146,9.817192,9.264238,8.713099,10.5695715,12.427858,14.284332,16.142618,17.999092,18.537542,19.074179,19.612629,20.149265,20.687716,18.671701,16.6575,14.643299,12.627284,10.613083,9.38752,8.161958,6.9382076,5.712645,4.4870825,3.1618068,3.2143826,3.2669585,3.3195345,3.3721104,3.4246864,3.6295512,3.834416,4.0392804,4.2441454,4.4508233,8.87989,13.308958,17.73984,22.17072,26.599787,28.128115,29.654629,31.182957,32.709473,34.237797,33.541622,32.847256,32.152893,31.456715,30.762348,33.084755,35.407158,37.729565,40.051968,42.374374,36.46593,30.555672,24.645412,18.735155,12.824898,11.155159,9.48542,7.8156815,6.14413,4.4743915,4.942136,5.40988,5.8776245,6.345369,6.813113,6.9944096,7.177519,7.360628,7.5419245,7.7250338,7.895452,8.06587,8.234476,8.404895,8.575313,7.6778965,6.78048,5.883064,4.985647,4.0882306,4.702825,5.317419,5.9320135,6.548421,7.1630154,7.993352,8.821876,9.652213,10.48255,11.312886,9.770056,8.227224,6.684393,5.143375,3.6005437,4.2024474,4.804351,5.408067,6.009971,6.6118746,6.2891674,5.9682727,5.6455655,5.3228583,5.0001507,4.365614,3.729264,3.094727,2.4601903,1.8256533,1.6026589,1.3796645,1.1566701,0.9354887,0.7124943,1.2708868,1.8274662,2.3858588,2.9424384,3.5008307,3.8017826,4.1045475,4.407312,4.710077,5.0128417,4.9203806,4.8279195,4.7354584,4.6429973,4.550536,4.4145637,4.2804046,4.1444325,4.0102735,3.874301,4.220577,4.5650396,4.9095025,5.2557783,5.600241,5.292038,4.985647,4.6774435,4.36924,4.062849,3.3829882,2.7031271,2.0232663,1.3415923,0.66173136,0.5747091,0.48768693,0.40066472,0.31182957,0.22480737,0.59283876,0.96087015,1.3270886,1.69512,2.0631514,3.5117085,4.9620786,6.412449,7.8628187,9.313189,9.1500225,8.9868555,8.825501,8.662335,8.499168,7.6017523,6.7043357,5.806919,4.9095025,4.0120864,3.6549325,3.2977788,2.9406252,2.5816586,2.2245052,2.474694,2.7248828,2.9750717,3.2252605,3.4754493,3.1871881,2.9007401,2.612479,2.324218,2.03777,2.1519866,2.268016,2.382233,2.4982624,2.612479,2.70494,2.7974012,2.8898623,2.9823234,3.0747845,3.3793623,3.6857529,3.9903307,4.2949085,4.599486,4.209699,3.8199122,3.4301252,3.0403383,2.6505513,2.5308957,2.4094272,2.2897718,2.1701162,2.0504606,2.2952106,2.5399606,2.7847104,3.0294604,3.2742105,3.4953918,3.7147603,3.9341288,4.15531,4.3746786,4.882308,5.389938,5.8975673,6.4051967,6.9128265,6.7442207,6.5774283,6.4106355,6.24203,6.0752378,7.3570023,8.640579,9.922344,11.204109,12.487686,13.225562,13.961625,14.699501,15.437376,16.175253,14.623356,13.069647,11.517752,9.965856,8.412147,9.398398,10.382836,11.367275,12.351714,13.337966,13.189302,13.042453,12.895603,12.74694,12.60009,10.988366,9.374829,7.763106,6.149569,4.537845,4.749962,4.9620786,5.1741953,5.388125,5.600241,7.783048,9.964043,12.14685,14.329657,16.512463,14.603414,12.692551,10.781689,8.872639,6.9617763,5.9320135,4.902251,3.872488,2.8427253,1.8129625,3.926877,6.0426044,8.158332,10.272246,12.387974,12.244749,12.103338,11.9601145,11.81689,11.675479,12.835775,13.994258,15.154554,16.31485,17.475147,18.167698,18.86025,19.552801,20.245354,20.937904,17.864933,14.791962,11.720803,8.647832,5.57486,5.034597,4.494334,3.9540713,3.4156215,2.8753586,2.6016014,2.3296568,2.0577126,1.7857682,1.5120108,1.3996071,1.2872034,1.1747998,1.062396,0.9499924,1.0605831,1.1693609,1.2799516,1.3905423,1.49932,1.2853905,1.0696479,0.8557183,0.6399758,0.42423326,0.47318324,0.52032024,0.56745726,0.61459434,0.66173136,0.65810543,0.6526665,0.64722764,0.6417888,0.63816285,0.8448406,1.0533313,1.260009,1.4666867,1.6751775,1.9598125,2.2444477,2.5308957,2.8155308,3.100166,2.9442513,2.7901495,2.6342347,2.4801328,2.324218,1.8981718,1.4703126,1.0424535,0.61459434,0.18673515,0.16497959,0.14322405,0.11965553,0.09789998,0.07433146,0.46411842,0.8557183,1.2455053,1.6352923,2.0250793,1.6207886,1.214685,0.8103943,0.40429065,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.43511102,0.87022203,1.305333,1.7404441,2.175555,2.220879,2.2643902,2.3097143,2.3550384,2.4003625,2.9442513,3.489953,4.0356545,4.5795436,5.125245,4.274966,3.4246864,2.5744069,1.7241274,0.87566096,0.7469406,0.6200332,0.49312583,0.36440548,0.2374981,0.2229944,0.20667773,0.19217403,0.17767033,0.16316663,0.14322405,0.12328146,0.10333887,0.08339628,0.06164073,0.07070554,0.07795739,0.08520924,0.092461094,0.099712946,0.092461094,0.08520924,0.07795739,0.07070554,0.06164073,0.08339628,0.10333887,0.12328146,0.14322405,0.16316663,1.6008459,3.0367124,4.4743915,5.9120708,7.3497505,5.8866897,4.4254417,2.962381,1.49932,0.038072214,0.034446288,0.032633327,0.030820364,0.027194439,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.29732585,0.5946517,0.8919776,1.1893034,1.4866294,3.3304121,5.1723824,7.0143523,8.858135,10.700105,12.099712,13.499319,14.90074,16.300346,17.699953,16.215137,14.730321,13.245504,11.760688,10.275872,9.402024,8.529989,7.6579537,6.784106,5.9120708,7.2844834,8.656897,10.029309,11.401722,12.774135,12.697989,12.620032,12.542075,12.464118,12.387974,11.111648,9.837135,8.562622,7.28811,6.011784,6.167699,6.3218007,6.4777155,6.6318173,6.787732,6.0824895,5.377247,4.6720047,3.966762,3.2633326,8.31062,13.357908,18.405195,23.452484,28.499771,22.814322,17.130684,11.445232,5.7597823,0.07433146,2.563529,5.049101,7.5382986,10.025683,12.513068,11.434355,10.357455,9.280556,8.201842,7.124943,7.915395,8.705847,9.494485,10.284937,11.075388,10.752681,10.429974,10.107266,9.784559,9.461852,8.841819,8.221786,7.6017523,6.981719,6.3616858,5.090799,3.8180993,2.5453994,1.2726997,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.032633327,0.03988518,0.047137026,0.054388877,0.06164073,0.09064813,0.11784257,0.14503701,0.17223145,0.19942589,0.22480737,0.25018883,0.2755703,0.2991388,0.3245203,0.2991388,0.2755703,0.25018883,0.22480737,0.19942589,0.27738327,0.35534066,0.43329805,0.5094425,0.5873999,0.8466535,1.1077201,1.3669738,1.6280404,1.887294,2.561716,3.2379513,3.9123733,4.5867953,5.2630305,4.2477713,3.2325122,2.2172532,1.2019942,0.18673515,2.1157274,4.0429068,5.9700856,7.897265,9.824444,11.559449,13.294455,15.02946,16.764465,18.49947,18.717026,18.934582,19.152136,19.369692,19.587248,20.294304,21.003172,21.710226,22.417282,23.124338,24.507627,25.889105,27.272396,28.655687,30.037165,29.101675,28.168,27.232512,26.297022,25.363346,22.720047,20.076748,17.43526,14.791962,12.1504755,14.055899,15.95951,17.864933,19.770357,21.675781,23.213173,24.750565,26.287958,27.82535,29.362741,27.410181,25.45762,23.50506,21.5525,19.59994,17.4407,15.279649,13.12041,10.959359,8.80012,7.51473,6.2293396,4.945762,3.6603715,2.374981,2.9442513,3.5153344,4.0846047,4.655688,5.224958,5.230397,5.235836,5.239462,5.2449007,5.2503395,5.618371,5.9845896,6.352621,6.720652,7.0868707,7.6398244,8.192778,8.745731,9.296872,9.849826,10.052877,10.255929,10.457169,10.66022,10.863272,10.419096,9.976733,9.53437,9.092008,8.649645,9.097446,9.545248,9.99305,10.440851,10.88684,10.370146,9.851639,9.334945,8.81825,8.299743,10.09095,11.880343,13.669738,15.459132,17.25034,17.87581,18.49947,19.124943,19.750414,20.375887,18.332678,16.289469,14.248073,12.2048645,10.161655,8.849071,7.5364857,6.2257137,4.9131284,3.6005437,3.0258346,3.0856624,3.1454902,3.2053177,3.2651455,3.3249733,3.6077955,3.8906176,4.171627,4.454449,4.7372713,8.444779,12.152288,15.859797,19.567305,23.274813,25.29808,27.319532,29.3428,31.364252,33.38752,33.09563,32.801933,32.510044,32.21816,31.924458,33.28962,34.65478,36.01994,37.3851,38.750263,33.53437,28.320288,23.104395,17.890314,12.674421,11.019187,9.365765,7.71053,6.055295,4.40006,5.1941376,5.9900284,6.7859187,7.5799966,8.375887,8.729415,9.084756,9.440096,9.795437,10.150778,10.118144,10.085511,10.052877,10.020245,9.987611,8.859948,7.7322855,6.604623,5.47696,4.349297,5.272095,6.1948934,7.117691,8.040489,8.963287,9.458226,9.953164,10.448103,10.943042,11.437981,9.9422865,8.448405,6.9527116,5.4570174,3.9631362,4.9983377,6.0317264,7.066928,8.10213,9.137331,8.685904,8.232663,7.7794223,7.327995,6.874754,5.8848767,4.894999,3.9051213,2.9152439,1.9253663,1.6842422,1.4449311,1.2056202,0.9644961,0.72518504,1.2672608,1.8093367,2.3532255,2.8953013,3.437377,3.7347028,4.0320287,4.329355,4.6266804,4.9258194,4.8170414,4.710077,4.603112,4.494334,4.3873696,4.2477713,4.1081734,3.966762,3.827164,3.6875658,3.8670492,4.0483456,4.227829,4.407312,4.5867953,4.307599,4.028403,3.7473936,3.4681973,3.1871881,2.7430124,2.2970235,1.8528478,1.4068589,0.96268314,0.8375887,0.7124943,0.5873999,0.46230546,0.33721104,0.54570174,0.7523795,0.96087015,1.167548,1.3742256,2.3876717,3.3993049,4.4127507,5.424384,6.43783,6.688019,6.9382076,7.1865835,7.4367723,7.686961,6.972654,6.258347,5.542227,4.8279195,4.1117992,3.8833659,3.6531196,3.4228733,3.1926272,2.962381,3.0747845,3.1871881,3.299592,3.4119956,3.5243993,3.2506418,2.9750717,2.6995013,2.4257438,2.1501737,2.2607644,2.3695421,2.4801328,2.5907235,2.6995013,2.8445382,2.9895754,3.1346123,3.2796493,3.4246864,3.7691493,4.115425,4.459888,4.804351,5.1506267,4.615803,4.079166,3.5443418,3.009518,2.474694,2.420305,2.3641033,2.3097143,2.2553256,2.1991236,2.4928236,2.7847104,3.0784104,3.3702974,3.6621845,3.7927177,3.923251,4.0519714,4.1825047,4.313038,4.8678045,5.422571,5.977338,6.532104,7.0868707,6.793171,6.497658,6.202145,5.906632,5.612932,6.642695,7.6724577,8.70222,9.731983,10.761745,12.337211,13.912675,15.488139,17.06179,18.637255,17.065416,15.491765,13.919927,12.348088,10.774437,11.439794,12.105151,12.770509,13.435865,14.09941,14.034143,13.97069,13.905423,13.840157,13.77489,12.06164,10.3502035,8.636953,6.925517,5.2122674,4.949388,4.688321,4.4254417,4.162562,3.8996825,6.2674117,8.63514,11.00287,13.370599,15.738328,14.097597,12.456866,10.817947,9.177217,7.5382986,6.3308654,5.123432,3.9141862,2.7067533,1.49932,4.3855567,7.26998,10.154404,13.04064,15.925063,14.7683935,13.60991,12.45324,11.294757,10.138086,11.802386,13.466686,15.132799,16.797098,18.463211,19.806616,21.151834,22.497053,23.842272,25.187489,20.997732,16.807976,12.618219,8.42665,4.2368937,3.8017826,3.3666716,2.9333735,2.4982624,2.0631514,1.9471219,1.8329052,1.7168756,1.6026589,1.4866294,1.3996071,1.3125849,1.2255627,1.1367276,1.0497054,1.0895905,1.1294757,1.1693609,1.209246,1.2491312,1.064209,0.8792868,0.69436467,0.5094425,0.3245203,0.3770962,0.42967212,0.48224804,0.53482395,0.5873999,0.55476654,0.52213323,0.4894999,0.45686656,0.42423326,0.58014804,0.73424983,0.8901646,1.0442665,1.2001812,1.8909199,2.5798457,3.2705846,3.9595103,4.650249,4.1045475,3.5606585,3.0149567,2.469255,1.9253663,1.5899682,1.2545701,0.91917205,0.5855869,0.25018883,0.2229944,0.19579996,0.16679256,0.13959812,0.11240368,0.36077955,0.6073425,0.8557183,1.1022812,1.3506571,1.0805258,0.8103943,0.5402629,0.27013144,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.45324063,0.90466833,1.357909,1.8093367,2.2625773,2.1302311,1.9978848,1.8655385,1.7331922,1.6008459,1.9670644,2.335096,2.7031271,3.0693457,3.437377,3.000453,2.561716,2.124792,1.6878681,1.2491312,1.0533313,0.8557183,0.65810543,0.4604925,0.26287958,0.2520018,0.24293698,0.23205921,0.2229944,0.21211663,0.18310922,0.15228885,0.12328146,0.092461094,0.06164073,0.06707962,0.072518505,0.07795739,0.08339628,0.0870222,0.08339628,0.07795739,0.072518505,0.06707962,0.06164073,0.092461094,0.12328146,0.15228885,0.18310922,0.21211663,1.7368182,3.2633326,4.788034,6.3127356,7.837437,6.2746634,4.7118897,3.149116,1.5881553,0.025381476,0.027194439,0.030820364,0.032633327,0.034446288,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.42785916,0.8557183,1.2817645,1.7096237,2.137483,3.832603,5.527723,7.2228427,8.917963,10.613083,11.874905,13.136727,14.400362,15.662184,16.92582,15.885179,14.844538,13.80571,12.76507,11.724429,10.622148,9.519867,8.417585,7.315304,6.2130227,7.2029004,8.192778,9.182655,10.172533,11.162411,11.176914,11.193231,11.207735,11.222239,11.236742,9.900589,8.562622,7.224656,5.8866897,4.550536,4.844236,5.139749,5.4352617,5.730775,6.0244746,5.3428006,4.6593137,3.97764,3.294153,2.612479,7.4911613,12.368031,17.2449,22.121769,27.000452,21.621391,16.245958,10.866898,5.4896507,0.11240368,2.2879589,4.461701,6.637256,8.812811,10.988366,10.065568,9.142771,8.219973,7.2971745,6.3743763,6.58468,6.794984,7.0052876,7.215591,7.424082,7.473032,7.520169,7.567306,7.614443,7.66158,7.3316207,7.0016613,6.6717024,6.341743,6.011784,4.8097897,3.6077955,2.4058013,1.2019942,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.04169814,0.047137026,0.052575916,0.058014803,0.06164073,0.09789998,0.13234627,0.16679256,0.2030518,0.2374981,0.26287958,0.28826106,0.31182957,0.33721104,0.36259252,0.3245203,0.28826106,0.25018883,0.21211663,0.17585737,0.3100166,0.44417584,0.58014804,0.71430725,0.85027945,1.1022812,1.3542831,1.6080978,1.8600996,2.1121013,2.4003625,2.6868105,2.9750717,3.2633326,3.5497808,2.864481,2.179181,1.4956942,0.8103943,0.12509441,2.759329,5.3953767,8.029612,10.665659,13.299893,15.040338,16.78078,18.519413,20.259857,22.000301,21.244295,20.490103,19.734098,18.979906,18.225714,18.82943,19.43496,20.04049,20.644205,21.249735,22.705544,24.15954,25.615349,27.069344,28.525154,27.747393,26.969631,26.19187,25.415922,24.63816,22.154404,19.672457,17.190512,14.706753,12.224807,14.407614,16.59042,18.773228,20.954222,23.137028,24.975372,26.811903,28.650248,30.486778,32.325123,30.539354,28.7554,26.969631,25.185677,23.399908,20.584377,17.770658,14.955129,12.139598,9.325879,7.9607186,6.5955577,5.230397,3.8652363,2.5000753,3.5679104,4.6357455,5.7017674,6.7696023,7.837437,7.795739,7.752228,7.71053,7.667019,7.6253204,7.931711,8.239915,8.548119,8.854509,9.162713,10.272246,11.381779,12.493125,13.602658,14.712192,14.422117,14.132043,13.8419695,13.551895,13.261822,12.368031,11.472427,10.576823,9.683033,8.78743,9.090195,9.39296,9.695724,9.9966755,10.29944,9.817192,9.334945,8.852696,8.370448,7.8882003,9.610515,11.332829,13.055143,14.777458,16.499773,17.212267,17.92476,18.637255,19.34975,20.062244,17.99184,15.921437,13.852847,11.782444,9.712041,8.312433,6.9128265,5.5132194,4.1117992,2.712192,2.8880494,2.955129,3.0222087,3.0892882,3.1581807,3.2252605,3.584227,3.9450066,4.305786,4.664753,5.0255322,8.009668,10.995618,13.979754,16.965704,19.94984,22.468046,24.984438,27.502642,30.020847,32.53724,32.64783,32.756607,32.8672,32.97779,33.08838,33.494484,33.9024,34.310318,34.718235,35.124336,30.604622,26.084906,21.56519,17.045475,12.525759,10.885027,9.244296,7.605378,5.964647,4.325729,5.4479527,6.5701766,7.6924005,8.814624,9.936848,10.46442,10.991992,11.519565,12.047136,12.574709,12.340837,12.105151,11.869466,11.635593,11.399909,10.042,8.685904,7.327995,5.9700856,4.612177,5.8431783,7.072367,8.303369,9.5325575,10.761745,10.9230995,11.082641,11.242181,11.401722,11.563075,10.114518,8.667774,7.219217,5.772473,4.325729,5.7924156,7.2591023,8.727602,10.194288,11.662788,11.080828,10.497053,9.915092,9.333132,8.749357,7.404139,6.060734,4.7155156,3.3702974,2.0250793,1.7676386,1.5101979,1.2527572,0.99531645,0.73787576,1.2654479,1.79302,2.3205922,2.8481643,3.3757362,3.6676233,3.9595103,4.25321,4.5450974,4.836984,4.7155156,4.592234,4.4707656,4.347484,4.2242026,4.079166,3.9341288,3.7890918,3.6458678,3.5008307,3.5153344,3.529838,3.5443418,3.5606585,3.5751622,3.3231604,3.0693457,2.817344,2.565342,2.3133402,2.1030366,1.892733,1.6824293,1.4721256,1.261822,1.1004683,0.93730164,0.774135,0.61278135,0.44961473,0.49675176,0.54570174,0.59283876,0.6399758,0.6871128,1.261822,1.8383441,2.4130533,2.9877625,3.5624714,4.2242026,4.8877473,5.5494785,6.2130227,6.874754,6.341743,5.810545,5.277534,4.744523,4.213325,4.1099863,4.006647,3.9051213,3.8017826,3.7002566,3.6748753,3.6494937,3.6241121,3.6005437,3.5751622,3.3122826,3.049403,2.7883365,2.525457,2.2625773,2.3677292,2.472881,2.5780327,2.6831846,2.7883365,2.9841363,3.1817493,3.3793623,3.576975,3.774588,4.160749,4.5450974,4.9294453,5.315606,5.6999545,5.0200934,4.3402324,3.6603715,2.9805105,2.3006494,2.3097143,2.3205922,2.3296568,2.3405347,2.3495996,2.6904364,3.0294604,3.3702974,3.7093215,4.0501585,4.0900435,4.1299286,4.169814,4.209699,4.249584,4.853301,5.4552045,6.057108,6.6608243,7.262728,6.8403077,6.4178877,5.995467,5.573047,5.1506267,5.9283876,6.7043357,7.4820967,8.259857,9.037619,11.450671,13.861912,16.274965,18.688019,21.099258,19.507477,17.915697,16.322102,14.730321,13.136727,13.483003,13.827466,14.171928,14.518205,14.862667,14.880796,14.897114,14.915243,14.9333725,14.94969,13.136727,11.325577,9.512614,7.699652,5.8866897,5.1506267,4.4127507,3.6748753,2.9369993,2.1991236,4.751775,7.304426,9.857078,12.409729,14.96238,13.591781,12.222994,10.852394,9.481794,8.113008,6.7279043,5.3428006,3.9576974,2.572594,1.1874905,4.842423,8.497355,12.152288,15.80722,19.462152,17.290224,15.118295,12.944552,10.772624,8.600695,10.770811,12.939114,15.10923,17.279346,19.449463,21.447348,23.445232,25.443117,27.439188,29.437073,24.130531,18.822178,13.515636,8.207282,2.9007401,2.570781,2.2408218,1.9108626,1.5809034,1.2491312,1.2926424,1.3343405,1.3778516,1.4195497,1.4630609,1.3996071,1.3379664,1.2745126,1.2128719,1.1494182,1.1204109,1.0895905,1.0605831,1.0297627,1.0007553,0.8448406,0.69073874,0.53482395,0.38072214,0.22480737,0.28282216,0.34083697,0.39703882,0.4550536,0.51306844,0.45324063,0.39159992,0.33177215,0.27194437,0.21211663,0.3154555,0.4169814,0.52032024,0.62184614,0.72518504,1.8202144,2.9152439,4.0102735,5.105303,6.200332,5.2648435,4.329355,3.395679,2.4601903,1.5247015,1.2817645,1.0406405,0.79770356,0.55476654,0.31182957,0.27919623,0.24837588,0.21574254,0.18310922,0.15047589,0.25562772,0.36077955,0.46411842,0.56927025,0.6744221,0.5402629,0.40429065,0.27013144,0.13415924,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.46955732,0.93911463,1.4104849,1.8800422,2.3495996,2.039583,1.7295663,1.4195497,1.1095331,0.7995165,0.9898776,1.1802386,1.3705997,1.5591478,1.7495089,1.7241274,1.7005589,1.6751775,1.649796,1.6244144,1.357909,1.0895905,0.823085,0.55476654,0.28826106,0.28282216,0.27738327,0.27194437,0.26831847,0.26287958,0.2229944,0.18310922,0.14322405,0.10333887,0.06164073,0.065266654,0.06707962,0.07070554,0.072518505,0.07433146,0.072518505,0.07070554,0.06707962,0.065266654,0.06164073,0.10333887,0.14322405,0.18310922,0.2229944,0.26287958,1.8746033,3.48814,5.0998635,6.7134004,8.325124,6.6626377,5.0001507,3.3376641,1.6751775,0.012690738,0.01994259,0.027194439,0.034446288,0.04169814,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.55839247,1.114972,1.6733645,2.229944,2.7883365,4.3347936,5.883064,7.4295206,8.977791,10.524248,11.650098,12.774135,13.899984,15.025834,16.14987,15.555219,14.960567,14.364102,13.769451,13.174799,11.842272,10.509744,9.177217,7.844689,6.5121617,7.119504,7.7268467,8.334189,8.943344,9.550687,9.657652,9.764616,9.873394,9.980359,10.087324,8.6877165,7.28811,5.8866897,4.4870825,3.0874753,3.5225863,3.9576974,4.3928084,4.8279195,5.2630305,4.603112,3.9431937,3.2832751,2.6233568,1.9616255,6.6698895,11.378153,16.084604,20.792868,25.49932,20.430275,15.359419,10.290376,5.219519,0.15047589,2.0123885,3.874301,5.7380266,7.5999393,9.461852,8.694968,7.9280853,7.159389,6.392506,5.6256227,5.2557783,4.8841214,4.514277,4.1444325,3.774588,4.1933823,4.610364,5.027345,5.4443264,5.863121,5.823236,5.7833505,5.7416525,5.7017674,5.661882,4.5305934,3.397492,2.2643902,1.1331016,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.052575916,0.054388877,0.058014803,0.059827764,0.06164073,0.10515183,0.14684997,0.19036107,0.23205921,0.2755703,0.2991388,0.3245203,0.34990177,0.37528324,0.40066472,0.34990177,0.2991388,0.25018883,0.19942589,0.15047589,0.34264994,0.53482395,0.726998,0.91917205,1.1131591,1.357909,1.6026589,1.8474089,2.0921588,2.3369088,2.2371957,2.137483,2.03777,1.938057,1.8383441,1.4830034,1.1276628,0.77232206,0.4169814,0.06164073,3.4047437,6.7478466,10.09095,13.43224,16.775343,18.519413,20.265295,22.009365,23.755249,25.49932,23.771564,22.045626,20.317871,18.590118,16.862366,17.364555,17.866747,18.37075,18.87294,19.375132,20.903458,22.429974,23.9583,25.484816,27.013142,26.393108,25.773077,25.153044,24.53301,23.912977,21.59057,19.268166,16.94576,14.623356,12.299138,14.759329,17.219519,19.679708,22.139898,24.60009,26.737572,28.875055,31.012537,33.15002,35.287502,33.67034,32.053177,30.434202,28.81704,27.199877,23.729868,20.259857,16.789846,13.319836,9.849826,8.404895,6.9599633,5.5150323,4.070101,2.6251698,4.1897564,5.754343,7.320743,8.885329,10.449916,10.359268,10.270433,10.179785,10.089137,10.000301,10.246864,10.49524,10.741803,10.990179,11.236742,12.904668,14.572594,16.240519,17.906631,19.574556,18.79317,18.00997,17.22677,16.445383,15.662184,14.315152,12.968122,11.619277,10.272246,8.925215,9.082943,9.24067,9.398398,9.554313,9.712041,9.264238,8.81825,8.370448,7.9226465,7.474845,9.130079,10.785315,12.440549,14.095784,15.749206,16.550535,17.350052,18.149569,18.949085,19.750414,17.652817,15.555219,13.457622,11.3600235,9.262425,7.7757964,6.2873545,4.800725,3.3122826,1.8256533,2.7502642,2.8245957,2.9007401,2.9750717,3.049403,3.1255474,3.5624714,3.9993954,4.4381323,4.8750563,5.3119802,7.574558,9.837135,12.099712,14.362289,16.624866,19.63801,22.649342,25.662485,28.675629,31.68696,32.200027,32.713097,33.224354,33.73742,34.25049,33.69935,33.15002,32.600693,32.049553,31.500225,27.674873,23.849524,20.024172,16.200634,12.375282,10.750868,9.12464,7.500226,5.8758116,4.249584,5.6999545,7.1503243,8.600695,10.049252,11.499621,12.199425,12.899229,13.600845,14.300649,15.000452,14.561715,14.124791,13.687867,13.24913,12.812206,11.225864,9.637709,8.049554,6.4632115,4.8750563,6.412449,7.949841,9.487233,11.024626,12.562017,12.387974,12.212116,12.038072,11.862214,11.6881695,10.28675,8.887142,7.4875355,6.0879283,4.688321,6.588306,8.488291,10.388275,12.28826,14.188245,13.475751,12.763257,12.050762,11.338268,10.625773,8.925215,7.224656,5.524097,3.825351,2.124792,1.8492218,1.5754645,1.2998942,1.0243238,0.7505665,1.261822,1.7748904,2.2879589,2.7992141,3.3122826,3.6005437,3.8869917,4.175253,4.461701,4.749962,4.612177,4.4743915,4.3366065,4.2006345,4.062849,3.9123733,3.7618973,3.6132345,3.4627585,3.3122826,3.1618068,3.0131438,2.8626678,2.712192,2.561716,2.3369088,2.1121013,1.887294,1.6624867,1.4376793,1.4630609,1.4866294,1.5120108,1.5373923,1.5627737,1.3633479,1.162109,0.96268314,0.76325727,0.5620184,0.44961473,0.33721104,0.22480737,0.11240368,0.0,0.13778515,0.2755703,0.41335547,0.5493277,0.6871128,1.7621996,2.8372865,3.9123733,4.98746,6.0625467,5.712645,5.3627434,5.0128417,4.6629395,4.313038,4.3366065,4.361988,4.3873696,4.4127507,4.4381323,4.274966,4.1117992,3.9504454,3.787279,3.6241121,3.3757362,3.1255474,2.8753586,2.6251698,2.374981,2.474694,2.5744069,2.6741197,2.7756457,2.8753586,3.1255474,3.3757362,3.6241121,3.874301,4.12449,4.550536,4.974769,5.4008155,5.825049,6.249282,5.424384,4.599486,3.774588,2.94969,2.124792,2.1991236,2.275268,2.3495996,2.4257438,2.5000753,2.8880494,3.2742105,3.6621845,4.0501585,4.4381323,4.3873696,4.3366065,4.2876563,4.2368937,4.1879435,4.836984,5.487838,6.1368785,6.787732,7.4367723,6.887445,6.338117,5.7869763,5.237649,4.688321,5.2122674,5.7380266,6.261973,6.787732,7.311678,10.56232,13.812962,17.06179,20.312433,23.563074,21.949537,20.337814,18.724277,17.112555,15.50083,15.524399,15.54978,15.575162,15.600543,15.624111,15.725637,15.825351,15.925063,16.024776,16.124489,14.211814,12.300951,10.388275,8.4756,6.5629244,5.3500524,4.137181,2.9243085,1.7132497,0.50037766,3.2379513,5.975525,8.713099,11.450671,14.188245,13.087777,11.9873085,10.88684,9.788185,8.6877165,7.124943,5.562169,3.9993954,2.4366217,0.87566096,5.2992897,9.724731,14.150173,18.575615,22.999243,19.812056,16.624866,13.437678,10.25049,7.063302,9.737422,12.411542,15.087475,17.763407,20.437527,23.088078,25.736816,28.387367,31.03792,33.686657,27.26333,20.838192,14.413053,7.987913,1.5627737,1.3379664,1.1131591,0.8883517,0.66173136,0.43692398,0.63816285,0.8375887,1.0370146,1.2382535,1.4376793,1.3996071,1.3633479,1.3252757,1.2872034,1.2491312,1.1494182,1.0497054,0.9499924,0.85027945,0.7505665,0.62547207,0.50037766,0.37528324,0.25018883,0.12509441,0.18673515,0.25018883,0.31182957,0.37528324,0.43692398,0.34990177,0.26287958,0.17585737,0.0870222,0.0,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,1.7495089,3.2506418,4.749962,6.249282,7.750415,6.4251394,5.0998635,3.774588,2.4493124,1.1258497,0.97537386,0.824898,0.6744221,0.52575916,0.37528324,0.33721104,0.2991388,0.26287958,0.22480737,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.48768693,0.97537386,1.4630609,1.9507477,2.4366217,1.9507477,1.4630609,0.97537386,0.48768693,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.44961473,0.8375887,1.2255627,1.6117238,1.9996977,1.6624867,1.3252757,0.9880646,0.6508536,0.31182957,0.31182957,0.31182957,0.31182957,0.31182957,0.31182957,0.26287958,0.21211663,0.16316663,0.11240368,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.11240368,0.16316663,0.21211663,0.26287958,0.31182957,2.0123885,3.7129474,5.411693,7.112252,8.812811,7.0506115,5.2884116,3.5243993,1.7621996,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.6871128,1.3742256,2.0631514,2.7502642,3.437377,4.836984,6.2365913,7.6380115,9.037619,10.437225,11.42529,12.413355,13.399607,14.387671,15.375735,15.22526,15.074784,14.924308,14.775645,14.625169,13.062395,11.499621,9.936848,8.374074,6.813113,7.037921,7.262728,7.4875355,7.7123427,7.93715,8.138389,8.337815,8.537241,8.736667,8.937905,7.474845,6.011784,4.550536,3.0874753,1.6244144,2.2009366,2.7756457,3.350355,3.925064,4.499773,3.8616104,3.2252605,2.5870976,1.9507477,1.3125849,5.8504305,10.386462,14.924308,19.462152,23.999998,19.237347,14.474693,9.712041,4.949388,0.18673515,1.7368182,3.2869012,4.836984,6.3870673,7.93715,7.324369,6.7134004,6.1006193,5.487838,4.8750563,3.925064,2.9750717,2.0250793,1.0750868,0.12509441,0.9119202,1.7005589,2.4873846,3.2742105,4.062849,4.313038,4.5632267,4.8116026,5.0617914,5.3119802,4.249584,3.1871881,2.124792,1.062396,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.11240368,0.16316663,0.21211663,0.26287958,0.31182957,0.33721104,0.36259252,0.387974,0.41335547,0.43692398,0.37528324,0.31182957,0.25018883,0.18673515,0.12509441,0.37528324,0.62547207,0.87566096,1.1258497,1.3742256,1.6117238,1.8492218,2.08672,2.324218,2.561716,2.0758421,1.5881553,1.1004683,0.61278135,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,4.0501585,8.100317,12.1504755,16.200634,20.250792,22.000301,23.74981,25.49932,27.25064,29.000149,26.300648,23.599335,20.899832,18.20033,15.50083,15.899682,16.300346,16.699198,17.099863,17.500528,19.099562,20.700407,22.29944,23.900286,25.49932,25.037014,24.574707,24.112402,23.650097,23.187792,21.024927,18.862062,16.699198,14.538147,12.375282,15.112856,17.85043,20.588003,23.325577,26.06315,28.499771,30.938206,33.37483,35.81145,38.249886,36.799515,35.349144,33.90059,32.45022,30.999847,26.875357,22.750868,18.624565,14.500074,10.375585,8.849071,7.324369,5.7996674,4.274966,2.7502642,4.8134155,6.874754,8.937905,10.999244,13.062395,12.92461,12.786825,12.650853,12.513068,12.375282,12.562017,12.750566,12.937301,13.125849,13.312584,15.537089,17.763407,19.987913,22.212418,24.436922,23.16241,21.887897,20.611572,19.337059,18.062546,16.262274,14.462003,12.661731,10.863272,9.063,9.07569,9.088382,9.099259,9.11195,9.12464,8.713099,8.299743,7.8882003,7.474845,7.063302,8.649645,10.2378,11.825955,13.412297,15.000452,15.8869915,16.775343,17.661882,18.550234,19.436771,17.31198,15.187187,13.062395,10.937603,8.812811,7.2373466,5.661882,4.0882306,2.5127661,0.93730164,2.6505513,2.7067533,2.764768,2.8227828,2.8807976,2.9369993,3.3249733,3.7129474,4.099108,4.4870825,4.8750563,7.309865,9.744674,12.179482,14.614291,17.0491,19.844688,22.640276,25.435865,28.229641,31.025229,31.329807,31.634384,31.940775,32.245354,32.54993,32.172832,31.795738,31.416828,31.039732,30.662636,26.940624,23.216799,19.494787,15.772775,12.050762,10.484363,8.919776,7.3551893,5.7906027,4.2242026,5.7017674,7.179332,8.656897,10.13446,11.612025,12.35534,13.096842,13.840157,14.581658,15.324973,14.935185,14.545399,14.155612,13.765825,13.374225,11.989121,10.605831,9.220728,7.835624,6.450521,7.512917,8.575313,9.637709,10.700105,11.762501,11.700861,11.637406,11.575767,11.512312,11.450671,10.29944,9.1500225,8.000604,6.849373,5.6999545,7.1956487,8.689529,10.185224,11.680918,13.174799,12.650853,12.125093,11.599335,11.075388,10.549629,9.202598,7.855567,6.506723,5.1596913,3.8126602,3.5080826,3.2016919,2.8971143,2.5925364,2.2879589,2.619731,2.953316,3.2850883,3.6168604,3.9504454,4.329355,4.710077,5.090799,5.469708,5.8504305,5.560356,5.2702823,4.9802084,4.690134,4.40006,4.1970086,3.9957695,3.7927177,3.589666,3.386614,3.198066,3.007705,2.817344,2.6269827,2.4366217,2.2081885,1.9779422,1.7476959,1.5174497,1.2872034,1.3542831,1.4231756,1.4902552,1.5573349,1.6244144,1.7803292,1.9344311,2.0903459,2.2444477,2.4003625,2.2045624,2.0105755,1.8147756,1.6207886,1.4249886,1.2491312,1.0750868,0.89922947,0.72518504,0.5493277,1.8945459,3.2397642,4.5849824,5.9302006,7.2754188,7.0125394,6.7496595,6.48678,6.2257137,5.962834,5.9120708,5.863121,5.812358,5.763408,5.712645,5.3428006,4.972956,4.603112,4.233268,3.8616104,3.5969179,3.3322253,3.0675328,2.8028402,2.5381477,2.6269827,2.7176309,2.808279,2.8971143,2.9877625,3.245203,3.5026438,3.7600844,4.017525,4.274966,4.5849824,4.894999,5.2050157,5.5150323,5.825049,5.0744824,4.325729,3.5751622,2.8245957,2.0758421,2.231757,2.3894846,2.5472124,2.70494,2.8626678,3.149116,3.437377,3.7256382,4.0120864,4.3003473,4.2894692,4.2804046,4.269527,4.2604623,4.249584,4.7282066,5.2050157,5.6818247,6.1604466,6.637256,6.209397,5.7833505,5.3554916,4.9276323,4.499773,5.4570174,6.414262,7.3733187,8.330563,9.287807,12.117842,14.947877,17.77791,20.607946,23.43798,22.042,20.647831,19.25185,17.857681,16.4617,16.427254,16.392807,16.358362,16.322102,16.287657,16.193382,16.097294,16.003021,15.906934,15.812659,14.567154,13.321649,12.077957,10.832452,9.5869465,7.9280853,6.2674117,4.606738,2.9478772,1.2872034,3.8108473,6.3326783,8.854509,11.378153,13.899984,12.665357,11.430729,10.194288,8.9596615,7.7250338,6.4269524,5.130684,3.832603,2.5345216,1.2382535,4.940323,8.642392,12.344462,16.048346,19.750414,16.972956,14.195497,11.418038,8.640579,5.863121,8.120259,10.377398,12.634536,14.891675,17.150625,19.465778,21.77912,24.094273,26.409426,28.724579,23.236742,17.750717,12.262879,6.775041,1.2872034,1.1530442,1.017072,0.88291276,0.7469406,0.61278135,0.73424983,0.8575313,0.9808127,1.1022812,1.2255627,1.2128719,1.2001812,1.1874905,1.1747998,1.162109,1.0497054,0.93730164,0.824898,0.7124943,0.6000906,0.50219065,0.40429065,0.30820364,0.21030366,0.11240368,0.22480737,0.33721104,0.44961473,0.5620184,0.6744221,0.5402629,0.40429065,0.27013144,0.13415924,0.0,0.08520924,0.17041849,0.25562772,0.34083697,0.42423326,1.5827163,2.7393866,3.8978696,5.0545397,6.2130227,5.3428006,4.4725785,3.6023567,2.7321346,1.8619126,1.7132497,1.5627737,1.4122978,1.261822,1.1131591,0.91917205,0.726998,0.53482395,0.34264994,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.45324063,0.90466833,1.357909,1.8093367,2.2625773,1.8093367,1.357909,0.90466833,0.45324063,0.0,0.15591478,0.3100166,0.46411842,0.6200332,0.774135,1.3125849,1.8492218,2.3876717,2.9243085,3.4627585,3.1146698,2.7683938,2.420305,2.0722163,1.7241274,1.4304274,1.1349145,0.83940166,0.54570174,0.25018883,0.21211663,0.17585737,0.13778515,0.099712946,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.25925365,0.45686656,0.6544795,0.8520924,1.0497054,2.467442,3.8851788,5.3029156,6.720652,8.138389,6.530291,4.9221935,3.3140955,1.7078108,0.099712946,0.092461094,0.08520924,0.07795739,0.07070554,0.06164073,0.052575916,0.04169814,0.032633327,0.02175555,0.012690738,0.6508536,1.2872034,1.9253663,2.561716,3.199879,4.445384,5.6890764,6.9345818,8.180087,9.425592,10.852394,12.279196,13.70781,15.134612,16.563227,15.917811,15.272397,14.626982,13.98338,13.337966,12.070704,10.801631,9.53437,8.267109,6.9998484,7.155763,7.309865,7.46578,7.6198816,7.7757964,7.9081426,8.040489,8.172835,8.3051815,8.437528,7.0506115,5.661882,4.274966,2.8880494,1.49932,2.0069497,2.514579,3.0222087,3.529838,4.0374675,3.576975,3.1182957,2.657803,2.1973107,1.7368182,5.9320135,10.127209,14.322405,18.5176,22.712795,18.43239,14.151986,9.871581,5.5929894,1.3125849,2.7974012,4.2822175,5.767034,7.25185,8.736667,7.8628187,6.987158,6.11331,5.237649,4.361988,3.5552197,2.7466383,1.93987,1.1331016,0.3245203,0.99531645,1.6642996,2.335096,3.005892,3.6748753,4.0846047,4.494334,4.9058766,5.315606,5.7253356,4.5867953,3.4500678,2.3133402,1.1747998,0.038072214,0.045324065,0.052575916,0.059827764,0.06707962,0.07433146,0.07795739,0.07977036,0.08339628,0.08520924,0.0870222,0.13415924,0.18310922,0.23024625,0.27738327,0.3245203,0.33721104,0.34990177,0.36259252,0.37528324,0.387974,0.35171473,0.31726846,0.28282216,0.24837588,0.21211663,0.46955732,0.726998,0.98443866,1.2418793,1.49932,1.6171626,1.7350051,1.8528478,1.9706904,2.08672,1.6896812,1.2926424,0.89560354,0.49675176,0.099712946,0.11421664,0.13053331,0.14503701,0.15954071,0.17585737,4.347484,8.519112,12.692551,16.864178,21.037619,22.462606,23.887594,25.312584,26.737572,28.162561,25.71325,23.262123,20.81281,18.363499,15.912373,15.810846,15.707508,15.604169,15.502643,15.399304,16.650248,17.89938,19.150324,20.399454,21.650398,21.512613,21.374828,21.237043,21.099258,20.963285,19.641636,18.3218,17.001963,15.682126,14.362289,16.728207,19.092308,21.458225,23.822329,26.188244,28.378304,30.56655,32.75842,34.946667,37.136726,36.328144,35.51775,34.707355,33.89696,33.08838,28.686506,24.28826,19.888199,15.488139,11.088079,9.804502,8.5227375,7.2391596,5.957395,4.6756306,6.4777155,8.2798,10.081885,11.885782,13.687867,13.446743,13.207433,12.968122,12.726997,12.487686,12.692551,12.897416,13.102281,13.307145,13.512011,15.212569,16.913128,18.611874,20.312433,22.01299,21.82807,21.643147,21.458225,21.273302,21.08838,18.782291,16.478018,14.171928,11.867653,9.563377,9.5525,9.541622,9.5325575,9.52168,9.512614,9.244296,8.977791,8.709473,8.442966,8.174648,9.441909,10.710983,11.978244,13.245504,14.512766,15.245202,15.977639,16.710075,17.442513,18.17495,16.026588,13.880041,11.731681,9.585134,7.4367723,6.1803894,4.9221935,3.6658103,2.4076142,1.1494182,2.5508385,2.5907235,2.6306088,2.6704938,2.7103791,2.7502642,3.0874753,3.4246864,3.7618973,4.099108,4.4381323,7.0451727,9.652213,12.259253,14.868106,17.475147,20.053179,22.629398,25.207432,27.785465,30.361685,30.459585,30.557484,30.655384,30.753284,30.849371,30.644506,30.439642,30.234777,30.029913,29.825047,26.204561,22.585888,18.9654,15.344915,11.724429,10.21967,8.714911,7.210152,5.7053933,4.2006345,5.7053933,7.210152,8.714911,10.21967,11.724429,12.509441,13.294455,14.079468,14.86448,15.649493,15.306843,14.964193,14.623356,14.280706,13.938056,12.754191,11.57214,10.390089,9.208037,8.024173,8.613385,9.200785,9.788185,10.375585,10.962985,11.011934,11.062697,11.111648,11.162411,11.213174,10.312131,9.412902,8.511859,7.61263,6.7134004,7.802991,8.892582,9.982172,11.071762,12.163166,11.8241415,11.486931,11.14972,10.812509,10.475298,9.479981,8.484665,7.4893484,6.495845,5.5005283,5.1651306,4.8297324,4.494334,4.160749,3.825351,3.97764,4.1299286,4.2822175,4.4345064,4.5867953,5.0599785,5.5331616,6.004532,6.4777155,6.9508986,6.506723,6.0643597,5.621997,5.179634,4.7372713,4.4816437,4.227829,3.972201,3.7183862,3.4627585,3.2325122,3.002266,2.7720199,2.5417736,2.3133402,2.077655,1.84197,1.6080978,1.3724127,1.1367276,1.2473183,1.357909,1.4666867,1.5772774,1.6878681,2.1973107,2.7067533,3.2180085,3.727451,4.2368937,3.9595103,3.682127,3.4047437,3.1273603,2.8499773,2.3622901,1.8746033,1.3869164,0.89922947,0.41335547,2.0268922,3.6422417,5.2575917,6.872941,8.488291,8.312433,8.138389,7.9625316,7.7866745,7.61263,7.4875355,7.362441,7.2373466,7.112252,6.987158,6.4106355,5.8323007,5.2557783,4.6774435,4.099108,3.8199122,3.540716,3.2597067,2.9805105,2.6995013,2.7792716,2.8608549,2.9406252,3.0203958,3.100166,3.3648586,3.6295512,3.8942437,4.160749,4.4254417,4.6194286,4.8152285,5.009216,5.2050157,5.4008155,4.7245803,4.0501585,3.3757362,2.6995013,2.0250793,2.2643902,2.5055144,2.7448254,2.9841363,3.2252605,3.4119956,3.6005437,3.787279,3.975827,4.162562,4.1933823,4.2223897,4.25321,4.2822175,4.313038,4.6176157,4.9221935,5.2267714,5.5331616,5.8377395,5.5331616,5.2267714,4.9221935,4.6176157,4.313038,5.7017674,7.0923095,8.482852,9.873394,11.262123,13.673364,16.08279,18.492218,20.901646,23.312885,22.13446,20.957848,19.77942,18.60281,17.424383,17.330109,17.235836,17.139748,17.045475,16.949387,16.659313,16.36924,16.079165,15.789091,15.50083,14.922495,14.34416,13.767638,13.189302,12.612781,10.504305,8.397643,6.2891674,4.1825047,2.0758421,4.3819304,6.6898317,8.997733,11.3056345,13.611723,12.242936,10.872336,9.501737,8.13295,6.7623506,5.730775,4.6973863,3.6658103,2.6324217,1.6008459,4.5795436,7.560054,10.540565,13.519262,16.499773,14.132043,11.764315,9.396585,7.0306687,4.6629395,6.5030966,8.343254,10.183411,12.021755,13.861912,15.841667,17.823235,19.80299,21.782745,23.7625,19.211964,14.663241,10.112705,5.562169,1.0116332,0.968122,0.922798,0.8774739,0.8321498,0.7868258,0.8321498,0.8774739,0.922798,0.968122,1.0116332,1.0243238,1.0370146,1.0497054,1.062396,1.0750868,0.9499924,0.824898,0.69980353,0.5747091,0.44961473,0.38072214,0.3100166,0.23931105,0.17041849,0.099712946,0.26287958,0.42423326,0.5873999,0.7505665,0.9119202,0.7306239,0.5475147,0.36440548,0.18310922,0.0,0.11965553,0.23931105,0.36077955,0.48043507,0.6000906,1.4159238,2.229944,3.045777,3.8597972,4.6756306,4.2604623,3.8452935,3.4301252,3.0149567,2.5997884,2.4493124,2.3006494,2.1501737,1.9996977,1.8492218,1.502946,1.1548572,0.80676836,0.4604925,0.11240368,0.09064813,0.06707962,0.045324065,0.02175555,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.4169814,0.83577573,1.2527572,1.6697385,2.08672,1.6697385,1.2527572,0.83577573,0.4169814,0.0,0.29732585,0.5946517,0.8919776,1.1893034,1.4866294,2.175555,2.8626678,3.5497808,4.2368937,4.9258194,4.5668526,4.209699,3.8525455,3.4953918,3.1382382,2.5472124,1.9579996,1.3669738,0.7777609,0.18673515,0.16316663,0.13778515,0.11240368,0.0870222,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.40791658,0.7523795,1.0968424,1.4431182,1.7875811,2.9224956,4.0574102,5.1923246,6.3272395,7.462154,6.009971,4.557788,3.105605,1.651609,0.19942589,0.17223145,0.14503701,0.11784257,0.09064813,0.06164073,0.054388877,0.047137026,0.03988518,0.032633327,0.025381476,0.61278135,1.2001812,1.7875811,2.374981,2.962381,4.0519714,5.141562,6.2329655,7.322556,8.412147,10.279498,12.14685,14.014201,15.883366,17.750717,16.610363,15.47001,14.329657,13.189302,12.050762,11.077202,10.1054535,9.131892,8.160145,7.1883965,7.271793,7.3570023,7.4422116,7.5274205,7.61263,7.6778965,7.743163,7.806617,7.8718834,7.93715,6.624565,5.3119802,3.9993954,2.6868105,1.3742256,1.8147756,2.2553256,2.6958754,3.1346123,3.5751622,3.29234,3.009518,2.7266958,2.4456866,2.1628644,6.01541,9.867955,13.720501,17.573046,21.425592,17.627436,13.829279,10.032935,6.2347784,2.4366217,3.8579843,5.277534,6.697084,8.116633,9.537996,8.399456,7.262728,6.1241875,4.98746,3.8507326,3.1853752,2.520018,1.8546607,1.1893034,0.52575916,1.0768998,1.6298534,2.182807,2.7357605,3.2869012,3.8579843,4.4272547,4.9983377,5.567608,6.1368785,4.9258194,3.7129474,2.5000753,1.2872034,0.07433146,0.07795739,0.07977036,0.08339628,0.08520924,0.0870222,0.092461094,0.09789998,0.10333887,0.10696479,0.11240368,0.15772775,0.2030518,0.24837588,0.291887,0.33721104,0.33721104,0.33721104,0.33721104,0.33721104,0.33721104,0.32995918,0.32270733,0.3154555,0.30820364,0.2991388,0.5656443,0.83033687,1.0950294,1.3597219,1.6244144,1.6226015,1.6207886,1.6171626,1.6153497,1.6117238,1.305333,0.99712944,0.69073874,0.3825351,0.07433146,0.13053331,0.18492219,0.23931105,0.2955129,0.34990177,4.64481,8.939718,13.234627,17.529535,21.824444,22.924911,24.025381,25.125849,26.224504,27.324972,25.124035,22.924911,20.725788,18.52485,16.325727,15.720199,15.114669,14.50914,13.905423,13.299893,14.200936,15.100165,15.999394,16.900436,17.799667,17.988214,18.17495,18.361685,18.550234,18.736969,18.260159,17.78335,17.304728,16.827919,16.349297,18.341742,20.334188,22.328447,24.31908,26.31334,28.255022,30.196705,32.1402,34.081882,36.02538,35.85496,35.684544,35.514126,35.34552,35.1751,30.49947,25.825651,21.15002,16.474392,11.800573,10.7599325,9.719293,8.680465,7.6398244,6.599184,8.1420145,9.684846,11.227677,12.770509,14.313339,13.97069,13.628039,13.28539,12.9427395,12.60009,12.823084,13.044266,13.267261,13.490254,13.713249,14.888049,16.062849,17.237648,18.412449,19.587248,20.491917,21.398397,22.303066,23.207733,24.112402,21.30231,18.492218,15.682126,12.872034,10.061942,10.029309,9.9966755,9.965856,9.933222,9.900589,9.7773075,9.655839,9.5325575,9.409276,9.287807,10.234174,11.182353,12.130532,13.0769,14.025079,14.603414,15.179935,15.758271,16.334793,16.913128,14.743011,12.572895,10.40278,8.232663,6.0625467,5.121619,4.1825047,3.2415771,2.3024626,1.3633479,2.4493124,2.472881,2.4946365,2.518205,2.5399606,2.561716,2.8499773,3.1382382,3.4246864,3.7129474,3.9993954,6.78048,9.5597515,12.340837,15.120108,17.89938,20.259857,22.620335,24.980812,27.339476,29.699953,29.589363,29.480585,29.369993,29.259403,29.150625,29.117992,29.08536,29.052725,29.020092,28.98746,25.470312,21.953163,18.434204,14.917056,11.399909,9.954978,8.510046,7.065115,5.620184,4.175253,5.7072062,7.2391596,8.772926,10.304879,11.836833,12.665357,13.492067,14.320591,15.147303,15.975826,15.680313,15.384801,15.089288,14.795588,14.500074,13.519262,12.540262,11.559449,10.58045,9.599637,9.712041,9.824444,9.936848,10.049252,10.161655,10.324821,10.487988,10.649343,10.812509,10.975676,10.324821,9.675781,9.024928,8.375887,7.7250338,8.410334,9.0956335,9.77912,10.46442,11.14972,10.999244,10.850581,10.700105,10.549629,10.399154,9.757364,9.115576,8.471974,7.8301854,7.1883965,6.8221784,6.4577727,6.093367,5.727149,5.3627434,5.335549,5.3083544,5.279347,5.2521524,5.224958,5.7906027,6.354434,6.9200783,7.4857225,8.049554,7.454902,6.8602505,6.265599,5.669134,5.0744824,4.7680917,4.459888,4.1516843,3.8452935,3.53709,3.2669585,2.9968271,2.7266958,2.4583774,2.1882458,1.9471219,1.7078108,1.4666867,1.2273756,0.9880646,1.1403534,1.2926424,1.4449311,1.5972201,1.7495089,2.6142921,3.4808881,4.345671,5.2104545,6.0752378,5.714458,5.3554916,4.994712,4.6357455,4.274966,3.4754493,2.675933,1.8746033,1.0750868,0.2755703,2.1592383,4.0447197,5.9302006,7.8156815,9.699349,9.612328,9.525306,9.438283,9.349448,9.262425,9.063,8.861761,8.662335,8.46291,8.26167,7.476658,6.6916447,5.906632,5.121619,4.3366065,4.0429068,3.7473936,3.4518807,3.1581807,2.8626678,2.9333735,3.002266,3.0729716,3.141864,3.2125697,3.484514,3.7582715,4.0302157,4.3021603,4.574105,4.655688,4.7354584,4.8152285,4.894999,4.974769,4.3746786,3.774588,3.1744974,2.5744069,1.9743162,2.2970235,2.619731,2.9424384,3.2651455,3.587853,3.6748753,3.7618973,3.8507326,3.9377546,4.024777,4.0954823,4.164375,4.2350807,4.305786,4.3746786,4.507025,4.6393714,4.7717175,4.9058766,5.038223,4.855114,4.6720047,4.4907084,4.307599,4.12449,5.9483304,7.7703576,9.592385,11.4144125,13.238253,15.227073,17.217705,19.208338,21.197159,23.187792,22.226921,21.267864,20.306993,19.347937,18.387066,18.232965,18.07705,17.922949,17.767033,17.612932,17.127058,16.642996,16.157122,15.673061,15.187187,15.277836,15.366671,15.457319,15.547967,15.636803,13.082338,10.527874,7.9715962,5.4171324,2.8626678,4.954827,7.0469856,9.140957,11.233116,13.325275,11.820516,10.315757,8.809185,7.304426,5.7996674,5.032784,4.265901,3.4972048,2.7303216,1.9616255,4.220577,6.4777155,8.734854,10.991992,13.24913,11.292944,9.334945,7.3769445,5.4207582,3.4627585,4.8841214,6.3072968,7.7304726,9.151835,10.57501,12.219368,13.865538,15.509895,17.154251,18.800423,15.187187,11.575767,7.9625316,4.349297,0.73787576,0.78319985,0.82671094,0.872035,0.91735905,0.96268314,0.9300498,0.8974165,0.86478317,0.8321498,0.7995165,0.8375887,0.87566096,0.9119202,0.9499924,0.9880646,0.85027945,0.7124943,0.5747091,0.43692398,0.2991388,0.2574407,0.21574254,0.17223145,0.13053331,0.0870222,0.2991388,0.51306844,0.72518504,0.93730164,1.1494182,0.91917205,0.69073874,0.4604925,0.23024625,0.0,0.15591478,0.3100166,0.46411842,0.6200332,0.774135,1.2473183,1.7205015,2.1918716,2.665055,3.1382382,3.1781235,3.2180085,3.2578938,3.2977788,3.3376641,3.1871881,3.0367124,2.8880494,2.7375734,2.5870976,2.084907,1.5827163,1.0805258,0.57833505,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.09064813,0.06707962,0.045324065,0.02175555,0.0,0.3825351,0.7650702,1.1476053,1.5301404,1.9126755,1.5301404,1.1476053,0.7650702,0.3825351,0.0,0.4405499,0.8792868,1.3198367,1.7603867,2.1991236,3.0367124,3.874301,4.7118897,5.5494785,6.3870673,6.0208488,5.6528172,5.2847857,4.9167547,4.550536,3.6658103,2.7792716,1.8945459,1.0098201,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.55476654,1.0478923,1.5392052,2.032331,2.525457,3.3775494,4.229642,5.081734,5.9356394,6.787732,5.4896507,4.1933823,2.8953013,1.5972201,0.2991388,0.2520018,0.20486477,0.15772775,0.11059072,0.06164073,0.058014803,0.052575916,0.047137026,0.04169814,0.038072214,0.5747091,1.1131591,1.649796,2.1882458,2.7248828,3.6603715,4.59586,5.529536,6.4650245,7.400513,9.708415,12.0145035,14.322405,16.630306,18.938208,17.302916,15.667623,14.0323305,12.397038,10.761745,10.085511,9.407463,8.729415,8.05318,7.3751316,7.3896356,7.404139,7.420456,7.4349594,7.4494634,7.4476504,7.4458375,7.4422116,7.440398,7.4367723,6.200332,4.9620786,3.7256382,2.4873846,1.2491312,1.6226015,1.9942589,2.3677292,2.7393866,3.1128569,3.007705,2.902553,2.7974012,2.6922495,2.5870976,6.096993,9.606889,13.116784,16.62668,20.138388,16.82248,13.508384,10.192475,6.876567,3.5624714,4.9167547,6.2728505,7.6271334,8.98323,10.337513,8.937905,7.5382986,6.1368785,4.7372713,3.3376641,2.8155308,2.2933977,1.7694515,1.2473183,0.72518504,1.1602961,1.5954071,2.030518,2.465629,2.9007401,3.6295512,4.360175,5.090799,5.81961,6.550234,5.2630305,3.975827,2.6868105,1.3996071,0.11240368,0.11059072,0.10696479,0.10515183,0.10333887,0.099712946,0.10696479,0.11421664,0.12328146,0.13053331,0.13778515,0.1794833,0.2229944,0.26469254,0.30820364,0.34990177,0.33721104,0.3245203,0.31182957,0.2991388,0.28826106,0.30820364,0.32814622,0.3480888,0.3680314,0.387974,0.65991837,0.9318628,1.2056202,1.4775645,1.7495089,1.6280404,1.504759,1.3832904,1.260009,1.1367276,0.91917205,0.7016165,0.48587397,0.26831847,0.05076295,0.14503701,0.23931105,0.33539808,0.42967212,0.52575916,4.942136,9.360326,13.778516,18.194893,22.613083,23.387217,24.163166,24.9373,25.71325,26.487383,24.536636,22.5877,20.636953,18.688019,16.73727,15.62955,14.521831,13.41411,12.308203,11.200482,11.74981,12.299138,12.850279,13.399607,13.9507475,14.462003,14.975071,15.488139,15.999394,16.512463,16.87687,17.243088,17.607492,17.971897,18.338116,19.957092,21.57788,23.196856,24.817644,26.43662,28.13174,29.82686,31.52198,33.217102,34.91222,35.38178,35.85315,36.322704,36.792263,37.26182,32.31243,27.363045,22.411844,17.462456,12.513068,11.715364,10.917661,10.119957,9.322253,8.52455,9.808127,11.089892,12.371656,13.655234,14.936998,14.492823,14.046834,13.602658,13.15667,12.712494,12.951805,13.192928,13.43224,13.673364,13.912675,14.561715,15.212569,15.861609,16.512463,17.163317,19.157576,21.153646,23.147905,25.142164,27.138237,23.822329,20.50642,17.192324,13.878228,10.56232,10.507931,10.451729,10.397341,10.342952,10.28675,10.310318,10.332074,10.355642,10.377398,10.399154,11.028252,11.655537,12.282822,12.910107,13.537392,13.959812,14.382232,14.804652,15.227073,15.649493,13.457622,11.263937,9.072064,6.880193,4.688321,4.064662,3.442816,2.819157,2.1973107,1.5754645,2.3495996,2.3550384,2.3604772,2.3641033,2.3695421,2.374981,2.612479,2.8499773,3.0874753,3.3249733,3.5624714,6.5157876,9.467291,12.420607,15.372109,18.325426,20.468348,22.609457,24.752378,26.8953,29.038221,28.719141,28.401873,28.084604,27.767334,27.450066,27.589664,27.729263,27.870674,28.010271,28.14987,24.73425,21.32044,17.904818,14.489197,11.075388,9.690285,8.3051815,6.9200783,5.5349746,4.1498713,5.710832,7.26998,8.830941,10.390089,11.949236,12.819458,13.68968,14.559902,15.430124,16.300346,16.051971,15.805408,15.557032,15.310469,15.062093,14.284332,13.508384,12.730623,11.952863,11.175101,10.812509,10.449916,10.087324,9.724731,9.362139,9.637709,9.91328,10.1870365,10.462607,10.738177,10.337513,9.936848,9.537996,9.137331,8.736667,9.017676,9.296872,9.577881,9.857078,10.138086,10.174346,10.212419,10.25049,10.28675,10.324821,10.034748,9.744674,9.4546,9.164526,8.874452,8.479226,8.0858135,7.690587,7.2953615,6.9001355,6.6916447,6.484967,6.2782893,6.069799,5.863121,6.5194135,7.177519,7.835624,8.491917,9.1500225,8.403082,7.654328,6.9073873,6.1604466,5.411693,5.0527267,4.691947,4.3329806,3.972201,3.6132345,3.303218,2.9932013,2.6831846,2.373168,2.0631514,1.8184015,1.5718386,1.3270886,1.0823387,0.8375887,1.0333886,1.2273756,1.4231756,1.6171626,1.8129625,3.0330863,4.25321,5.473334,6.6916447,7.911769,7.4694057,7.027043,6.58468,6.1423173,5.6999545,4.5867953,3.4754493,2.3622901,1.2491312,0.13778515,2.2915847,4.4471974,6.60281,8.758422,10.912222,10.912222,10.912222,10.912222,10.912222,10.912222,10.636651,10.362894,10.087324,9.811753,9.537996,8.544493,7.552802,6.5592985,5.567608,4.574105,4.265901,3.9558845,3.6458678,3.3358512,3.0258346,3.0856624,3.1454902,3.2053177,3.2651455,3.3249733,3.6041696,3.8851788,4.164375,4.445384,4.7245803,4.690134,4.655688,4.6194286,4.5849824,4.550536,4.024777,3.5008307,2.9750717,2.4493124,1.9253663,2.3296568,2.7357605,3.1400511,3.5443418,3.9504454,3.9377546,3.925064,3.9123733,3.8996825,3.8869917,3.9975824,4.1081734,4.216951,4.327542,4.4381323,4.3982472,4.358362,4.3166637,4.2767787,4.2368937,4.177066,4.117238,4.0574102,3.9975824,3.9377546,6.19308,8.446592,10.701918,12.957244,15.212569,16.782595,18.352621,19.922646,21.492672,23.062696,22.319382,21.57788,20.834566,20.093063,19.34975,19.13582,18.920078,18.704334,18.490406,18.274662,17.5948,16.914942,16.23508,15.555219,14.875358,15.633177,16.389181,17.147,17.904818,18.662638,15.660371,12.658105,9.654026,6.6517596,3.6494937,5.527723,7.404139,9.282369,11.160598,13.037014,11.398096,9.757364,8.116633,6.4777155,4.836984,4.3347936,3.832603,3.3304121,2.8282216,2.324218,3.8597972,5.3953767,6.930956,8.464723,10.000301,8.452031,6.9055743,5.3573046,3.8108473,2.2625773,3.2669585,4.273153,5.277534,6.281915,7.28811,8.597069,9.907841,11.2168,12.527572,13.838344,11.162411,8.488291,5.812358,3.1382382,0.46230546,0.5982776,0.7324369,0.8684091,1.0025684,1.1367276,1.0279498,0.91735905,0.80676836,0.6979906,0.5873999,0.6508536,0.7124943,0.774135,0.8375887,0.89922947,0.7505665,0.6000906,0.44961473,0.2991388,0.15047589,0.13415924,0.11965553,0.10515183,0.09064813,0.07433146,0.33721104,0.6000906,0.8629702,1.1258497,1.3869164,1.1095331,0.8321498,0.55476654,0.27738327,0.0,0.19036107,0.38072214,0.56927025,0.75963134,0.9499924,1.0805258,1.209246,1.3397794,1.4703126,1.6008459,2.0957847,2.5907235,3.0856624,3.5806012,4.07554,3.925064,3.774588,3.6241121,3.4754493,3.3249733,2.666868,2.0105755,1.35247,0.69436467,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.3480888,0.69436467,1.0424535,1.3905423,1.7368182,1.3905423,1.0424535,0.69436467,0.3480888,0.0,0.581961,1.1657349,1.7476959,2.3296568,2.911618,3.8996825,4.8877473,5.8758116,6.8620634,7.850128,7.473032,7.0941224,6.717026,6.33993,5.962834,4.782595,3.6023567,2.422118,1.2418793,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.70342946,1.3415923,1.983381,2.6233568,3.2633326,3.832603,4.401873,4.972956,5.542227,6.11331,4.9693303,3.827164,2.6849976,1.5428312,0.40066472,0.33177215,0.26469254,0.19761293,0.13053331,0.06164073,0.059827764,0.058014803,0.054388877,0.052575916,0.05076295,0.53663695,1.0243238,1.5120108,1.9996977,2.4873846,3.2669585,4.0483456,4.8279195,5.6074934,6.3870673,9.135518,11.882156,14.630608,17.377247,20.125698,17.995466,15.865235,13.735004,11.6047735,9.474543,9.092008,8.709473,8.326937,7.944402,7.5618668,7.507478,7.453089,7.3968873,7.3424983,7.28811,7.217404,7.1466985,7.077806,7.0071006,6.9382076,5.774286,4.612177,3.4500678,2.2879589,1.1258497,1.4304274,1.7350051,2.039583,2.3441606,2.6505513,2.72307,2.7955883,2.8681068,2.9406252,3.0131438,6.1803894,9.347635,12.514881,15.682126,18.849373,16.017525,13.185677,10.352016,7.520169,4.688321,5.977338,7.268167,8.557183,9.848013,11.137029,9.474543,7.8120556,6.149569,4.4870825,2.8245957,2.4456866,2.0649643,1.6842422,1.305333,0.9246109,1.2418793,1.5591478,1.8782293,2.1954978,2.5127661,3.4029307,4.2930956,5.18326,6.071612,6.9617763,5.600241,4.2368937,2.8753586,1.5120108,0.15047589,0.14322405,0.13415924,0.12690738,0.11965553,0.11240368,0.12328146,0.13234627,0.14322405,0.15228885,0.16316663,0.2030518,0.24293698,0.28282216,0.32270733,0.36259252,0.33721104,0.31182957,0.28826106,0.26287958,0.2374981,0.28463513,0.33177215,0.38072214,0.42785916,0.4749962,0.7541924,1.0352017,1.3143979,1.5954071,1.8746033,1.6316663,1.3905423,1.1476053,0.90466833,0.66173136,0.53482395,0.40791658,0.27919623,0.15228885,0.025381476,0.15954071,0.2955129,0.42967212,0.5656443,0.69980353,5.239462,9.77912,14.320591,18.86025,23.399908,23.849524,24.299137,24.750565,25.20018,25.649796,23.949236,22.25049,20.54993,18.849373,17.150625,15.540715,13.930804,12.31908,10.710983,9.099259,9.300498,9.499924,9.699349,9.900589,10.100015,10.937603,11.775192,12.612781,13.45037,14.287958,15.495391,16.702824,17.910257,19.117691,20.325123,21.572441,22.81976,24.067078,25.314396,26.561714,28.010271,29.457016,30.905573,32.352318,33.800873,34.910408,36.01994,37.129475,38.240818,39.350353,34.125393,28.900436,23.675478,18.45052,13.225562,12.670795,12.114216,11.559449,11.004683,10.449916,11.472427,12.494938,13.517449,14.53996,15.56247,15.014956,14.467442,13.919927,13.372412,12.824898,13.082338,13.339779,13.597219,13.85466,14.112101,14.237195,14.362289,14.487384,14.612478,14.737573,17.823235,20.907085,23.992746,27.076595,30.162258,26.342346,22.522434,18.702522,14.882609,11.062697,10.98474,10.906783,10.830639,10.752681,10.674724,10.843329,11.010121,11.176914,11.34552,11.512312,11.820516,12.126906,12.43511,12.743314,13.049705,13.318023,13.584529,13.852847,14.119352,14.387671,12.172231,9.956791,7.743163,5.527723,3.3122826,3.007705,2.7031271,2.3967366,2.0921588,1.7875811,2.2498865,2.2371957,2.2245052,2.2118144,2.1991236,2.1882458,2.374981,2.561716,2.7502642,2.9369993,3.1255474,6.249282,9.374829,12.500377,15.625924,18.749659,20.675026,22.600391,24.525759,26.44931,28.374678,27.85073,27.324972,26.799213,26.275267,25.749508,26.06315,26.374979,26.68681,27.000452,27.31228,23.999998,20.687716,17.375433,14.06315,10.750868,9.425592,8.100317,6.775041,5.4497657,4.12449,5.712645,7.3008003,8.887142,10.475298,12.06164,12.975373,13.887294,14.799213,15.712947,16.624866,16.425442,16.224201,16.024776,15.825351,15.624111,15.049402,14.474693,13.899984,13.325275,12.750566,11.912977,11.075388,10.2378,9.400211,8.562622,8.950596,9.336758,9.724731,10.112705,10.500679,10.3502035,10.199727,10.049252,9.900589,9.750113,9.625018,9.499924,9.374829,9.249735,9.12464,9.349448,9.574255,9.800876,10.025683,10.25049,10.312131,10.375585,10.437225,10.500679,10.56232,10.138086,9.712041,9.287807,8.861761,8.437528,8.049554,7.663393,7.2754188,6.887445,6.4994707,7.250037,8.000604,8.749357,9.499924,10.25049,9.349448,8.450218,7.549176,6.6499467,5.750717,5.337362,4.9258194,4.512464,4.099108,3.6875658,3.3376641,2.9877625,2.6378605,2.2879589,1.938057,1.6878681,1.4376793,1.1874905,0.93730164,0.6871128,0.9246109,1.162109,1.3996071,1.6371052,1.8746033,3.4500678,5.0255322,6.599184,8.174648,9.750113,9.224354,8.700407,8.174648,7.650702,7.124943,5.6999545,4.274966,2.8499773,1.4249886,0.0,2.4257438,4.8496747,7.2754188,9.699349,12.125093,12.212116,12.299138,12.387974,12.474996,12.562017,12.212116,11.862214,11.512312,11.162411,10.812509,9.612328,8.412147,7.211965,6.011784,4.8116026,4.4870825,4.162562,3.8380418,3.5117085,3.1871881,3.2379513,3.2869012,3.3376641,3.386614,3.437377,3.7256382,4.0120864,4.3003473,4.5867953,4.8750563,4.7245803,4.574105,4.4254417,4.274966,4.12449,3.6748753,3.2252605,2.7756457,2.324218,1.8746033,2.3622901,2.8499773,3.3376641,3.825351,4.313038,4.2006345,4.0882306,3.975827,3.8616104,3.7492065,3.8996825,4.0501585,4.2006345,4.349297,4.499773,4.2876563,4.07554,3.8616104,3.6494937,3.437377,3.5008307,3.5624714,3.6241121,3.6875658,3.7492065,6.43783,9.12464,11.813264,14.500074,17.186886,18.338116,19.487535,20.636953,21.788185,22.937603,22.411844,21.887897,21.362139,20.838192,20.312433,20.036863,19.763105,19.487535,19.211964,18.938208,18.062546,17.186886,16.313038,15.437376,14.561715,15.986704,17.411694,18.836681,20.26167,21.686659,18.238403,14.788336,11.338268,7.8882003,4.4381323,6.1006193,7.763106,9.425592,11.088079,12.750566,10.975676,9.200785,7.424082,5.6491914,3.874301,3.636803,3.3993049,3.1618068,2.9243085,2.6868105,3.5008307,4.313038,5.125245,5.9374523,6.7496595,5.612932,4.4743915,3.3376641,2.1991236,1.062396,1.649796,2.2371957,2.8245957,3.4119956,3.9993954,4.974769,5.9501433,6.925517,7.900891,8.874452,7.137634,5.4008155,3.6621845,1.9253663,0.18673515,0.41335547,0.63816285,0.8629702,1.0877775,1.3125849,1.1258497,0.93730164,0.7505665,0.5620184,0.37528324,0.46230546,0.5493277,0.63816285,0.72518504,0.8122072,0.6508536,0.48768693,0.3245203,0.16316663,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.37528324,0.6871128,1.0007553,1.3125849,1.6244144,1.2998942,0.97537386,0.6508536,0.3245203,0.0,0.22480737,0.44961473,0.6744221,0.89922947,1.1258497,0.9119202,0.69980353,0.48768693,0.2755703,0.06164073,1.0134461,1.9616255,2.913431,3.8616104,4.8116026,4.6629395,4.512464,4.361988,4.213325,4.062849,3.2506418,2.4366217,1.6244144,0.8122072,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.31182957,0.62547207,0.93730164,1.2491312,1.5627737,1.2491312,0.93730164,0.62547207,0.31182957,0.0,0.72518504,1.4503701,2.175555,2.9007401,3.6241121,4.762653,5.89938,7.037921,8.174648,9.313189,8.925215,8.537241,8.149267,7.763106,7.3751316,5.89938,4.4254417,2.94969,1.4757515,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.85027945,1.6371052,2.4257438,3.2125697,3.9993954,4.2876563,4.574105,4.8623657,5.1506267,5.4370747,4.4508233,3.4627585,2.474694,1.4866294,0.50037766,0.41335547,0.3245203,0.2374981,0.15047589,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.50037766,0.93730164,1.3742256,1.8129625,2.2498865,2.8753586,3.5008307,4.12449,4.749962,5.375434,8.562622,11.74981,14.936998,18.124187,21.313189,18.688019,16.062849,13.437678,10.812509,8.187339,8.100317,8.013294,7.9244595,7.837437,7.750415,7.6253204,7.500226,7.3751316,7.250037,7.124943,6.987158,6.849373,6.7134004,6.5756154,6.43783,5.3500524,4.262275,3.1744974,2.08672,1.0007553,1.2382535,1.4757515,1.7132497,1.9507477,2.1882458,2.4366217,2.6868105,2.9369993,3.1871881,3.437377,6.261973,9.086569,11.912977,14.737573,17.562168,15.212569,12.862969,10.511557,8.161958,5.812358,7.037921,8.26167,9.487233,10.712796,11.938358,10.012992,8.087626,6.16226,4.2368937,2.3133402,2.0758421,1.8383441,1.6008459,1.3633479,1.1258497,1.3252757,1.5247015,1.7241274,1.9253663,2.124792,3.1744974,4.2242026,5.275721,6.3254266,7.3751316,5.9374523,4.499773,3.0620937,1.6244144,0.18673515,0.17585737,0.16316663,0.15047589,0.13778515,0.12509441,0.13778515,0.15047589,0.16316663,0.17585737,0.18673515,0.22480737,0.26287958,0.2991388,0.33721104,0.37528324,0.33721104,0.2991388,0.26287958,0.22480737,0.18673515,0.26287958,0.33721104,0.41335547,0.48768693,0.5620184,0.85027945,1.1367276,1.4249886,1.7132497,1.9996977,1.6371052,1.2745126,0.9119202,0.5493277,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.17585737,0.34990177,0.52575916,0.69980353,0.87566096,5.538601,10.199727,14.862667,19.525606,24.186733,24.311829,24.436922,24.562017,24.68711,24.812206,23.361835,21.913279,20.462908,19.012539,17.562168,15.4500675,13.337966,11.224051,9.11195,6.9998484,6.849373,6.70071,6.550234,6.399758,6.249282,7.413204,8.575313,9.737422,10.899531,12.06164,14.112101,16.162561,18.213022,20.26167,22.31213,23.187792,24.06164,24.9373,25.812962,26.68681,27.88699,29.087172,30.287354,31.487534,32.687714,34.437225,36.186733,37.938053,39.687565,41.437073,35.936543,30.437828,24.9373,19.438585,13.938056,13.6244135,13.312584,13.000754,12.687112,12.375282,13.136727,13.899984,14.663241,15.4246855,16.187943,15.537089,14.888049,14.237195,13.588155,12.937301,13.212872,13.486629,13.762199,14.037769,14.313339,13.912675,13.512011,13.113158,12.712494,12.311829,16.487082,20.662334,24.837587,29.01284,33.18809,28.862364,24.536636,20.212719,15.8869915,11.563075,11.463363,11.361836,11.262123,11.162411,11.062697,11.374527,11.6881695,11.999999,12.311829,12.625471,12.612781,12.60009,12.5873995,12.574709,12.562017,12.674421,12.786825,12.899229,13.011633,13.125849,10.88684,8.649645,6.412449,4.175253,1.938057,1.9507477,1.9616255,1.9743162,1.987007,1.9996977,2.3876717,2.4003625,2.4130533,2.4257438,2.4366217,2.4493124,2.5526514,2.6541772,2.7575161,2.8608549,2.962381,5.9447045,8.927028,11.909351,14.891675,17.87581,19.922646,21.96948,24.018127,26.064962,28.111797,27.430124,26.746637,26.064962,25.38329,24.699802,25.082336,25.464872,25.847408,26.229942,26.612478,23.075388,19.538298,15.999394,12.462305,8.925215,7.8882003,6.849373,5.812358,4.7753434,3.738329,5.1198063,6.5030966,7.8845744,9.267865,10.649343,11.689982,12.730623,13.769451,14.810091,15.850732,15.821725,15.79453,15.767336,15.740141,15.712947,15.431937,15.152741,14.871732,14.592536,14.313339,13.172986,12.032633,10.89228,9.751925,8.613385,8.939718,9.267865,9.594198,9.922344,10.25049,9.976733,9.704789,9.432844,9.1609,8.887142,8.660522,8.432089,8.205468,7.9770355,7.750415,7.989726,8.23085,8.470161,8.709473,8.950596,9.354887,9.759177,10.165281,10.5695715,10.975676,11.077202,11.18054,11.282066,11.385405,11.486931,11.466989,11.447045,11.427103,11.407161,11.3872175,11.30926,11.233116,11.155159,11.077202,10.999244,9.945912,8.890768,7.835624,6.78048,5.7253356,5.2467136,4.7699046,4.2930956,3.8144734,3.3376641,3.1182957,2.8971143,2.6777458,2.4583774,2.2371957,2.2825198,2.327844,2.373168,2.4166791,2.4620032,2.5870976,2.712192,2.8372865,2.962381,3.0874753,4.6266804,6.167699,7.706904,9.247922,10.7871275,9.960417,9.131892,8.3051815,7.476658,6.6499467,5.3246713,3.9993954,2.6741197,1.3506571,0.025381476,2.3423476,4.6593137,6.978093,9.295059,11.612025,11.9601145,12.308203,12.654479,13.002567,13.3506565,13.009819,12.670795,12.329959,11.989121,11.650098,10.484363,9.32044,8.154706,6.9907837,5.825049,5.389938,4.954827,4.519716,4.0846047,3.6494937,3.5951047,3.540716,3.484514,3.4301252,3.3757362,3.7056956,4.0356545,4.365614,4.695573,5.0255322,4.893186,4.76084,4.6266804,4.494334,4.361988,3.9377546,3.5117085,3.0874753,2.663242,2.2371957,2.7266958,3.2180085,3.7075086,4.1970086,4.688321,4.507025,4.327542,4.1480584,3.966762,3.787279,3.9558845,4.122677,4.2894692,4.458075,4.6248674,4.499773,4.3746786,4.249584,4.12449,3.9993954,3.9903307,3.9794528,3.9703882,3.9595103,3.9504454,6.497658,9.04487,11.592083,14.139296,16.68832,17.932013,19.177519,20.423023,21.666716,22.912222,22.264994,21.617765,20.97054,20.32331,19.67427,19.75948,19.844688,19.929897,20.015106,20.100317,18.82943,17.560356,16.289469,15.020395,13.749508,14.86448,15.979452,17.094423,18.209396,19.324368,16.29672,13.270886,10.243238,7.215591,4.1879435,5.5857377,6.981719,8.379513,9.7773075,11.175101,9.935035,8.694968,7.454902,6.2148356,4.974769,4.8696175,4.764466,4.6593137,4.554162,4.4508233,4.9693303,5.4896507,6.009971,6.530291,7.0506115,6.0770507,5.105303,4.1317415,3.159994,2.1882458,2.474694,2.762955,3.049403,3.3376641,3.6241121,4.439945,5.2557783,6.069799,6.885632,7.699652,6.338117,4.974769,3.6132345,2.2498865,0.8883517,1.1040943,1.3216497,1.5392052,1.7567607,1.9743162,1.7277533,1.4793775,1.2328146,0.98443866,0.73787576,0.83033687,0.922798,1.015259,1.1077201,1.2001812,0.9644961,0.7306239,0.4949388,0.25925365,0.025381476,0.045324065,0.065266654,0.08520924,0.10515183,0.12509441,0.5148814,0.90466833,1.2944553,1.6842422,2.0758421,1.845596,1.6153497,1.3851035,1.1548572,0.9246109,1.0497054,1.1747998,1.2998942,1.4249886,1.550083,1.3651608,1.1802386,0.99531645,0.8103943,0.62547207,1.3796645,2.13567,2.8898623,3.6458678,4.40006,4.1879435,3.975827,3.7618973,3.5497808,3.3376641,2.6704938,2.0033236,1.3343405,0.6671702,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03988518,0.07977036,0.11965553,0.15954071,0.19942589,0.15954071,0.11965553,0.07977036,0.03988518,0.0,0.25018883,0.50037766,0.7505665,1.0007553,1.2491312,1.0007553,0.7505665,0.50037766,0.25018883,0.0,0.58014804,1.1602961,1.7404441,2.3205922,2.9007401,3.8380418,4.7753434,5.712645,6.6499467,7.5872483,7.304426,7.021604,6.740595,6.4577727,6.1749506,5.42801,4.6792564,3.9323158,3.1853752,2.4366217,1.9598125,1.4830034,1.0043813,0.5275721,0.05076295,0.052575916,0.054388877,0.058014803,0.059827764,0.06164073,0.072518505,0.08339628,0.092461094,0.10333887,0.11240368,0.8194591,1.5283275,2.2353828,2.9424384,3.6494937,3.8507326,4.0501585,4.249584,4.4508233,4.650249,3.8054085,2.960568,2.1157274,1.2708868,0.42423326,0.35171473,0.27919623,0.20667773,0.13415924,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.41335547,0.76325727,1.1131591,1.4630609,1.8129625,2.3695421,2.9279346,3.484514,4.0429068,4.599486,7.135821,9.670342,12.2048645,14.739386,17.27572,15.250641,13.225562,11.200482,9.175404,7.1503243,7.1648283,7.179332,7.1956487,7.210152,7.224656,7.0868707,6.9508986,6.813113,6.6753283,6.5375433,6.640882,6.742408,6.8457465,6.947273,7.0506115,5.8323007,4.615803,3.397492,2.179181,0.96268314,1.260009,1.5573349,1.8546607,2.1519866,2.4493124,2.6052272,2.759329,2.9152439,3.0693457,3.2252605,6.169512,9.115576,12.059827,15.005891,17.950142,16.739084,15.529838,14.320591,13.109532,11.900287,11.735307,11.570327,11.405348,11.240368,11.075388,9.2606125,7.4458375,5.6292486,3.8144734,1.9996977,1.8093367,1.6207886,1.4304274,1.2400664,1.0497054,1.2473183,1.4449311,1.6425442,1.840157,2.03777,3.350355,4.6629395,5.975525,7.28811,8.600695,6.9182653,5.235836,3.5515938,1.8691645,0.18673515,0.17767033,0.16679256,0.15772775,0.14684997,0.13778515,0.15228885,0.16679256,0.18310922,0.19761293,0.21211663,0.23024625,0.24837588,0.26469254,0.28282216,0.2991388,0.27013144,0.23931105,0.21030366,0.1794833,0.15047589,0.24474995,0.34083697,0.43511102,0.5293851,0.62547207,0.82671094,1.0297627,1.2328146,1.4358664,1.6371052,1.3397794,1.0424535,0.7451276,0.44780177,0.15047589,0.24474995,0.34083697,0.43511102,0.5293851,0.62547207,1.1421664,1.6606737,2.1773682,2.6958754,3.2125697,7.1031876,10.991992,14.882609,18.771414,22.662033,22.872335,23.08264,23.292944,23.503246,23.711737,22.049252,20.386765,18.724277,17.06179,15.399304,13.517449,11.635593,9.751925,7.8700705,5.9882154,5.826862,5.667321,5.5077806,5.3482394,5.186886,6.298232,7.407765,8.517298,9.626831,10.738177,13.029762,15.32316,17.614744,19.908142,22.199726,22.75812,23.3147,23.87309,24.42967,24.988064,26.083092,27.178122,28.273151,29.368181,30.463211,32.265297,34.06738,35.869465,37.67155,39.47545,34.77806,30.080675,25.381475,20.685904,15.986704,15.544341,15.101978,14.6596155,14.217253,13.77489,14.376793,14.98051,15.582414,16.184317,16.788034,16.117237,15.448255,14.777458,14.106662,13.437678,13.637105,13.838344,14.037769,14.237195,14.436621,13.961625,13.486629,13.011633,12.536636,12.06164,16.450823,20.838192,25.225561,29.61293,34.0003,30.457771,26.915243,23.372713,19.830185,16.287657,16.177065,16.068287,15.957697,15.847106,15.738328,14.960567,14.182806,13.4050455,12.627284,11.849524,12.203052,12.554766,12.908294,13.260008,13.611723,13.318023,13.022511,12.726997,12.433297,12.137785,10.067381,7.996978,5.9265747,3.8579843,1.7875811,1.8582866,1.9271792,1.9978848,2.0667772,2.137483,2.525457,2.561716,2.5997884,2.6378605,2.6741197,2.712192,2.7303216,2.7466383,2.764768,2.7828975,2.7992141,5.6401267,8.479226,11.320138,14.159238,17.00015,19.170267,21.340382,23.510498,25.680614,27.85073,27.009516,26.170115,25.330713,24.489498,23.650097,24.103338,24.554766,25.008005,25.459433,25.912674,22.150776,18.387066,14.625169,10.863272,7.0995617,6.350808,5.600241,4.8496747,4.099108,3.350355,4.5269675,5.7053933,6.882006,8.0604315,9.237044,10.4045925,11.57214,12.739688,13.907236,15.074784,15.219821,15.364858,15.509895,15.654932,15.799969,15.814472,15.83079,15.845293,15.859797,15.8743,14.432995,12.989877,11.546759,10.1054535,8.662335,8.930654,9.197159,9.465478,9.731983,10.000301,9.605076,9.20985,8.814624,8.419398,8.024173,7.6942134,7.364254,7.0342946,6.7043357,6.3743763,6.630004,6.885632,7.1394467,7.3950744,7.650702,8.397643,9.144584,9.893337,10.640278,11.3872175,12.018129,12.647227,13.278138,13.907236,14.538147,14.884423,15.2325115,15.580601,15.926876,16.274965,15.3702965,14.465629,13.559147,12.654479,11.74981,10.540565,9.329506,8.120259,6.9092,5.6999545,5.1578784,4.615803,4.071914,3.529838,2.9877625,2.8971143,2.808279,2.7176309,2.6269827,2.5381477,2.8771715,3.2180085,3.5570326,3.8978696,4.2368937,4.249584,4.262275,4.274966,4.2876563,4.3003473,5.805106,7.309865,8.814624,10.319383,11.8241415,10.694666,9.56519,8.435715,7.304426,6.1749506,4.949388,3.7256382,2.5000753,1.2745126,0.05076295,2.2607644,4.4707656,6.680767,8.890768,11.10077,11.708113,12.3154545,12.922797,13.53014,14.137483,13.807523,13.477564,13.147605,12.817645,12.487686,11.358211,10.226922,9.097446,7.9679704,6.836682,6.2927933,5.7470913,5.2032027,4.6575007,4.1117992,3.9522583,3.7927177,3.633177,3.4718235,3.3122826,3.6857529,4.0574102,4.4308805,4.802538,5.1741953,5.0599785,4.945762,4.8297324,4.7155156,4.599486,4.2006345,3.7999697,3.3993049,3.000453,2.5997884,3.092914,3.584227,4.077353,4.5704784,5.0617914,4.8152285,4.5668526,4.3202896,4.071914,3.825351,4.0102735,4.195195,4.3801174,4.5650396,4.749962,4.7118897,4.6756306,4.6375585,4.599486,4.5632267,4.4798307,4.3982472,4.314851,4.233268,4.1498713,6.5574856,8.9651,11.372714,13.780329,16.187943,17.527721,18.867502,20.207281,21.54706,22.886839,22.118143,21.347635,20.577126,19.806616,19.03792,19.482096,19.928085,20.372261,20.818249,21.262424,19.598125,17.932013,16.267714,14.601601,12.937301,13.742256,14.547212,15.352167,16.157122,16.962078,14.356851,11.753436,9.14821,6.542982,3.9377546,5.0708566,6.202145,7.3352466,8.4683485,9.599637,8.894395,8.189152,7.4857225,6.78048,6.0752378,6.1024323,6.1296263,6.156821,6.185828,6.2130227,6.439643,6.6680765,6.8946967,7.12313,7.3497505,6.542982,5.7344007,4.9276323,4.120864,3.3122826,3.299592,3.2869012,3.2742105,3.2633326,3.2506418,3.9051213,4.559601,5.2158933,5.870373,6.5248523,5.5367875,4.550536,3.5624714,2.5744069,1.5881553,1.7966459,2.0069497,2.2172532,2.427557,2.6378605,2.3296568,2.0232663,1.7150626,1.4068589,1.1004683,1.1983683,1.2944553,1.3923552,1.4902552,1.5881553,1.2799516,0.97174793,0.6653573,0.35715362,0.05076295,0.07795739,0.10515183,0.13234627,0.15954071,0.18673515,0.6544795,1.1222239,1.5899682,2.0577126,2.525457,2.3894846,2.2553256,2.1193533,1.9851941,1.8492218,1.8746033,1.8999848,1.9253663,1.9507477,1.9743162,1.8165885,1.6606737,1.502946,1.3452182,1.1874905,1.7476959,2.3079014,2.8681068,3.4283123,3.9867048,3.7129474,3.437377,3.1618068,2.8880494,2.612479,2.0903459,1.5682126,1.0442665,0.52213323,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.04169814,0.08520924,0.12690738,0.17041849,0.21211663,0.17041849,0.12690738,0.08520924,0.04169814,0.0,0.18673515,0.37528324,0.5620184,0.7505665,0.93730164,0.7505665,0.5620184,0.37528324,0.18673515,0.0,0.43511102,0.87022203,1.305333,1.7404441,2.175555,2.913431,3.6494937,4.3873696,5.125245,5.863121,5.6854506,5.5077806,5.33011,5.1524396,4.974769,4.954827,4.934884,4.914942,4.894999,4.8750563,3.9069343,2.9406252,1.9725033,1.0043813,0.038072214,0.04169814,0.047137026,0.052575916,0.058014803,0.06164073,0.08339628,0.10333887,0.12328146,0.14322405,0.16316663,0.7904517,1.4177368,2.0450218,2.6723068,3.299592,3.4119956,3.5243993,3.636803,3.7492065,3.8616104,3.159994,2.4583774,1.7549478,1.0533313,0.34990177,0.291887,0.23568514,0.17767033,0.11965553,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.3245203,0.5873999,0.85027945,1.1131591,1.3742256,1.8655385,2.3550384,2.8445382,3.3358512,3.825351,5.7072062,7.5890613,9.47273,11.354585,13.238253,11.813264,10.388275,8.963287,7.5382986,6.11331,6.2293396,6.347182,6.4650245,6.582867,6.70071,6.550234,6.399758,6.249282,6.1006193,5.9501433,6.2927933,6.635443,6.978093,7.320743,7.663393,6.3145485,4.9675174,3.6204863,2.2716422,0.9246109,1.2817645,1.6407311,1.9978848,2.3550384,2.712192,2.7720199,2.8318477,2.8916752,2.953316,3.0131438,6.0770507,9.142771,12.20849,15.272397,18.338116,18.26741,18.196705,18.127813,18.057108,17.988214,16.432693,14.877171,13.321649,11.7679405,10.212419,8.508233,6.8022356,5.0980506,3.392053,1.6878681,1.5446441,1.403233,1.260009,1.1167849,0.97537386,1.1693609,1.3651608,1.5591478,1.7549478,1.9507477,3.5243993,5.0998635,6.6753283,8.2507925,9.824444,7.897265,5.9700856,4.0429068,2.1157274,0.18673515,0.1794833,0.17223145,0.16497959,0.15772775,0.15047589,0.16679256,0.18492219,0.2030518,0.21936847,0.2374981,0.23568514,0.23205921,0.23024625,0.22662032,0.22480737,0.2030518,0.1794833,0.15772775,0.13415924,0.11240368,0.22662032,0.34264994,0.45686656,0.5728962,0.6871128,0.80495536,0.922798,1.0406405,1.1566701,1.2745126,1.0424535,0.8103943,0.57833505,0.3444629,0.11240368,0.34083697,0.56745726,0.79589057,1.0225109,1.2491312,2.1102884,2.9696326,3.83079,4.690134,5.5494785,8.667774,11.784257,14.902553,18.019035,21.137331,21.432844,21.728357,22.022057,22.31757,22.613083,20.736666,18.862062,16.98746,15.112856,13.238253,11.584831,9.933222,8.2798,6.628191,4.974769,4.804351,4.6357455,4.465327,4.2949085,4.12449,5.18326,6.240217,7.2971745,8.354132,9.412902,11.947423,14.481945,17.01828,19.552801,22.087322,22.326633,22.567759,22.80707,23.048193,23.287504,24.277382,25.26726,26.257137,27.247015,28.236893,30.093367,31.948027,33.80269,35.65735,37.51201,33.617764,29.723522,25.827465,21.933222,18.037165,17.464268,16.893185,16.32029,15.747393,15.174497,15.616859,16.059223,16.503399,16.94576,17.388124,16.697386,16.006647,15.31772,14.626982,13.938056,14.06315,14.188245,14.313339,14.436621,14.561715,14.012388,13.46306,12.91192,12.362592,11.813264,16.41275,21.012236,25.613535,30.213022,34.812508,32.053177,29.292036,26.532707,23.773378,21.012236,20.89258,20.772924,20.653269,20.531801,20.412146,18.544794,16.677443,14.810091,12.9427395,11.075388,11.793322,12.509441,13.227375,13.945308,14.663241,13.959812,13.258195,12.554766,11.853149,11.14972,9.247922,7.344311,5.4425135,3.540716,1.6371052,1.7658255,1.892733,2.0196402,2.1483607,2.275268,2.663242,2.7248828,2.7883365,2.8499773,2.911618,2.9750717,2.907992,2.8390994,2.7720199,2.70494,2.6378605,5.335549,8.033237,10.730926,13.426801,16.124489,18.417887,20.70947,23.002869,25.294455,27.587852,26.590723,25.59178,24.59465,23.59752,22.600391,23.122524,23.644657,24.166792,24.690737,25.212872,21.224354,17.237648,13.24913,9.262425,5.275721,4.8116026,4.349297,3.8869917,3.4246864,2.962381,3.9341288,4.9076896,5.8794374,6.8529987,7.8247466,9.119202,10.41547,11.709926,13.00438,14.300649,14.617917,14.935185,15.252454,15.569723,15.8869915,16.197008,16.507025,16.817041,17.127058,17.437075,15.693004,13.947122,12.203052,10.457169,8.713099,8.919776,9.128266,9.334945,9.541622,9.750113,9.231606,8.714911,8.198216,7.6797094,7.1630154,6.7297173,6.298232,5.864934,5.431636,5.0001507,5.2702823,5.540414,5.810545,6.0806766,6.350808,7.440398,8.529989,9.619579,10.70917,11.800573,12.957244,14.115726,15.272397,16.43088,17.58755,18.301857,19.017977,19.732285,20.448404,21.162712,19.42952,17.698141,15.964949,14.231756,12.500377,11.135216,9.770056,8.404895,7.039734,5.674573,5.06723,4.459888,3.8525455,3.245203,2.6378605,2.6777458,2.7176309,2.7575161,2.7974012,2.8372865,3.4718235,4.1081734,4.74271,5.377247,6.011784,5.9120708,5.812358,5.712645,5.612932,5.5132194,6.981719,8.452031,9.922344,11.392657,12.862969,11.430729,9.9966755,8.564435,7.132195,5.6999545,4.5759177,3.4500678,2.324218,1.2001812,0.07433146,2.1773682,4.2804046,6.3834414,8.484665,10.587702,11.454298,12.322706,13.189302,14.057712,14.924308,14.6052265,14.284332,13.965251,13.644357,13.325275,12.230246,11.135216,10.040187,8.945157,7.850128,7.1956487,6.539356,5.8848767,5.230397,4.574105,4.309412,4.0447197,3.780027,3.5153344,3.2506418,3.6658103,4.079166,4.494334,4.9095025,5.3246713,5.2267714,5.130684,5.032784,4.934884,4.836984,4.461701,4.0882306,3.7129474,3.3376641,2.962381,3.4573197,3.9522583,4.4471974,4.942136,5.4370747,5.121619,4.8079767,4.4925213,4.177066,3.8616104,4.064662,4.267714,4.4707656,4.6720047,4.8750563,4.9258194,4.974769,5.0255322,5.0744824,5.125245,4.9693303,4.8152285,4.6593137,4.505212,4.349297,6.6173134,8.885329,11.153346,13.419549,15.687565,17.121618,18.557486,19.993351,21.427404,22.863272,21.96948,21.077503,20.185526,19.291735,18.399757,19.204712,20.009668,20.814623,21.61958,22.424534,20.36501,18.305483,16.244144,14.184619,12.125093,12.620032,13.114971,13.60991,14.104849,14.599788,12.416981,10.234174,8.05318,5.870373,3.6875658,4.554162,5.422571,6.2891674,7.157576,8.024173,7.855567,7.6851482,7.51473,7.344311,7.175706,7.3352466,7.494787,7.654328,7.8156815,7.9752226,7.909956,7.844689,7.7794223,7.7141557,7.650702,7.0071006,6.3653116,5.7217097,5.0799212,4.4381323,4.12449,3.8126602,3.5008307,3.1871881,2.8753586,3.3702974,3.8652363,4.360175,4.855114,5.3500524,4.7372713,4.12449,3.5117085,2.9007401,2.2879589,2.4891977,2.6922495,2.8953013,3.0983531,3.299592,2.9333735,2.565342,2.1973107,1.8292793,1.4630609,1.5645868,1.6679256,1.7694515,1.8727903,1.9743162,1.5954071,1.214685,0.83577573,0.4550536,0.07433146,0.11059072,0.14503701,0.1794833,0.21574254,0.25018883,0.79589057,1.3397794,1.8854811,2.42937,2.9750717,2.9351864,2.8953013,2.855416,2.8155308,2.7756457,2.6995013,2.6251698,2.5508385,2.474694,2.4003625,2.269829,2.1392958,2.0105755,1.8800422,1.7495089,2.1157274,2.4801328,2.8445382,3.2107568,3.5751622,3.2379513,2.9007401,2.561716,2.2245052,1.887294,1.5101979,1.1331016,0.7541924,0.3770962,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.045324065,0.09064813,0.13415924,0.1794833,0.22480737,0.1794833,0.13415924,0.09064813,0.045324065,0.0,0.12509441,0.25018883,0.37528324,0.50037766,0.62547207,0.50037766,0.37528324,0.25018883,0.12509441,0.0,0.29007402,0.58014804,0.87022203,1.1602961,1.4503701,1.987007,2.525457,3.0620937,3.6005437,4.137181,4.064662,3.9921436,3.919625,3.8471067,3.774588,4.4816437,5.1905117,5.8975673,6.604623,7.311678,5.8540564,4.3982472,2.9406252,1.4830034,0.025381476,0.032633327,0.03988518,0.047137026,0.054388877,0.06164073,0.092461094,0.12328146,0.15228885,0.18310922,0.21211663,0.75963134,1.3071461,1.8546607,2.4021754,2.94969,2.9750717,3.000453,3.0258346,3.049403,3.0747845,2.514579,1.9543737,1.3941683,0.83577573,0.2755703,0.23205921,0.19036107,0.14684997,0.10515183,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.2374981,0.41335547,0.5873999,0.76325727,0.93730164,1.3597219,1.7821422,2.2045624,2.6269827,3.049403,4.2804046,5.5095935,6.740595,7.9697833,9.200785,8.374074,7.549176,6.7242785,5.89938,5.0744824,5.295664,5.5150323,5.7344007,5.955582,6.1749506,6.011784,5.8504305,5.6872635,5.524097,5.3627434,5.9447045,6.526665,7.1104393,7.6924005,8.274362,6.796797,5.319232,3.8416677,2.3641033,0.8883517,1.305333,1.7223145,2.1392958,2.5580902,2.9750717,2.9406252,2.904366,2.8699198,2.8354735,2.7992141,5.9845896,9.169965,12.35534,15.540715,18.724277,19.795738,20.865387,21.935034,23.004683,24.07433,21.13008,18.185827,15.239763,12.295512,9.349448,7.754041,6.1604466,4.5650396,2.9696326,1.3742256,1.2799516,1.1856775,1.0895905,0.99531645,0.89922947,1.0932164,1.2853905,1.4775645,1.6697385,1.8619126,3.7002566,5.5367875,7.3751316,9.211663,11.050007,8.8780775,6.7043357,4.5324063,2.3604772,0.18673515,0.18310922,0.17767033,0.17223145,0.16679256,0.16316663,0.18310922,0.2030518,0.2229944,0.24293698,0.26287958,0.23931105,0.21755551,0.19579996,0.17223145,0.15047589,0.13415924,0.11965553,0.10515183,0.09064813,0.07433146,0.21030366,0.3444629,0.48043507,0.61459434,0.7505665,0.78319985,0.81583315,0.8466535,0.8792868,0.9119202,0.7451276,0.57833505,0.40972954,0.24293698,0.07433146,0.43511102,0.79589057,1.1548572,1.5156367,1.8746033,3.0784104,4.2804046,5.482399,6.684393,7.8882003,10.232361,12.578335,14.922495,17.266655,19.612629,19.993351,20.372261,20.752983,21.131891,21.512613,19.424082,17.33736,15.250641,13.162108,11.075388,9.652213,8.23085,6.8076744,5.384499,3.9631362,3.7818398,3.6023567,3.4228733,3.24339,3.0620937,4.068288,5.0726695,6.0770507,7.083245,8.087626,10.865085,13.642544,16.420002,19.19746,21.97492,21.896961,21.820818,21.74286,21.664904,21.586945,22.471672,23.35821,24.242935,25.12766,26.012386,27.919624,29.82686,31.73591,33.643147,35.550385,32.45747,29.364555,26.27164,23.18054,20.087626,19.384195,18.682579,17.97915,17.277533,16.575916,16.856926,17.139748,17.422571,17.705393,17.988214,17.277533,16.566853,15.857984,15.147303,14.436621,14.487384,14.538147,14.587097,14.63786,14.68681,14.06315,13.437678,12.812206,12.186734,11.563075,16.374678,21.188093,25.999697,30.813112,35.624714,33.646774,31.670643,29.692701,27.71476,25.736816,25.608097,25.477564,25.34703,25.21831,25.087776,22.12902,19.17208,16.215137,13.258195,10.29944,11.381779,12.465931,13.548269,14.630608,15.712947,14.601601,13.492067,12.382534,11.273002,10.161655,8.42665,6.6916447,4.95664,3.2234476,1.4866294,1.6733645,1.8582866,2.0432088,2.228131,2.4130533,2.7992141,2.8880494,2.9750717,3.0620937,3.149116,3.2379513,3.0856624,2.9333735,2.7792716,2.6269827,2.474694,5.029158,7.5854354,10.139899,12.694364,15.250641,17.665508,20.080374,22.49524,24.910107,27.324972,26.170115,25.015257,23.860401,22.705544,21.550686,22.141712,22.73455,23.327389,23.920229,24.513067,20.299742,16.08823,11.874905,7.66158,3.4500678,3.2742105,3.100166,2.9243085,2.7502642,2.5744069,3.343103,4.1099863,4.876869,5.6455655,6.412449,7.835624,9.256987,10.680162,12.103338,13.524701,14.014201,14.505513,14.995013,15.484513,15.975826,16.579542,17.185072,17.790602,18.394318,18.999847,16.953012,14.904366,12.857531,10.810696,8.762048,8.910711,9.057561,9.2044115,9.353074,9.499924,8.859948,8.219973,7.5799966,6.9400206,6.300045,5.765221,5.230397,4.695573,4.160749,3.6241121,3.9105604,4.195195,4.4798307,4.764466,5.049101,6.4831543,7.915395,9.347635,10.779876,12.212116,13.898171,15.582414,17.266655,18.952711,20.636953,21.719292,22.80163,23.885782,24.96812,26.050459,23.490557,20.930653,18.37075,15.810846,13.24913,11.729868,10.210606,8.689529,7.170267,5.6491914,4.9783955,4.305786,3.633177,2.960568,2.2879589,2.4583774,2.6269827,2.7974012,2.9678197,3.1382382,4.068288,4.9983377,5.9283876,6.8566246,7.7866745,7.574558,7.362441,7.1503243,6.9382076,6.7242785,8.160145,9.594198,11.030065,12.464118,13.899984,12.164979,10.429974,8.694968,6.9599633,5.224958,4.2006345,3.1744974,2.1501737,1.1258497,0.099712946,2.0957847,4.0900435,6.0843024,8.080374,10.074633,11.202296,12.329959,13.457622,14.585284,15.712947,15.40293,15.092914,14.782897,14.47288,14.162864,13.102281,12.0416975,10.982927,9.922344,8.861761,8.096691,7.3316207,6.5683637,5.803293,5.038223,4.668379,4.2967215,3.926877,3.5570326,3.1871881,3.6458678,4.102734,4.559601,5.0182805,5.475147,5.3953767,5.315606,5.235836,5.1542525,5.0744824,4.7245803,4.3746786,4.024777,3.6748753,3.3249733,3.8217251,4.3202896,4.8170414,5.315606,5.812358,5.429823,5.047288,4.664753,4.2822175,3.8996825,4.120864,4.3402324,4.559601,4.780782,5.0001507,5.137936,5.275721,5.411693,5.5494785,5.6872635,5.4606433,5.23221,5.0055895,4.7771564,4.550536,6.677141,8.805559,10.932164,13.060582,15.187187,16.717327,18.247469,19.777609,21.307749,22.837889,21.82263,20.807371,19.792112,18.776854,17.763407,18.92733,20.093063,21.256987,22.422722,23.586643,21.131891,18.677141,16.22239,13.767638,11.312886,11.497808,11.682731,11.867653,12.052575,12.237497,10.477111,8.716724,6.9581504,5.197764,3.437377,4.0392804,4.6429973,5.2449007,5.846804,6.450521,6.814926,7.179332,7.5455503,7.909956,8.274362,8.568061,8.859948,9.151835,9.445535,9.737422,9.380268,9.023115,8.664148,8.306994,7.949841,7.473032,6.9944096,6.5176005,6.0407915,5.562169,4.949388,4.3384194,3.7256382,3.1128569,2.5000753,2.8354735,3.1708715,3.5044568,3.8398547,4.175253,3.9377546,3.7002566,3.4627585,3.2252605,2.9877625,3.1817493,3.3775494,3.5733492,3.7673361,3.9631362,3.5352771,3.1074178,2.6795588,2.2516994,1.8256533,1.9326181,2.039583,2.1483607,2.2553256,2.3622901,1.9108626,1.4576219,1.0043813,0.5529536,0.099712946,0.14322405,0.18492219,0.22662032,0.27013144,0.31182957,0.9354887,1.5573349,2.179181,2.8028402,3.4246864,3.4808881,3.5352771,3.589666,3.6458678,3.7002566,3.5243993,3.350355,3.1744974,3.000453,2.8245957,2.72307,2.619731,2.518205,2.4148662,2.3133402,2.4819458,2.6523643,2.8227828,2.9932013,3.1618068,2.762955,2.3622901,1.9616255,1.5627737,1.162109,0.9300498,0.6979906,0.46411842,0.23205921,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.047137026,0.09427405,0.14322405,0.19036107,0.2374981,0.19036107,0.14322405,0.09427405,0.047137026,0.0,0.06164073,0.12509441,0.18673515,0.25018883,0.31182957,0.25018883,0.18673515,0.12509441,0.06164073,0.0,0.14503701,0.29007402,0.43511102,0.58014804,0.72518504,1.062396,1.3996071,1.7368182,2.0758421,2.4130533,2.4456866,2.47832,2.5091403,2.5417736,2.5744069,4.0102735,5.4443264,6.880193,8.314246,9.750113,7.802991,5.8558693,3.9069343,1.9598125,0.012690738,0.02175555,0.032633327,0.04169814,0.052575916,0.06164073,0.10333887,0.14322405,0.18310922,0.2229944,0.26287958,0.7306239,1.1983683,1.6642996,2.132044,2.5997884,2.5381477,2.474694,2.4130533,2.3495996,2.2879589,1.8691645,1.452183,1.0352017,0.61822027,0.19942589,0.17223145,0.14503701,0.11784257,0.09064813,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.15047589,0.2374981,0.3245203,0.41335547,0.50037766,0.8557183,1.209246,1.5645868,1.9199274,2.275268,2.8517902,3.4301252,4.006647,4.5849824,5.163317,4.936697,4.7118897,4.4870825,4.262275,4.0374675,4.360175,4.6828823,5.0055895,5.328297,5.6491914,5.475147,5.2992897,5.125245,4.949388,4.7753434,5.5984282,6.4197006,7.2427855,8.06587,8.887142,7.2790446,5.67276,4.064662,2.4583774,0.85027945,1.3270886,1.8057107,2.2825198,2.759329,3.2379513,3.1074178,2.9768846,2.8481643,2.7176309,2.5870976,5.8921285,9.197159,12.50219,15.80722,19.112251,21.322252,23.532255,25.742256,27.952257,30.162258,25.827465,21.492672,17.157877,12.823084,8.488291,7.0016613,5.516845,4.0320287,2.5472124,1.062396,1.015259,0.968122,0.91917205,0.872035,0.824898,1.015259,1.2056202,1.3941683,1.5845293,1.7748904,3.874301,5.975525,8.074935,10.174346,12.27557,9.857078,7.440398,5.0219064,2.6052272,0.18673515,0.18492219,0.18310922,0.1794833,0.17767033,0.17585737,0.19761293,0.21936847,0.24293698,0.26469254,0.28826106,0.24474995,0.2030518,0.15954071,0.11784257,0.07433146,0.06707962,0.059827764,0.052575916,0.045324065,0.038072214,0.19217403,0.3480888,0.50219065,0.65810543,0.8122072,0.75963134,0.7070554,0.6544795,0.60190356,0.5493277,0.44780177,0.3444629,0.24293698,0.13959812,0.038072214,0.5293851,1.0225109,1.5156367,2.0069497,2.5000753,4.0447197,5.5893636,7.135821,8.680465,10.225109,11.7969475,13.370599,14.942437,16.514277,18.087927,18.552046,19.017977,19.482096,19.948027,20.412146,18.111496,15.812659,13.512011,11.213174,8.912524,7.7195945,6.526665,5.335549,4.1426196,2.94969,2.759329,2.570781,2.38042,2.1900587,1.9996977,2.953316,3.9051213,4.856927,5.810545,6.7623506,9.782746,12.803142,15.821725,18.84212,21.862516,21.46729,21.072063,20.676838,20.283426,19.888199,20.667774,21.447348,22.226921,23.008308,23.787882,25.747694,27.707508,29.66732,31.627132,33.586945,31.297173,29.0074,26.71763,24.427858,22.138086,21.304123,20.471973,19.639824,18.807674,17.975525,18.096992,18.220274,18.341742,18.465023,18.588305,17.857681,17.127058,16.398247,15.667623,14.936998,14.911617,14.888049,14.862667,14.837286,14.811904,14.112101,13.412297,12.712494,12.012691,11.312886,16.338419,21.36395,26.38767,31.41139,36.43692,35.24218,34.047436,32.852695,31.657953,30.463211,30.321798,30.182201,30.042603,29.903006,29.761593,25.715061,21.666716,17.620184,13.573651,9.525306,10.97205,12.420607,13.867351,15.314095,16.762651,15.245202,13.727753,12.210303,10.692853,9.175404,7.607191,6.0389786,4.4725785,2.904366,1.3379664,1.5809034,1.8220274,2.0649643,2.3079014,2.5508385,2.9369993,3.049403,3.1618068,3.2742105,3.386614,3.5008307,3.2633326,3.0258346,2.7883365,2.5508385,2.3133402,4.7245803,7.137634,9.550687,11.961927,14.37498,16.913128,19.449463,21.98761,24.525759,27.062092,25.749508,24.436922,23.124338,21.811752,20.499168,21.162712,21.824444,22.487988,23.14972,23.813263,19.375132,14.936998,10.500679,6.0625467,1.6244144,1.7368182,1.8492218,1.9616255,2.0758421,2.1882458,2.7502642,3.3122826,3.874301,4.4381323,5.0001507,6.550234,8.100317,9.6504,11.200482,12.750566,13.412297,14.075842,14.737573,15.399304,16.062849,16.962078,17.863121,18.76235,19.663393,20.562622,18.213022,15.863422,13.512011,11.162411,8.812811,8.899834,8.9868555,9.07569,9.162713,9.249735,8.488291,7.7250338,6.9617763,6.200332,5.4370747,4.800725,4.162562,3.5243993,2.8880494,2.2498865,2.5508385,2.8499773,3.149116,3.4500678,3.7492065,5.524097,7.3008003,9.07569,10.850581,12.625471,14.837286,17.0491,19.262728,21.474543,23.68817,25.136726,26.587097,28.037466,29.487837,30.938206,27.54978,24.163166,20.774738,17.388124,13.999697,12.32452,10.649343,8.974165,7.3008003,5.6256227,4.8877473,4.1498713,3.4119956,2.6741197,1.938057,2.2371957,2.5381477,2.8372865,3.1382382,3.437377,4.6629395,5.8866897,7.112252,8.337815,9.563377,9.237044,8.912524,8.588004,8.26167,7.93715,9.336758,10.738177,12.137785,13.537392,14.936998,12.899229,10.863272,8.825501,6.787732,4.749962,3.825351,2.9007401,1.9743162,1.0497054,0.12509441,2.0123885,3.8996825,5.7869763,7.6742706,9.563377,10.950294,12.337211,13.72594,15.112856,16.499773,16.200634,15.899682,15.600543,15.299591,15.000452,13.974316,12.949992,11.925668,10.899531,9.875207,8.999546,8.125698,7.250037,6.3743763,5.5005283,5.0255322,4.550536,4.07554,3.6005437,3.1255474,3.6241121,4.12449,4.6248674,5.125245,5.6256227,5.562169,5.5005283,5.4370747,5.375434,5.3119802,4.98746,4.6629395,4.3366065,4.0120864,3.6875658,4.1879435,4.688321,5.186886,5.6872635,6.187641,5.7380266,5.2884116,4.836984,4.3873696,3.9377546,4.175253,4.4127507,4.650249,4.8877473,5.125245,5.3500524,5.57486,5.7996674,6.0244746,6.249282,5.9501433,5.6491914,5.3500524,5.049101,4.749962,6.736969,8.725789,10.712796,12.699803,14.68681,16.313038,17.937452,19.561867,21.188093,22.812508,21.675781,20.537241,19.400513,18.261972,17.125244,18.649946,20.174648,21.699348,23.225864,24.750565,21.900587,19.050611,16.200634,13.3506565,10.500679,10.375585,10.25049,10.125396,10.000301,9.875207,8.537241,7.1992745,5.863121,4.5251546,3.1871881,3.5243993,3.8616104,4.2006345,4.537845,4.8750563,5.774286,6.6753283,7.574558,8.4756,9.374829,9.800876,10.225109,10.649343,11.075388,11.499621,10.850581,10.199727,9.550687,8.899834,8.2507925,7.93715,7.6253204,7.311678,6.9998484,6.688019,5.774286,4.8623657,3.9504454,3.0367124,2.124792,2.3006494,2.474694,2.6505513,2.8245957,3.000453,3.1382382,3.2742105,3.4119956,3.5497808,3.6875658,3.874301,4.062849,4.249584,4.4381323,4.6248674,4.137181,3.6494937,3.1618068,2.6741197,2.1882458,2.3006494,2.4130533,2.525457,2.6378605,2.7502642,2.2245052,1.7005589,1.1747998,0.6508536,0.12509441,0.17585737,0.22480737,0.2755703,0.3245203,0.37528324,1.0750868,1.7748904,2.474694,3.1744974,3.874301,4.024777,4.175253,4.325729,4.4743915,4.6248674,4.349297,4.07554,3.7999697,3.5243993,3.2506418,3.1744974,3.100166,3.0258346,2.94969,2.8753586,2.8499773,2.8245957,2.7992141,2.7756457,2.7502642,2.2879589,1.8256533,1.3633479,0.89922947,0.43692398,0.34990177,0.26287958,0.17585737,0.0870222,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13778515,0.2755703,0.41335547,0.5493277,0.6871128,0.824898,0.96268314,1.1004683,1.2382535,1.3742256,3.53709,5.6999545,7.8628187,10.025683,12.186734,9.750113,7.311678,4.8750563,2.4366217,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.11240368,0.16316663,0.21211663,0.26287958,0.31182957,0.69980353,1.0877775,1.4757515,1.8619126,2.2498865,2.0994108,1.9507477,1.8002719,1.649796,1.49932,1.2255627,0.9499924,0.6744221,0.40066472,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.34990177,0.63816285,0.9246109,1.2128719,1.49932,1.4249886,1.3506571,1.2745126,1.2001812,1.1258497,1.49932,1.8746033,2.2498865,2.6251698,3.000453,3.4246864,3.8507326,4.274966,4.699199,5.125245,4.936697,4.749962,4.5632267,4.3746786,4.1879435,5.2503395,6.3127356,7.3751316,8.437528,9.499924,7.763106,6.0244746,4.2876563,2.5508385,0.8122072,1.3506571,1.887294,2.4257438,2.962381,3.5008307,3.2742105,3.049403,2.8245957,2.5997884,2.374981,5.7996674,9.224354,12.650853,16.075539,19.500225,22.85058,26.199121,29.549477,32.899834,36.250187,30.52485,24.799515,19.074179,13.3506565,7.6253204,6.249282,4.8750563,3.5008307,2.124792,0.7505665,0.7505665,0.7505665,0.7505665,0.7505665,0.7505665,0.93730164,1.1258497,1.3125849,1.49932,1.6878681,4.0501585,6.412449,8.774739,11.137029,13.499319,10.837891,8.174648,5.5132194,2.8499773,0.18673515,0.18673515,0.18673515,0.18673515,0.18673515,0.18673515,0.21211663,0.2374981,0.26287958,0.28826106,0.31182957,0.25018883,0.18673515,0.12509441,0.06164073,0.0,0.0,0.0,0.0,0.0,0.0,0.17585737,0.34990177,0.52575916,0.69980353,0.87566096,0.73787576,0.6000906,0.46230546,0.3245203,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.62547207,1.2491312,1.8746033,2.5000753,3.1255474,5.0128417,6.9001355,8.78743,10.674724,12.562017,13.363347,14.162864,14.96238,15.761897,16.563227,17.112555,17.661882,18.213022,18.76235,19.311678,16.800724,14.287958,11.775192,9.262425,6.7496595,5.7869763,4.8242936,3.8616104,2.9007401,1.938057,1.7368182,1.5373923,1.3379664,1.1367276,0.93730164,1.8383441,2.7375734,3.636803,4.537845,5.4370747,8.700407,11.961927,15.22526,18.48678,21.750113,21.037619,20.325123,19.612629,18.900135,18.187641,18.862062,19.538298,20.212719,20.887142,21.563377,23.575766,25.588154,27.600542,29.61293,31.625319,30.136877,28.650248,27.161806,25.675177,24.186733,23.22405,22.26318,21.300497,20.337814,19.375132,19.337059,19.3008,19.262728,19.224655,19.188396,18.43783,17.687263,16.936697,16.187943,15.437376,15.337664,15.23795,15.138238,15.036712,14.936998,14.162864,13.386916,12.612781,11.836833,11.062697,16.300346,21.537996,26.775644,32.01148,37.24913,36.837585,36.424232,36.012688,35.599335,35.18779,35.037315,34.88684,34.738174,34.5877,34.437225,29.299288,24.161352,19.025229,13.887294,8.749357,10.56232,12.375282,14.188245,15.999394,17.812357,15.8869915,13.961625,12.038072,10.112705,8.187339,6.787732,5.388125,3.9867048,2.5870976,1.1874905,1.4866294,1.7875811,2.08672,2.3876717,2.6868105,2.9007401,2.9968271,3.094727,3.1926272,3.290527,3.386614,3.159994,2.9333735,2.70494,2.47832,2.2498865,4.6230545,6.9944096,9.367578,11.740746,14.112101,16.7554,19.396887,22.040186,24.681673,27.324972,25.704184,24.085207,22.464418,20.845444,19.224655,19.52742,19.830185,20.13295,20.435715,20.736666,17.23221,13.727753,10.223296,6.717026,3.2125697,3.0657198,2.9170568,2.770207,2.6233568,2.474694,3.2524548,4.0302157,4.8079767,5.5857377,6.3616858,7.614443,8.8672,10.119957,11.372714,12.625471,13.390542,14.155612,14.920682,15.685752,16.450823,17.025532,17.60024,18.17495,18.749659,19.324368,17.369995,15.415621,13.4594345,11.50506,9.550687,9.697536,9.844387,9.99305,10.139899,10.28675,9.644961,9.003172,8.3595705,7.7177815,7.07418,6.6644506,6.2547207,5.844991,5.4352617,5.0255322,5.4407005,5.8558693,6.2692246,6.684393,7.0995617,8.074935,9.050309,10.025683,10.999244,11.974618,14.222692,16.470764,18.717026,20.9651,23.213173,24.944551,26.677744,28.410936,30.142317,31.875507,29.589363,27.305029,25.020697,22.73455,20.450218,17.589363,14.730321,11.869466,9.010424,6.149569,5.3953767,4.6393714,3.8851788,3.1291735,2.374981,2.6233568,2.8699198,3.1182957,3.3648586,3.6132345,4.8152285,6.017223,7.219217,8.423024,9.625018,9.247922,8.870826,8.491917,8.1148205,7.7377243,9.175404,10.613083,12.050762,13.486629,14.924308,13.15667,11.390844,9.623205,7.855567,6.0879283,4.9276323,3.7673361,2.6070402,1.4467441,0.28826106,3.4283123,6.5665503,9.708415,12.848466,15.986704,15.925063,15.863422,15.799969,15.738328,15.674874,14.96238,14.249886,13.537392,12.824898,12.112403,11.552197,10.991992,10.431787,9.871581,9.313189,8.392203,7.473032,6.552047,5.632875,4.7118897,4.2930956,3.872488,3.4518807,3.0330863,2.612479,3.1654327,3.7183862,4.269527,4.8224807,5.375434,5.282973,5.1905117,5.0980506,5.0055895,4.9131284,4.650249,4.3873696,4.12449,3.8616104,3.6005437,4.0483456,4.494334,4.942136,5.389938,5.8377395,5.516845,5.197764,4.876869,4.557788,4.2368937,4.4508233,4.6629395,4.8750563,5.087173,5.2992897,5.620184,5.9392653,6.26016,6.5792413,6.9001355,6.5955577,6.2891674,5.9845896,5.6800117,5.375434,6.9744673,8.575313,10.174346,11.775192,13.374225,15.547967,17.719896,19.891825,22.065567,24.237497,23.43798,22.63665,21.837133,21.037619,20.238102,20.87445,21.512613,22.150776,22.787127,23.42529,20.629702,17.835926,15.040338,12.244749,9.449161,9.287807,9.12464,8.963287,8.80012,8.636953,7.4331465,6.2275267,5.0219064,3.8180993,2.612479,2.8699198,3.1273603,3.3848011,3.6422417,3.8996825,4.6973863,5.4950895,6.2927933,7.0904965,7.8882003,8.23085,8.571687,8.914337,9.256987,9.599637,9.325879,9.050309,8.774739,8.499168,8.225411,8.080374,7.935337,7.7903004,7.645263,7.500226,6.5030966,5.504154,4.507025,3.5098956,2.5127661,2.5744069,2.6378605,2.6995013,2.762955,2.8245957,3.1926272,3.5606585,3.926877,4.2949085,4.6629395,4.710077,4.7572136,4.804351,4.853301,4.900438,4.5469103,4.195195,3.8416677,3.489953,3.1382382,3.2651455,3.392053,3.5207734,3.6476808,3.774588,3.2651455,2.7557032,2.2444477,1.7350051,1.2255627,1.260009,1.2944553,1.3307146,1.3651608,1.3996071,1.9199274,2.4402475,2.960568,3.4808881,3.9993954,4.1970086,4.3946214,4.592234,4.7898474,4.98746,4.748149,4.507025,4.267714,4.028403,3.787279,3.7401419,3.6930048,3.6458678,3.5969179,3.5497808,3.343103,3.1346123,2.9279346,2.7194438,2.5127661,2.079468,1.647983,1.214685,0.78319985,0.34990177,0.27919623,0.21030366,0.13959812,0.07070554,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.15772775,0.3154555,0.47318324,0.630911,0.7868258,0.726998,0.6671702,0.6073425,0.5475147,0.48768693,0.38978696,0.291887,0.19579996,0.09789998,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.11059072,0.21936847,0.32995918,0.4405499,0.5493277,0.65991837,0.7705091,0.8792868,0.9898776,1.1004683,2.8409123,4.5795436,6.319988,8.0604315,9.800876,7.846502,5.8957543,3.9431937,1.9906329,0.038072214,0.11784257,0.19761293,0.27738327,0.35715362,0.43692398,0.41335547,0.387974,0.36259252,0.33721104,0.31182957,0.678048,1.0424535,1.4068589,1.7730774,2.137483,1.983381,1.8274662,1.6733645,1.5174497,1.3633479,1.114972,0.8684091,0.6200332,0.37165734,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.32270733,0.581961,0.8430276,1.1022812,1.3633479,1.2726997,1.1820517,1.0932164,1.0025684,0.9119202,1.2273756,1.5428312,1.8582866,2.1719291,2.4873846,2.8717327,3.2578938,3.6422417,4.028403,4.4127507,4.209699,4.006647,3.8054085,3.6023567,3.3993049,4.2804046,5.1596913,6.0407915,6.9200783,7.799365,6.688019,5.57486,4.461701,3.350355,2.2371957,2.810092,3.3829882,3.9558845,4.5269675,5.0998635,5.0074024,4.914942,4.8224807,4.7300196,4.6375585,7.703278,10.767185,13.832905,16.89681,19.96253,22.078259,24.192173,26.3079,28.421814,30.537542,25.885479,21.233418,16.579542,11.927481,7.2754188,6.1731377,5.0708566,3.966762,2.864481,1.7621996,1.5573349,1.35247,1.1476053,0.94274056,0.73787576,0.88472575,1.0333886,1.1802386,1.3270886,1.4757515,3.346729,5.219519,7.0923095,8.9651,10.837891,8.780178,6.722465,4.664753,2.6070402,0.5493277,0.5420758,0.53482395,0.5275721,0.52032024,0.51306844,0.46411842,0.4169814,0.36984438,0.32270733,0.2755703,0.21936847,0.16497959,0.11059072,0.054388877,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.15954071,0.30820364,0.4550536,0.60190356,0.7505665,0.629098,0.5094425,0.38978696,0.27013144,0.15047589,0.15047589,0.15047589,0.15047589,0.15047589,0.15047589,1.0424535,1.9344311,2.8282216,3.720199,4.612177,6.169512,7.7268467,9.284182,10.843329,12.400664,13.008006,13.615349,14.222692,14.830034,15.437376,15.589665,15.741954,15.894243,16.048346,16.200634,14.046834,11.894848,9.742861,7.590874,5.4370747,5.0799212,4.7227674,4.365614,4.006647,3.6494937,3.1128569,2.5744069,2.03777,1.49932,0.96268314,1.7168756,2.472881,3.2270734,3.9830787,4.7372713,7.4367723,10.138086,12.837588,15.537089,18.236591,17.85043,17.462456,17.074482,16.68832,16.300346,16.956638,17.614744,18.27285,18.929142,19.587248,21.19172,22.798004,24.402477,26.006948,27.613234,26.349598,25.087776,23.82414,22.562319,21.300497,20.675026,20.049553,19.424082,18.800423,18.17495,18.610062,19.045172,19.480284,19.915394,20.350506,19.387821,18.425138,17.462456,16.499773,15.537089,15.528025,15.517147,15.508082,15.497204,15.488139,14.487384,13.486629,12.487686,11.486931,10.487988,14.880796,19.273605,23.6646,28.05741,32.45022,32.930653,33.409275,33.88971,34.370144,34.85058,34.964798,35.080826,35.19504,35.309258,35.42529,30.392506,25.35972,20.326937,15.295965,10.263181,11.630155,12.9971285,14.365915,15.732889,17.099863,15.06028,13.018885,10.979301,8.939718,6.9001355,5.805106,4.710077,3.6150475,2.520018,1.4249886,1.6207886,1.8147756,2.0105755,2.2045624,2.4003625,2.8626678,2.9442513,3.0276475,3.1092308,3.1926272,3.2742105,3.056655,2.8409123,2.6233568,2.4058013,2.1882458,4.519716,6.8529987,9.184468,11.517752,13.849221,16.597672,19.34431,22.092762,24.839401,27.587852,25.660673,23.73168,21.8045,19.877321,17.950142,17.892128,17.834112,17.77791,17.719896,17.661882,15.089288,12.516694,9.944099,7.3733187,4.800725,4.3928084,3.9848917,3.576975,3.1708715,2.762955,3.7546456,4.748149,5.7398396,6.733343,7.7250338,8.680465,9.634083,10.589515,11.544946,12.500377,13.366973,14.235382,15.101978,15.970387,16.836983,17.087172,17.33736,17.58755,17.837738,18.087927,16.526966,14.967819,13.406858,11.847711,10.28675,10.49524,10.701918,10.910409,11.117086,11.325577,10.801631,10.279498,9.757364,9.235231,8.713099,8.529989,8.34688,8.165584,7.9824743,7.799365,8.330563,8.859948,9.389333,9.920531,10.449916,10.625773,10.799818,10.975676,11.14972,11.325577,13.608097,15.890617,18.173138,20.455656,22.738176,24.752378,26.766579,28.782595,30.796795,32.81281,31.630758,30.446894,29.264841,28.08279,26.90074,22.854206,18.809486,14.764768,10.720048,6.6753283,5.903006,5.130684,4.358362,3.584227,2.811905,3.007705,3.2016919,3.397492,3.5932918,3.787279,4.9675174,6.147756,7.327995,8.508233,9.686659,9.256987,8.827314,8.397643,7.9679704,7.5382986,9.012237,10.487988,11.961927,13.437678,14.911617,13.415923,11.918416,10.419096,8.921589,7.4258947,6.0299134,4.6357455,3.2397642,1.845596,0.44961473,4.842423,9.235231,13.628039,18.020847,22.411844,20.899832,19.387821,17.87581,16.361988,14.849977,13.724127,12.60009,11.47424,10.3502035,9.224354,9.130079,9.035806,8.939718,8.845445,8.749357,7.7848616,6.8203654,5.8558693,4.88956,3.925064,3.5606585,3.1944401,2.8300345,2.465629,2.0994108,2.70494,3.3104696,3.9141862,4.519716,5.125245,5.0019636,4.880495,4.7572136,4.6357455,4.512464,4.313038,4.1117992,3.9123733,3.7129474,3.5117085,3.9069343,4.3021603,4.6973863,5.092612,5.487838,5.297477,5.1071157,4.9167547,4.7282066,4.537845,4.7245803,4.9131284,5.0998635,5.2865987,5.475147,5.8903155,6.305484,6.720652,7.135821,7.549176,7.2391596,6.929143,6.6191263,6.3091097,6.000906,7.211965,8.424837,9.637709,10.850581,12.06164,14.782897,17.50234,20.221785,22.94304,25.662485,25.20018,24.737875,24.27557,23.813263,23.349146,23.100769,22.85058,22.600391,22.350203,22.100014,19.360628,16.619429,13.880041,11.1406555,8.399456,8.200029,8.000604,7.799365,7.5999393,7.400513,6.3272395,5.2557783,4.1825047,3.1092308,2.03777,2.2154403,2.3931105,2.570781,2.7466383,2.9243085,3.6204863,4.314851,5.009216,5.7053933,6.399758,6.6608243,6.9200783,7.179332,7.440398,7.699652,7.799365,7.900891,8.000604,8.100317,8.200029,8.221786,8.245354,8.267109,8.290678,8.312433,7.230095,6.147756,5.0654173,3.9830787,2.9007401,2.8499773,2.7992141,2.7502642,2.6995013,2.6505513,3.247016,3.8452935,4.441758,5.040036,5.638314,5.5458527,5.4533916,5.3591175,5.2666564,5.1741953,4.95664,4.740897,4.5233417,4.305786,4.0882306,4.229642,4.3728657,4.514277,4.6575007,4.800725,4.305786,3.8108473,3.3140955,2.819157,2.324218,2.3441606,2.3641033,2.3858588,2.4058013,2.4257438,2.764768,3.105605,3.444629,3.785466,4.12449,4.36924,4.615803,4.860553,5.105303,5.3500524,5.145188,4.940323,4.7354584,4.5305934,4.325729,4.305786,4.2858434,4.265901,4.2441454,4.2242026,3.834416,3.444629,3.054842,2.665055,2.275268,1.8727903,1.4703126,1.067835,0.6653573,0.26287958,0.21030366,0.15772775,0.10515183,0.052575916,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.3154555,0.629098,0.9445535,1.260009,1.5754645,1.405046,1.2346275,1.064209,0.89560354,0.72518504,0.58014804,0.43511102,0.29007402,0.14503701,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0,0.0,0.0,0.0,0.0,0.08339628,0.16497959,0.24837588,0.32995918,0.41335547,0.4949388,0.57833505,0.65991837,0.7433147,0.824898,2.1429217,3.4591327,4.7771564,6.09518,7.413204,5.9447045,4.478018,3.009518,1.5428312,0.07433146,0.2229944,0.36984438,0.5166943,0.6653573,0.8122072,0.7124943,0.61278135,0.51306844,0.41335547,0.31182957,0.6544795,0.99712944,1.3397794,1.6824293,2.0250793,1.8655385,1.7041848,1.5446441,1.3851035,1.2255627,1.0043813,0.7850128,0.5656443,0.3444629,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.2955129,0.5275721,0.75963134,0.9916905,1.2255627,1.1204109,1.015259,0.9101072,0.80495536,0.69980353,0.9554313,1.209246,1.4648738,1.7205015,1.9743162,2.3205922,2.665055,3.009518,3.3557937,3.7002566,3.482701,3.2651455,3.04759,2.8300345,2.612479,3.3104696,4.006647,4.704638,5.4026284,6.1006193,5.612932,5.125245,4.6375585,4.1498713,3.6621845,4.269527,4.876869,5.484212,6.093367,6.70071,6.740595,6.78048,6.8203654,6.8602505,6.9001355,9.605076,12.310016,15.014956,17.719896,20.424837,21.305937,22.185223,23.06451,23.94561,24.824896,21.244295,17.665508,14.084907,10.504305,6.925517,6.09518,5.2648435,4.4345064,3.6041696,2.7756457,2.3641033,1.9543737,1.5446441,1.1349145,0.72518504,0.8321498,0.93911463,1.0478923,1.1548572,1.261822,2.6451125,4.02659,5.40988,6.793171,8.174648,6.722465,5.2702823,3.8180993,2.3641033,0.9119202,0.8974165,0.88291276,0.8665961,0.8520924,0.8375887,0.7179332,0.5982776,0.47680917,0.35715362,0.2374981,0.19036107,0.14322405,0.09427405,0.047137026,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.14503701,0.26469254,0.38434806,0.5058166,0.62547207,0.52213323,0.42060733,0.31726846,0.21574254,0.11240368,0.15047589,0.18673515,0.22480737,0.26287958,0.2991388,1.4594349,2.619731,3.780027,4.940323,6.1006193,7.327995,8.55537,9.782746,11.010121,12.237497,12.652666,13.067834,13.483003,13.898171,14.313339,14.066776,13.822026,13.577277,13.332527,13.087777,11.294757,9.501737,7.71053,5.91751,4.12449,4.3728657,4.6194286,4.8678045,5.1143675,5.3627434,4.4870825,3.6132345,2.7375734,1.8619126,0.9880646,1.5972201,2.2081885,2.817344,3.4283123,4.0374675,6.1749506,8.312433,10.449916,12.5873995,14.724882,14.663241,14.599788,14.538147,14.474693,14.413053,15.053028,15.693004,16.33298,16.972956,17.612932,18.809486,20.007854,21.20441,22.402779,23.599335,22.562319,21.525305,20.48829,19.449463,18.412449,18.124187,17.837738,17.549479,17.26303,16.97477,17.883062,18.789545,19.697838,20.60432,21.512613,20.337814,19.163015,17.988214,16.813416,15.636803,15.718386,15.798156,15.877926,15.957697,16.037468,14.811904,13.588155,12.362592,11.137029,9.91328,13.4594345,17.007402,20.55537,24.101524,27.649492,29.021906,30.394318,31.766731,33.139145,34.51337,34.892277,35.273,35.65191,36.03263,36.413353,31.483908,26.556276,21.630457,16.702824,11.775192,12.697989,13.620788,14.541773,15.464571,16.38737,14.231756,12.077957,9.922344,7.7667317,5.612932,4.8224807,4.0320287,3.2415771,2.4529383,1.6624867,1.7531348,1.84197,1.9326181,2.0232663,2.1121013,2.8245957,2.8916752,2.960568,3.0276475,3.094727,3.1618068,2.955129,2.7466383,2.5399606,2.333283,2.124792,4.41819,6.7097745,9.003172,11.294757,13.588155,16.439945,19.291735,22.145338,24.997128,27.85073,25.615349,23.379965,21.144583,18.9092,16.67563,16.256836,15.839854,15.422873,15.004078,14.587097,12.948178,11.307447,9.666717,8.027799,6.3870673,5.719897,5.0527267,4.3855567,3.7183862,3.049403,4.256836,5.464269,6.6717024,7.8791356,9.088382,9.744674,10.40278,11.060884,11.717177,12.375282,13.345218,14.315152,15.285088,16.255022,17.224958,17.150625,17.074482,17.00015,16.92582,16.849674,15.685752,14.520018,13.354282,12.19036,11.024626,11.292944,11.559449,11.827768,12.094274,12.362592,11.9601145,11.557636,11.155159,10.752681,10.3502035,10.395528,10.440851,10.484363,10.529687,10.57501,11.220426,11.86584,12.509441,13.154857,13.800271,13.174799,12.549327,11.925668,11.300196,10.674724,12.99169,15.310469,17.627436,19.9444,22.26318,24.560204,26.857227,29.154251,31.453089,33.75011,33.67034,33.590572,33.5108,33.42922,33.349445,28.120863,22.890465,17.660069,12.429671,7.1992745,6.4106355,5.620184,4.8297324,4.0392804,3.2506418,3.392053,3.5352771,3.6766882,3.8199122,3.9631362,5.1198063,6.2782893,7.4349594,8.59163,9.750113,9.267865,8.785617,8.303369,7.819308,7.3370595,8.849071,10.362894,11.874905,13.386916,14.90074,13.673364,12.444175,11.2168,9.989424,8.762048,7.132195,5.5023413,3.872488,2.2426348,0.61278135,6.256534,11.9021,17.547665,23.19323,28.836983,25.874601,22.912222,19.94984,16.98746,14.025079,12.487686,10.950294,9.412902,7.8755093,6.338117,6.7079616,7.077806,7.4476504,7.817495,8.187339,7.177519,6.167699,5.1578784,4.1480584,3.1382382,2.8282216,2.518205,2.2081885,1.8981718,1.5881553,2.2444477,2.902553,3.5606585,4.216951,4.8750563,4.7227674,4.5704784,4.41819,4.264088,4.1117992,3.975827,3.8380418,3.7002566,3.5624714,3.4246864,3.7673361,4.1099863,4.4526362,4.795286,5.137936,5.0781083,5.0182805,4.95664,4.896812,4.836984,5.0001507,5.163317,5.3246713,5.487838,5.6491914,6.1604466,6.6698895,7.179332,7.690587,8.200029,7.8845744,7.569119,7.2554765,6.9400206,6.624565,7.4494634,8.274362,9.099259,9.924157,10.750868,14.017827,17.284784,20.551744,23.820515,27.087475,26.96238,26.837286,26.71219,26.587097,26.462002,25.325274,24.186733,23.050007,21.913279,20.774738,18.08974,15.404743,12.719746,10.034748,7.3497505,7.112252,6.874754,6.637256,6.399758,6.16226,5.223145,4.2822175,3.343103,2.4021754,1.4630609,1.5591478,1.6570477,1.7549478,1.8528478,1.9507477,2.5417736,3.1346123,3.727451,4.3202896,4.9131284,5.090799,5.2666564,5.4443264,5.621997,5.7996674,6.2746634,6.7496595,7.224656,7.699652,8.174648,8.365009,8.55537,8.745731,8.934279,9.12464,7.957093,6.789545,5.621997,4.454449,3.2869012,3.1255474,2.962381,2.7992141,2.6378605,2.474694,3.303218,4.1299286,4.95664,5.7851634,6.6118746,6.379815,6.147756,5.915697,5.6818247,5.4497657,5.368182,5.2847857,5.2032027,5.1198063,5.038223,5.1941376,5.351866,5.5095935,5.667321,5.825049,5.3446136,4.8641787,4.3855567,3.9051213,3.4246864,3.4301252,3.435564,3.43919,3.444629,3.4500678,3.6096084,3.7691493,3.930503,4.0900435,4.249584,4.5432844,4.835171,5.127058,5.4207582,5.712645,5.542227,5.371808,5.2032027,5.032784,4.8623657,4.8696175,4.876869,4.8841214,4.893186,4.900438,4.327542,3.7546456,3.1817493,2.610666,2.03777,1.6642996,1.2926424,0.91917205,0.5475147,0.17585737,0.13959812,0.10515183,0.07070554,0.034446288,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.47318324,0.9445535,1.4177368,1.8909199,2.3622901,2.0830941,1.8020848,1.5228885,1.2418793,0.96268314,0.7705091,0.57833505,0.38434806,0.19217403,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.0,0.0,0.0,0.0,0.0,0.054388877,0.11059072,0.16497959,0.21936847,0.2755703,0.32995918,0.38434806,0.4405499,0.4949388,0.5493277,1.4449311,2.3405347,3.2343252,4.1299286,5.0255322,4.0429068,3.0602808,2.077655,1.0950294,0.11240368,0.32814622,0.5420758,0.75781834,0.97174793,1.1874905,1.0116332,0.8375887,0.66173136,0.48768693,0.31182957,0.6327239,0.95180535,1.2726997,1.5917811,1.9126755,1.7476959,1.5827163,1.4177368,1.2527572,1.0877775,0.89560354,0.7016165,0.5094425,0.31726846,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.26831847,0.47318324,0.678048,0.88291276,1.0877775,0.968122,0.8466535,0.726998,0.6073425,0.48768693,0.68167394,0.8774739,1.0732739,1.2672608,1.4630609,1.7676386,2.0722163,2.3767939,2.6831846,2.9877625,2.7557032,2.521831,2.2897718,2.0577126,1.8256533,2.3405347,2.855416,3.3702974,3.8851788,4.40006,4.537845,4.6756306,4.8116026,4.949388,5.087173,5.730775,6.3725634,7.0143523,7.6579537,8.299743,8.471974,8.644206,8.81825,8.990481,9.162713,11.506873,13.852847,16.197008,18.542982,20.887142,20.531801,20.178274,19.822933,19.467592,19.112251,16.604925,14.097597,11.59027,9.082943,6.5756154,6.017223,5.4606433,4.902251,4.345671,3.787279,3.1726844,2.5580902,1.9416829,1.3270886,0.7124943,0.7795739,0.8466535,0.9155461,0.9826257,1.0497054,1.9416829,2.8354735,3.727451,4.6194286,5.5132194,4.664753,3.8180993,2.9696326,2.1229792,1.2745126,1.2527572,1.2291887,1.2074331,1.1856775,1.162109,0.969935,0.7777609,0.5855869,0.39159992,0.19942589,0.15954071,0.11965553,0.07977036,0.03988518,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.13053331,0.2229944,0.3154555,0.40791658,0.50037766,0.41516843,0.32995918,0.24474995,0.15954071,0.07433146,0.15047589,0.22480737,0.2991388,0.37528324,0.44961473,1.8782293,3.3050308,4.7318325,6.1604466,7.5872483,8.484665,9.382081,10.279498,11.176914,12.07433,12.297325,12.52032,12.743314,12.964496,13.1874895,12.545701,11.9021,11.26031,10.616709,9.97492,8.54268,7.1104393,5.678199,4.2459583,2.811905,3.6658103,4.517903,5.369995,6.2220874,7.07418,5.863121,4.650249,3.437377,2.2245052,1.0116332,1.4775645,1.9416829,2.4076142,2.8717327,3.3376641,4.9131284,6.48678,8.062244,9.637709,11.213174,11.47424,11.73712,11.999999,12.262879,12.525759,13.147605,13.769451,14.39311,15.014956,15.636803,16.427254,17.217705,18.008158,18.796797,19.587248,18.77504,17.962833,17.150625,16.338419,15.524399,15.575162,15.624111,15.674874,15.725637,15.774588,17.154251,18.53573,19.915394,21.29506,22.674723,21.287807,19.899076,18.512161,17.125244,15.738328,15.906934,16.077353,16.24777,16.41819,16.586794,15.138238,13.687867,12.237497,10.7871275,9.336758,12.039885,14.743011,17.444326,20.147453,22.85058,25.114971,27.37936,29.645565,31.909954,34.174343,34.81976,35.465176,36.110588,36.75419,37.399605,32.577126,27.754644,22.932163,18.109684,13.287203,13.765825,14.242634,14.719443,15.198066,15.674874,13.4050455,11.135216,8.865387,6.5955577,4.325729,3.8398547,3.3557937,2.8699198,2.3858588,1.8999848,1.8854811,1.8691645,1.8546607,1.840157,1.8256533,2.7883365,2.8390994,2.8916752,2.9442513,2.9968271,3.049403,2.8517902,2.6541772,2.4583774,2.2607644,2.0631514,4.314851,6.5665503,8.820063,11.071762,13.325275,16.282217,19.239159,22.197914,25.154856,28.111797,25.570024,23.028252,20.484665,17.94289,15.399304,14.623356,13.845595,13.067834,12.290073,11.512312,10.805257,10.098202,9.389333,8.682278,7.9752226,7.0469856,6.1205616,5.1923246,4.264088,3.3376641,4.76084,6.1822023,7.605378,9.026741,10.449916,10.810696,11.169662,11.530442,11.889409,12.250188,13.321649,14.394923,15.468197,16.539658,17.612932,17.212267,16.813416,16.41275,16.012085,15.613234,14.842725,14.072216,13.301706,12.5330105,11.762501,12.090648,12.416981,12.745127,13.073273,13.399607,13.116784,12.835775,12.552953,12.270131,11.9873085,12.259253,12.5330105,12.804955,13.0769,13.3506565,14.110288,14.869919,15.62955,16.389181,17.150625,15.725637,14.300649,12.87566,11.450671,10.025683,12.377095,14.730321,17.081734,19.43496,21.788185,24.36803,26.947876,29.527721,32.107567,34.687412,35.709923,36.732433,37.754948,38.77746,39.79997,33.385708,26.969631,20.55537,14.139296,7.7250338,6.9182653,6.109684,5.3029156,4.494334,3.6875658,3.778214,3.8670492,3.9576974,4.0483456,4.137181,5.272095,6.4070096,7.5419245,8.676839,9.811753,9.27693,8.7421055,8.207282,7.6724577,7.137634,8.6877165,10.2378,11.787883,13.337966,14.888049,13.930804,12.971747,12.0145035,11.057259,10.100015,8.234476,6.3707504,4.505212,2.6396735,0.774135,7.6724577,14.568967,21.46729,28.365612,35.262123,30.849371,26.438433,22.025682,17.612932,13.200181,11.249433,9.300498,7.3497505,5.4008155,3.4500678,4.2858434,5.1198063,5.955582,6.789545,7.6253204,6.5701766,5.5150323,4.459888,3.4047437,2.3495996,2.0957847,1.840157,1.5845293,1.3307146,1.0750868,1.7857682,2.4946365,3.2053177,3.9141862,4.6248674,4.441758,4.2604623,4.077353,3.8942437,3.7129474,3.636803,3.5624714,3.48814,3.4119956,3.3376641,3.6277382,3.917812,4.207886,4.49796,4.788034,4.856927,4.9276323,4.9983377,5.06723,5.137936,5.275721,5.411693,5.5494785,5.6872635,5.825049,6.430578,7.0342946,7.6398244,8.245354,8.8508835,8.529989,8.210908,7.890013,7.569119,7.250037,7.686961,8.125698,8.562622,8.999546,9.438283,13.252756,17.06723,20.883516,24.697989,28.512463,28.724579,28.936695,29.150625,29.362741,29.574858,27.54978,25.5247,23.49962,21.474543,19.449463,16.820667,14.190058,11.559449,8.930654,6.300045,6.0244746,5.750717,5.475147,5.199577,4.9258194,4.117238,3.3104696,2.5018883,1.69512,0.8883517,0.90466833,0.922798,0.93911463,0.9572442,0.97537386,1.4648738,1.9543737,2.4456866,2.9351864,3.4246864,3.5207734,3.6150475,3.7093215,3.8054085,3.8996825,4.749962,5.600241,6.450521,7.3008003,8.149267,8.508233,8.865387,9.222541,9.579695,9.936848,8.685904,7.4331465,6.1803894,4.9276323,3.6748753,3.3993049,3.1255474,2.8499773,2.5744069,2.3006494,3.3576066,4.4145637,5.473334,6.530291,7.5872483,7.215591,6.8421206,6.4704633,6.096993,5.7253356,5.7779117,5.8304877,5.883064,5.9356394,5.9882154,6.1604466,6.3326783,6.5049095,6.677141,6.849373,6.3852544,5.919323,5.4552045,4.989273,4.5251546,4.514277,4.505212,4.494334,4.4852695,4.4743915,4.454449,4.4345064,4.4145637,4.3946214,4.3746786,4.7155156,5.0545397,5.3953767,5.7344007,6.0752378,5.9392653,5.805106,5.669134,5.5349746,5.4008155,5.4352617,5.469708,5.504154,5.540414,5.57486,4.8206677,4.064662,3.3104696,2.5544643,1.8002719,1.4576219,1.114972,0.77232206,0.42967212,0.0870222,0.07070554,0.052575916,0.034446288,0.018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.630911,1.260009,1.8909199,2.520018,3.149116,2.759329,2.3695421,1.9797552,1.5899682,1.2001812,0.96087015,0.7197462,0.48043507,0.23931105,0.0,0.03988518,0.07977036,0.11965553,0.15954071,0.19942589,0.15954071,0.11965553,0.07977036,0.03988518,0.0,0.0,0.0,0.0,0.0,0.0,0.027194439,0.054388877,0.08339628,0.11059072,0.13778515,0.16497959,0.19217403,0.21936847,0.24837588,0.2755703,0.7469406,1.2201238,1.693307,2.1646774,2.6378605,2.1392958,1.6425442,1.1457924,0.64722764,0.15047589,0.43329805,0.71430725,0.99712944,1.2799516,1.5627737,1.3125849,1.062396,0.8122072,0.5620184,0.31182957,0.6091554,0.90829426,1.2056202,1.502946,1.8002719,1.6298534,1.4594349,1.2908293,1.1204109,0.9499924,0.7850128,0.6200332,0.4550536,0.29007402,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.23931105,0.4169814,0.5946517,0.77232206,0.9499924,0.81583315,0.67986095,0.54570174,0.40972954,0.2755703,0.40972954,0.54570174,0.67986095,0.81583315,0.9499924,1.214685,1.4793775,1.745883,2.0105755,2.275268,2.0268922,1.7803292,1.5319533,1.2853905,1.0370146,1.3705997,1.7023718,2.034144,2.3677292,2.6995013,3.4627585,4.2242026,4.98746,5.750717,6.5121617,7.1902094,7.8682575,8.544493,9.222541,9.900589,10.205167,10.509744,10.8143215,11.120712,11.42529,13.410484,15.3956785,17.380873,19.364254,21.349447,19.75948,18.169512,16.579542,14.989574,13.399607,11.965553,10.529687,9.0956335,7.6597667,6.2257137,5.9392653,5.65463,5.369995,5.08536,4.800725,3.9794528,3.159994,2.3405347,1.5192627,0.69980353,0.726998,0.7541924,0.78319985,0.8103943,0.8375887,1.2400664,1.6425442,2.0450218,2.4474995,2.8499773,2.6070402,2.3659163,2.1229792,1.8800422,1.6371052,1.6080978,1.5772774,1.54827,1.5174497,1.4866294,1.2219368,0.9572442,0.69255173,0.42785916,0.16316663,0.13053331,0.09789998,0.065266654,0.032633327,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.11421664,0.1794833,0.24474995,0.3100166,0.37528324,0.30820364,0.23931105,0.17223145,0.10515183,0.038072214,0.15047589,0.26287958,0.37528324,0.48768693,0.6000906,2.2952106,3.9903307,5.6854506,7.380571,9.07569,9.643148,10.210606,10.778063,11.34552,11.912977,11.941984,11.972805,12.001812,12.032633,12.06164,11.022813,9.982172,8.943344,7.902704,6.8620634,5.7906027,4.7173285,3.6458678,2.572594,1.49932,2.956942,4.4145637,5.8721857,7.3298078,8.78743,7.2373466,5.6872635,4.137181,2.5870976,1.0370146,1.357909,1.6769904,1.9978848,2.3169663,2.6378605,3.6494937,4.6629395,5.674573,6.688019,7.699652,8.287052,8.874452,9.461852,10.049252,10.636651,11.242181,11.847711,12.45324,13.056956,13.662486,14.045021,14.427556,14.810091,15.192626,15.575162,14.9877615,14.400362,13.812962,13.225562,12.638163,13.024323,13.412297,13.800271,14.188245,14.574407,16.427254,18.280102,20.13295,21.983984,23.836832,22.237799,20.636953,19.03792,17.437075,15.838041,16.097294,16.358362,16.617615,16.87687,17.137936,15.462758,13.7875805,12.112403,10.437225,8.762048,10.620335,12.4786215,14.335095,16.191568,18.049856,21.208036,24.366217,27.522585,30.678953,33.837135,34.747242,35.65735,36.567455,37.477562,38.38767,33.67034,28.951199,24.235683,19.518354,14.799213,14.831847,14.86448,14.897114,14.929747,14.96238,12.576522,10.192475,7.806617,5.422571,3.0367124,2.857229,2.6777458,2.4982624,2.3169663,2.137483,2.0178273,1.8981718,1.7767034,1.6570477,1.5373923,2.7502642,2.7883365,2.8245957,2.8626678,2.9007401,2.9369993,2.7502642,2.561716,2.374981,2.1882458,1.9996977,4.213325,6.4251394,8.636953,10.850581,13.062395,16.124489,19.186583,22.25049,25.312584,28.374678,25.5247,22.674723,19.824745,16.97477,14.124791,12.988064,11.849524,10.712796,9.574255,8.437528,8.662335,8.887142,9.11195,9.336758,9.563377,8.375887,7.1883965,5.999093,4.8116026,3.6241121,5.2630305,6.9001355,8.537241,10.174346,11.813264,11.874905,11.938358,11.999999,12.06164,12.125093,13.299893,14.474693,15.649493,16.824293,18.000906,17.27572,16.550535,15.825351,15.100165,14.37498,13.999697,13.6244135,13.24913,12.87566,12.500377,12.888351,13.274512,13.662486,14.05046,14.436621,14.275268,14.112101,13.9507475,13.7875805,13.6244135,14.124791,14.625169,15.125546,15.624111,16.124489,17.00015,17.87581,18.749659,19.62532,20.499168,18.274662,16.050158,13.825653,11.599335,9.374829,11.762501,14.150173,16.537846,18.925516,21.313189,24.175856,27.03671,29.89938,32.762047,35.624714,37.749508,39.8743,42.000904,44.125698,46.25049,38.65055,31.05061,23.45067,15.850732,8.2507925,7.4258947,6.599184,5.774286,4.949388,4.12449,4.162562,4.2006345,4.2368937,4.274966,4.313038,5.424384,6.5375433,7.650702,8.762048,9.875207,9.287807,8.700407,8.113008,7.5256076,6.9382076,8.52455,10.112705,11.700861,13.287203,14.875358,14.188245,13.499319,12.812206,12.125093,11.437981,9.336758,7.2373466,5.137936,3.0367124,0.93730164,9.086569,17.237648,25.386915,33.537994,41.687263,35.825954,29.962833,24.099712,18.236591,12.375282,10.012992,7.650702,5.2865987,2.9243085,0.5620184,1.8619126,3.1618068,4.461701,5.763408,7.063302,5.962834,4.8623657,3.7618973,2.663242,1.5627737,1.3633479,1.162109,0.96268314,0.76325727,0.5620184,1.3252757,2.08672,2.8499773,3.6132345,4.3746786,4.162562,3.9504454,3.738329,3.5243993,3.3122826,3.299592,3.2869012,3.2742105,3.2633326,3.2506418,3.48814,3.7256382,3.9631362,4.2006345,4.4381323,4.6375585,4.836984,5.038223,5.237649,5.4370747,5.5494785,5.661882,5.774286,5.8866897,6.000906,6.70071,7.400513,8.100317,8.80012,9.499924,9.175404,8.8508835,8.52455,8.200029,7.8755093,7.9244595,7.9752226,8.024173,8.074935,8.125698,12.487686,16.849674,21.213474,25.575462,29.93745,30.486778,31.03792,31.587248,32.13839,32.687714,29.774284,26.862667,23.949236,21.037619,18.124187,15.54978,12.975373,10.399154,7.8247466,5.2503395,4.936697,4.6248674,4.313038,3.9993954,3.6875658,3.0131438,2.3369088,1.6624867,0.9880646,0.31182957,0.25018883,0.18673515,0.12509441,0.06164073,0.0,0.387974,0.774135,1.162109,1.550083,1.938057,1.9507477,1.9616255,1.9743162,1.987007,1.9996977,3.2252605,4.4508233,5.674573,6.9001355,8.125698,8.649645,9.175404,9.699349,10.225109,10.750868,9.412902,8.074935,6.736969,5.4008155,4.062849,3.6748753,3.2869012,2.9007401,2.5127661,2.124792,3.4119956,4.699199,5.9882154,7.2754188,8.562622,8.049554,7.5382986,7.02523,6.5121617,6.000906,6.187641,6.3743763,6.5629244,6.7496595,6.9382076,7.124943,7.311678,7.500226,7.686961,7.8755093,7.4258947,6.9744673,6.5248523,6.0752378,5.6256227,5.600241,5.57486,5.5494785,5.524097,5.5005283,5.2992897,5.0998635,4.900438,4.699199,4.499773,4.8877473,5.275721,5.661882,6.049856,6.43783,6.338117,6.2384043,6.1368785,6.037165,5.9374523,6.000906,6.0625467,6.1241875,6.187641,6.249282,5.3119802,4.3746786,3.437377,2.5000753,1.5627737,1.2491312,0.93730164,0.62547207,0.31182957,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.7868258,1.5754645,2.3622901,3.149116,3.9377546,3.437377,2.9369993,2.4366217,1.938057,1.4376793,1.1494182,0.8629702,0.5747091,0.28826106,0.0,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,0.2374981,0.22480737,0.21211663,0.19942589,0.18673515,0.53663695,0.8883517,1.2382535,1.5881553,1.938057,1.6117238,1.2872034,0.96268314,0.63816285,0.31182957,0.5873999,0.8629702,1.1367276,1.4122978,1.6878681,1.5120108,1.3379664,1.162109,0.9880646,0.8122072,0.6744221,0.53663695,0.40066472,0.26287958,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.21211663,0.36259252,0.51306844,0.66173136,0.8122072,0.66173136,0.51306844,0.36259252,0.21211663,0.06164073,0.13778515,0.21211663,0.28826106,0.36259252,0.43692398,0.66173136,0.8883517,1.1131591,1.3379664,1.5627737,1.2998942,1.0370146,0.774135,0.51306844,0.25018883,0.40066472,0.5493277,0.69980353,0.85027945,1.0007553,2.3876717,3.774588,5.163317,6.550234,7.93715,8.649645,9.362139,10.074633,10.7871275,11.499621,11.938358,12.375282,12.812206,13.24913,13.687867,15.312282,16.936697,18.562923,20.187338,21.811752,18.987158,16.162561,13.337966,10.511557,7.686961,7.324369,6.9617763,6.599184,6.2365913,5.8758116,5.863121,5.8504305,5.8377395,5.825049,5.812358,4.788034,3.7618973,2.7375734,1.7132497,0.6871128,0.6744221,0.66173136,0.6508536,0.63816285,0.62547207,0.53663695,0.44961473,0.36259252,0.2755703,0.18673515,0.5493277,0.9119202,1.2745126,1.6371052,1.9996977,1.9616255,1.9253663,1.887294,1.8492218,1.8129625,1.4757515,1.1367276,0.7995165,0.46230546,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.099712946,0.13778515,0.17585737,0.21211663,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.15047589,0.2991388,0.44961473,0.6000906,0.7505665,2.712192,4.6756306,6.637256,8.600695,10.56232,10.799818,11.037316,11.274815,11.512312,11.74981,11.586644,11.42529,11.262123,11.10077,10.937603,9.499924,8.062244,6.624565,5.186886,3.7492065,3.0367124,2.324218,1.6117238,0.89922947,0.18673515,2.2498865,4.313038,6.3743763,8.437528,10.500679,8.611572,6.7242785,4.836984,2.94969,1.062396,1.2382535,1.4122978,1.5881553,1.7621996,1.938057,2.3876717,2.8372865,3.2869012,3.738329,4.1879435,5.0998635,6.011784,6.925517,7.837437,8.749357,9.336758,9.924157,10.51337,11.10077,11.6881695,11.662788,11.637406,11.612025,11.586644,11.563075,11.200482,10.837891,10.475298,10.112705,9.750113,10.475298,11.200482,11.925668,12.650853,13.374225,15.700256,18.024473,20.350506,22.674723,25.000753,23.187792,21.374828,19.561867,17.750717,15.937754,16.287657,16.637558,16.98746,17.33736,17.687263,15.787278,13.887294,11.9873085,10.087324,8.187339,9.200785,10.212419,11.225864,12.237497,13.24913,17.301102,21.351261,25.399607,29.449764,33.499924,34.67472,35.84952,37.024323,38.199123,39.375732,34.761745,30.149569,25.537392,20.925215,16.313038,15.899682,15.488139,15.074784,14.663241,14.249886,11.74981,9.249735,6.7496595,4.249584,1.7495089,1.8746033,1.9996977,2.124792,2.2498865,2.374981,2.1501737,1.9253663,1.7005589,1.4757515,1.2491312,2.712192,2.8046532,2.8971143,2.9895754,3.0820365,3.1744974,2.9732587,2.770207,2.5671551,2.3641033,2.1628644,4.4272547,6.6916447,8.957849,11.222239,13.486629,16.213324,18.938208,21.66309,24.387972,27.112856,24.598276,22.081884,19.567305,17.052727,14.538147,13.232814,11.927481,10.622148,9.316814,8.013294,8.145641,8.2779875,8.410334,8.54268,8.675026,7.549176,6.4251394,5.2992897,4.175253,3.049403,4.5342193,6.0208488,7.5056653,8.990481,10.475298,10.410031,10.344765,10.279498,10.2142315,10.150778,11.651911,13.154857,14.657803,16.160748,17.661882,16.940323,16.21695,15.495391,14.772019,14.05046,13.45037,12.850279,12.250188,11.650098,11.050007,11.49237,11.934732,12.377095,12.819458,13.261822,13.339779,13.417736,13.495693,13.571837,13.649796,13.979754,14.309713,14.639673,14.969632,15.299591,15.676687,16.055597,16.432693,16.80979,17.186886,15.484513,13.782142,12.07977,10.377398,8.675026,11.030065,13.385102,15.740141,18.095179,20.450218,22.620335,24.790451,26.960567,29.130682,31.300798,32.858135,34.41547,35.972805,37.53014,39.087475,32.72035,26.353224,19.984287,13.617162,7.250037,6.5701766,5.8903155,5.2104545,4.5305934,3.8507326,4.0030212,4.15531,4.307599,4.459888,4.612177,5.859495,7.1068134,8.355945,9.603263,10.850581,10.275872,9.699349,9.12464,8.549932,7.9752226,8.870826,9.764616,10.66022,11.555823,12.449615,12.5873995,12.725184,12.862969,13.000754,13.136727,11.535881,9.933222,8.330563,6.7279043,5.125245,11.512312,17.89938,24.28826,30.675327,37.062393,32.379513,27.698442,23.01556,18.332678,13.649796,11.432542,9.215289,6.9980354,4.780782,2.561716,3.442816,4.322103,5.2032027,6.0824895,6.9617763,5.9447045,4.9276323,3.9105604,2.8916752,1.8746033,1.6624867,1.4503701,1.2382535,1.0243238,0.8122072,1.4376793,2.0631514,2.6868105,3.3122826,3.9377546,3.8616104,3.787279,3.7129474,3.636803,3.5624714,3.5570326,3.5534067,3.5479677,3.5425289,3.53709,3.7492065,3.9631362,4.175253,4.3873696,4.599486,4.8496747,5.0998635,5.3500524,5.600241,5.8504305,6.011784,6.1749506,6.338117,6.4994707,6.6626377,7.364254,8.067683,8.7693,9.47273,10.174346,9.77912,9.385707,8.990481,8.595256,8.200029,8.7693,9.340384,9.909654,10.480737,11.050007,15.167245,19.284483,23.403534,27.520773,31.63801,31.817493,31.996977,32.178272,32.357758,32.53724,29.362741,26.188244,23.011934,19.837437,16.66294,14.665054,12.66717,10.669285,8.673213,6.6753283,6.19308,5.710832,5.2267714,4.744523,4.262275,3.491766,2.72307,1.9525607,1.1820517,0.41335547,0.34264994,0.27194437,0.2030518,0.13234627,0.06164073,0.36077955,0.65810543,0.9554313,1.2527572,1.550083,1.7096237,1.8691645,2.030518,2.1900587,2.3495996,3.5642843,4.780782,5.995467,7.210152,8.424837,8.667774,8.910711,9.151835,9.394773,9.637709,8.452031,7.268167,6.0824895,4.896812,3.7129474,3.4953918,3.2778363,3.0602808,2.8427253,2.6251698,3.6077955,4.590421,5.573047,6.5556726,7.5382986,7.1956487,6.8529987,6.510349,6.167699,5.825049,6.017223,6.209397,6.4033837,6.5955577,6.787732,6.9545245,7.12313,7.2899227,7.456715,7.6253204,7.2355337,6.8457465,6.454147,6.0643597,5.674573,5.620184,5.565795,5.5095935,5.4552045,5.4008155,5.375434,5.3500524,5.3246713,5.2992897,5.275721,5.4932766,5.710832,5.9283876,6.14413,6.3616858,6.2293396,6.096993,5.964647,5.8323007,5.6999545,5.8558693,6.009971,6.165886,6.319988,6.4759026,6.008158,5.540414,5.0726695,4.604925,4.137181,3.4500678,2.762955,2.0758421,1.3869164,0.69980353,0.56020546,0.42060733,0.27919623,0.13959812,0.0,0.07977036,0.15954071,0.23931105,0.3208944,0.40066472,0.3208944,0.23931105,0.15954071,0.07977036,0.0,0.7650702,1.5301404,2.2952106,3.0602808,3.825351,3.9631362,4.099108,4.2368937,4.3746786,4.512464,4.0900435,3.6676233,3.245203,2.8227828,2.4003625,2.2952106,2.1900587,2.084907,1.9797552,1.8746033,1.5101979,1.1457924,0.7795739,0.41516843,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.047137026,0.058014803,0.06707962,0.07795739,0.0870222,0.11421664,0.14322405,0.17041849,0.19761293,0.22480737,0.21755551,0.21030366,0.2030518,0.19579996,0.18673515,0.4604925,0.7324369,1.0043813,1.2781386,1.550083,1.3017071,1.0551442,0.80676836,0.56020546,0.31182957,0.5275721,0.7433147,0.9572442,1.1729867,1.3869164,1.2491312,1.1131591,0.97537386,0.8375887,0.69980353,0.5855869,0.46955732,0.35534066,0.23931105,0.12509441,0.11421664,0.10515183,0.09427405,0.08520924,0.07433146,0.07433146,0.07433146,0.07433146,0.07433146,0.07433146,0.072518505,0.07070554,0.06707962,0.065266654,0.06164073,0.28826106,0.51306844,0.73787576,0.96268314,1.1874905,0.96268314,0.73787576,0.51306844,0.28826106,0.06164073,0.14503701,0.22662032,0.3100166,0.39159992,0.4749962,0.65810543,0.83940166,1.0225109,1.2056202,1.3869164,1.1548572,0.922798,0.69073874,0.45686656,0.22480737,0.3444629,0.46411842,0.5855869,0.70524246,0.824898,2.182807,3.540716,4.896812,6.2547207,7.61263,8.105756,8.597069,9.090195,9.583321,10.074633,10.390089,10.705544,11.019187,11.334642,11.650098,12.975373,14.300649,15.625924,16.949387,18.274662,15.992143,13.709623,11.427103,9.144584,6.8620634,6.5230393,6.1822023,5.8431783,5.5023413,5.163317,5.317419,5.473334,5.6274357,5.7833505,5.9374523,4.9693303,4.0030212,3.0348995,2.0667772,1.1004683,1.0007553,0.89922947,0.7995165,0.69980353,0.6000906,0.52575916,0.44961473,0.37528324,0.2991388,0.22480737,0.73424983,1.2455053,1.7549478,2.2643902,2.7756457,2.5272698,2.280707,2.032331,1.7857682,1.5373923,1.2491312,0.96268314,0.6744221,0.387974,0.099712946,0.10333887,0.10515183,0.10696479,0.11059072,0.11240368,0.12690738,0.14322405,0.15772775,0.17223145,0.18673515,0.19036107,0.19217403,0.19579996,0.19761293,0.19942589,0.15954071,0.11965553,0.07977036,0.03988518,0.0,0.20486477,0.40972954,0.61459434,0.8194591,1.0243238,2.8481643,4.670192,6.492219,8.314246,10.138086,10.31757,10.497053,10.6783495,10.857833,11.037316,10.779876,10.522435,10.264994,10.007553,9.750113,8.582565,7.415017,6.247469,5.0799212,3.9123733,3.3793623,2.8481643,2.3151531,1.7821422,1.2491312,2.9732587,4.695573,6.4178877,8.140202,9.862516,8.412147,6.9617763,5.5132194,4.062849,2.612479,2.6976883,2.7828975,2.8681068,2.953316,3.0367124,3.2796493,3.5225863,3.7655232,4.006647,4.249584,5.1723824,6.09518,7.017978,7.9407763,8.861761,9.342196,9.822631,10.303066,10.781689,11.262123,10.937603,10.613083,10.28675,9.96223,9.637709,9.385707,9.131892,8.87989,8.627889,8.375887,9.0956335,9.815379,10.535126,11.254871,11.974618,14.333282,16.690134,19.046986,21.40565,23.7625,22.283123,20.801933,19.322556,17.843178,16.361988,16.702824,17.04185,17.382685,17.721708,18.062546,16.499773,14.936998,13.374225,11.813264,10.25049,10.827013,11.405348,11.98187,12.5602045,13.136727,16.447197,19.757666,23.068136,26.376793,29.687262,31.143072,32.59707,34.052876,35.50687,36.96268,32.615196,28.267712,23.920229,19.572744,15.22526,14.904366,14.585284,14.26439,13.945308,13.6244135,11.392657,9.159087,6.92733,4.695573,2.4620032,2.3876717,2.3133402,2.2371957,2.1628644,2.08672,2.030518,1.9725033,1.9144884,1.8582866,1.8002719,2.6741197,2.8227828,2.9696326,3.1182957,3.2651455,3.4119956,3.1944401,2.9768846,2.759329,2.5417736,2.324218,4.6429973,6.9599633,9.27693,11.595709,13.912675,16.300346,18.688019,21.07569,23.463362,25.84922,23.67004,21.490858,19.309864,17.130684,14.94969,13.477564,12.005438,10.533313,9.059374,7.5872483,7.6271334,7.667019,7.706904,7.746789,7.7866745,6.7242785,5.661882,4.599486,3.53709,2.474694,3.8072214,5.139749,6.472276,7.804804,9.137331,8.945157,8.752983,8.560809,8.366822,8.174648,10.00574,11.83502,13.664299,15.495391,17.32467,16.604925,15.885179,15.165432,14.445685,13.724127,12.899229,12.07433,11.249433,10.424535,9.599637,10.098202,10.594954,11.091705,11.59027,12.087022,12.40429,12.7233715,13.04064,13.357908,13.675177,13.834718,13.994258,14.155612,14.315152,14.474693,14.355038,14.235382,14.115726,13.994258,13.874602,12.694364,11.514126,10.3357,9.155461,7.9752226,10.297627,12.620032,14.942437,17.264843,19.587248,21.064812,22.542377,24.019941,25.497505,26.97507,27.964949,28.954826,29.944702,30.93458,31.924458,26.790148,21.655838,16.519714,11.385405,6.249282,5.714458,5.179634,4.64481,4.1099863,3.5751622,3.8416677,4.1099863,4.3783045,4.64481,4.9131284,6.294606,7.6778965,9.059374,10.442664,11.8241415,11.262123,10.700105,10.138086,9.574255,9.012237,9.215289,9.418341,9.619579,9.822631,10.025683,10.988366,11.949236,12.91192,13.874602,14.837286,13.7331915,12.627284,11.5231905,10.417283,9.313189,13.938056,18.562923,23.187792,27.812658,32.437527,28.934883,25.43224,21.929596,18.426952,14.924308,12.852092,10.779876,8.70766,6.635443,4.5632267,5.0219064,5.482399,5.942891,6.4033837,6.8620634,5.9283876,4.992899,4.0574102,3.1219215,2.1882458,1.9616255,1.7368182,1.5120108,1.2872034,1.062396,1.550083,2.03777,2.525457,3.0131438,3.5008307,3.5624714,3.6241121,3.6875658,3.7492065,3.8126602,3.8144734,3.8180993,3.8199122,3.8217251,3.825351,4.0120864,4.2006345,4.3873696,4.574105,4.762653,5.0617914,5.3627434,5.661882,5.962834,6.261973,6.4759026,6.688019,6.9001355,7.112252,7.324369,8.029612,8.734854,9.440096,10.145339,10.850581,10.384649,9.920531,9.4546,8.990481,8.52455,9.6141405,10.705544,11.795135,12.884725,13.974316,17.846804,21.719292,25.59178,29.464268,33.336758,33.14821,32.957848,32.767487,32.577126,32.386765,28.949387,25.512009,22.074633,18.637255,15.199879,13.780329,12.360779,10.939416,9.519867,8.100317,7.4476504,6.794984,6.1423173,5.4896507,4.836984,3.972201,3.1074178,2.2426348,1.3778516,0.51306844,0.43511102,0.35715362,0.27919623,0.2030518,0.12509441,0.33177215,0.5402629,0.7469406,0.9554313,1.162109,1.4703126,1.7767034,2.084907,2.3931105,2.6995013,3.9051213,5.1107416,6.3145485,7.520169,8.725789,8.685904,8.644206,8.604321,8.564435,8.52455,7.4929743,6.4595857,5.42801,4.3946214,3.3630457,3.3140955,3.2669585,3.2198215,3.1726844,3.1255474,3.8017826,4.4798307,5.1578784,5.8341136,6.5121617,6.33993,6.167699,5.995467,5.823236,5.6491914,5.846804,6.0444174,6.24203,6.439643,6.637256,6.784106,6.932769,7.079619,7.228282,7.3751316,7.0451727,6.7152133,6.3852544,6.055295,5.7253356,5.6401267,5.5549173,5.469708,5.384499,5.2992897,5.4497657,5.600241,5.750717,5.89938,6.049856,6.096993,6.14413,6.19308,6.240217,6.2873545,6.1223745,5.957395,5.7924156,5.6274357,5.462456,5.710832,5.957395,6.205771,6.452334,6.70071,6.7025228,6.7043357,6.7079616,6.7097745,6.7134004,5.6491914,4.5867953,3.5243993,2.4620032,1.3996071,1.1204109,0.83940166,0.56020546,0.27919623,0.0,0.15954071,0.3208944,0.48043507,0.6399758,0.7995165,0.6399758,0.48043507,0.3208944,0.15954071,0.0,0.7433147,1.4848163,2.228131,2.9696326,3.7129474,4.4870825,5.2630305,6.037165,6.813113,7.5872483,7.0306687,6.472276,5.915697,5.3573046,4.800725,4.539658,4.2804046,4.019338,3.7600844,3.5008307,2.819157,2.1392958,1.4594349,0.7795739,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.09427405,0.11421664,0.13415924,0.15410182,0.17585737,0.1794833,0.18492219,0.19036107,0.19579996,0.19942589,0.19761293,0.19579996,0.19217403,0.19036107,0.18673515,0.3825351,0.57833505,0.77232206,0.968122,1.162109,0.9916905,0.823085,0.6526665,0.48224804,0.31182957,0.46774435,0.62184614,0.7777609,0.9318628,1.0877775,0.9880646,0.8883517,0.7868258,0.6871128,0.5873999,0.4949388,0.40247768,0.3100166,0.21755551,0.12509441,0.11784257,0.11059072,0.10333887,0.09427405,0.0870222,0.0870222,0.0870222,0.0870222,0.0870222,0.0870222,0.08339628,0.07795739,0.072518505,0.06707962,0.06164073,0.36259252,0.66173136,0.96268314,1.261822,1.5627737,1.261822,0.96268314,0.66173136,0.36259252,0.06164073,0.15228885,0.24293698,0.33177215,0.4224203,0.51306844,0.6526665,0.79226464,0.9318628,1.0732739,1.2128719,1.0098201,0.80676836,0.6055295,0.40247768,0.19942589,0.29007402,0.38072214,0.46955732,0.56020546,0.6508536,1.9779422,3.3050308,4.632119,5.959208,7.28811,7.560054,7.8319983,8.105756,8.3777,8.649645,8.841819,9.035806,9.22798,9.420154,9.612328,10.636651,11.662788,12.687112,13.713249,14.737573,12.9971285,11.256684,9.518054,7.7776093,6.037165,5.719897,5.4026284,5.08536,4.7680917,4.4508233,4.7717175,5.0944247,5.4171324,5.7398396,6.0625467,5.1524396,4.2423325,3.3322253,2.422118,1.5120108,1.3252757,1.1367276,0.9499924,0.76325727,0.5747091,0.51306844,0.44961473,0.387974,0.3245203,0.26287958,0.91917205,1.5772774,2.2353828,2.8916752,3.5497808,3.092914,2.6342347,2.1773682,1.7205015,1.261822,1.0243238,0.7868258,0.5493277,0.31182957,0.07433146,0.10515183,0.13415924,0.16497959,0.19579996,0.22480737,0.24293698,0.25925365,0.27738327,0.2955129,0.31182957,0.27919623,0.24837588,0.21574254,0.18310922,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.25925365,0.52032024,0.7795739,1.0406405,1.2998942,2.9823234,4.664753,6.347182,8.029612,9.712041,9.835322,9.956791,10.080072,10.203354,10.324821,9.973107,9.619579,9.267865,8.914337,8.562622,7.665206,6.7677894,5.870373,4.972956,4.07554,3.7220123,3.3702974,3.0167696,2.665055,2.3133402,3.6948178,5.0781083,6.4595857,7.842876,9.224354,8.212721,7.1992745,6.187641,5.1741953,4.162562,4.157123,4.1516843,4.1480584,4.1426196,4.137181,4.171627,4.207886,4.2423325,4.2767787,4.313038,5.2449007,6.1767635,7.1104393,8.042302,8.974165,9.347635,9.719293,10.092763,10.46442,10.837891,10.212419,9.5869465,8.963287,8.337815,7.7123427,7.569119,7.4277077,7.2844834,7.1430726,6.9998484,7.7141557,8.430276,9.144584,9.860703,10.57501,12.964496,15.355793,17.745277,20.134762,22.524246,21.376642,20.229036,19.083244,17.935638,16.788034,17.117992,17.447952,17.77791,18.10787,18.43783,17.212267,15.986704,14.762955,13.537392,12.311829,12.455053,12.598277,12.739688,12.882912,13.024323,15.595104,18.165886,20.734854,23.305634,25.874601,27.609608,29.344612,31.079618,32.81462,34.54963,30.466837,26.384045,22.303066,18.220274,14.137483,13.910862,13.682428,13.455809,13.227375,13.000754,11.035503,9.070251,7.1050005,5.139749,3.1744974,2.9007401,2.6251698,2.3495996,2.0758421,1.8002719,1.9108626,2.0196402,2.1302311,2.2408218,2.3495996,2.6378605,2.8390994,3.0421512,3.245203,3.4482548,3.6494937,3.4174345,3.1853752,2.953316,2.7194438,2.4873846,4.856927,7.228282,9.597824,11.967366,14.336908,16.38737,18.43783,20.48829,22.536938,24.587399,22.741802,20.89802,19.052423,17.206827,15.363045,13.722314,12.083396,10.442664,8.801933,7.1630154,7.1104393,7.057863,7.0052876,6.9527116,6.9001355,5.89938,4.900438,3.8996825,2.9007401,1.8999848,3.0802233,4.2604623,5.4407005,6.6191263,7.799365,7.4802837,7.159389,6.8403077,6.5194135,6.200332,8.357758,10.515183,12.672608,14.830034,16.98746,16.269526,15.553406,14.835473,14.117539,13.399607,12.349901,11.300196,10.25049,9.200785,8.149267,8.70222,9.255174,9.808127,10.359268,10.912222,11.470614,12.027194,12.585587,13.142166,13.700559,13.68968,13.680615,13.669738,13.660673,13.649796,13.033388,12.415168,11.7969475,11.18054,10.56232,9.904215,9.247922,8.589817,7.931711,7.2754188,9.56519,11.854962,14.144734,16.434505,18.724277,19.50929,20.294304,21.079315,21.864328,22.649342,23.071762,23.494183,23.916603,24.340836,24.763256,20.859947,16.958452,13.055143,9.151835,5.2503395,4.860553,4.4707656,4.079166,3.6893787,3.299592,3.682127,4.064662,4.4471974,4.8297324,5.2122674,6.7297173,8.247167,9.764616,11.282066,12.799516,12.250188,11.700861,11.14972,10.600392,10.049252,9.5597515,9.070251,8.580752,8.089439,7.5999393,9.38752,11.175101,12.962683,14.750263,16.537846,15.930502,15.32316,14.715817,14.106662,13.499319,16.361988,19.224655,22.087322,24.949991,27.812658,25.490253,23.167849,20.845444,18.523039,16.200634,14.271642,12.344462,10.417283,8.490104,6.5629244,6.60281,6.642695,6.68258,6.722465,6.7623506,5.910258,5.0581656,4.2042603,3.3521678,2.5000753,2.2625773,2.0250793,1.7875811,1.550083,1.3125849,1.6624867,2.0123885,2.3622901,2.712192,3.0620937,3.2633326,3.4627585,3.6621845,3.8616104,4.062849,4.071914,4.082792,4.0918565,4.102734,4.1117992,4.274966,4.4381323,4.599486,4.762653,4.9258194,5.275721,5.6256227,5.975525,6.3254266,6.6753283,6.9382076,7.1992745,7.462154,7.7250338,7.987913,8.694968,9.402024,10.110892,10.817947,11.525003,10.990179,10.455356,9.920531,9.385707,8.8508835,10.460794,12.070704,13.680615,15.290526,16.900436,20.528175,24.1541,27.78184,31.409576,35.037315,34.477108,33.916904,33.356697,32.798306,32.238102,28.537844,24.837587,21.137331,17.437075,13.736817,12.895603,12.052575,11.209548,10.368333,9.525306,8.70222,7.8791356,7.057863,6.2347784,5.411693,4.4526362,3.491766,2.5327086,1.5718386,0.61278135,0.5275721,0.44236287,0.35715362,0.27194437,0.18673515,0.3045777,0.4224203,0.5402629,0.65810543,0.774135,1.2291887,1.6842422,2.1392958,2.5943494,3.049403,4.2441454,5.4407005,6.635443,7.8301854,9.024928,8.70222,8.379513,8.056806,7.7340984,7.413204,6.532104,5.6528172,4.7717175,3.8924308,3.0131438,3.1346123,3.2578938,3.3793623,3.5026438,3.6241121,3.9975824,4.36924,4.74271,5.1143675,5.487838,5.484212,5.482399,5.480586,5.47696,5.475147,5.678199,5.8794374,6.0824895,6.285541,6.48678,6.6155005,6.742408,6.869315,6.9980354,7.124943,6.8548117,6.58468,6.3145485,6.0444174,5.774286,5.660069,5.5458527,5.429823,5.315606,5.199577,5.524097,5.8504305,6.1749506,6.4994707,6.825804,6.7025228,6.5792413,6.4577727,6.3344913,6.2130227,6.01541,5.8177967,5.620184,5.422571,5.224958,5.565795,5.904819,6.245656,6.58468,6.925517,7.3968873,7.8700705,8.343254,8.814624,9.287807,7.850128,6.412449,4.974769,3.53709,2.0994108,1.6806163,1.260009,0.83940166,0.42060733,0.0,0.23931105,0.48043507,0.7197462,0.96087015,1.2001812,0.96087015,0.7197462,0.48043507,0.23931105,0.0,0.7197462,1.4394923,2.1592383,2.8807976,3.6005437,5.0128417,6.4251394,7.837437,9.249735,10.662033,9.969481,9.27693,8.584378,7.891826,7.1992745,6.784106,6.3707504,5.955582,5.540414,5.125245,4.1299286,3.1346123,2.1392958,1.1457924,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.14322405,0.17223145,0.2030518,0.23205921,0.26287958,0.24474995,0.22662032,0.21030366,0.19217403,0.17585737,0.17767033,0.1794833,0.18310922,0.18492219,0.18673515,0.3045777,0.4224203,0.5402629,0.65810543,0.774135,0.68167394,0.58921283,0.49675176,0.40429065,0.31182957,0.40791658,0.50219065,0.5982776,0.69255173,0.7868258,0.72518504,0.66173136,0.6000906,0.53663695,0.4749962,0.40429065,0.33539808,0.26469254,0.19579996,0.12509441,0.11965553,0.11421664,0.11059072,0.10515183,0.099712946,0.099712946,0.099712946,0.099712946,0.099712946,0.099712946,0.092461094,0.08520924,0.07795739,0.07070554,0.06164073,0.43692398,0.8122072,1.1874905,1.5627737,1.938057,1.5627737,1.1874905,0.8122072,0.43692398,0.06164073,0.15954071,0.2574407,0.35534066,0.45324063,0.5493277,0.64722764,0.7451276,0.8430276,0.93911463,1.0370146,0.86478317,0.69255173,0.52032024,0.3480888,0.17585737,0.23568514,0.2955129,0.35534066,0.41516843,0.4749962,1.7730774,3.0693457,4.367427,5.6655083,6.9617763,7.0143523,7.066928,7.119504,7.17208,7.224656,7.2953615,7.364254,7.4349594,7.5056653,7.574558,8.299743,9.024928,9.750113,10.475298,11.200482,10.002114,8.805559,7.607191,6.4106355,5.2122674,4.9167547,4.6230545,4.327542,4.0320287,3.738329,4.227829,4.7173285,5.2068286,5.6981416,6.187641,5.335549,4.4816437,3.6295512,2.7774587,1.9253663,1.649796,1.3742256,1.1004683,0.824898,0.5493277,0.50037766,0.44961473,0.40066472,0.34990177,0.2991388,1.1059072,1.9108626,2.715818,3.5207734,4.325729,3.6567454,2.9895754,2.322405,1.6552348,0.9880646,0.7995165,0.61278135,0.42423326,0.2374981,0.05076295,0.10696479,0.16497959,0.2229944,0.27919623,0.33721104,0.35715362,0.3770962,0.39703882,0.4169814,0.43692398,0.36984438,0.30276474,0.23568514,0.16679256,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.3154555,0.629098,0.9445535,1.260009,1.5754645,3.1182957,4.6593137,6.202145,7.744976,9.287807,9.353074,9.418341,9.481794,9.547061,9.612328,9.164526,8.716724,8.270736,7.8229337,7.3751316,6.7478466,6.1205616,5.4932766,4.8641787,4.2368937,4.064662,3.8924308,3.720199,3.5479677,3.3757362,4.41819,5.4606433,6.5030966,7.5455503,8.588004,8.013294,7.4367723,6.8620634,6.2873545,5.712645,5.618371,5.522284,5.42801,5.331923,5.237649,5.0654173,4.893186,4.7191415,4.5469103,4.3746786,5.317419,6.26016,7.2029004,8.145641,9.088382,9.353074,9.617766,9.882459,10.147152,10.411844,9.487233,8.562622,7.6380115,6.7134004,5.7869763,5.754343,5.7217097,5.6890764,5.658256,5.6256227,6.3344913,7.0451727,7.755854,8.464723,9.175404,11.597522,14.01964,16.441757,18.865688,21.287807,20.471973,19.657953,18.84212,18.0281,17.212267,17.533161,17.852243,18.173138,18.492218,18.813112,17.92476,17.038223,16.14987,15.263332,14.37498,14.083094,13.789393,13.497506,13.20562,12.91192,14.743011,16.57229,18.403383,20.232662,22.061941,24.077955,26.092157,28.108171,30.122374,32.136574,28.320288,24.50219,20.68409,16.867804,13.049705,12.915545,12.779573,12.645414,12.509441,12.375282,10.676537,8.979604,7.2826705,5.5857377,3.8869917,3.4119956,2.9369993,2.4620032,1.987007,1.5120108,1.789394,2.0667772,2.3441606,2.6233568,2.9007401,2.5997884,2.857229,3.1146698,3.3721104,3.6295512,3.8869917,3.6404288,3.392053,3.1454902,2.8971143,2.6505513,5.0726695,7.494787,9.916905,12.340837,14.762955,16.474392,18.187641,19.90089,21.612328,23.325577,21.815378,20.305182,18.794983,17.284784,15.774588,13.967064,12.15954,10.352016,8.544493,6.736969,6.591932,6.446895,6.301858,6.156821,6.011784,5.0744824,4.137181,3.199879,2.2625773,1.3252757,2.3532255,3.3793623,4.407312,5.4352617,6.4632115,6.01541,5.567608,5.1198063,4.6720047,4.2242026,6.7097745,9.195346,11.680918,14.164677,16.650248,15.934128,15.219821,14.505513,13.789393,13.075087,11.800573,10.524248,9.249735,7.9752226,6.70071,7.308052,7.915395,8.5227375,9.130079,9.737422,10.535126,11.332829,12.130532,12.928236,13.724127,13.544643,13.36516,13.185677,13.00438,12.824898,11.709926,10.594954,9.479981,8.365009,7.250037,7.115878,6.979906,6.8457465,6.7097745,6.5756154,8.832754,11.089892,13.347031,15.604169,17.863121,17.955582,18.048042,18.140503,18.232965,18.325426,18.18039,18.035353,17.890314,17.745277,17.60024,14.929747,12.259253,9.590572,6.9200783,4.249584,4.004834,3.7600844,3.5153344,3.2705846,3.0258346,3.5225863,4.019338,4.517903,5.0146546,5.5132194,7.1648283,8.81825,10.469859,12.123281,13.77489,13.238253,12.699803,12.163166,11.624716,11.088079,9.904215,8.722163,7.5401115,6.35806,5.1741953,7.7866745,10.399154,13.013446,15.625924,18.236591,18.127813,18.017221,17.906631,17.797853,17.687263,18.787731,19.888199,20.986855,22.087322,23.187792,22.045626,20.901646,19.75948,18.617313,17.475147,15.693004,13.910862,12.126906,10.344765,8.562622,8.1819,7.802991,7.422269,7.0433598,6.6626377,5.8921285,5.121619,4.3529234,3.5824142,2.811905,2.561716,2.3133402,2.0631514,1.8129625,1.5627737,1.7748904,1.987007,2.1991236,2.4130533,2.6251698,2.962381,3.299592,3.636803,3.975827,4.313038,4.329355,4.347484,4.365614,4.3819304,4.40006,4.537845,4.6756306,4.8116026,4.949388,5.087173,5.487838,5.8866897,6.2873545,6.688019,7.0868707,7.400513,7.7123427,8.024173,8.337815,8.649645,9.360326,10.069194,10.779876,11.490557,12.199425,11.595709,10.990179,10.384649,9.77912,9.175404,11.3056345,13.434052,15.564283,17.694515,19.824745,23.207733,26.590723,29.971897,33.354885,36.737873,35.807823,34.877773,33.947723,33.017673,32.087624,28.124489,24.163166,20.20003,16.236893,12.27557,12.010877,11.744371,11.479679,11.214987,10.950294,9.956791,8.9651,7.9715962,6.979906,5.9882154,4.933071,3.877927,2.8227828,1.7676386,0.7124943,0.6200332,0.5275721,0.43511102,0.34264994,0.25018883,0.27738327,0.3045777,0.33177215,0.36077955,0.387974,0.9898776,1.5917811,2.1954978,2.7974012,3.3993049,4.5849824,5.77066,6.9545245,8.140202,9.325879,8.72035,8.1148205,7.509291,6.9055743,6.300045,5.573047,4.844236,4.117238,3.39024,2.663242,2.955129,3.247016,3.540716,3.832603,4.12449,4.1933823,4.2604623,4.327542,4.3946214,4.461701,4.6303062,4.797099,4.9657044,5.132497,5.2992897,5.5077806,5.714458,5.922949,6.1296263,6.338117,6.445082,6.552047,6.6608243,6.7677894,6.874754,6.6644506,6.454147,6.245656,6.035352,5.825049,5.6800117,5.5349746,5.389938,5.2449007,5.0998635,5.600241,6.1006193,6.599184,7.0995617,7.5999393,7.308052,7.0143523,6.722465,6.430578,6.1368785,5.906632,5.678199,5.4479527,5.217706,4.98746,5.4207582,5.8522434,6.285541,6.717026,7.1503243,8.093065,9.035806,9.976733,10.919474,11.862214,10.049252,8.238102,6.4251394,4.612177,2.7992141,2.2408218,1.6806163,1.1204109,0.56020546,0.0,0.3208944,0.6399758,0.96087015,1.2799516,1.6008459,1.2799516,0.96087015,0.6399758,0.3208944,0.0,0.6979906,1.3941683,2.0921588,2.7901495,3.48814,5.5367875,7.5872483,9.637709,11.6881695,13.736817,12.910107,12.083396,11.254871,10.428161,9.599637,9.030367,8.459284,7.890013,7.320743,6.7496595,5.4407005,4.1299286,2.819157,1.5101979,0.19942589,0.15954071,0.11965553,0.07977036,0.03988518,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.19036107,0.23024625,0.27013144,0.3100166,0.34990177,0.3100166,0.27013144,0.23024625,0.19036107,0.15047589,0.15772775,0.16497959,0.17223145,0.1794833,0.18673515,0.22662032,0.26831847,0.30820364,0.3480888,0.387974,0.37165734,0.35715362,0.34264994,0.32814622,0.31182957,0.3480888,0.3825351,0.4169814,0.45324063,0.48768693,0.46230546,0.43692398,0.41335547,0.387974,0.36259252,0.3154555,0.26831847,0.21936847,0.17223145,0.12509441,0.12328146,0.11965553,0.11784257,0.11421664,0.11240368,0.11240368,0.11240368,0.11240368,0.11240368,0.11240368,0.10333887,0.092461094,0.08339628,0.072518505,0.06164073,0.51306844,0.96268314,1.4122978,1.8619126,2.3133402,1.8619126,1.4122978,0.96268314,0.51306844,0.06164073,0.16679256,0.27194437,0.3770962,0.48224804,0.5873999,0.6417888,0.6979906,0.7523795,0.80676836,0.8629702,0.7197462,0.57833505,0.43511102,0.291887,0.15047589,0.1794833,0.21030366,0.23931105,0.27013144,0.2991388,1.5682126,2.8354735,4.102734,5.369995,6.637256,6.4704633,6.301858,6.1350656,5.9682727,5.7996674,5.7470913,5.6945157,5.6419396,5.5893636,5.5367875,5.962834,6.3870673,6.813113,7.2373466,7.663393,7.0071006,6.352621,5.6981416,5.041849,4.3873696,4.115425,3.8416677,3.5697234,3.2977788,3.0258346,3.682127,4.3402324,4.9983377,5.65463,6.3127356,5.516845,4.7227674,3.926877,3.1327994,2.3369088,1.9743162,1.6117238,1.2491312,0.8883517,0.52575916,0.48768693,0.44961473,0.41335547,0.37528324,0.33721104,1.2908293,2.2426348,3.1944401,4.1480584,5.0998635,4.2223897,3.3449159,2.467442,1.5899682,0.7124943,0.5747091,0.43692398,0.2991388,0.16316663,0.025381476,0.11059072,0.19579996,0.27919623,0.36440548,0.44961473,0.47318324,0.4949388,0.5166943,0.5402629,0.5620184,0.4604925,0.35715362,0.25562772,0.15228885,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.36984438,0.73968875,1.1095331,1.4793775,1.8492218,3.2524548,4.655688,6.057108,7.460341,8.861761,8.870826,8.8780775,8.885329,8.892582,8.899834,8.357758,7.8156815,7.271793,6.7297173,6.187641,5.8304877,5.473334,5.1143675,4.7572136,4.40006,4.407312,4.4145637,4.421816,4.4308805,4.4381323,5.139749,5.8431783,6.544795,7.2482243,7.949841,7.8120556,7.6742706,7.5382986,7.400513,7.262728,7.077806,6.892884,6.7079616,6.5230393,6.338117,5.957395,5.576673,5.197764,4.8170414,4.4381323,5.389938,6.341743,7.2953615,8.247167,9.200785,9.3567,9.514427,9.672155,9.829884,9.987611,8.762048,7.5382986,6.3127356,5.087173,3.8616104,3.9395678,4.017525,4.0954823,4.171627,4.249584,4.954827,5.660069,6.3653116,7.0705543,7.7757964,10.230548,12.685299,15.140051,17.5948,20.049553,19.567305,19.085056,18.60281,18.120562,17.638313,17.94833,18.258347,18.568363,18.87838,19.188396,18.637255,18.087927,17.536787,16.98746,16.438131,15.709321,14.982323,14.255324,13.528327,12.799516,13.89092,14.98051,16.0701,17.15969,18.24928,20.544493,22.839703,25.134912,27.430124,29.725334,26.171928,22.620335,19.066927,15.515334,11.961927,11.920229,11.876718,11.83502,11.793322,11.74981,10.319383,8.888955,7.460341,6.0299134,4.599486,3.925064,3.2506418,2.5744069,1.8999848,1.2255627,1.6697385,2.1157274,2.5599031,3.004079,3.4500678,2.561716,2.8753586,3.1871881,3.5008307,3.8126602,4.12449,3.8616104,3.6005437,3.3376641,3.0747845,2.811905,5.2865987,7.763106,10.2378,12.712494,15.187187,16.563227,17.937452,19.311678,20.687716,22.061941,20.887142,19.712341,18.537542,17.362743,16.187943,14.211814,12.237497,10.263181,8.287052,6.3127356,6.0752378,5.8377395,5.600241,5.3627434,5.125245,4.249584,3.3757362,2.5000753,1.6244144,0.7505665,1.6244144,2.5000753,3.3757362,4.249584,5.125245,4.550536,3.975827,3.3993049,2.8245957,2.2498865,5.0617914,7.8755093,10.687414,13.499319,16.313038,15.600543,14.888049,14.175554,13.46306,12.750566,11.249433,9.750113,8.2507925,6.7496595,5.2503395,5.9120708,6.5756154,7.2373466,7.900891,8.562622,9.599637,10.636651,11.675479,12.712494,13.749508,13.399607,13.049705,12.699803,12.349901,11.999999,10.388275,8.774739,7.1630154,5.5494785,3.9377546,4.325729,4.7118897,5.0998635,5.487838,5.8758116,8.100317,10.324821,12.549327,14.775645,17.00015,16.400059,15.799969,15.199879,14.599788,13.999697,13.287203,12.574709,11.862214,11.14972,10.437225,8.999546,7.5618668,6.1241875,4.688321,3.2506418,3.149116,3.049403,2.94969,2.8499773,2.7502642,3.3630457,3.975827,4.5867953,5.199577,5.812358,7.5999393,9.38752,11.175101,12.962683,14.750263,14.224504,13.700559,13.174799,12.650853,12.125093,10.25049,8.375887,6.4994707,4.6248674,2.7502642,6.187641,9.625018,13.062395,16.499773,19.93715,20.325123,20.713097,21.099258,21.487232,21.875206,21.211662,20.54993,19.888199,19.224655,18.562923,18.599184,18.637255,18.675327,18.7134,18.749659,17.112555,15.475449,13.838344,12.199425,10.56232,9.762803,8.963287,8.161958,7.362441,6.5629244,5.8758116,5.186886,4.499773,3.8126602,3.1255474,2.8626678,2.5997884,2.3369088,2.0758421,1.8129625,1.887294,1.9616255,2.03777,2.1121013,2.1882458,2.663242,3.1382382,3.6132345,4.0882306,4.5632267,4.5867953,4.612177,4.6375585,4.6629395,4.688321,4.800725,4.9131284,5.0255322,5.137936,5.2503395,5.6999545,6.149569,6.599184,7.0506115,7.500226,7.8628187,8.225411,8.588004,8.950596,9.313189,10.025683,10.738177,11.450671,12.163166,12.87566,12.199425,11.525003,10.850581,10.174346,9.499924,12.1504755,14.799213,17.449764,20.100317,22.750868,25.887293,29.025532,32.161957,35.300194,38.43662,37.136726,35.83683,34.536938,33.23704,31.93715,27.712946,23.48693,19.262728,15.036712,10.812509,11.124338,11.437981,11.74981,12.06164,12.375282,11.213174,10.049252,8.887142,7.7250338,6.5629244,5.411693,4.262275,3.1128569,1.9616255,0.8122072,0.7124943,0.61278135,0.51306844,0.41335547,0.31182957,0.25018883,0.18673515,0.12509441,0.06164073,0.0,0.7505665,1.49932,2.2498865,3.000453,3.7492065,4.9258194,6.1006193,7.2754188,8.450218,9.625018,8.736667,7.850128,6.9617763,6.0752378,5.186886,4.612177,4.0374675,3.4627585,2.8880494,2.3133402,2.7756457,3.2379513,3.7002566,4.162562,4.6248674,4.3873696,4.1498713,3.9123733,3.6748753,3.437377,3.774588,4.1117992,4.4508233,4.788034,5.125245,5.337362,5.5494785,5.763408,5.975525,6.187641,6.2746634,6.3616858,6.450521,6.5375433,6.624565,6.4759026,6.3254266,6.1749506,6.0244746,5.8758116,5.6999545,5.52591,5.3500524,5.1741953,5.0001507,5.674573,6.350808,7.02523,7.699652,8.375887,7.911769,7.4494634,6.987158,6.5248523,6.0625467,5.7996674,5.5367875,5.275721,5.0128417,4.749962,5.275721,5.7996674,6.3254266,6.849373,7.3751316,8.78743,10.199727,11.612025,13.024323,14.436621,12.250188,10.061942,7.8755093,5.6872635,3.5008307,2.7992141,2.0994108,1.3996071,0.69980353,0.0,0.40066472,0.7995165,1.2001812,1.6008459,1.9996977,1.6008459,1.2001812,0.7995165,0.40066472,0.0,0.6744221,1.3506571,2.0250793,2.6995013,3.3757362,6.0625467,8.749357,11.437981,14.124791,16.811602,15.850732,14.888049,13.925365,12.962683,11.999999,11.274815,10.549629,9.824444,9.099259,8.375887,6.7496595,5.125245,3.5008307,1.8746033,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.2374981,0.28826106,0.33721104,0.387974,0.43692398,0.37528324,0.31182957,0.25018883,0.18673515,0.12509441,0.13778515,0.15047589,0.16316663,0.17585737,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.06164073,0.12509441,0.18673515,0.25018883,0.31182957,0.28826106,0.26287958,0.2374981,0.21211663,0.18673515,0.19942589,0.21211663,0.22480737,0.2374981,0.25018883,0.22480737,0.19942589,0.17585737,0.15047589,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.5873999,1.1131591,1.6371052,2.1628644,2.6868105,2.1628644,1.6371052,1.1131591,0.5873999,0.06164073,0.17585737,0.28826106,0.40066472,0.51306844,0.62547207,0.63816285,0.6508536,0.66173136,0.6744221,0.6871128,0.5747091,0.46230546,0.34990177,0.2374981,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,1.3633479,2.5997884,3.8380418,5.0744824,6.3127356,5.924762,5.5367875,5.1506267,4.762653,4.3746786,4.2006345,4.024777,3.8507326,3.6748753,3.5008307,3.6241121,3.7492065,3.874301,3.9993954,4.12449,4.0120864,3.8996825,3.787279,3.6748753,3.5624714,3.3122826,3.0620937,2.811905,2.561716,2.3133402,3.1382382,3.9631362,4.788034,5.612932,6.43783,5.6999545,4.9620786,4.2242026,3.48814,2.7502642,2.3006494,1.8492218,1.3996071,0.9499924,0.50037766,0.4749962,0.44961473,0.42423326,0.40066472,0.37528324,1.4757515,2.5744069,3.6748753,4.7753434,5.8758116,4.788034,3.7002566,2.612479,1.5247015,0.43692398,0.34990177,0.26287958,0.17585737,0.0870222,0.0,0.11240368,0.22480737,0.33721104,0.44961473,0.5620184,0.5873999,0.61278135,0.63816285,0.66173136,0.6871128,0.5493277,0.41335547,0.2755703,0.13778515,0.0,0.0,0.0,0.0,0.0,0.0,0.42423326,0.85027945,1.2745126,1.7005589,2.124792,3.388427,4.650249,5.9120708,7.175706,8.437528,8.386765,8.337815,8.287052,8.238102,8.187339,7.549176,6.9128265,6.2746634,5.638314,5.0001507,4.9131284,4.8242936,4.7372713,4.650249,4.5632267,4.749962,4.936697,5.125245,5.3119802,5.5005283,5.863121,6.2257137,6.588306,6.9490857,7.311678,7.61263,7.911769,8.212721,8.511859,8.812811,8.537241,8.26167,7.987913,7.7123427,7.4367723,6.849373,6.261973,5.674573,5.087173,4.499773,5.462456,6.4251394,7.3878226,8.350506,9.313189,9.362139,9.412902,9.461852,9.512614,9.563377,8.036863,6.5121617,4.98746,3.4627585,1.938057,2.124792,2.3133402,2.5000753,2.6868105,2.8753586,3.5751622,4.274966,4.974769,5.674573,6.3743763,8.861761,11.350959,13.838344,16.325727,18.813112,18.662638,18.512161,18.361685,18.213022,18.062546,18.361685,18.662638,18.961775,19.262728,19.561867,19.34975,19.137632,18.925516,18.7134,18.49947,17.33736,16.175253,15.013144,13.849221,12.687112,13.037014,13.386916,13.736817,14.0867195,14.436621,17.01284,19.587248,22.163467,24.737875,27.31228,24.025381,20.736666,17.449764,14.162864,10.874149,10.924912,10.975676,11.024626,11.075388,11.124338,9.96223,8.80012,7.6380115,6.4759026,5.3119802,4.4381323,3.5624714,2.6868105,1.8129625,0.93730164,1.550083,2.1628644,2.7756457,3.386614,3.9993954,2.5870976,2.817344,3.04759,3.2778363,3.5080826,3.738329,3.4700103,3.2016919,2.9351864,2.666868,2.4003625,4.5849824,6.7696023,8.954222,11.1406555,13.325275,14.78471,16.244144,17.705393,19.164827,20.624262,19.585434,18.544794,17.504154,16.465326,15.4246855,13.397794,11.370901,9.342196,7.315304,5.2865987,5.06723,4.847862,4.6266804,4.407312,4.1879435,3.5207734,2.8517902,2.18462,1.5174497,0.85027945,1.5446441,2.2408218,2.9351864,3.6295512,4.325729,3.972201,3.6204863,3.2669585,2.9152439,2.561716,4.9258194,7.28811,9.6504,12.012691,14.37498,13.820213,13.265448,12.710681,12.154101,11.599335,10.2958145,8.990481,7.6851482,6.379815,5.0744824,5.7833505,6.490406,7.1974616,7.9045167,8.613385,9.365765,10.118144,10.870523,11.622903,12.375282,12.0145035,11.655537,11.294757,10.93579,10.57501,9.275117,7.9752226,6.6753283,5.375434,4.07554,4.6230545,5.1705694,5.718084,6.265599,6.813113,8.780178,10.747242,12.714307,14.683184,16.650248,16.030214,15.410182,14.790149,14.170115,13.550082,12.810393,12.070704,11.329204,10.589515,9.849826,8.557183,7.264541,5.9718986,4.6792564,3.386614,3.4156215,3.442816,3.4700103,3.4972048,3.5243993,3.8597972,4.195195,4.5305934,4.8641787,5.199577,6.6644506,8.129324,9.594198,11.060884,12.525759,12.449615,12.375282,12.299138,12.224807,12.1504755,10.161655,8.174648,6.187641,4.2006345,2.2118144,5.0255322,7.837437,10.649343,13.46306,16.274965,17.163317,18.049856,18.938208,19.824745,20.713097,20.840004,20.966911,21.095633,21.22254,21.349447,20.55537,19.75948,18.9654,18.169512,17.375433,15.979452,14.585284,13.189302,11.795135,10.399154,9.702975,9.004985,8.306994,7.610817,6.9128265,6.09518,5.277534,4.459888,3.6422417,2.8245957,2.7176309,2.610666,2.5018883,2.3949237,2.2879589,2.4021754,2.518205,2.6324217,2.7466383,2.8626678,3.299592,3.738329,4.175253,4.612177,5.049101,5.0146546,4.9802084,4.945762,4.9095025,4.8750563,4.985647,5.0944247,5.2050157,5.315606,5.424384,5.7797246,6.1350656,6.490406,6.8457465,7.1992745,7.5781837,7.95528,8.3323765,8.709473,9.088382,9.73017,10.371959,11.015561,11.65735,12.299138,12.143224,11.985496,11.827768,11.67004,11.512312,13.822026,16.13174,18.443268,20.752983,23.062696,24.92461,26.788336,28.650248,30.51216,32.374073,31.541924,30.709774,29.877623,29.045473,28.213324,24.529385,20.847258,17.16513,13.483003,9.800876,9.842574,9.884272,9.927783,9.969481,10.012992,9.063,8.113008,7.1630154,6.2130227,5.2630305,4.3547363,3.4482548,2.5399606,1.6316663,0.72518504,0.6744221,0.62547207,0.5747091,0.52575916,0.4749962,0.46411842,0.4550536,0.44417584,0.43511102,0.42423326,1.2128719,1.9996977,2.7883365,3.5751622,4.361988,5.4370747,6.5121617,7.5872483,8.662335,9.737422,9.697536,9.657652,9.617766,9.577881,9.537996,8.597069,7.6579537,6.717026,5.7779117,4.836984,4.6357455,4.4326935,4.229642,4.028403,3.825351,3.7473936,3.6694362,3.5932918,3.5153344,3.437377,3.8054085,4.171627,4.539658,4.9076896,5.275721,5.3428006,5.40988,5.47696,5.5458527,5.612932,5.727149,5.8431783,5.957395,6.071612,6.187641,6.0244746,5.863121,5.6999545,5.5367875,5.375434,5.186886,5.0001507,4.8116026,4.6248674,4.4381323,5.0998635,5.7615952,6.4251394,7.0868707,7.750415,7.5854354,7.420456,7.2554765,7.0904965,6.925517,6.7442207,6.5647373,6.3852544,6.205771,6.0244746,6.5194135,7.0143523,7.509291,8.00423,8.499168,10.047439,11.595709,13.142166,14.690435,16.236893,13.671551,11.108022,8.54268,5.977338,3.4119956,2.7303216,2.0468347,1.3651608,0.68167394,0.0,0.3208944,0.6399758,0.96087015,1.2799516,1.6008459,1.3216497,1.0442665,0.7668832,0.4894999,0.21211663,1.8909199,3.5679104,5.2449007,6.921891,8.600695,10.422722,12.244749,14.066776,15.890617,17.712645,17.092611,16.472578,15.852545,15.2325115,14.612478,13.622601,12.632723,11.642846,10.652968,9.663091,8.239915,6.816739,5.3953767,3.972201,2.5508385,2.3205922,2.0903459,1.8600996,1.6298534,1.3996071,1.1494182,0.89922947,0.6508536,0.40066472,0.15047589,0.19036107,0.23024625,0.27013144,0.3100166,0.34990177,0.30276474,0.25562772,0.20667773,0.15954071,0.11240368,0.11965553,0.12690738,0.13415924,0.14322405,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.054388877,0.11059072,0.16497959,0.21936847,0.2755703,0.25562772,0.23568514,0.21574254,0.19579996,0.17585737,0.18673515,0.19942589,0.21211663,0.22480737,0.2374981,0.2229944,0.20667773,0.19217403,0.17767033,0.16316663,0.15772775,0.15228885,0.14684997,0.14322405,0.13778515,0.13778515,0.13778515,0.13778515,0.13778515,0.13778515,0.13415924,0.13234627,0.13053331,0.12690738,0.12509441,0.6000906,1.0750868,1.550083,2.0250793,2.5000753,2.0123885,1.5247015,1.0370146,0.5493277,0.06164073,0.1794833,0.29732585,0.41516843,0.533011,0.6508536,0.6653573,0.67986095,0.69436467,0.7106813,0.72518504,0.6091554,0.4949388,0.38072214,0.26469254,0.15047589,0.14684997,0.14503701,0.14322405,0.13959812,0.13778515,1.4304274,2.72307,4.0157123,5.3083544,6.599184,6.004532,5.40988,4.8152285,4.220577,3.6241121,3.484514,3.3449159,3.2053177,3.0657198,2.9243085,3.007705,3.0892882,3.1726844,3.254268,3.3376641,3.2506418,3.1618068,3.0747845,2.9877625,2.9007401,2.7031271,2.5055144,2.3079014,2.1102884,1.9126755,2.8608549,3.8072214,4.7554007,5.7017674,6.6499467,5.844991,5.040036,4.2350807,3.4301252,2.6251698,2.5345216,2.4456866,2.3550384,2.2643902,2.175555,1.8075237,1.4394923,1.0732739,0.70524246,0.33721104,1.3977941,2.4565642,3.5171473,4.5777307,5.638314,4.5867953,3.53709,2.4873846,1.4376793,0.387974,0.33721104,0.28826106,0.2374981,0.18673515,0.13778515,0.3480888,0.55839247,0.7668832,0.97718686,1.1874905,1.062396,0.93730164,0.8122072,0.6871128,0.5620184,0.44961473,0.33721104,0.22480737,0.11240368,0.0,0.0,0.0,0.0,0.0,0.0,0.5946517,1.1893034,1.7857682,2.38042,2.9750717,4.0030212,5.029158,6.057108,7.0850577,8.113008,8.096691,8.082188,8.067683,8.05318,8.036863,7.4820967,6.92733,6.3725634,5.8177967,5.2630305,5.2122674,5.163317,5.1125546,5.0617914,5.0128417,5.034597,5.0581656,5.0799212,5.101677,5.125245,5.812358,6.4994707,7.1883965,7.8755093,8.562622,8.595256,8.627889,8.660522,8.693155,8.725789,8.564435,8.404895,8.245354,8.0858135,7.9244595,7.440398,6.9545245,6.4704633,5.9845896,5.5005283,6.2746634,7.0506115,7.8247466,8.600695,9.374829,9.518054,9.659465,9.802689,9.944099,10.087324,8.898021,7.706904,6.5176005,5.328297,4.137181,4.49796,4.856927,5.217706,5.576673,5.9374523,6.5973706,7.2572894,7.9172077,8.577126,9.237044,10.964798,12.692551,14.420304,16.148058,17.87581,18.093367,18.310923,18.526665,18.74422,18.961775,19.17208,19.382383,19.592686,19.80299,20.013294,19.610817,19.208338,18.80586,18.403383,17.999092,16.784407,15.569723,14.355038,13.140353,11.925668,12.52032,13.114971,13.709623,14.304275,14.90074,17.114367,19.329807,21.545248,23.760687,25.974316,23.002869,20.02961,17.058165,14.084907,11.111648,10.955733,10.798005,10.640278,10.48255,10.324821,9.293246,8.259857,7.228282,6.1948934,5.163317,4.307599,3.4518807,2.5979755,1.742257,0.8883517,1.5101979,2.132044,2.7557032,3.3775494,3.9993954,2.612479,2.759329,2.907992,3.054842,3.2016919,3.350355,3.0765975,2.8046532,2.5327086,2.2607644,1.987007,3.8833659,5.7779117,7.6724577,9.567003,11.463363,13.008006,14.55265,16.097294,17.64194,19.186583,18.281914,17.377247,16.472578,15.567909,14.663241,12.581961,10.502492,8.423024,6.341743,4.262275,4.059223,3.8579843,3.6549325,3.4518807,3.2506418,2.7901495,2.3296568,1.8691645,1.4104849,0.9499924,1.4648738,1.9797552,2.4946365,3.009518,3.5243993,3.395679,3.2651455,3.1346123,3.005892,2.8753586,4.788034,6.70071,8.613385,10.524248,12.436923,12.039885,11.642846,11.245807,10.846955,10.449916,9.340384,8.23085,7.119504,6.009971,4.900438,5.6528172,6.4051967,7.157576,7.909956,8.662335,9.130079,9.597824,10.065568,10.533313,10.999244,10.629399,10.259555,9.88971,9.519867,9.1500225,8.161958,7.175706,6.187641,5.199577,4.213325,4.9203806,5.6274357,6.3344913,7.0433598,7.750415,9.460039,11.169662,12.879286,14.590723,16.300346,15.660371,15.020395,14.380419,13.740443,13.100468,12.331772,11.564888,10.798005,10.029309,9.262425,8.1148205,6.967215,5.81961,4.6720047,3.5243993,3.680314,3.834416,3.9903307,4.1444325,4.3003473,4.358362,4.4145637,4.4725785,4.5305934,4.5867953,5.730775,6.872941,8.015107,9.157274,10.29944,10.674724,11.050007,11.42529,11.800573,12.175857,10.074633,7.9752226,5.8758116,3.774588,1.6751775,3.8616104,6.049856,8.238102,10.424535,12.612781,13.999697,15.386614,16.775343,18.16226,19.549175,20.468348,21.385706,22.303066,23.220425,24.137783,22.509743,20.881702,19.255476,17.627436,15.999394,14.848164,13.695119,12.542075,11.390844,10.2378,9.643148,9.046683,8.452031,7.85738,7.262728,6.3145485,5.368182,4.420003,3.4718235,2.525457,2.572594,2.619731,2.666868,2.715818,2.762955,2.9170568,3.0729716,3.2270734,3.3829882,3.53709,3.9377546,4.3366065,4.7372713,5.137936,5.5367875,5.4425135,5.3482394,5.2521524,5.1578784,5.0617914,5.1705694,5.277534,5.384499,5.4932766,5.600241,5.859495,6.1205616,6.379815,6.640882,6.9001355,7.2917356,7.6851482,8.076748,8.470161,8.861761,9.434657,10.007553,10.58045,11.153346,11.724429,12.085209,12.444175,12.804955,13.165734,13.524701,15.495391,17.464268,19.43496,21.40565,23.374527,23.961926,24.549326,25.136726,25.724127,26.31334,25.94712,25.582714,25.21831,24.85209,24.487686,21.347635,18.207582,15.067532,11.927481,8.78743,8.560809,8.3323765,8.105756,7.877322,7.650702,6.9128265,6.1749506,5.4370747,4.699199,3.9631362,3.2977788,2.6324217,1.9670644,1.3017071,0.63816285,0.63816285,0.63816285,0.63816285,0.63816285,0.63816285,0.67986095,0.72337204,0.7650702,0.80676836,0.85027945,1.6751775,2.5000753,3.3249733,4.1498713,4.974769,5.9501433,6.925517,7.900891,8.874452,9.849826,10.656594,11.465176,12.271944,13.080525,13.887294,12.581961,11.27844,9.973107,8.667774,7.362441,6.495845,5.6274357,4.76084,3.8924308,3.0258346,3.1074178,3.1908143,3.2723975,3.3557937,3.437377,3.834416,4.233268,4.6303062,5.027345,5.424384,5.3482394,5.2702823,5.1923246,5.1143675,5.038223,5.179634,5.3228583,5.464269,5.6074934,5.750717,5.57486,5.4008155,5.224958,5.049101,4.8750563,4.6756306,4.4743915,4.274966,4.07554,3.874301,4.5251546,5.1741953,5.825049,6.4759026,7.124943,7.2572894,7.3896356,7.5219817,7.654328,7.7866745,7.690587,7.592687,7.494787,7.3968873,7.3008003,7.764919,8.23085,8.694968,9.1609,9.625018,11.307447,12.989877,14.672306,16.354736,18.037165,15.094727,12.152288,9.20985,6.2674117,3.3249733,2.659616,1.9942589,1.3307146,0.6653573,0.0,0.23931105,0.48043507,0.7197462,0.96087015,1.2001812,1.0442665,0.8901646,0.73424983,0.58014804,0.42423326,3.105605,5.7851634,8.464723,11.144281,13.825653,14.782897,15.740141,16.697386,17.654629,18.611874,18.33449,18.057108,17.779724,17.50234,17.224958,15.970387,14.715817,13.4594345,12.2048645,10.950294,9.73017,8.510046,7.2899227,6.069799,4.8496747,4.439945,4.0302157,3.6204863,3.2107568,2.7992141,2.2625773,1.7241274,1.1874905,0.6508536,0.11240368,0.14322405,0.17223145,0.2030518,0.23205921,0.26287958,0.23024625,0.19761293,0.16497959,0.13234627,0.099712946,0.10333887,0.10515183,0.10696479,0.11059072,0.11240368,0.09064813,0.06707962,0.045324065,0.02175555,0.0,0.047137026,0.09427405,0.14322405,0.19036107,0.2374981,0.2229944,0.20667773,0.19217403,0.17767033,0.16316663,0.17585737,0.18673515,0.19942589,0.21211663,0.22480737,0.21936847,0.21574254,0.21030366,0.20486477,0.19942589,0.19036107,0.1794833,0.17041849,0.15954071,0.15047589,0.15047589,0.15047589,0.15047589,0.15047589,0.15047589,0.15772775,0.16497959,0.17223145,0.1794833,0.18673515,0.61278135,1.0370146,1.4630609,1.887294,2.3133402,1.8619126,1.4122978,0.96268314,0.51306844,0.06164073,0.18492219,0.30820364,0.42967212,0.5529536,0.6744221,0.69255173,0.7106813,0.726998,0.7451276,0.76325727,0.64541465,0.5275721,0.40972954,0.291887,0.17585737,0.17041849,0.16497959,0.15954071,0.15410182,0.15047589,1.4975071,2.8445382,4.1933823,5.540414,6.887445,6.0843024,5.282973,4.4798307,3.6766882,2.8753586,2.770207,2.665055,2.5599031,2.4547513,2.3495996,2.3894846,2.42937,2.469255,2.5091403,2.5508385,2.4873846,2.4257438,2.3622901,2.3006494,2.2371957,2.0921588,1.9471219,1.8020848,1.6570477,1.5120108,2.5816586,3.6531196,4.7227674,5.7924156,6.8620634,5.9900284,5.1179934,4.2441454,3.3721104,2.5000753,2.770207,3.0403383,3.3104696,3.5806012,3.8507326,3.1400511,2.42937,1.7205015,1.0098201,0.2991388,1.3198367,2.3405347,3.3594196,4.3801174,5.4008155,4.3873696,3.3757362,2.3622901,1.3506571,0.33721104,0.3245203,0.31182957,0.2991388,0.28826106,0.2755703,0.581961,0.8901646,1.1983683,1.504759,1.8129625,1.5373923,1.261822,0.9880646,0.7124943,0.43692398,0.34990177,0.26287958,0.17585737,0.0870222,0.0,0.0,0.0,0.0,0.0,0.0,0.7650702,1.5301404,2.2952106,3.0602808,3.825351,4.6176157,5.40988,6.202145,6.9944096,7.7866745,7.806617,7.8283725,7.8483152,7.8682575,7.8882003,7.415017,6.9418335,6.4704633,5.99728,5.524097,5.5132194,5.5005283,5.487838,5.475147,5.462456,5.319232,5.177821,5.034597,4.893186,4.749962,5.763408,6.775041,7.7866745,8.80012,9.811753,9.577881,9.342196,9.108324,8.872639,8.636953,8.59163,8.548119,8.502794,8.457471,8.412147,8.029612,7.647076,7.264541,6.882006,6.4994707,7.0868707,7.6742706,8.26167,8.849071,9.438283,9.672155,9.907841,10.141713,10.377398,10.613083,9.757364,8.901647,8.047741,7.192023,6.338117,6.869315,7.402326,7.935337,8.4683485,8.999546,9.619579,10.239613,10.859646,11.479679,12.099712,13.067834,14.035956,15.002265,15.970387,16.936697,17.522284,18.10787,18.691645,19.277231,19.862818,19.982473,20.102129,20.221785,20.343254,20.462908,19.87007,19.277231,18.684393,18.093367,17.500528,16.233267,14.964193,13.696932,12.429671,11.162411,12.001812,12.843027,13.682428,14.521831,15.363045,17.217705,19.072367,20.927027,22.781689,24.63816,21.980358,19.322556,16.664753,14.006948,11.349146,10.98474,10.620335,10.254116,9.88971,9.525306,8.62245,7.7195945,6.816739,5.915697,5.0128417,4.177066,3.343103,2.5073273,1.6733645,0.8375887,1.4703126,2.1030366,2.7357605,3.3666716,3.9993954,2.6378605,2.7031271,2.7683938,2.8318477,2.8971143,2.962381,2.6849976,2.4076142,2.1302311,1.8528478,1.5754645,3.1799364,4.784408,6.390693,7.995165,9.599637,11.22949,12.859344,14.489197,16.120863,17.750717,16.980207,16.209698,15.439189,14.670493,13.899984,11.7679405,9.635896,7.502039,5.369995,3.2379513,3.053029,2.8681068,2.6831846,2.4982624,2.3133402,2.0595255,1.8075237,1.5555218,1.3017071,1.0497054,1.3851035,1.7205015,2.0558996,2.3894846,2.7248828,2.817344,2.909805,3.002266,3.094727,3.1871881,4.650249,6.11331,7.574558,9.037619,10.500679,10.259555,10.020245,9.77912,9.539809,9.300498,8.384952,7.4694057,6.5556726,5.6401267,4.7245803,5.522284,6.319988,7.117691,7.915395,8.713099,8.894395,9.077503,9.2606125,9.441909,9.625018,9.244296,8.865387,8.484665,8.105756,7.7250338,7.0506115,6.3743763,5.6999545,5.0255322,4.349297,5.217706,6.0843024,6.9527116,7.819308,8.6877165,10.139899,11.592083,13.044266,14.498261,15.950445,15.290526,14.630608,13.97069,13.310771,12.650853,11.854962,11.060884,10.264994,9.469104,8.675026,7.6724577,6.6698895,5.667321,4.664753,3.6621845,3.9450066,4.227829,4.510651,4.7916603,5.0744824,4.855114,4.6357455,4.4145637,4.195195,3.975827,4.795286,5.614745,6.434204,7.2554765,8.074935,8.899834,9.724731,10.549629,11.374527,12.199425,9.987611,7.7757964,5.562169,3.350355,1.1367276,2.6995013,4.262275,5.825049,7.3878226,8.950596,10.837891,12.725184,14.612478,16.499773,18.387066,20.094877,21.802689,23.510498,25.21831,26.924307,24.46593,22.00574,19.54555,17.08536,14.625169,13.715062,12.804955,11.894848,10.98474,10.074633,9.583321,9.090195,8.597069,8.105756,7.61263,6.53573,5.4570174,4.3801174,3.303218,2.2245052,2.427557,2.6306088,2.8318477,3.0348995,3.2379513,3.4319382,3.6277382,3.8217251,4.017525,4.213325,4.574105,4.936697,5.2992897,5.661882,6.0244746,5.870373,5.714458,5.560356,5.4044414,5.2503395,5.3554916,5.4606433,5.565795,5.669134,5.774286,5.9392653,6.104245,6.2692246,6.434204,6.599184,7.0071006,7.415017,7.8229337,8.23085,8.636953,9.139144,9.643148,10.145339,10.64753,11.14972,12.027194,12.904668,13.782142,14.6596155,15.537089,17.166943,18.796797,20.428463,22.058315,23.68817,22.999243,22.31213,21.625017,20.937904,20.250792,20.352318,20.455656,20.557182,20.660522,20.762047,18.165886,15.567909,12.969934,10.371959,7.7757964,7.2772317,6.78048,6.281915,5.7851634,5.2865987,4.762653,4.2368937,3.7129474,3.1871881,2.663242,2.2408218,1.8184015,1.3941683,0.97174793,0.5493277,0.6000906,0.6508536,0.69980353,0.7505665,0.7995165,0.89560354,0.9898776,1.0841516,1.1802386,1.2745126,2.137483,3.000453,3.8634233,4.7245803,5.5875506,6.4632115,7.3370595,8.212721,9.088382,9.96223,11.617464,13.272699,14.927934,16.583168,18.238403,16.566853,14.897114,13.227375,11.557636,9.8878975,8.355945,6.8221784,5.290225,3.7582715,2.2245052,2.467442,2.7103791,2.953316,3.1944401,3.437377,3.8652363,4.2930956,4.7191415,5.147001,5.57486,5.351866,5.130684,4.9076896,4.6846952,4.461701,4.632119,4.802538,4.972956,5.143375,5.3119802,5.125245,4.936697,4.749962,4.5632267,4.3746786,4.162562,3.9504454,3.738329,3.5243993,3.3122826,3.9504454,4.5867953,5.224958,5.863121,6.4994707,6.929143,7.360628,7.7903004,8.219973,8.649645,8.63514,8.620637,8.604321,8.589817,8.575313,9.010424,9.445535,9.880646,10.315757,10.750868,12.567456,14.385859,16.202446,18.020847,19.837437,16.517902,13.198368,9.87702,6.5574856,3.2379513,2.5907235,1.9416829,1.2944553,0.64722764,0.0,0.15954071,0.3208944,0.48043507,0.6399758,0.7995165,0.7668832,0.73424983,0.7016165,0.67079616,0.63816285,4.3202896,8.002417,11.684544,15.368484,19.050611,19.143072,19.235533,19.327993,19.420456,19.512917,19.578182,19.641636,19.706903,19.77217,19.837437,18.318174,16.797098,15.277836,13.75676,12.237497,11.220426,10.203354,9.184468,8.167397,7.1503243,6.5592985,5.9700856,5.3808727,4.7898474,4.2006345,3.3757362,2.5508385,1.7241274,0.89922947,0.07433146,0.09427405,0.11421664,0.13415924,0.15410182,0.17585737,0.15772775,0.13959812,0.12328146,0.10515183,0.0870222,0.08520924,0.08339628,0.07977036,0.07795739,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.03988518,0.07977036,0.11965553,0.15954071,0.19942589,0.19036107,0.1794833,0.17041849,0.15954071,0.15047589,0.16316663,0.17585737,0.18673515,0.19942589,0.21211663,0.21755551,0.2229944,0.22662032,0.23205921,0.2374981,0.2229944,0.20667773,0.19217403,0.17767033,0.16316663,0.16316663,0.16316663,0.16316663,0.16316663,0.16316663,0.1794833,0.19761293,0.21574254,0.23205921,0.25018883,0.62547207,1.0007553,1.3742256,1.7495089,2.124792,1.7132497,1.2998942,0.8883517,0.4749962,0.06164073,0.19036107,0.31726846,0.44417584,0.5728962,0.69980353,0.7197462,0.73968875,0.75963134,0.7795739,0.7995165,0.67986095,0.56020546,0.4405499,0.3208944,0.19942589,0.19217403,0.18492219,0.17767033,0.17041849,0.16316663,1.5645868,2.9678197,4.36924,5.772473,7.175706,6.164073,5.1542525,4.1444325,3.1346123,2.124792,2.0540867,1.9851941,1.9144884,1.845596,1.7748904,1.7730774,1.7694515,1.7676386,1.7658255,1.7621996,1.7241274,1.6878681,1.649796,1.6117238,1.5754645,1.4830034,1.3905423,1.2980812,1.2056202,1.1131591,2.3042755,3.4972048,4.690134,5.883064,7.07418,6.1350656,5.1941376,4.255023,3.3140955,2.374981,3.005892,3.63499,4.265901,4.894999,5.52591,4.4725785,3.4192474,2.3677292,1.3143979,0.26287958,1.2418793,2.222692,3.2016919,4.1825047,5.163317,4.1879435,3.2125697,2.2371957,1.261822,0.28826106,0.31182957,0.33721104,0.36259252,0.387974,0.41335547,0.81764615,1.2219368,1.6280404,2.032331,2.4366217,2.0123885,1.5881553,1.162109,0.73787576,0.31182957,0.25018883,0.18673515,0.12509441,0.06164073,0.0,0.0,0.0,0.0,0.0,0.0,0.9354887,1.8691645,2.8046532,3.7401419,4.6756306,5.23221,5.7906027,6.347182,6.9055743,7.462154,7.518356,7.572745,7.6271334,7.6833353,7.7377243,7.3479376,6.9581504,6.5683637,6.1767635,5.7869763,5.812358,5.8377395,5.863121,5.8866897,5.9120708,5.6056805,5.297477,4.989273,4.6828823,4.3746786,5.712645,7.0506115,8.386765,9.724731,11.062697,10.560507,10.058316,9.554313,9.052122,8.549932,8.620637,8.689529,8.760235,8.829127,8.899834,8.620637,8.339628,8.0604315,7.7794223,7.500226,7.900891,8.299743,8.700407,9.099259,9.499924,9.82807,10.154404,10.48255,10.810696,11.137029,10.616709,10.098202,9.577881,9.057561,8.537241,9.242483,9.947725,10.652968,11.358211,12.06164,12.6417885,13.221936,13.802084,14.382232,14.96238,15.170871,15.377548,15.584227,15.792717,15.999394,16.953012,17.904818,18.858437,19.810242,20.762047,20.792868,20.821875,20.852695,20.881702,20.912523,20.129324,19.347937,18.564737,17.78335,17.00015,15.680313,14.3604765,13.04064,11.720803,10.399154,11.485118,12.569269,13.655234,14.739386,15.825351,17.319231,18.814926,20.31062,21.8045,23.300196,20.957848,18.6155,16.273151,13.930804,11.586644,11.015561,10.442664,9.869768,9.296872,8.725789,7.951654,7.179332,6.4070096,5.634688,4.8623657,4.0483456,3.2325122,2.4166791,1.6026589,0.7868258,1.4304274,2.0722163,2.715818,3.3576066,3.9993954,2.663242,2.6451125,2.6269827,2.610666,2.5925364,2.5744069,2.2933977,2.0105755,1.7277533,1.4449311,1.162109,2.47832,3.7927177,5.1071157,6.4233265,7.7377243,9.452786,11.16785,12.882912,14.597975,16.313038,15.676687,15.0421505,14.407614,13.773077,13.136727,10.952107,8.767487,6.582867,4.3982472,2.2118144,2.0450218,1.8782293,1.7096237,1.5428312,1.3742256,1.3307146,1.2853905,1.2400664,1.1947423,1.1494182,1.305333,1.4594349,1.6153497,1.7694515,1.9253663,2.2408218,2.5544643,2.8699198,3.1853752,3.5008307,4.512464,5.524097,6.5375433,7.549176,8.562622,8.479226,8.397643,8.314246,8.232663,8.149267,7.4295206,6.7097745,5.9900284,5.2702823,4.550536,5.391751,6.2347784,7.077806,7.9208336,8.762048,8.660522,8.557183,8.455658,8.352319,8.2507925,7.859193,7.4694057,7.079619,6.6898317,6.300045,5.9374523,5.57486,5.2122674,4.8496747,4.4870825,5.5150323,6.542982,7.570932,8.597069,9.625018,10.81976,12.0145035,13.209246,14.405801,15.600543,14.920682,14.240821,13.559147,12.879286,12.199425,11.378153,10.555068,9.731983,8.910711,8.087626,7.230095,6.3725634,5.5150323,4.6575007,3.7999697,4.209699,4.6194286,5.029158,5.4407005,5.8504305,5.351866,4.855114,4.358362,3.8597972,3.3630457,3.8597972,4.358362,4.855114,5.351866,5.8504305,7.124943,8.399456,9.675781,10.950294,12.224807,9.900589,7.574558,5.2503395,2.9243085,0.6000906,1.5373923,2.474694,3.4119956,4.349297,5.2884116,7.6742706,10.061942,12.449615,14.837286,17.224958,19.72322,22.21967,24.717932,27.214382,29.712645,26.420303,23.127964,19.835623,16.543283,13.24913,12.581961,11.91479,11.24762,10.58045,9.91328,9.52168,9.131892,8.7421055,8.352319,7.9625316,6.755099,5.5476656,4.3402324,3.1327994,1.9253663,2.2825198,2.6396735,2.9968271,3.3557937,3.7129474,3.9468195,4.1825047,4.41819,4.652062,4.8877473,5.2122674,5.5367875,5.863121,6.187641,6.5121617,6.298232,6.0824895,5.866747,5.6528172,5.4370747,5.540414,5.6419396,5.7452784,5.846804,5.9501433,6.0208488,6.089741,6.1604466,6.2293396,6.300045,6.722465,7.1448855,7.567306,7.989726,8.412147,8.845445,9.27693,9.710228,10.141713,10.57501,11.969179,13.36516,14.759329,16.15531,17.549479,18.840307,20.129324,21.420153,22.70917,23.999998,22.038374,20.074934,18.11331,16.14987,14.188245,14.757515,15.326786,15.897869,16.467138,17.038223,14.982323,12.928236,10.872336,8.81825,6.7623506,5.995467,5.2267714,4.459888,3.6930048,2.9243085,2.612479,2.3006494,1.987007,1.6751775,1.3633479,1.1820517,1.0025684,0.823085,0.6417888,0.46230546,0.5620184,0.66173136,0.76325727,0.8629702,0.96268314,1.1095331,1.258196,1.405046,1.551896,1.7005589,2.5997884,3.5008307,4.40006,5.2992897,6.200332,6.9744673,7.750415,8.52455,9.300498,10.074633,12.578335,15.080223,17.582111,20.085812,22.5877,20.551744,18.5176,16.481644,14.447499,12.413355,10.2142315,8.01692,5.81961,3.6222992,1.4249886,1.8274662,2.229944,2.6324217,3.0348995,3.437377,3.8942437,4.3529234,4.8097897,5.2666564,5.7253356,5.3573046,4.989273,4.6230545,4.255023,3.8869917,4.0846047,4.2822175,4.4798307,4.6774435,4.8750563,4.6756306,4.4743915,4.274966,4.07554,3.874301,3.6494937,3.4246864,3.199879,2.9750717,2.7502642,3.3757362,3.9993954,4.6248674,5.2503395,5.8758116,6.60281,7.3298078,8.056806,8.785617,9.512614,9.579695,9.646774,9.715667,9.782746,9.849826,10.254116,10.66022,11.06451,11.470614,11.874905,13.827466,15.780026,17.732588,19.685148,21.637709,17.939264,14.242634,10.54419,6.8475595,3.149116,2.520018,1.8909199,1.260009,0.629098,0.0,0.07977036,0.15954071,0.23931105,0.3208944,0.40066472,0.4894999,0.58014804,0.67079616,0.75963134,0.85027945,5.5349746,10.21967,14.904366,19.590874,24.27557,23.503246,22.729113,21.956789,21.184467,20.412146,20.820063,21.22798,21.635895,22.042,22.449915,20.664148,18.880192,17.094423,15.310469,13.524701,12.710681,11.894848,11.080828,10.264994,9.449161,8.680465,7.909956,7.1394467,6.3707504,5.600241,4.4870825,3.3757362,2.2625773,1.1494182,0.038072214,0.047137026,0.058014803,0.06707962,0.07795739,0.0870222,0.08520924,0.08339628,0.07977036,0.07795739,0.07433146,0.06707962,0.059827764,0.052575916,0.045324065,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.032633327,0.065266654,0.09789998,0.13053331,0.16316663,0.15772775,0.15228885,0.14684997,0.14322405,0.13778515,0.15047589,0.16316663,0.17585737,0.18673515,0.19942589,0.21574254,0.23024625,0.24474995,0.25925365,0.2755703,0.25562772,0.23568514,0.21574254,0.19579996,0.17585737,0.17585737,0.17585737,0.17585737,0.17585737,0.17585737,0.2030518,0.23024625,0.2574407,0.28463513,0.31182957,0.63816285,0.96268314,1.2872034,1.6117238,1.938057,1.5627737,1.1874905,0.8122072,0.43692398,0.06164073,0.19579996,0.32814622,0.4604925,0.59283876,0.72518504,0.7469406,0.7705091,0.79226464,0.81583315,0.8375887,0.71430725,0.59283876,0.46955732,0.3480888,0.22480737,0.21574254,0.20486477,0.19579996,0.18492219,0.17585737,1.6334792,3.0892882,4.5469103,6.004532,7.462154,6.245656,5.027345,3.8108473,2.5925364,1.3742256,1.3397794,1.305333,1.2708868,1.2346275,1.2001812,1.1548572,1.1095331,1.064209,1.020698,0.97537386,0.96268314,0.9499924,0.93730164,0.9246109,0.9119202,0.872035,0.8321498,0.79226464,0.7523795,0.7124943,2.0268922,3.343103,4.6575007,5.9718986,7.28811,6.2801023,5.272095,4.264088,3.2578938,2.2498865,3.2397642,4.229642,5.219519,6.209397,7.1992745,5.805106,4.410938,3.0149567,1.6207886,0.22480737,1.1657349,2.1048496,3.045777,3.9848917,4.9258194,3.9867048,3.049403,2.1121013,1.1747998,0.2374981,0.2991388,0.36259252,0.42423326,0.48768693,0.5493277,1.0533313,1.5555218,2.0577126,2.5599031,3.0620937,2.4873846,1.9126755,1.3379664,0.76325727,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.0,0.0,0.0,0.0,0.0,1.1059072,2.2100015,3.3159087,4.420003,5.524097,5.846804,6.169512,6.492219,6.814926,7.137634,7.228282,7.317117,7.407765,7.4966,7.5872483,7.2808576,6.972654,6.6644506,6.35806,6.049856,6.11331,6.1749506,6.2384043,6.300045,6.3616858,5.8903155,5.4171324,4.945762,4.4725785,3.9993954,5.661882,7.324369,8.9868555,10.649343,12.311829,11.543133,10.772624,10.002114,9.233418,8.46291,8.647832,8.832754,9.017676,9.202598,9.38752,9.20985,9.03218,8.854509,8.676839,8.499168,8.713099,8.925215,9.137331,9.349448,9.563377,9.982172,10.40278,10.823386,11.242181,11.662788,11.477866,11.292944,11.108022,10.9230995,10.738177,11.615651,12.493125,13.370599,14.248073,15.125546,15.66581,16.20426,16.744522,17.284784,17.825048,17.272095,16.719141,16.168001,15.6150465,15.062093,16.38193,17.701767,19.023417,20.343254,21.66309,21.603262,21.541622,21.481794,21.421967,21.362139,20.39039,19.41683,18.445082,17.473333,16.499773,15.127359,13.754947,12.382534,11.010121,9.637709,10.968424,12.297325,13.628039,14.956942,16.287657,17.422571,18.557486,19.6924,20.827314,21.962229,19.935337,17.906631,15.879739,13.852847,11.8241415,11.044568,10.264994,9.48542,8.705847,7.9244595,7.2826705,6.639069,5.99728,5.3554916,4.7118897,3.917812,3.1219215,2.327844,1.5319533,0.73787576,1.3905423,2.0432088,2.6958754,3.346729,3.9993954,2.6868105,2.5870976,2.4873846,2.3876717,2.2879589,2.1882458,1.8999848,1.6117238,1.3252757,1.0370146,0.7505665,1.7748904,2.7992141,3.825351,4.8496747,5.8758116,7.6742706,9.474543,11.274815,13.075087,14.875358,14.37498,13.874602,13.374225,12.87566,12.375282,10.138086,7.900891,5.661882,3.4246864,1.1874905,1.0370146,0.8883517,0.73787576,0.5873999,0.43692398,0.6000906,0.76325727,0.9246109,1.0877775,1.2491312,1.2255627,1.2001812,1.1747998,1.1494182,1.1258497,1.6624867,2.1991236,2.7375734,3.2742105,3.8126602,4.3746786,4.936697,5.5005283,6.0625467,6.624565,6.70071,6.775041,6.849373,6.925517,6.9998484,6.4759026,5.9501433,5.424384,4.900438,4.3746786,5.2630305,6.149569,7.037921,7.9244595,8.812811,8.424837,8.036863,7.650702,7.262728,6.874754,6.4759026,6.0752378,5.674573,5.275721,4.8750563,4.8242936,4.7753434,4.7245803,4.6756306,4.6248674,5.812358,6.9998484,8.187339,9.374829,10.56232,11.499621,12.436923,13.374225,14.313339,15.250641,14.5508375,13.849221,13.149418,12.449615,11.74981,10.899531,10.049252,9.200785,8.350506,7.500226,6.787732,6.0752378,5.3627434,4.650249,3.9377546,4.4743915,5.0128417,5.5494785,6.0879283,6.624565,5.8504305,5.0744824,4.3003473,3.5243993,2.7502642,2.9243085,3.100166,3.2742105,3.4500678,3.6241121,5.3500524,7.07418,8.80012,10.524248,12.250188,9.811753,7.3751316,4.936697,2.5000753,0.06164073,0.37528324,0.6871128,1.0007553,1.3125849,1.6244144,4.512464,7.400513,10.28675,13.174799,16.062849,19.34975,22.63665,25.925365,29.212267,32.49917,28.374678,24.250187,20.125698,15.999394,11.874905,11.450671,11.024626,10.600392,10.174346,9.750113,9.461852,9.175404,8.887142,8.600695,8.312433,6.9744673,5.638314,4.3003473,2.962381,1.6244144,2.137483,2.6505513,3.1618068,3.6748753,4.1879435,4.461701,4.7372713,5.0128417,5.2865987,5.562169,5.8504305,6.1368785,6.4251394,6.7134004,6.9998484,6.7242785,6.450521,6.1749506,5.89938,5.6256227,5.7253356,5.825049,5.924762,6.0244746,6.1241875,6.1006193,6.0752378,6.049856,6.0244746,6.000906,6.43783,6.874754,7.311678,7.750415,8.187339,8.549932,8.912524,9.275117,9.637709,10.000301,11.912977,13.825653,15.738328,17.64919,19.561867,20.511858,21.461851,22.411844,23.361835,24.311829,21.07569,17.837738,14.599788,11.361836,8.125698,9.162713,10.199727,11.236742,12.27557,13.312584,11.800573,10.28675,8.774739,7.262728,5.750717,4.7118897,3.6748753,2.6378605,1.6008459,0.5620184,0.46230546,0.36259252,0.26287958,0.16316663,0.06164073,0.12509441,0.18673515,0.25018883,0.31182957,0.37528324,0.52575916,0.6744221,0.824898,0.97537386,1.1258497,1.3252757,1.5247015,1.7241274,1.9253663,2.124792,3.0620937,3.9993954,4.936697,5.8758116,6.813113,7.4875355,8.161958,8.838193,9.512614,10.1870365,13.537392,16.887747,20.238102,23.588457,26.936998,24.536636,22.138086,19.737724,17.33736,14.936998,12.07433,9.213476,6.350808,3.48814,0.62547207,1.1874905,1.7495089,2.3133402,2.8753586,3.437377,3.925064,4.4127507,4.900438,5.388125,5.8758116,5.3627434,4.8496747,4.3366065,3.825351,3.3122826,3.53709,3.7618973,3.9867048,4.213325,4.4381323,4.2242026,4.0120864,3.7999697,3.587853,3.3757362,3.1382382,2.9007401,2.663242,2.4257438,2.1882458,2.7992141,3.4119956,4.024777,4.6375585,5.2503395,6.2746634,7.3008003,8.325124,9.349448,10.375585,10.524248,10.674724,10.825199,10.975676,11.124338,11.499621,11.874905,12.250188,12.625471,13.000754,15.087475,17.174194,19.262728,21.349447,23.43798,19.36244,15.2869005,11.213174,7.137634,3.0620937,2.4493124,1.8383441,1.2255627,0.61278135,0.0,0.0,0.0,0.0,0.0,0.0,0.21211663,0.42423326,0.63816285,0.85027945,1.062396,6.7496595,12.436923,18.126,23.813263,29.500526,27.861609,26.224504,24.587399,22.950293,21.313189,22.061941,22.812508,23.563074,24.311829,25.062395,23.011934,20.963285,18.912827,16.862366,14.811904,14.199123,13.588155,12.975373,12.362592,11.74981,10.799818,9.849826,8.899834,7.949841,6.9998484,5.600241,4.2006345,2.7992141,1.3996071,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.13778515,0.15047589,0.16316663,0.17585737,0.18673515,0.21211663,0.2374981,0.26287958,0.28826106,0.31182957,0.28826106,0.26287958,0.2374981,0.21211663,0.18673515,0.18673515,0.18673515,0.18673515,0.18673515,0.18673515,0.22480737,0.26287958,0.2991388,0.33721104,0.37528324,0.6508536,0.9246109,1.2001812,1.4757515,1.7495089,1.4122978,1.0750868,0.73787576,0.40066472,0.06164073,0.19942589,0.33721104,0.4749962,0.61278135,0.7505665,0.774135,0.7995165,0.824898,0.85027945,0.87566096,0.7505665,0.62547207,0.50037766,0.37528324,0.25018883,0.2374981,0.22480737,0.21211663,0.19942589,0.18673515,1.7005589,3.2125697,4.7245803,6.2384043,7.750415,6.3254266,4.900438,3.4754493,2.0504606,0.62547207,0.62547207,0.62547207,0.62547207,0.62547207,0.62547207,0.53663695,0.44961473,0.36259252,0.2755703,0.18673515,0.19942589,0.21211663,0.22480737,0.2374981,0.25018883,0.26287958,0.2755703,0.28826106,0.2991388,0.31182957,1.7495089,3.1871881,4.6248674,6.0625467,7.500226,6.4251394,5.3500524,4.274966,3.199879,2.124792,3.4754493,4.8242936,6.1749506,7.5256076,8.874452,7.137634,5.4008155,3.6621845,1.9253663,0.18673515,1.0877775,1.987007,2.8880494,3.787279,4.688321,3.787279,2.8880494,1.987007,1.0877775,0.18673515,0.28826106,0.387974,0.48768693,0.5873999,0.6871128,1.2872034,1.887294,2.4873846,3.0874753,3.6875658,2.962381,2.2371957,1.5120108,0.7868258,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,1.2745126,2.5508385,3.825351,5.0998635,6.3743763,6.4632115,6.550234,6.637256,6.7242785,6.813113,6.9382076,7.063302,7.1883965,7.311678,7.4367723,7.211965,6.987158,6.7623506,6.5375433,6.3127356,6.412449,6.5121617,6.6118746,6.7134004,6.813113,6.1749506,5.5367875,4.900438,4.262275,3.6241121,5.612932,7.5999393,9.5869465,11.575767,13.562773,12.525759,11.486931,10.449916,9.412902,8.375887,8.675026,8.974165,9.275117,9.574255,9.875207,9.800876,9.724731,9.6504,9.574255,9.499924,9.525306,9.550687,9.574255,9.599637,9.625018,10.138086,10.649343,11.162411,11.675479,12.186734,12.337211,12.487686,12.638163,12.786825,12.937301,13.987006,15.036712,16.08823,17.137936,18.187641,18.688019,19.186583,19.68696,20.187338,20.687716,19.375132,18.062546,16.749962,15.437376,14.124791,15.812659,17.500528,19.188396,20.87445,22.562319,22.411844,22.26318,22.112705,21.962229,21.811752,20.649643,19.487535,18.325426,17.163317,15.999394,14.574407,13.149418,11.724429,10.29944,8.874452,10.449916,12.025381,13.600845,15.174497,16.749962,17.52591,18.300045,19.074179,19.850128,20.624262,18.912827,17.199575,15.488139,13.77489,12.06164,11.075388,10.087324,9.099259,8.113008,7.124943,6.6118746,6.1006193,5.5875506,5.0744824,4.5632267,3.787279,3.0131438,2.2371957,1.4630609,0.6871128,1.3506571,2.0123885,2.6741197,3.3376641,3.9993954,2.374981,2.2825198,2.1900587,2.0975976,2.0051367,1.9126755,1.6552348,1.3977941,1.1403534,0.88291276,0.62547207,1.6878681,2.7502642,3.8126602,4.8750563,5.9374523,8.027799,10.118144,12.206677,14.297023,16.38737,15.805408,15.221634,14.639673,14.057712,13.475751,11.030065,8.584378,6.1405044,3.6948178,1.2491312,1.2654479,1.2799516,1.2944553,1.310772,1.3252757,1.261822,1.2001812,1.1367276,1.0750868,1.0116332,1.0043813,0.99712944,0.9898776,0.9826257,0.97537386,1.5881553,2.1991236,2.811905,3.4246864,4.0374675,4.782595,5.527723,6.2728505,7.017978,7.763106,7.755854,7.746789,7.7395372,7.7322855,7.7250338,7.0451727,6.3653116,5.6854506,5.0055895,4.325729,5.045475,5.765221,6.484967,7.2047133,7.9244595,8.392203,8.859948,9.327692,9.795437,10.263181,9.570629,8.8780775,8.185526,7.4929743,6.8004227,7.2572894,7.7141557,8.172835,8.629702,9.088382,10.549629,12.012691,13.475751,14.936998,16.400059,16.171627,15.945006,15.718386,15.489952,15.263332,14.567154,13.872789,13.176612,12.482247,11.787883,10.995618,10.203354,9.409276,8.617011,7.8247466,7.1267557,6.430578,5.732588,5.034597,4.3366065,4.6176157,4.896812,5.177821,5.4570174,5.7380266,5.1107416,4.4816437,3.8543584,3.2270734,2.5997884,3.0403383,3.4808881,3.919625,4.360175,4.800725,6.1006193,7.400513,8.700407,10.000301,11.300196,9.155461,7.0107265,4.8641787,2.7194438,0.5747091,0.7650702,0.9554313,1.1457924,1.3343405,1.5247015,4.517903,7.509291,10.502492,13.495693,16.487082,18.515787,20.542679,22.56957,24.598276,26.625168,24.69255,22.759932,20.827314,18.894695,16.962078,15.250641,13.537392,11.8241415,10.112705,8.399456,8.080374,7.75948,7.440398,7.119504,6.8004227,5.774286,4.749962,3.7256382,2.6995013,1.6751775,2.1719291,2.6704938,3.1672456,3.6658103,4.162562,4.7554007,5.3482394,5.9392653,6.532104,7.124943,7.1466985,7.170267,7.192023,7.215591,7.2373466,6.965402,6.6916447,6.4197006,6.147756,5.8758116,6.189454,6.5049095,6.8203654,7.135821,7.4494634,7.2826705,7.115878,6.947273,6.78048,6.6118746,6.9744673,7.3370595,7.699652,8.062244,8.424837,8.890768,9.354887,9.820818,10.284937,10.750868,12.67986,14.610665,16.539658,18.470463,20.399454,20.535427,20.669586,20.80556,20.939718,21.07569,18.314548,15.555219,12.794077,10.034748,7.2754188,8.370448,9.465478,10.560507,11.655537,12.750566,11.3056345,9.860703,8.415772,6.970841,5.524097,4.7227674,3.919625,3.1182957,2.3151531,1.5120108,1.2400664,0.968122,0.69436467,0.4224203,0.15047589,0.36440548,0.58014804,0.79589057,1.0098201,1.2255627,1.1856775,1.1457924,1.1040943,1.064209,1.0243238,1.1602961,1.2944553,1.4304274,1.5645868,1.7005589,2.5073273,3.3140955,4.122677,4.9294453,5.7380266,6.836682,7.93715,9.037619,10.138086,11.236742,14.817343,18.397943,21.976732,25.557333,29.137934,26.597975,24.058014,21.518053,18.978092,16.438131,13.45037,10.462607,7.474845,4.4870825,1.49932,1.8129625,2.124792,2.4366217,2.7502642,3.0620937,4.0483456,5.032784,6.017223,7.0016613,7.987913,7.0052876,6.0226617,5.040036,4.0574102,3.0747845,3.4246864,3.774588,4.12449,4.4743915,4.8242936,4.590421,4.3547363,4.120864,3.8851788,3.6494937,3.5153344,3.3793623,3.245203,3.1092308,2.9750717,3.5515938,4.1299286,4.708264,5.2847857,5.863121,6.794984,7.7268467,8.660522,9.592385,10.524248,10.440851,10.355642,10.270433,10.185224,10.100015,11.588457,13.075087,14.561715,16.050158,17.536787,17.779724,18.022661,18.265598,18.506721,18.749659,15.754644,12.75963,9.764616,6.7696023,3.774588,3.0203958,2.2643902,1.5101979,0.7541924,0.0,0.0,0.0,0.0,0.0,0.0,0.17041849,0.34083697,0.5094425,0.67986095,0.85027945,5.5132194,10.174346,14.837286,19.500225,24.163166,22.749054,21.336756,19.92446,18.512161,17.099863,17.859495,18.619125,19.38057,20.140202,20.899832,19.090496,17.279346,15.47001,13.660673,11.849524,11.470614,11.089892,10.70917,10.330261,9.949538,9.380268,8.809185,8.239915,7.6706448,7.0995617,5.6800117,4.2604623,2.8390994,1.4195497,0.0,0.0,0.0,0.0,0.0,0.0,0.15591478,0.3100166,0.46411842,0.6200332,0.774135,0.62184614,0.46955732,0.31726846,0.16497959,0.012690738,0.014503701,0.018129626,0.01994259,0.02175555,0.025381476,0.04169814,0.059827764,0.07795739,0.09427405,0.11240368,0.11240368,0.11240368,0.11240368,0.11240368,0.11240368,0.12328146,0.13234627,0.14322405,0.15228885,0.16316663,0.19217403,0.2229944,0.2520018,0.28282216,0.31182957,0.291887,0.27194437,0.2520018,0.23205921,0.21211663,0.21755551,0.2229944,0.22662032,0.23205921,0.2374981,0.2755703,0.31182957,0.34990177,0.387974,0.42423326,0.83033687,1.2346275,1.6407311,2.0450218,2.4493124,1.9706904,1.4902552,1.0098201,0.5293851,0.05076295,0.18492219,0.3208944,0.4550536,0.58921283,0.72518504,0.7523795,0.7795739,0.80676836,0.83577573,0.8629702,0.7433147,0.62184614,0.50219065,0.3825351,0.26287958,0.24837588,0.23205921,0.21755551,0.2030518,0.18673515,1.8129625,3.437377,5.0617914,6.688019,8.312433,6.755099,5.197764,3.6404288,2.0830941,0.52575916,0.6200332,0.71430725,0.8103943,0.90466833,1.0007553,0.8375887,0.6744221,0.51306844,0.34990177,0.18673515,0.29007402,0.39159992,0.4949388,0.5982776,0.69980353,0.8122072,0.9246109,1.0370146,1.1494182,1.261822,2.3876717,3.5117085,4.6375585,5.763408,6.887445,5.8540564,4.8224807,3.7890918,2.7575161,1.7241274,2.808279,3.8906176,4.972956,6.055295,7.137634,5.7470913,4.358362,2.9678197,1.5772774,0.18673515,1.0043813,1.8220274,2.6396735,3.4573197,4.274966,3.4500678,2.6251698,1.8002719,0.97537386,0.15047589,0.4949388,0.83940166,1.1856775,1.5301404,1.8746033,2.0957847,2.3151531,2.5345216,2.7557032,2.9750717,2.3894846,1.8057107,1.2201238,0.6345369,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,1.0424535,2.084907,3.1273603,4.169814,5.2122674,5.6473784,6.0824895,6.5176005,6.9527116,7.3878226,7.344311,7.3026133,7.2591023,7.217404,7.175706,7.115878,7.0542374,6.9944096,6.9345818,6.874754,6.78048,6.684393,6.590119,6.495845,6.399758,6.1405044,5.8794374,5.620184,5.3591175,5.0998635,7.0052876,8.910711,10.8143215,12.719746,14.625169,13.457622,12.290073,11.122525,9.954978,8.78743,9.070251,9.353074,9.635896,9.916905,10.199727,10.1326475,10.065568,9.9966755,9.929596,9.862516,9.815379,9.768243,9.719293,9.672155,9.625018,10.110892,10.594954,11.080828,11.564888,12.050762,12.500377,12.949992,13.399607,13.849221,14.300649,15.781839,17.264843,18.747847,20.229036,21.71204,22.344765,22.977488,23.610212,24.242935,24.87566,23.327389,21.77912,20.232662,18.684393,17.137936,18.446894,19.757666,21.068438,22.377398,23.68817,23.816889,23.947422,24.077955,24.206676,24.33721,22.886839,21.43647,19.987913,18.537542,17.087172,15.680313,14.271642,12.864782,11.457924,10.049252,10.991992,11.934732,12.877473,13.820213,14.762955,15.62955,16.49796,17.364555,18.232965,19.099562,17.660069,16.220575,14.779271,13.339779,11.900287,10.845142,9.789998,8.734854,7.6797094,6.624565,6.2347784,5.844991,5.4552045,5.0654173,4.6756306,3.8597972,3.045777,2.229944,1.4159238,0.6000906,1.1222239,1.6443571,2.1683033,2.6904364,3.2125697,2.0631514,1.9779422,1.892733,1.8075237,1.7223145,1.6371052,1.4104849,1.1820517,0.9554313,0.726998,0.50037766,1.6008459,2.6995013,3.7999697,4.900438,6.000906,8.379513,10.7599325,13.140353,15.520773,17.89938,17.235836,16.570478,15.905121,15.239763,14.574407,11.922042,9.269678,6.6173134,3.9649491,1.3125849,1.4920682,1.6733645,1.8528478,2.032331,2.2118144,1.9253663,1.6371052,1.3506571,1.062396,0.774135,0.7850128,0.79589057,0.80495536,0.81583315,0.824898,1.5120108,2.1991236,2.8880494,3.5751622,4.262275,5.1905117,6.1169357,7.0451727,7.9734097,8.899834,8.809185,8.72035,8.629702,8.540867,8.450218,7.614443,6.78048,5.9447045,5.1107416,4.274966,4.8279195,5.3808727,5.9320135,6.484967,7.037921,8.3595705,9.683033,11.004683,12.328146,13.649796,12.665357,11.680918,10.694666,9.710228,8.725789,9.690285,10.654781,11.619277,12.585587,13.550082,15.2869005,17.025532,18.76235,20.499168,22.237799,20.845444,19.453089,18.060734,16.668379,15.27421,14.585284,13.894546,13.20562,12.514881,11.8241415,11.089892,10.355642,9.619579,8.885329,8.149267,7.4675927,6.7859187,6.1024323,5.4207582,4.7372713,4.76084,4.782595,4.804351,4.8279195,4.8496747,4.36924,3.8906176,3.4101827,2.9297476,2.4493124,3.1545548,3.8597972,4.5650396,5.2702823,5.975525,6.849373,7.7250338,8.600695,9.474543,10.3502035,8.497355,6.644508,4.7916603,2.9406252,1.0877775,1.1548572,1.2219368,1.2908293,1.357909,1.4249886,4.5233417,7.6198816,10.718235,13.8147745,16.913128,17.680012,18.446894,19.21559,19.982473,20.749357,21.010424,21.269676,21.530745,21.789997,22.049252,19.050611,16.050158,13.049705,10.049252,7.0506115,6.697084,6.345369,5.9918413,5.6401267,5.2865987,4.574105,3.8616104,3.149116,2.4366217,1.7241274,2.2081885,2.6904364,3.1726844,3.6549325,4.137181,5.047288,5.957395,6.867502,7.7776093,8.6877165,8.444779,8.201842,7.9607186,7.7177815,7.474845,7.2047133,6.9345818,6.6644506,6.394319,6.1241875,6.6553855,7.1847706,7.7141557,8.245354,8.774739,8.464723,8.154706,7.844689,7.5346723,7.224656,7.512917,7.799365,8.087626,8.375887,8.662335,9.229793,9.79725,10.364707,10.932164,11.499621,13.446743,15.3956785,17.3428,19.289923,21.237043,20.557182,19.877321,19.19746,18.5176,17.837738,15.555219,13.272699,10.990179,8.70766,6.4251394,7.5781837,8.729415,9.882459,11.035503,12.186734,10.810696,9.432844,8.054993,6.677141,5.2992897,4.7318325,4.164375,3.5969179,3.0294604,2.4620032,2.0178273,1.5718386,1.1276628,0.68167394,0.2374981,0.6055295,0.97174793,1.3397794,1.7078108,2.0758421,1.845596,1.6153497,1.3851035,1.1548572,0.9246109,0.99531645,1.064209,1.1349145,1.2056202,1.2745126,1.9525607,2.6306088,3.3068438,3.9848917,4.6629395,6.187641,7.7123427,9.237044,10.761745,12.28826,16.097294,19.908142,23.717176,27.528025,31.337059,28.6575,25.977942,23.29657,20.61701,17.937452,14.824595,11.711739,8.600695,5.487838,2.374981,2.4366217,2.5000753,2.561716,2.6251698,2.6868105,4.169814,5.6528172,7.135821,8.617011,10.100015,8.647832,7.1956487,5.7416525,4.2894692,2.8372865,3.3122826,3.787279,4.262275,4.7372713,5.2122674,4.954827,4.6973863,4.439945,4.1825047,3.925064,3.8924308,3.8597972,3.827164,3.7945306,3.7618973,4.305786,4.847862,5.389938,5.9320135,6.4759026,7.315304,8.154706,8.99592,9.835322,10.674724,10.355642,10.034748,9.715667,9.394773,9.07569,11.675479,14.275268,16.875055,19.474844,22.074633,20.471973,18.869314,17.266655,15.66581,14.06315,12.14685,10.232361,8.317872,6.401571,4.4870825,3.589666,2.6922495,1.794833,0.8974165,0.0,0.0,0.0,0.0,0.0,0.0,0.12690738,0.25562772,0.3825351,0.5094425,0.63816285,4.274966,7.911769,11.5503845,15.187187,18.825804,17.6365,16.450823,15.263332,14.075842,12.888351,13.657047,14.427556,15.198066,15.966762,16.73727,15.167245,13.597219,12.027194,10.457169,8.887142,8.740293,8.59163,8.444779,8.29793,8.149267,7.9607186,7.7703576,7.5799966,7.3896356,7.1992745,5.7597823,4.3202896,2.8807976,1.4394923,0.0,0.0,0.0,0.0,0.0,0.0,0.29732585,0.5946517,0.8919776,1.1893034,1.4866294,1.1947423,0.90285534,0.6091554,0.31726846,0.025381476,0.030820364,0.034446288,0.03988518,0.045324065,0.05076295,0.059827764,0.07070554,0.07977036,0.09064813,0.099712946,0.099712946,0.099712946,0.099712946,0.099712946,0.099712946,0.10696479,0.11421664,0.12328146,0.13053331,0.13778515,0.17223145,0.20667773,0.24293698,0.27738327,0.31182957,0.29732585,0.28282216,0.26831847,0.2520018,0.2374981,0.24837588,0.2574407,0.26831847,0.27738327,0.28826106,0.3245203,0.36259252,0.40066472,0.43692398,0.4749962,1.0098201,1.5446441,2.079468,2.6142921,3.149116,2.5272698,1.9054236,1.2817645,0.65991837,0.038072214,0.17041849,0.30276474,0.43511102,0.56745726,0.69980353,0.7306239,0.75963134,0.7904517,0.8194591,0.85027945,0.73424983,0.6200332,0.5058166,0.38978696,0.2755703,0.2574407,0.23931105,0.2229944,0.20486477,0.18673515,1.9253663,3.6621845,5.4008155,7.137634,8.874452,7.1847706,5.4950895,3.8054085,2.1157274,0.42423326,0.61459434,0.80495536,0.99531645,1.1856775,1.3742256,1.1367276,0.89922947,0.66173136,0.42423326,0.18673515,0.38072214,0.5728962,0.7650702,0.9572442,1.1494182,1.3633479,1.5754645,1.7875811,1.9996977,2.2118144,3.0258346,3.8380418,4.650249,5.462456,6.2746634,5.2847857,4.2949085,3.3050308,2.3151531,1.3252757,2.1392958,2.955129,3.7691493,4.5849824,5.4008155,4.3565493,3.3159087,2.2716422,1.2291887,0.18673515,0.922798,1.6570477,2.3931105,3.1273603,3.8616104,3.1128569,2.3622901,1.6117238,0.8629702,0.11240368,0.70342946,1.2926424,1.8818551,2.472881,3.0620937,2.902553,2.7430124,2.5816586,2.422118,2.2625773,1.8165885,1.3724127,0.92823684,0.48224804,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.8103943,1.6207886,2.42937,3.2397642,4.0501585,4.8333583,5.614745,6.397945,7.179332,7.9625316,7.752228,7.5419245,7.3316207,7.12313,6.9128265,7.017978,7.12313,7.228282,7.3316207,7.4367723,7.1466985,6.8566246,6.5683637,6.2782893,5.9882154,6.104245,6.2220874,6.33993,6.4577727,6.5756154,8.397643,10.21967,12.0416975,13.865538,15.687565,14.389484,13.093216,11.795135,10.497053,9.200785,9.465478,9.73017,9.994863,10.259555,10.524248,10.46442,10.4045925,10.344765,10.284937,10.225109,10.1054535,9.985798,9.864329,9.744674,9.625018,10.081885,10.540565,10.997431,11.454298,11.912977,12.661731,13.412297,14.162864,14.911617,15.662184,17.578485,19.492973,21.407463,23.32195,25.238253,26.003323,26.768393,27.53165,28.29672,29.06179,27.279648,25.497505,23.715364,21.933222,20.149265,21.082941,22.014805,22.946667,23.880342,24.812206,25.221935,25.631664,26.043207,26.452936,26.862667,25.124035,23.387217,21.650398,19.911768,18.17495,16.784407,15.3956785,14.005136,12.6145935,11.225864,11.535881,11.845898,12.154101,12.464118,12.774135,13.735004,14.695875,15.654932,16.615803,17.57486,16.40731,15.239763,14.072216,12.904668,11.73712,10.614896,9.492672,8.370448,7.2482243,6.1241875,5.857682,5.5893636,5.3228583,5.0545397,4.788034,3.9323158,3.0765975,2.222692,1.3669738,0.51306844,0.89560354,1.2781386,1.6606737,2.0432088,2.4257438,1.7495089,1.6733645,1.5954071,1.5174497,1.4394923,1.3633479,1.1657349,0.968122,0.7705091,0.5728962,0.37528324,1.5120108,2.6505513,3.787279,4.9258194,6.0625467,8.733041,11.401722,14.072216,16.74271,19.413204,18.66445,17.91751,17.170568,16.421816,15.674874,12.815832,9.954978,7.0941224,4.2350807,1.3742256,1.7205015,2.0649643,2.4094272,2.7557032,3.100166,2.5870976,2.0758421,1.5627737,1.0497054,0.53663695,0.5656443,0.59283876,0.6200332,0.64722764,0.6744221,1.4376793,2.1991236,2.962381,3.7256382,4.4870825,5.5966153,6.7079616,7.817495,8.927028,10.038374,9.864329,9.692098,9.519867,9.347635,9.175404,8.185526,7.1956487,6.205771,5.2140803,4.2242026,4.610364,4.994712,5.3808727,5.765221,6.149569,8.326937,10.504305,12.683486,14.860854,17.038223,15.760084,14.481945,13.20562,11.927481,10.649343,12.123281,13.595407,15.067532,16.539658,18.011784,20.024172,22.038374,24.050762,26.06315,28.075539,25.517448,22.959358,20.40308,17.84499,15.2869005,14.603414,13.918114,13.232814,12.547514,11.862214,11.184166,10.507931,9.829884,9.151835,8.4756,7.806617,7.1394467,6.472276,5.805106,5.137936,4.902251,4.668379,4.4326935,4.1970086,3.9631362,3.6295512,3.2977788,2.9641938,2.6324217,2.3006494,3.2705846,4.2405195,5.2104545,6.1803894,7.1503243,7.5999393,8.049554,8.499168,8.950596,9.400211,7.83925,6.2801023,4.7191415,3.159994,1.6008459,1.5446441,1.4902552,1.4358664,1.3796645,1.3252757,4.5269675,7.7304726,10.932164,14.13567,17.33736,16.844234,16.352922,15.859797,15.366671,14.875358,17.328297,19.77942,22.23236,24.685299,27.138237,22.85058,18.562923,14.275268,9.987611,5.6999545,5.315606,4.9294453,4.5450974,4.160749,3.774588,3.3757362,2.9750717,2.5744069,2.175555,1.7748904,2.2426348,2.7103791,3.1781235,3.6458678,4.1117992,5.3391747,6.5683637,7.795739,9.023115,10.25049,9.742861,9.235231,8.727602,8.219973,7.7123427,7.4458375,7.177519,6.9092,6.642695,6.3743763,7.119504,7.8646317,8.609759,9.354887,10.100015,9.646774,9.195346,8.7421055,8.290678,7.837437,8.049554,8.26167,8.4756,8.6877165,8.899834,9.570629,10.239613,10.910409,11.579392,12.250188,14.21544,16.18069,18.145943,20.10938,22.074633,20.580751,19.085056,17.589363,16.095482,14.599788,12.79589,10.990179,9.184468,7.380571,5.57486,6.784106,7.995165,9.2044115,10.41547,11.624716,10.315757,9.004985,7.6942134,6.3852544,5.0744824,4.74271,4.409125,4.077353,3.7455807,3.4119956,2.7955883,2.1773682,1.5591478,0.94274056,0.3245203,0.8448406,1.3651608,1.8854811,2.4058013,2.9243085,2.5055144,2.084907,1.6642996,1.2455053,0.824898,0.83033687,0.83577573,0.83940166,0.8448406,0.85027945,1.3977941,1.9453088,2.4928236,3.0403383,3.587853,5.5367875,7.4875355,9.438283,11.3872175,13.337966,17.377247,21.416527,25.45762,29.4969,33.537994,30.717026,27.89787,25.076899,22.257742,19.436771,16.200634,12.962683,9.724731,6.48678,3.2506418,3.0620937,2.8753586,2.6868105,2.5000753,2.3133402,4.2930956,6.2728505,8.252605,10.232361,12.212116,10.290376,8.366822,6.445082,4.5233417,2.5997884,3.199879,3.7999697,4.40006,5.0001507,5.600241,5.319232,5.040036,4.76084,4.4798307,4.2006345,4.269527,4.3402324,4.409125,4.4798307,4.550536,5.0581656,5.565795,6.073425,6.5792413,7.0868707,7.835624,8.582565,9.329506,10.078259,10.825199,10.270433,9.715667,9.159087,8.604321,8.049554,11.762501,15.475449,19.188396,22.89953,26.612478,23.164223,19.717781,16.269526,12.823084,9.374829,8.539054,7.705091,6.869315,6.035352,5.199577,4.160749,3.1201086,2.079468,1.0406405,0.0,0.0,0.0,0.0,0.0,0.0,0.08520924,0.17041849,0.25562772,0.34083697,0.42423326,3.0385253,5.6491914,8.26167,10.874149,13.486629,12.525759,11.563075,10.600392,9.637709,8.675026,9.4546,10.234174,11.015561,11.795135,12.574709,11.243994,9.915092,8.584378,7.2554765,5.924762,6.009971,6.09518,6.1803894,6.265599,6.350808,6.539356,6.7297173,6.9200783,7.1104393,7.3008003,5.8395524,4.3801174,2.9206827,1.4594349,0.0,0.0,0.0,0.0,0.0,0.0,0.4405499,0.8792868,1.3198367,1.7603867,2.1991236,1.7676386,1.3343405,0.90285534,0.46955732,0.038072214,0.045324065,0.052575916,0.059827764,0.06707962,0.07433146,0.07795739,0.07977036,0.08339628,0.08520924,0.0870222,0.0870222,0.0870222,0.0870222,0.0870222,0.0870222,0.092461094,0.09789998,0.10333887,0.10696479,0.11240368,0.15228885,0.19217403,0.23205921,0.27194437,0.31182957,0.30276474,0.291887,0.28282216,0.27194437,0.26287958,0.27738327,0.291887,0.30820364,0.32270733,0.33721104,0.37528324,0.41335547,0.44961473,0.48768693,0.52575916,1.1893034,1.8546607,2.520018,3.1853752,3.8507326,3.0856624,2.3205922,1.5555218,0.7904517,0.025381476,0.15410182,0.28463513,0.41516843,0.54570174,0.6744221,0.7070554,0.73968875,0.77232206,0.80495536,0.8375887,0.726998,0.61822027,0.5076295,0.39703882,0.28826106,0.26831847,0.24837588,0.22662032,0.20667773,0.18673515,2.03777,3.8869917,5.7380266,7.5872483,9.438283,7.614443,5.7924156,3.9703882,2.1483607,0.3245203,0.6091554,0.89560354,1.1802386,1.4648738,1.7495089,1.4376793,1.1258497,0.8122072,0.50037766,0.18673515,0.46955732,0.7523795,1.0352017,1.3180238,1.6008459,1.9126755,2.2245052,2.5381477,2.8499773,3.1618068,3.6621845,4.162562,4.6629395,5.163317,5.661882,4.7155156,3.7673361,2.819157,1.8727903,0.9246109,1.4721256,2.0196402,2.5671551,3.1146698,3.6621845,2.9678197,2.2716422,1.5772774,0.88291276,0.18673515,0.83940166,1.4920682,2.1447346,2.7974012,3.4500678,2.7756457,2.0994108,1.4249886,0.7505665,0.07433146,0.9101072,1.745883,2.5798457,3.4156215,4.249584,3.7093215,3.1708715,2.6306088,2.0903459,1.550083,1.2455053,0.93911463,0.6345369,0.32995918,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.57833505,1.1548572,1.7331922,2.3097143,2.8880494,4.017525,5.147001,6.2782893,7.407765,8.537241,8.160145,7.783048,7.404139,7.027043,6.6499467,6.9200783,7.1902094,7.460341,7.7304726,8.000604,7.51473,7.0306687,6.544795,6.060734,5.57486,6.069799,6.5647373,7.059676,7.554615,8.049554,9.789998,11.530442,13.270886,15.009518,16.749962,15.32316,13.894546,12.467744,11.040942,9.612328,9.860703,10.107266,10.355642,10.602205,10.850581,10.798005,10.745429,10.692853,10.640278,10.587702,10.395528,10.203354,10.009366,9.817192,9.625018,10.05469,10.484363,10.915848,11.34552,11.775192,12.824898,13.874602,14.924308,15.975826,17.025532,19.373318,21.719292,24.067078,26.414865,28.762651,29.660069,30.557484,31.4549,32.352318,33.249733,31.231907,29.214079,27.198065,25.180237,23.16241,23.717176,24.271942,24.82671,25.38329,25.938055,26.626982,27.31772,28.006645,28.697384,29.388123,27.363045,25.337965,23.312885,21.287807,19.262728,17.890314,16.517902,15.14549,13.773077,12.400664,12.077957,11.755249,11.432542,11.109835,10.7871275,11.840459,12.891977,13.945308,14.996826,16.050158,15.154554,14.260764,13.36516,12.469557,11.575767,10.384649,9.195346,8.00423,6.814926,5.6256227,5.480586,5.335549,5.1905117,5.045475,4.900438,4.004834,3.1092308,2.2154403,1.3198367,0.42423326,0.6671702,0.9101072,1.1530442,1.3941683,1.6371052,1.4376793,1.3669738,1.2980812,1.2273756,1.1566701,1.0877775,0.91917205,0.7523795,0.5855869,0.4169814,0.25018883,1.4249886,2.5997884,3.774588,4.949388,6.1241875,9.084756,12.045323,15.005891,17.964645,20.925215,20.094877,19.26454,18.434204,17.60568,16.775343,13.70781,10.640278,7.572745,4.505212,1.4376793,1.9471219,2.4583774,2.9678197,3.4772623,3.9867048,3.2506418,2.5127661,1.7748904,1.0370146,0.2991388,0.3444629,0.38978696,0.43511102,0.48043507,0.52575916,1.3633479,2.1991236,3.0367124,3.874301,4.7118897,6.004532,7.2971745,8.589817,9.882459,11.175101,10.919474,10.665659,10.410031,10.154404,9.900589,8.754796,7.610817,6.4650245,5.319232,4.175253,4.3928084,4.610364,4.8279195,5.045475,5.2630305,8.294304,11.327391,14.3604765,17.39175,20.424837,18.85481,17.284784,15.71476,14.144734,12.574709,14.554463,16.534218,18.515787,20.495543,22.475298,24.763256,27.049402,29.33736,31.625319,33.913277,30.189453,26.467442,22.745428,19.021603,15.299591,14.61973,13.939869,13.260008,12.580148,11.900287,11.280253,10.66022,10.040187,9.420154,8.80012,8.147454,7.494787,6.8421206,6.189454,5.5367875,5.045475,4.552349,4.059223,3.5679104,3.0747845,2.8898623,2.70494,2.520018,2.335096,2.1501737,3.3848011,4.6194286,5.8558693,7.0904965,8.325124,8.350506,8.375887,8.399456,8.424837,8.450218,7.1829576,5.915697,4.646623,3.3793623,2.1121013,1.9344311,1.7567607,1.5790904,1.403233,1.2255627,4.5324063,7.83925,11.147907,14.454751,17.761595,16.010273,14.257137,12.5058155,10.752681,8.999546,13.644357,18.289167,22.93579,27.580599,32.22541,26.65055,21.07569,15.499017,9.924157,4.349297,3.9323158,3.5153344,3.0983531,2.6795588,2.2625773,2.175555,2.08672,1.9996977,1.9126755,1.8256533,2.277081,2.7303216,3.1817493,3.63499,4.0882306,5.632875,7.177519,8.722163,10.266808,11.813264,11.039129,10.266808,9.494485,8.722163,7.949841,7.6851482,7.420456,7.155763,6.889258,6.624565,7.5854354,8.544493,9.5053625,10.46442,11.42529,10.830639,10.234174,9.639522,9.04487,8.450218,8.588004,8.725789,8.861761,8.999546,9.137331,9.909654,10.681975,11.454298,12.22662,13.000754,14.982323,16.965704,18.947271,20.930653,22.912222,20.602507,18.292793,15.983078,13.673364,11.361836,10.034748,8.70766,7.380571,6.051669,4.7245803,5.9918413,7.2591023,8.528176,9.795437,11.062697,9.820818,8.577126,7.3352466,6.093367,4.8496747,4.751775,4.655688,4.557788,4.459888,4.361988,3.5733492,2.7828975,1.9924458,1.2019942,0.41335547,1.0841516,1.7567607,2.42937,3.101979,3.774588,3.1654327,2.5544643,1.9453088,1.3343405,0.72518504,0.6653573,0.6055295,0.54570174,0.48587397,0.42423326,0.8430276,1.260009,1.6769904,2.0957847,2.5127661,4.8877473,7.262728,9.637709,12.012691,14.387671,18.657198,22.926725,27.198065,31.467592,35.737118,32.778362,29.817795,26.857227,23.89666,20.937904,17.57486,14.211814,10.850581,7.4875355,4.12449,3.6875658,3.2506418,2.811905,2.374981,1.938057,4.4145637,6.892884,9.3693905,11.847711,14.324218,11.9329195,9.539809,7.1466985,4.7554007,2.3622901,3.0874753,3.8126602,4.537845,5.2630305,5.9882154,5.6854506,5.382686,5.0799212,4.7771564,4.4743915,4.646623,4.8206677,4.992899,5.1651306,5.337362,5.810545,6.281915,6.755099,7.228282,7.699652,8.355945,9.010424,9.664904,10.319383,10.975676,10.185224,9.394773,8.604321,7.8156815,7.02523,11.849524,16.67563,21.499924,26.324217,31.150324,25.856472,20.564434,15.272397,9.980359,4.688321,4.933071,5.177821,5.422571,5.667321,5.9120708,4.7300196,3.5479677,2.3641033,1.1820517,0.0,0.0,0.0,0.0,0.0,0.0,0.04169814,0.08520924,0.12690738,0.17041849,0.21211663,1.8002719,3.386614,4.974769,6.5629244,8.149267,7.413204,6.6753283,5.9374523,5.199577,4.461701,5.2521524,6.0426044,6.833056,7.6216946,8.412147,7.322556,6.2329655,5.143375,4.0519714,2.962381,3.2796493,3.5969179,3.9141862,4.233268,4.550536,5.1198063,5.6908894,6.26016,6.82943,7.400513,5.919323,4.439945,2.960568,1.4793775,0.0,0.0,0.0,0.0,0.0,0.0,0.581961,1.1657349,1.7476959,2.3296568,2.911618,2.3405347,1.7676386,1.1947423,0.62184614,0.05076295,0.059827764,0.07070554,0.07977036,0.09064813,0.099712946,0.09427405,0.09064813,0.08520924,0.07977036,0.07433146,0.07433146,0.07433146,0.07433146,0.07433146,0.07433146,0.07795739,0.07977036,0.08339628,0.08520924,0.0870222,0.13234627,0.17767033,0.2229944,0.26831847,0.31182957,0.30820364,0.30276474,0.29732585,0.291887,0.28826106,0.30820364,0.32814622,0.3480888,0.3680314,0.387974,0.42423326,0.46230546,0.50037766,0.53663695,0.5747091,1.3705997,2.1646774,2.960568,3.7546456,4.550536,3.6422417,2.7357605,1.8274662,0.91917205,0.012690738,0.13959812,0.26831847,0.39522585,0.52213323,0.6508536,0.6852999,0.7197462,0.7541924,0.7904517,0.824898,0.7197462,0.61459434,0.5094425,0.40429065,0.2991388,0.27738327,0.25562772,0.23205921,0.21030366,0.18673515,2.1501737,4.1117992,6.0752378,8.036863,10.000301,8.044115,6.089741,4.135368,2.179181,0.22480737,0.6055295,0.98443866,1.3651608,1.745883,2.124792,1.7368182,1.3506571,0.96268314,0.5747091,0.18673515,0.56020546,0.9318628,1.305333,1.6769904,2.0504606,2.4620032,2.8753586,3.2869012,3.7002566,4.1117992,4.3003473,4.4870825,4.6756306,4.8623657,5.049101,4.1444325,3.2397642,2.335096,1.4304274,0.52575916,0.80495536,1.0841516,1.3651608,1.6443571,1.9253663,1.5772774,1.2291887,0.88291276,0.53482395,0.18673515,0.75781834,1.3270886,1.8981718,2.467442,3.0367124,2.4366217,1.8383441,1.2382535,0.63816285,0.038072214,1.1167849,2.1973107,3.2778363,4.358362,5.4370747,4.517903,3.5969179,2.6777458,1.7567607,0.8375887,0.6726091,0.5076295,0.34264994,0.17767033,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.3444629,0.69073874,1.0352017,1.3796645,1.7241274,3.2016919,4.6792564,6.156821,7.6343856,9.11195,8.568061,8.02236,7.476658,6.932769,6.3870673,6.8221784,7.2572894,7.6924005,8.127511,8.562622,7.8827615,7.2029004,6.5230393,5.8431783,5.163317,6.035352,6.9073873,7.7794223,8.653271,9.525306,11.182353,12.839401,14.498261,16.15531,17.812357,16.255022,14.697688,13.140353,11.583018,10.025683,10.254116,10.484363,10.714609,10.944855,11.175101,11.129777,11.084454,11.039129,10.995618,10.950294,10.685601,10.420909,10.154404,9.88971,9.625018,10.027496,10.429974,10.832452,11.234929,11.637406,12.988064,14.336908,15.687565,17.038223,18.387066,21.168152,23.947422,26.726694,29.507778,32.287052,33.316814,34.346577,35.37815,36.407913,37.437675,35.184166,32.932465,30.680765,28.427254,26.175554,26.353224,26.530895,26.70675,26.884422,27.062092,28.032028,29.001963,29.971897,30.941832,31.911768,29.60024,27.2869,24.975372,22.662033,20.350506,18.99441,17.640125,16.285843,14.929747,13.575464,12.620032,11.664601,10.70917,9.755551,8.80012,9.945912,11.089892,12.235684,13.379663,14.525456,13.901797,13.279951,12.658105,12.034446,11.4126,10.154404,8.898021,7.6398244,6.3834414,5.125245,5.101677,5.0799212,5.0581656,5.034597,5.0128417,4.077353,3.141864,2.2081885,1.2726997,0.33721104,0.4405499,0.5420758,0.64541465,0.7469406,0.85027945,1.1258497,1.062396,1.0007553,0.93730164,0.87566096,0.8122072,0.6744221,0.53663695,0.40066472,0.26287958,0.12509441,1.3379664,2.5508385,3.7618973,4.974769,6.187641,9.438283,12.687112,15.937754,19.188396,22.437225,21.525305,20.613384,19.699652,18.787731,17.87581,14.599788,11.325577,8.049554,4.7753434,1.49932,2.175555,2.8499773,3.5243993,4.2006345,4.8750563,3.9123733,2.94969,1.987007,1.0243238,0.06164073,0.12509441,0.18673515,0.25018883,0.31182957,0.37528324,1.2872034,2.1991236,3.1128569,4.024777,4.936697,6.412449,7.8882003,9.362139,10.837891,12.311829,11.974618,11.637406,11.300196,10.962985,10.625773,9.325879,8.024173,6.7242785,5.424384,4.12449,4.175253,4.2242026,4.274966,4.325729,4.3746786,8.26167,12.1504755,16.037468,19.92446,23.813263,21.949537,20.087626,18.225714,16.361988,14.500074,16.98746,19.474844,21.962229,24.449614,26.936998,29.500526,32.062244,34.62577,37.18749,39.749203,34.86327,29.975523,25.087776,20.20003,15.312282,14.63786,13.961625,13.287203,12.612781,11.938358,11.374527,10.812509,10.25049,9.686659,9.12464,8.488291,7.850128,7.211965,6.5756154,5.9374523,5.186886,4.4381323,3.6875658,2.9369993,2.1882458,2.1501737,2.1121013,2.0758421,2.03777,1.9996977,3.5008307,5.0001507,6.4994707,8.000604,9.499924,9.099259,8.700407,8.299743,7.900891,7.500226,6.5248523,5.5494785,4.574105,3.6005437,2.6251698,2.324218,2.0250793,1.7241274,1.4249886,1.1258497,4.537845,7.949841,11.361836,14.775645,18.187641,15.174497,12.163166,9.1500225,6.1368785,3.1255474,9.96223,16.798912,23.637405,30.4759,37.312584,30.45052,23.588457,16.72458,9.862516,3.000453,2.5508385,2.0994108,1.649796,1.2001812,0.7505665,0.97537386,1.2001812,1.4249886,1.649796,1.8746033,2.3133402,2.7502642,3.1871881,3.6241121,4.062849,5.924762,7.7866745,9.6504,11.512312,13.374225,12.337211,11.300196,10.263181,9.224354,8.187339,7.9244595,7.663393,7.400513,7.137634,6.874754,8.049554,9.224354,10.399154,11.575767,12.750566,12.012691,11.274815,10.536939,9.800876,9.063,9.12464,9.188094,9.249735,9.313189,9.374829,10.25049,11.124338,11.999999,12.87566,13.749508,15.749206,17.750717,19.750414,21.750113,23.74981,20.624262,17.500528,14.37498,11.249433,8.125698,7.2754188,6.4251394,5.57486,4.7245803,3.874301,5.199577,6.5248523,7.850128,9.175404,10.500679,9.325879,8.149267,6.9744673,5.7996674,4.6248674,4.762653,4.900438,5.038223,5.1741953,5.3119802,4.349297,3.388427,2.4257438,1.4630609,0.50037766,1.3252757,2.1501737,2.9750717,3.7999697,4.6248674,3.825351,3.0258346,2.2245052,1.4249886,0.62547207,0.50037766,0.37528324,0.25018883,0.12509441,0.0,0.28826106,0.5747091,0.8629702,1.1494182,1.4376793,4.2368937,7.037921,9.837135,12.638163,15.437376,19.93715,24.436922,28.938509,33.438282,37.938053,34.83789,31.737722,28.637556,25.537392,22.437225,18.950897,15.462758,11.974618,8.488291,5.0001507,4.313038,3.625925,2.9369993,2.2498865,1.5627737,4.537845,7.512917,10.487988,13.46306,16.438131,13.575464,10.712796,7.850128,4.98746,2.124792,2.9750717,3.825351,4.6756306,5.52591,6.3743763,6.049856,5.7253356,5.4008155,5.0744824,4.749962,5.0255322,5.2992897,5.57486,5.8504305,6.1241875,6.5629244,6.9998484,7.4367723,7.8755093,8.312433,8.874452,9.438283,10.000301,10.56232,11.124338,10.100015,9.07569,8.049554,7.02523,6.000906,11.938358,17.873999,23.813263,29.750715,35.688168,28.548721,21.4129,14.275268,7.137634,0.0,1.3252757,2.6505513,3.975827,5.2992897,6.624565,5.2992897,3.975827,2.6505513,1.3252757,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.5620184,1.1258497,1.6878681,2.2498865,2.811905,2.3006494,1.7875811,1.2745126,0.76325727,0.25018883,1.0497054,1.8492218,2.6505513,3.4500678,4.249584,3.3993049,2.5508385,1.7005589,0.85027945,0.0,0.5493277,1.1004683,1.649796,2.1991236,2.7502642,3.7002566,4.650249,5.600241,6.550234,7.500226,5.999093,4.499773,3.000453,1.49932,0.0,0.0,0.0,0.0,0.0,0.0,0.72518504,1.4503701,2.175555,2.9007401,3.6241121,2.911618,2.1991236,1.4866294,0.774135,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.11240368,0.16316663,0.21211663,0.26287958,0.31182957,0.31182957,0.31182957,0.31182957,0.31182957,0.31182957,0.33721104,0.36259252,0.387974,0.41335547,0.43692398,0.4749962,0.51306844,0.5493277,0.5873999,0.62547207,1.550083,2.474694,3.3993049,4.325729,5.2503395,4.2006345,3.150929,2.0994108,1.0497054,0.0,0.12509441,0.25018883,0.37528324,0.50037766,0.62547207,0.66173136,0.69980353,0.73787576,0.774135,0.8122072,0.7124943,0.61278135,0.51306844,0.41335547,0.31182957,0.28826106,0.26287958,0.2374981,0.21211663,0.18673515,2.2625773,4.3366065,6.412449,8.488291,10.56232,8.4756,6.3870673,4.3003473,2.2118144,0.12509441,0.6000906,1.0750868,1.550083,2.0250793,2.5000753,2.03777,1.5754645,1.1131591,0.6508536,0.18673515,0.6508536,1.1131591,1.5754645,2.03777,2.5000753,3.0131438,3.5243993,4.0374675,4.550536,5.0617914,4.936697,4.8116026,4.688321,4.5632267,4.4381323,3.5751622,2.712192,1.8492218,0.9880646,0.12509441,0.13778515,0.15047589,0.16316663,0.17585737,0.18673515,0.18673515,0.18673515,0.18673515,0.18673515,0.18673515,0.6744221,1.162109,1.649796,2.137483,2.6251698,2.0994108,1.5754645,1.0497054,0.52575916,0.0,1.3252757,2.6505513,3.975827,5.2992897,6.624565,5.3246713,4.024777,2.7248828,1.4249886,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.11240368,0.22480737,0.33721104,0.44961473,0.5620184,2.3876717,4.213325,6.037165,7.8628187,9.686659,8.974165,8.26167,7.549176,6.836682,6.1241875,6.7242785,7.324369,7.9244595,8.52455,9.12464,8.2507925,7.3751316,6.4994707,5.6256227,4.749962,6.000906,7.250037,8.499168,9.750113,10.999244,12.574709,14.150173,15.725637,17.29929,18.874754,17.186886,15.50083,13.812962,12.125093,10.437225,10.649343,10.863272,11.075388,11.287505,11.499621,11.463363,11.42529,11.3872175,11.349146,11.312886,10.975676,10.636651,10.29944,9.96223,9.625018,10.000301,10.375585,10.750868,11.124338,11.499621,13.149418,14.799213,16.450823,18.100618,19.750414,22.962984,26.175554,29.388123,32.600693,35.813263,36.975372,38.13748,39.29959,40.4617,41.62562,39.138237,36.64904,34.161655,31.674269,29.186884,28.98746,28.788033,28.586794,28.387367,28.187943,29.437073,30.688017,31.93715,33.18809,34.437225,31.837437,29.237648,26.63786,24.03807,21.438282,20.100317,18.76235,17.424383,16.08823,14.750263,13.162108,11.573953,9.987611,8.399456,6.813113,8.049554,9.287807,10.524248,11.762501,13.000754,12.650853,12.299138,11.949236,11.599335,11.249433,9.924157,8.600695,7.2754188,5.9501433,4.6248674,4.7245803,4.8242936,4.9258194,5.0255322,5.125245,4.1498713,3.1744974,2.1991236,1.2255627,0.25018883,0.21211663,0.17585737,0.13778515,0.099712946,0.06164073,1.0007553,0.93911463,0.8792868,0.8194591,0.75963134,0.69980353,0.58921283,0.48043507,0.36984438,0.25925365,0.15047589,1.1421664,2.13567,3.1273603,4.120864,5.1125546,7.844689,10.576823,13.310771,16.042906,18.77504,18.590118,18.405195,18.220274,18.035353,17.85043,14.849977,11.849524,8.849071,5.8504305,2.8499773,3.0620937,3.2742105,3.48814,3.7002566,3.9123733,3.442816,2.9732587,2.5018883,2.032331,1.5627737,2.3079014,3.053029,3.7981565,4.5432844,5.2884116,5.3482394,5.408067,5.467895,5.527723,5.5875506,6.8983226,8.207282,9.518054,10.827013,12.137785,12.179482,12.222994,12.264692,12.308203,12.349901,11.512312,10.674724,9.837135,8.999546,8.161958,8.406708,8.653271,8.898021,9.142771,9.38752,11.952863,14.518205,17.081734,19.647076,22.212418,20.865387,19.518354,18.169512,16.82248,15.475449,17.857681,20.239914,22.622147,25.00438,27.386612,29.415318,31.44221,33.470917,35.497807,37.5247,33.530743,29.534973,25.539204,21.545248,17.549479,16.195194,14.840912,13.484816,12.130532,10.774437,10.504305,10.234174,9.965856,9.695724,9.425592,9.102885,8.780178,8.457471,8.134763,7.8120556,6.6753283,5.5367875,4.40006,3.2633326,2.124792,2.6378605,3.149116,3.6621845,4.175253,4.688321,5.620184,6.552047,7.4857225,8.417585,9.349448,8.725789,8.100317,7.474845,6.849373,6.2257137,5.520471,4.8152285,4.1099863,3.4047437,2.6995013,2.42937,2.1592383,1.889107,1.6207886,1.3506571,5.4443264,9.539809,13.635292,17.730774,21.824444,18.635443,15.444629,12.255627,9.064813,5.8758116,11.631968,17.389936,23.147905,28.905876,34.662033,28.894999,23.127964,17.359118,11.592083,5.825049,5.0726695,4.3202896,3.5679104,2.8155308,2.0631514,1.9978848,1.9326181,1.8673514,1.8020848,1.7368182,2.0595255,2.382233,2.70494,3.0276475,3.350355,4.8297324,6.3091097,7.7903004,9.269678,10.750868,9.929596,9.110137,8.290678,7.4694057,6.6499467,6.4795284,6.3091097,6.1405044,5.9700856,5.7996674,7.12313,8.444779,9.768243,11.089892,12.413355,11.958302,11.503247,11.048194,10.593141,10.138086,10.2378,10.337513,10.437225,10.536939,10.636651,11.459737,12.282822,13.1059065,13.927178,14.750263,16.322102,17.895754,19.467592,21.03943,22.613083,19.61988,16.628492,13.635292,10.642091,7.650702,7.115878,6.5792413,6.0444174,5.5095935,4.974769,6.009971,7.0451727,8.080374,9.115576,10.150778,9.142771,8.134763,7.1267557,6.1205616,5.1125546,5.473334,5.8323007,6.19308,6.552047,6.9128265,5.955582,4.9983377,4.0392804,3.0820365,2.124792,2.764768,3.4047437,4.0447197,4.6846952,5.3246713,4.365614,3.4047437,2.4456866,1.4848163,0.52575916,0.6671702,0.8103943,0.95180535,1.0950294,1.2382535,1.6824293,2.126605,2.572594,3.0167696,3.4627585,5.667321,7.8718834,10.078259,12.282822,14.487384,18.164072,21.842573,25.51926,29.197762,32.87445,30.688017,28.499771,26.311525,24.125093,21.936848,19.150324,16.361988,13.575464,10.7871275,8.000604,6.7623506,5.52591,4.2876563,3.049403,1.8129625,4.274966,6.736969,9.200785,11.662788,14.124791,11.795135,9.465478,7.135821,4.804351,2.474694,3.5352771,4.59586,5.65463,6.7152133,7.7757964,7.231908,6.6898317,6.147756,5.6056805,5.0617914,5.2865987,5.5132194,5.7380266,5.962834,6.187641,6.622752,7.057863,7.4929743,7.9280853,8.363196,9.115576,9.867955,10.620335,11.372714,12.125093,11.289318,10.455356,9.619579,8.785617,7.949841,12.097899,16.244144,20.392202,24.540262,28.68832,23.182352,17.678198,12.172231,6.6680765,1.162109,2.0758421,2.9877625,3.8996825,4.8134155,5.7253356,4.5795436,3.435564,2.2897718,1.1457924,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.15954071,0.20667773,0.25562772,0.30276474,0.34990177,0.73787576,1.1258497,1.5120108,1.8999848,2.2879589,1.8691645,1.452183,1.0352017,0.61822027,0.19942589,0.83940166,1.4793775,2.1193533,2.759329,3.3993049,2.7393866,2.079468,1.4195497,0.75963134,0.099712946,0.52032024,0.93911463,1.3597219,1.7803292,2.1991236,3.045777,3.8906176,4.7354584,5.580299,6.4251394,5.145188,3.8652363,2.5852847,1.305333,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.61278135,1.2255627,1.8383441,2.4493124,3.0620937,2.469255,1.8782293,1.2853905,0.69255173,0.099712946,0.10515183,0.11059072,0.11421664,0.11965553,0.12509441,0.26287958,0.40066472,0.53663695,0.6744221,0.8122072,0.75781834,0.7016165,0.64722764,0.59283876,0.53663695,0.44780177,0.35715362,0.26831847,0.17767033,0.0870222,0.12328146,0.15772775,0.19217403,0.22662032,0.26287958,0.2755703,0.28826106,0.2991388,0.31182957,0.3245203,0.3680314,0.40972954,0.45324063,0.4949388,0.53663695,0.5493277,0.5620184,0.5747091,0.5873999,0.6000906,1.5772774,2.5544643,3.531651,4.510651,5.487838,4.3982472,3.3068438,2.2172532,1.1276628,0.038072214,0.13959812,0.24293698,0.3444629,0.44780177,0.5493277,0.6055295,0.65991837,0.71430725,0.7705091,0.824898,0.7324369,0.6399758,0.5475147,0.4550536,0.36259252,0.32814622,0.291887,0.2574407,0.2229944,0.18673515,1.8909199,3.5932918,5.295664,6.9980354,8.700407,7.0016613,5.3047285,3.6077955,1.9108626,0.21211663,0.6852999,1.1566701,1.6298534,2.1030366,2.5744069,2.1229792,1.6697385,1.2183108,0.7650702,0.31182957,0.6544795,0.99712944,1.3397794,1.6824293,2.0250793,2.4583774,2.8898623,3.3231604,3.7546456,4.1879435,4.1281157,4.068288,4.006647,3.9468195,3.8869917,3.1346123,2.382233,1.6298534,0.8774739,0.12509441,0.13234627,0.13959812,0.14684997,0.15410182,0.16316663,0.17585737,0.18673515,0.19942589,0.21211663,0.22480737,0.65810543,1.0895905,1.5228885,1.9543737,2.3876717,1.9126755,1.4376793,0.96268314,0.48768693,0.012690738,1.1367276,2.2625773,3.388427,4.512464,5.638314,4.5305934,3.4228733,2.3151531,1.2074331,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.21574254,0.40429065,0.5946517,0.7850128,0.97537386,2.6034143,4.229642,5.857682,7.4857225,9.11195,8.72035,8.326937,7.935337,7.5419245,7.1503243,7.4694057,7.7903004,8.109382,8.430276,8.749357,7.842876,6.9345818,6.0281005,5.1198063,4.213325,5.411693,6.6118746,7.8120556,9.012237,10.212419,11.564888,12.917358,14.269829,15.622298,16.97477,15.700256,14.425743,13.149418,11.874905,10.600392,11.057259,11.514126,11.972805,12.429671,12.888351,12.9427395,12.9971285,13.05333,13.107719,13.162108,12.621845,12.083396,11.543133,11.00287,10.462607,10.491614,10.522435,10.553255,10.582263,10.613083,12.083396,13.551895,15.022208,16.492521,17.962833,21.13008,24.297325,27.464571,30.631815,33.800873,34.952106,36.10515,37.258194,38.409424,39.56247,36.884724,34.206978,31.529232,28.8533,26.175554,26.139294,26.104849,26.070402,26.034143,25.999697,27.252453,28.50521,29.757967,31.010725,32.26167,29.785162,27.306843,24.830336,22.352016,19.87551,18.5176,17.15969,15.801782,14.445685,13.087777,11.6881695,10.28675,8.887142,7.4875355,6.0879283,7.0451727,8.002417,8.9596615,9.916905,10.874149,10.863272,10.850581,10.837891,10.825199,10.812509,9.570629,8.326937,7.0850577,5.8431783,4.599486,4.5324063,4.465327,4.3982472,4.329355,4.262275,3.4555066,2.6469254,1.840157,1.0333886,0.22480737,0.19761293,0.17041849,0.14322405,0.11421664,0.0870222,0.87566096,0.81764615,0.75963134,0.7016165,0.64541465,0.5873999,0.5058166,0.4224203,0.34083697,0.2574407,0.17585737,0.9481794,1.7205015,2.4928236,3.2651455,4.0374675,6.2529078,8.466536,10.681975,12.897416,15.112856,15.654932,16.197008,16.740896,17.282972,17.825048,15.100165,12.375282,9.6504,6.925517,4.2006345,3.9504454,3.7002566,3.4500678,3.199879,2.94969,2.9732587,2.9950142,3.0167696,3.0403383,3.0620937,4.4907084,5.91751,7.344311,8.772926,10.199727,9.407463,8.615198,7.8229337,7.0306687,6.2384043,7.382384,8.528176,9.672155,10.817947,11.961927,12.384347,12.806767,13.229188,13.653421,14.075842,13.700559,13.325275,12.949992,12.574709,12.199425,12.639976,13.080525,13.519262,13.959812,14.400362,15.6422415,16.88412,18.127813,19.369692,20.613384,19.77942,18.947271,18.115122,17.282972,16.450823,18.727903,21.004984,23.282066,25.559147,27.838041,29.330109,30.822176,32.314243,33.808125,35.300194,32.198215,29.094423,25.992445,22.890465,19.786674,17.75253,15.718386,13.682428,11.648285,9.612328,9.635896,9.657652,9.679407,9.702975,9.724731,9.71748,9.710228,9.702975,9.695724,9.686659,8.161958,6.637256,5.1125546,3.587853,2.0631514,3.1255474,4.1879435,5.2503395,6.3127356,7.3751316,7.7395372,8.105756,8.470161,8.834567,9.200785,8.350506,7.500226,6.6499467,5.7996674,4.949388,4.514277,4.079166,3.6458678,3.2107568,2.7756457,2.5345216,2.2952106,2.0558996,1.8147756,1.5754645,6.352621,11.129777,15.906934,20.685904,25.46306,22.094576,18.727903,15.359419,11.992747,8.624263,13.301706,17.97915,22.658407,27.33585,32.013294,27.339476,22.66747,17.995466,13.321649,8.649645,7.5945,6.539356,5.484212,4.4308805,3.3757362,3.0203958,2.665055,2.3097143,1.9543737,1.6008459,1.8075237,2.0142014,2.222692,2.42937,2.6378605,3.7347028,4.8333583,5.9302006,7.027043,8.125698,7.5219817,6.9200783,6.3181744,5.714458,5.1125546,5.034597,4.95664,4.880495,4.802538,4.7245803,6.1948934,7.665206,9.135518,10.605831,12.07433,11.9021,11.729868,11.557636,11.385405,11.213174,11.349146,11.486931,11.624716,11.762501,11.900287,12.670795,13.439491,14.210001,14.98051,15.749206,16.894999,18.04079,19.18477,20.330563,21.474543,18.6155,15.754644,12.895603,10.034748,7.175706,6.9545245,6.735156,6.5157876,6.294606,6.0752378,6.8203654,7.5654926,8.31062,9.055748,9.800876,8.9596615,8.120259,7.2808576,6.439643,5.600241,6.1822023,6.7641635,7.3479376,7.9298983,8.511859,7.560054,6.6082487,5.65463,4.702825,3.7492065,4.2042603,4.6593137,5.1143675,5.569421,6.0244746,4.9058766,3.785466,2.665055,1.5446441,0.42423326,0.83577573,1.2455053,1.6552348,2.0649643,2.474694,3.0765975,3.680314,4.2822175,4.8841214,5.487838,7.0977483,8.70766,10.31757,11.927481,13.537392,16.392807,19.248224,22.101828,24.957243,27.812658,26.538147,25.26182,23.987309,22.712795,21.438282,19.34975,17.26303,15.174497,13.087777,10.999244,9.211663,7.4258947,5.638314,3.8507326,2.0631514,4.0120864,5.962834,7.911769,9.862516,11.813264,10.014805,8.21816,6.4197006,4.6230545,2.8245957,4.0954823,5.3645563,6.635443,7.9045167,9.175404,8.415772,7.654328,6.8946967,6.1350656,5.375434,5.5494785,5.7253356,5.89938,6.0752378,6.249282,6.68258,7.115878,7.5473633,7.9806614,8.412147,9.354887,10.297627,11.240368,12.183108,13.125849,12.480434,11.83502,11.189605,10.54419,9.900589,12.25744,14.614291,16.972956,19.329807,21.686659,17.81417,13.943495,10.069194,6.1967063,2.324218,2.8245957,3.3249733,3.825351,4.325729,4.8242936,3.8597972,2.8953013,1.9308052,0.9644961,0.0,0.045324065,0.09064813,0.13415924,0.1794833,0.22480737,0.3208944,0.41516843,0.5094425,0.6055295,0.69980353,0.9119202,1.1258497,1.3379664,1.550083,1.7621996,1.4394923,1.1167849,0.79589057,0.47318324,0.15047589,0.630911,1.1095331,1.5899682,2.0704033,2.5508385,2.079468,1.6099107,1.1403534,0.67079616,0.19942589,0.4894999,0.7795739,1.0696479,1.3597219,1.649796,2.3894846,3.1291735,3.870675,4.610364,5.3500524,4.2894692,3.2306993,2.1701162,1.1095331,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.50037766,1.0007553,1.49932,1.9996977,2.5000753,2.0268922,1.5555218,1.0823387,0.6091554,0.13778515,0.13415924,0.13234627,0.13053331,0.12690738,0.12509441,0.41335547,0.69980353,0.9880646,1.2745126,1.5627737,1.452183,1.3434052,1.2328146,1.1222239,1.0116332,0.8321498,0.6526665,0.47318324,0.291887,0.11240368,0.13234627,0.15228885,0.17223145,0.19217403,0.21211663,0.2374981,0.26287958,0.28826106,0.31182957,0.33721104,0.39703882,0.45686656,0.5166943,0.57833505,0.63816285,0.62547207,0.61278135,0.6000906,0.5873999,0.5747091,1.6044719,2.6342347,3.6658103,4.695573,5.7253356,4.594047,3.4645715,2.335096,1.2056202,0.07433146,0.15410182,0.23568514,0.3154555,0.39522585,0.4749962,0.5475147,0.6200332,0.69255173,0.7650702,0.8375887,0.7523795,0.6671702,0.581961,0.49675176,0.41335547,0.3680314,0.32270733,0.27738327,0.23205921,0.18673515,1.5174497,2.8481643,4.177066,5.5077806,6.836682,5.529536,4.2223897,2.9152439,1.6080978,0.2991388,0.7705091,1.2400664,1.7096237,2.179181,2.6505513,2.2081885,1.7658255,1.3216497,0.8792868,0.43692398,0.65991837,0.88291276,1.1059072,1.3270886,1.550083,1.9017978,2.2553256,2.6070402,2.960568,3.3122826,3.3177216,3.3231604,3.3267863,3.3322253,3.3376641,2.6940625,2.0522738,1.4104849,0.7668832,0.12509441,0.12690738,0.13053331,0.13234627,0.13415924,0.13778515,0.16316663,0.18673515,0.21211663,0.2374981,0.26287958,0.6399758,1.017072,1.3941683,1.7730774,2.1501737,1.7241274,1.2998942,0.87566096,0.44961473,0.025381476,0.9499924,1.8746033,2.7992141,3.7256382,4.650249,3.7347028,2.819157,1.9054236,0.9898776,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.31726846,0.5855869,0.8520924,1.1204109,1.3869164,2.817344,4.2477713,5.678199,7.1068134,8.537241,8.464723,8.392203,8.319685,8.247167,8.174648,8.214534,8.254418,8.294304,8.334189,8.375887,7.4349594,6.495845,5.5549173,4.615803,3.6748753,4.8242936,5.975525,7.124943,8.274362,9.425592,10.555068,11.684544,12.815832,13.945308,15.074784,14.211814,13.3506565,12.487686,11.624716,10.761745,11.465176,12.166792,12.870221,13.571837,14.275268,14.422117,14.57078,14.71763,14.86448,15.013144,14.269829,13.528327,12.785012,12.0416975,11.300196,10.98474,10.669285,10.355642,10.040187,9.724731,11.015561,12.304577,13.595407,14.884423,16.175253,19.297174,22.419096,25.54283,28.664751,31.786673,32.930653,34.07282,35.214985,36.35715,37.499317,34.633022,31.764917,28.89681,26.030518,23.16241,23.292944,23.421663,23.552197,23.68273,23.813263,25.067833,26.322403,27.576973,28.831545,30.087927,27.73289,25.37785,23.022812,20.667774,18.312735,16.934883,15.557032,14.17918,12.803142,11.42529,10.212419,8.999546,7.7866745,6.5756154,5.3627434,6.0407915,6.717026,7.3950744,8.073122,8.749357,9.07569,9.400211,9.724731,10.049252,10.375585,9.215289,8.054993,6.8946967,5.7344007,4.574105,4.3402324,4.1045475,3.870675,3.63499,3.3993049,2.759329,2.1193533,1.4793775,0.83940166,0.19942589,0.18310922,0.16497959,0.14684997,0.13053331,0.11240368,0.7505665,0.69436467,0.6399758,0.5855869,0.5293851,0.4749962,0.42060733,0.36440548,0.3100166,0.25562772,0.19942589,0.7523795,1.305333,1.8582866,2.4094272,2.962381,4.6593137,6.35806,8.054993,9.751925,11.450671,12.719746,13.990632,15.2597065,16.530592,17.799667,15.350354,12.899229,10.449916,8.000604,5.5494785,4.836984,4.12449,3.4119956,2.6995013,1.987007,2.5018883,3.0167696,3.531651,4.0483456,4.5632267,6.6717024,8.781991,10.89228,13.002567,15.112856,13.466686,11.822329,10.177972,8.531802,6.887445,7.8682575,8.847258,9.82807,10.80707,11.787883,12.589212,13.392355,14.195497,14.996826,15.799969,15.8869915,15.975826,16.062849,16.14987,16.236893,16.873243,17.50778,18.142317,18.776854,19.413204,19.333433,19.25185,19.17208,19.092308,19.012539,18.69527,18.378002,18.060734,17.741652,17.424383,19.598125,21.770054,23.941984,26.115726,28.287655,29.2449,30.202143,31.159388,32.11663,33.07569,30.865688,28.655687,26.445684,24.235683,22.025682,19.309864,16.59586,13.880041,11.164224,8.450218,8.765674,9.079316,9.394773,9.710228,10.025683,10.332074,10.640278,10.946668,11.254871,11.563075,9.6504,7.7377243,5.825049,3.9123733,1.9996977,3.6132345,5.224958,6.836682,8.450218,10.061942,9.860703,9.657652,9.4546,9.253361,9.050309,7.9752226,6.9001355,5.825049,4.749962,3.6748753,3.5098956,3.3449159,3.1799364,3.0149567,2.8499773,2.6396735,2.42937,2.220879,2.0105755,1.8002719,7.2591023,12.719746,18.18039,23.63922,29.099863,25.555521,22.009365,18.465023,14.920682,11.374527,14.973258,18.570175,22.167093,25.765823,29.362741,25.785767,22.206978,18.630003,15.053028,11.47424,10.118144,8.760235,7.402326,6.0444174,4.688321,4.0429068,3.397492,2.752077,2.1066625,1.4630609,1.5555218,1.647983,1.7404441,1.8329052,1.9253663,2.6396735,3.3557937,4.070101,4.784408,5.5005283,5.1143675,4.7300196,4.345671,3.9595103,3.5751622,3.589666,3.6041696,3.6204863,3.63499,3.6494937,5.2666564,6.885632,8.502794,10.119957,11.73712,11.847711,11.958302,12.067079,12.17767,12.28826,12.462305,12.638163,12.812206,12.988064,13.162108,13.880041,14.597975,15.3159075,16.032028,16.749962,17.467894,18.185827,18.901947,19.61988,20.337814,17.609306,14.882609,12.154101,9.427405,6.70071,6.794984,6.889258,6.985345,7.079619,7.175706,7.6307597,8.0858135,8.540867,8.994107,9.449161,8.778365,8.105756,7.4331465,6.7605376,6.0879283,6.892884,7.6978393,8.502794,9.30775,10.112705,9.164526,8.21816,7.26998,6.3218007,5.375434,5.6455655,5.915697,6.185828,6.454147,6.7242785,5.4443264,4.164375,2.8844235,1.6044719,0.3245203,1.0025684,1.6806163,2.3568513,3.0348995,3.7129474,4.4725785,5.23221,5.9918413,6.7532854,7.512917,8.528176,9.541622,10.556881,11.57214,12.5873995,14.61973,16.652061,18.684393,20.716722,22.749054,22.388275,22.025682,21.66309,21.300497,20.937904,19.549175,18.16226,16.775343,15.386614,13.999697,11.662788,9.325879,6.987158,4.650249,2.3133402,3.7492065,5.186886,6.624565,8.062244,9.499924,8.234476,6.970841,5.7053933,4.439945,3.1744974,4.655688,6.1350656,7.614443,9.0956335,10.57501,9.597824,8.620637,7.6416373,6.6644506,5.6872635,5.812358,5.9374523,6.0625467,6.187641,6.3127356,6.742408,7.17208,7.6017523,8.033237,8.46291,9.594198,10.7273,11.860401,12.99169,14.124791,13.669738,13.2146845,12.75963,12.304577,11.849524,12.416981,12.984438,13.551895,14.119352,14.68681,12.447801,10.20698,7.9679704,5.727149,3.48814,3.5751622,3.6621845,3.7492065,3.8380418,3.925064,3.1400511,2.3550384,1.5700256,0.7850128,0.0,0.06707962,0.13415924,0.2030518,0.27013144,0.33721104,0.48043507,0.62184614,0.7650702,0.90829426,1.0497054,1.0877775,1.1258497,1.162109,1.2001812,1.2382535,1.0098201,0.78319985,0.55476654,0.32814622,0.099712946,0.42060733,0.73968875,1.0605831,1.3796645,1.7005589,1.4195497,1.1403534,0.85934424,0.58014804,0.2991388,0.4604925,0.6200332,0.7795739,0.93911463,1.1004683,1.7350051,2.3695421,3.005892,3.6404288,4.274966,3.435564,2.5943494,1.7549478,0.9155461,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.387974,0.774135,1.162109,1.550083,1.938057,1.5845293,1.2328146,0.8792868,0.5275721,0.17585737,0.16497959,0.15410182,0.14503701,0.13415924,0.12509441,0.5620184,1.0007553,1.4376793,1.8746033,2.3133402,2.1483607,1.983381,1.8184015,1.651609,1.4866294,1.2183108,0.9481794,0.678048,0.40791658,0.13778515,0.14322405,0.14684997,0.15228885,0.15772775,0.16316663,0.19942589,0.2374981,0.2755703,0.31182957,0.34990177,0.42785916,0.5058166,0.581961,0.65991837,0.73787576,0.69980353,0.66173136,0.62547207,0.5873999,0.5493277,1.6316663,2.715818,3.7981565,4.880495,5.962834,4.7916603,3.6222992,2.4529383,1.2817645,0.11240368,0.17041849,0.22662032,0.28463513,0.34264994,0.40066472,0.4894999,0.58014804,0.67079616,0.75963134,0.85027945,0.77232206,0.69436467,0.61822027,0.5402629,0.46230546,0.40791658,0.35171473,0.29732585,0.24293698,0.18673515,1.1457924,2.1030366,3.0602808,4.017525,4.974769,4.0574102,3.1400511,2.222692,1.305333,0.387974,0.8557183,1.3216497,1.789394,2.2571385,2.7248828,2.2915847,1.8600996,1.4268016,0.99531645,0.5620184,0.6653573,0.7668832,0.87022203,0.97174793,1.0750868,1.3470312,1.6207886,1.892733,2.1646774,2.4366217,2.5073273,2.5780327,2.6469254,2.7176309,2.7883365,2.2553256,1.7223145,1.1893034,0.65810543,0.12509441,0.12328146,0.11965553,0.11784257,0.11421664,0.11240368,0.15047589,0.18673515,0.22480737,0.26287958,0.2991388,0.62184614,0.9445535,1.2672608,1.5899682,1.9126755,1.5373923,1.162109,0.7868258,0.41335547,0.038072214,0.76325727,1.4866294,2.2118144,2.9369993,3.6621845,2.9406252,2.2172532,1.4956942,0.77232206,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.42060733,0.7650702,1.1095331,1.455809,1.8002719,3.0330863,4.264088,5.4969025,6.7297173,7.9625316,8.210908,8.457471,8.705847,8.952409,9.200785,8.9596615,8.72035,8.479226,8.239915,8.000604,7.027043,6.055295,5.081734,4.1099863,3.1382382,4.2368937,5.337362,6.43783,7.5382986,8.636953,9.545248,10.451729,11.3600235,12.268318,13.174799,12.725184,12.27557,11.8241415,11.374527,10.924912,11.873092,12.819458,13.767638,14.715817,15.662184,15.903308,16.142618,16.38193,16.623055,16.862366,15.917811,14.973258,14.026892,13.082338,12.137785,11.477866,10.817947,10.15803,9.498111,8.838193,9.947725,11.057259,12.166792,13.278138,14.387671,17.464268,20.542679,23.619276,26.697687,29.774284,30.907387,32.04049,33.171776,34.30488,35.43798,32.379513,29.322857,26.264389,23.207733,20.149265,20.444778,20.740292,21.035805,21.329504,21.625017,22.883213,24.139597,25.397793,26.654177,27.912373,25.680614,23.447044,21.215288,18.981718,16.749962,15.352167,13.954373,12.556579,11.160598,9.762803,8.736667,7.7123427,6.688019,5.661882,4.6375585,5.034597,5.431636,5.8304877,6.2275267,6.624565,7.28811,7.949841,8.613385,9.275117,9.936848,8.859948,7.783048,6.7043357,5.6274357,4.550536,4.1480584,3.7455807,3.343103,2.9406252,2.5381477,2.0649643,1.5917811,1.1204109,0.64722764,0.17585737,0.16679256,0.15954071,0.15228885,0.14503701,0.13778515,0.62547207,0.5728962,0.52032024,0.46774435,0.41516843,0.36259252,0.33539808,0.30820364,0.27919623,0.2520018,0.22480737,0.55839247,0.8901646,1.2219368,1.5555218,1.887294,3.0675328,4.2477713,5.42801,6.6082487,7.7866745,9.784559,11.782444,13.780329,15.7782135,17.774284,15.600543,13.424988,11.249433,9.07569,6.9001355,5.7253356,4.550536,3.3757362,2.1991236,1.0243238,2.032331,3.0403383,4.0483456,5.0545397,6.0625467,8.854509,11.648285,14.440247,17.23221,20.024172,17.527721,15.02946,12.5330105,10.034748,7.5382986,8.352319,9.168152,9.982172,10.798005,11.612025,12.794077,13.9779415,15.159993,16.342045,17.524096,18.075237,18.624565,19.175705,19.725033,20.27436,21.104698,21.935034,22.765371,23.595709,24.424232,23.022812,21.61958,20.218159,18.814926,17.411694,17.609306,17.80692,18.004532,18.202145,18.399757,20.468348,22.535126,24.601902,26.670492,28.73727,29.15969,29.582111,30.00453,30.42695,30.849371,29.533161,28.215137,26.897114,25.579088,24.262878,20.867199,17.473333,14.077655,10.681975,7.28811,7.895452,8.502794,9.110137,9.71748,10.324821,10.946668,11.570327,12.192173,12.815832,13.437678,11.137029,8.838193,6.5375433,4.2368937,1.938057,4.099108,6.261973,8.424837,10.587702,12.750566,11.980057,11.209548,10.440851,9.670342,8.899834,7.5999393,6.300045,5.0001507,3.7002566,2.4003625,2.5055144,2.610666,2.715818,2.819157,2.9243085,2.7448254,2.565342,2.3858588,2.2045624,2.0250793,8.167397,14.309713,20.45203,26.594349,32.736664,29.014652,25.29264,21.57063,17.846804,14.124791,16.642996,19.15939,21.677593,24.195799,26.71219,24.230246,21.748299,19.26454,16.782595,14.300649,12.639976,10.979301,9.32044,7.6597667,5.999093,5.0654173,4.1299286,3.1944401,2.2607644,1.3252757,1.3017071,1.2799516,1.258196,1.2346275,1.2128719,1.5446441,1.8782293,2.2100015,2.5417736,2.8753586,2.7067533,2.5399606,2.373168,2.2045624,2.03777,2.1447346,2.2516994,2.3604772,2.467442,2.5744069,4.3402324,6.104245,7.8700705,9.635896,11.399909,11.793322,12.184921,12.578335,12.969934,13.363347,13.575464,13.7875805,13.999697,14.211814,14.425743,15.089288,15.754644,16.420002,17.08536,17.750717,18.04079,18.330864,18.619125,18.9092,19.199274,16.604925,14.010575,11.4144125,8.820063,6.2257137,6.635443,7.0451727,7.454902,7.8646317,8.274362,8.439341,8.604321,8.7693,8.934279,9.099259,8.595256,8.089439,7.5854354,7.079619,6.5756154,7.6017523,8.629702,9.657652,10.685601,11.711739,10.770811,9.82807,8.885329,7.9425893,6.9998484,7.0850577,7.170267,7.2554765,7.3406854,7.4258947,5.9845896,4.5450974,3.105605,1.6642996,0.22480737,1.1693609,2.1157274,3.0602808,4.004834,4.949388,5.866747,6.784106,7.703278,8.620637,9.537996,9.956791,10.377398,10.798005,11.2168,11.637406,12.846653,14.057712,15.266958,16.478018,17.687263,18.238403,18.787731,19.337059,19.888199,20.437527,19.750414,19.063301,18.374376,17.687263,17.00015,14.112101,11.225864,8.337815,5.4497657,2.561716,3.48814,4.4127507,5.337362,6.261973,7.1883965,6.454147,5.7217097,4.989273,4.256836,3.5243993,5.2140803,6.9055743,8.595256,10.284937,11.974618,10.779876,9.585134,8.39039,7.1956487,5.999093,6.0752378,6.149569,6.2257137,6.300045,6.3743763,6.8022356,7.230095,7.6579537,8.0858135,8.511859,9.835322,11.156972,12.480434,13.802084,15.125546,14.860854,14.594349,14.329657,14.064963,13.800271,12.576522,11.354585,10.1326475,8.910711,7.686961,7.079619,6.472276,5.864934,5.2575917,4.650249,4.325729,3.9993954,3.6748753,3.350355,3.0258346,2.420305,1.8147756,1.209246,0.6055295,0.0,0.09064813,0.1794833,0.27013144,0.36077955,0.44961473,0.6399758,0.83033687,1.020698,1.209246,1.3996071,1.261822,1.1258497,0.9880646,0.85027945,0.7124943,0.58014804,0.44780177,0.3154555,0.18310922,0.05076295,0.21030366,0.36984438,0.5293851,0.69073874,0.85027945,0.75963134,0.67079616,0.58014804,0.4894999,0.40066472,0.42967212,0.4604925,0.4894999,0.52032024,0.5493277,1.0805258,1.6099107,2.1392958,2.6704938,3.199879,2.5798457,1.9598125,1.3397794,0.7197462,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.2755703,0.5493277,0.824898,1.1004683,1.3742256,1.1421664,0.9101072,0.678048,0.44417584,0.21211663,0.19579996,0.17767033,0.15954071,0.14322405,0.12509441,0.7124943,1.2998942,1.887294,2.474694,3.0620937,2.8427253,2.6233568,2.4021754,2.182807,1.9616255,1.6026589,1.2418793,0.88291276,0.52213323,0.16316663,0.15228885,0.14322405,0.13234627,0.12328146,0.11240368,0.16316663,0.21211663,0.26287958,0.31182957,0.36259252,0.45686656,0.5529536,0.64722764,0.7433147,0.8375887,0.774135,0.7124943,0.6508536,0.5873999,0.52575916,1.6606737,2.7955883,3.930503,5.0654173,6.200332,4.989273,3.780027,2.570781,1.3597219,0.15047589,0.18492219,0.21936847,0.25562772,0.29007402,0.3245203,0.43329805,0.5402629,0.64722764,0.7541924,0.8629702,0.79226464,0.72337204,0.6526665,0.581961,0.51306844,0.44780177,0.3825351,0.31726846,0.2520018,0.18673515,0.77232206,1.357909,1.9416829,2.5272698,3.1128569,2.5852847,2.0577126,1.5301404,1.0025684,0.4749962,0.94092757,1.405046,1.8691645,2.335096,2.7992141,2.3767939,1.9543737,1.5319533,1.1095331,0.6871128,0.67079616,0.6526665,0.6345369,0.61822027,0.6000906,0.79226464,0.98443866,1.1766127,1.3705997,1.5627737,1.696933,1.8329052,1.9670644,2.1030366,2.2371957,1.8147756,1.3923552,0.969935,0.5475147,0.12509441,0.11784257,0.11059072,0.10333887,0.09427405,0.0870222,0.13778515,0.18673515,0.2374981,0.28826106,0.33721104,0.6055295,0.872035,1.1403534,1.4068589,1.6751775,1.3506571,1.0243238,0.69980353,0.37528324,0.05076295,0.5747091,1.1004683,1.6244144,2.1501737,2.6741197,2.1447346,1.6153497,1.0841516,0.55476654,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.52213323,0.9445535,1.3669738,1.789394,2.2118144,3.247016,4.2822175,5.317419,6.352621,7.3878226,7.95528,8.5227375,9.090195,9.657652,10.225109,9.704789,9.184468,8.664148,8.145641,7.6253204,6.6191263,5.614745,4.610364,3.6041696,2.5997884,3.6494937,4.699199,5.750717,6.8004227,7.850128,8.535428,9.220728,9.904215,10.589515,11.274815,11.236742,11.200482,11.162411,11.124338,11.088079,12.279196,13.472125,14.665054,15.857984,17.0491,17.382685,17.714457,18.048042,18.379814,18.7134,17.565794,16.41819,15.270584,14.122978,12.975373,11.969179,10.964798,9.960417,8.954222,7.949841,8.87989,9.80994,10.73999,11.67004,12.60009,15.633177,18.66445,21.697536,24.730623,27.761896,28.885933,30.008156,31.13038,32.252605,33.37483,30.127811,26.878983,23.631968,20.38495,17.137936,17.598429,18.057108,18.5176,18.978092,19.436771,20.696781,21.956789,23.216799,24.476809,25.736816,23.626528,21.518053,19.407764,17.297476,15.187187,13.769451,12.351714,10.93579,9.518054,8.100317,7.262728,6.4251394,5.5875506,4.749962,3.9123733,4.0302157,4.1480584,4.265901,4.3819304,4.499773,5.5005283,6.4994707,7.500226,8.499168,9.499924,8.504607,7.509291,6.5157876,5.520471,4.5251546,3.9540713,3.3848011,2.8155308,2.2444477,1.6751775,1.3705997,1.064209,0.75963134,0.4550536,0.15047589,0.15228885,0.15410182,0.15772775,0.15954071,0.16316663,0.50037766,0.44961473,0.40066472,0.34990177,0.2991388,0.25018883,0.25018883,0.25018883,0.25018883,0.25018883,0.25018883,0.36259252,0.4749962,0.5873999,0.69980353,0.8122072,1.4757515,2.137483,2.7992141,3.4627585,4.12449,6.849373,9.574255,12.300951,15.025834,17.750717,15.850732,13.9507475,12.050762,10.150778,8.2507925,6.6118746,4.974769,3.3376641,1.7005589,0.06164073,1.5627737,3.0620937,4.5632267,6.0625467,7.5618668,11.037316,14.512766,17.988214,21.461851,24.9373,21.586945,18.238403,14.888049,11.537694,8.187339,8.838193,9.487233,10.138086,10.7871275,11.437981,13.000754,14.561715,16.124489,17.687263,19.250036,20.26167,21.275116,22.286749,23.300196,24.311829,25.337965,26.36229,27.388426,28.41275,29.437073,26.71219,23.987309,21.262424,18.537542,15.812659,16.525154,17.237648,17.950142,18.662638,19.375132,21.336756,23.300196,25.26182,27.22526,29.186884,29.07448,28.962078,28.849674,28.73727,28.624866,28.200632,27.774588,27.350353,26.924307,26.500074,22.424534,18.350807,14.275268,10.199727,6.1241875,7.02523,7.9244595,8.825501,9.724731,10.625773,11.563075,12.500377,13.437678,14.37498,15.312282,12.625471,9.936848,7.250037,4.5632267,1.8746033,4.5867953,7.3008003,10.012992,12.725184,15.437376,14.09941,12.763257,11.42529,10.087324,8.749357,7.224656,5.6999545,4.175253,2.6505513,1.1258497,1.49932,1.8746033,2.2498865,2.6251698,3.000453,2.8499773,2.6995013,2.5508385,2.4003625,2.2498865,9.07569,15.899682,22.725487,29.549477,36.375282,32.475597,28.575916,24.674421,20.774738,16.875055,18.312735,19.750414,21.188093,22.625772,24.06164,22.674723,21.287807,19.899076,18.512161,17.125244,15.161806,13.200181,11.236742,9.275117,7.311678,6.0879283,4.8623657,3.636803,2.4130533,1.1874905,1.0497054,0.9119202,0.774135,0.63816285,0.50037766,0.44961473,0.40066472,0.34990177,0.2991388,0.25018883,0.2991388,0.34990177,0.40066472,0.44961473,0.50037766,0.69980353,0.89922947,1.1004683,1.2998942,1.49932,3.4119956,5.3246713,7.2373466,9.1500225,11.062697,11.73712,12.413355,13.087777,13.762199,14.436621,14.68681,14.936998,15.187187,15.437376,15.687565,16.300346,16.913128,17.52591,18.136877,18.749659,18.611874,18.475903,18.338116,18.20033,18.062546,15.600543,13.136727,10.674724,8.212721,5.750717,6.474089,7.1992745,7.9244595,8.649645,9.374829,9.249735,9.12464,8.999546,8.874452,8.749357,8.412147,8.074935,7.7377243,7.400513,7.063302,8.312433,9.561564,10.812509,12.06164,13.312584,12.375282,11.437981,10.500679,9.563377,8.624263,8.52455,8.424837,8.325124,8.225411,8.125698,6.5248523,4.9258194,3.3249733,1.7241274,0.12509441,1.3379664,2.5508385,3.7618973,4.974769,6.187641,7.262728,8.337815,9.412902,10.487988,11.563075,11.3872175,11.213174,11.037316,10.863272,10.687414,11.075388,11.463363,11.849524,12.237497,12.625471,14.0867195,15.54978,17.01284,18.475903,19.93715,19.94984,19.96253,19.975222,19.987913,20.000603,16.563227,13.125849,9.686659,6.249282,2.811905,3.2252605,3.636803,4.0501585,4.461701,4.8750563,4.6756306,4.4743915,4.274966,4.07554,3.874301,5.774286,7.6742706,9.574255,11.47424,13.374225,11.961927,10.549629,9.137331,7.7250338,6.3127356,6.338117,6.3616858,6.3870673,6.412449,6.43783,6.8620634,7.28811,7.7123427,8.138389,8.562622,10.074633,11.586644,13.100468,14.612478,16.124489,16.050158,15.975826,15.899682,15.825351,15.749206,12.737875,9.724731,6.7115874,3.7002566,0.6871128,1.7132497,2.7375734,3.7618973,4.788034,5.812358,5.0744824,4.3384194,3.6005437,2.8626678,2.124792,1.7005589,1.2745126,0.85027945,0.42423326,0.0,0.11240368,0.22480737,0.33721104,0.44961473,0.5620184,0.7995165,1.0370146,1.2745126,1.5120108,1.7495089,1.4376793,1.1258497,0.8122072,0.50037766,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.0,0.0,0.0,0.0,0.0,0.099712946,0.19942589,0.2991388,0.40066472,0.50037766,0.40066472,0.2991388,0.19942589,0.099712946,0.0,0.42423326,0.85027945,1.2745126,1.7005589,2.124792,1.7241274,1.3252757,0.9246109,0.52575916,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.16316663,0.3245203,0.48768693,0.6508536,0.8122072,0.69980353,0.5873999,0.4749962,0.36259252,0.25018883,0.22480737,0.19942589,0.17585737,0.15047589,0.12509441,0.8629702,1.6008459,2.3369088,3.0747845,3.8126602,3.53709,3.2633326,2.9877625,2.712192,2.4366217,1.987007,1.5373923,1.0877775,0.63816285,0.18673515,0.16316663,0.13778515,0.11240368,0.0870222,0.06164073,0.12509441,0.18673515,0.25018883,0.31182957,0.37528324,0.48768693,0.6000906,0.7124943,0.824898,0.93730164,0.85027945,0.76325727,0.6744221,0.5873999,0.50037766,1.6878681,2.8753586,4.062849,5.2503395,6.43783,5.186886,3.9377546,2.6868105,1.4376793,0.18673515,0.19942589,0.21211663,0.22480737,0.2374981,0.25018883,0.37528324,0.50037766,0.62547207,0.7505665,0.87566096,0.8122072,0.7505665,0.6871128,0.62547207,0.5620184,0.48768693,0.41335547,0.33721104,0.26287958,0.18673515,0.40066472,0.61278135,0.824898,1.0370146,1.2491312,1.1131591,0.97537386,0.8375887,0.69980353,0.5620184,1.0243238,1.4866294,1.9507477,2.4130533,2.8753586,2.4620032,2.0504606,1.6371052,1.2255627,0.8122072,0.6744221,0.53663695,0.40066472,0.26287958,0.12509441,0.2374981,0.34990177,0.46230546,0.5747091,0.6871128,0.8883517,1.0877775,1.2872034,1.4866294,1.6878681,1.3742256,1.062396,0.7505665,0.43692398,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.12509441,0.18673515,0.25018883,0.31182957,0.37528324,0.5873999,0.7995165,1.0116332,1.2255627,1.4376793,1.162109,0.8883517,0.61278135,0.33721104,0.06164073,0.387974,0.7124943,1.0370146,1.3633479,1.6878681,1.3506571,1.0116332,0.6744221,0.33721104,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.62547207,1.1258497,1.6244144,2.124792,2.6251698,3.4627585,4.3003473,5.137936,5.975525,6.813113,7.699652,8.588004,9.474543,10.362894,11.249433,10.449916,9.6504,8.849071,8.049554,7.250037,6.2130227,5.1741953,4.137181,3.100166,2.0631514,3.0620937,4.062849,5.0617914,6.0625467,7.063302,7.5256076,7.987913,8.450218,8.912524,9.374829,9.750113,10.125396,10.500679,10.874149,11.249433,12.687112,14.124791,15.56247,17.00015,18.43783,18.862062,19.288109,19.712341,20.136576,20.562622,19.211964,17.863121,16.512463,15.161806,13.812962,12.462305,11.111648,9.762803,8.412147,7.063302,7.8120556,8.562622,9.313189,10.061942,10.812509,13.800271,16.788034,19.775795,22.761745,25.749508,26.862667,27.975826,29.087172,30.20033,31.311676,27.8743,24.436922,20.999546,17.562168,14.124791,14.750263,15.375735,15.999394,16.624866,17.25034,18.512161,19.775795,21.037619,22.29944,23.563074,21.574255,19.587248,17.60024,15.613234,13.6244135,12.186734,10.749055,9.313189,7.8755093,6.43783,5.7869763,5.137936,4.4870825,3.8380418,3.1871881,3.0258346,2.8626678,2.6995013,2.5381477,2.374981,3.7129474,5.050914,6.3870673,7.7250338,9.063,8.149267,7.2373466,6.3254266,5.411693,4.499773,3.7618973,3.0240216,2.2879589,1.550083,0.8122072,0.6744221,0.53663695,0.40066472,0.26287958,0.12509441,0.13778515,0.15047589,0.16316663,0.17585737,0.18673515,0.50037766,0.44236287,0.38434806,0.32814622,0.27013144,0.21211663,0.25018883,0.28826106,0.3245203,0.36259252,0.40066472,0.72337204,1.0442665,1.3669738,1.6896812,2.0123885,2.4148662,2.817344,3.2198215,3.6222992,4.024777,6.9744673,9.924157,12.87566,15.825351,18.77504,16.421816,14.070402,11.717177,9.365765,7.0125394,7.518356,8.02236,8.528176,9.03218,9.537996,9.751925,9.967669,10.181598,10.397341,10.613083,13.599032,16.586794,19.574556,22.562319,25.550081,22.516994,19.485722,16.452635,13.419549,10.388275,10.975676,11.563075,12.1504755,12.737875,13.325275,14.501887,15.680313,16.856926,18.035353,19.211964,20.352318,21.492672,22.633024,23.773378,24.911919,26.046833,27.181747,28.316662,29.45339,30.588305,28.120863,25.653421,23.184166,20.716722,18.24928,18.361685,18.474089,18.588305,18.700708,18.813112,20.412146,22.01299,23.612024,25.212872,26.811903,26.844538,26.87717,26.909803,26.942436,26.97507,26.719442,26.465628,26.210001,25.954372,25.700558,22.399153,19.099562,15.799969,12.500377,9.200785,9.712041,10.225109,10.738177,11.249433,11.762501,12.40429,13.047892,13.68968,14.333282,14.975071,12.815832,10.654781,8.495543,6.3344913,4.175253,6.1006193,8.024173,9.949538,11.874905,13.800271,12.620032,11.439794,10.259555,9.079316,7.900891,6.9508986,6.000906,5.049101,4.099108,3.149116,3.8507326,4.550536,5.2503395,5.9501433,6.6499467,6.338117,6.0244746,5.712645,5.4008155,5.087173,10.874149,16.66294,22.449915,28.236893,34.02568,30.769602,27.515333,24.259253,21.004984,17.750717,19.117691,20.484665,21.851639,23.220425,24.587399,23.361835,22.138086,20.912523,19.68696,18.463211,16.006647,13.551895,11.097144,8.642392,6.187641,5.1542525,4.122677,3.0892882,2.0577126,1.0243238,0.89922947,0.774135,0.6508536,0.52575916,0.40066472,0.37165734,0.3444629,0.31726846,0.29007402,0.26287958,0.3154555,0.3680314,0.42060733,0.47318324,0.52575916,0.8122072,1.1004683,1.3869164,1.6751775,1.9616255,3.7256382,5.487838,7.250037,9.012237,10.774437,11.543133,12.310016,13.0769,13.845595,14.612478,14.802839,14.9932,15.181748,15.372109,15.56247,16.148058,16.731833,17.31742,17.903006,18.48678,18.16226,17.837738,17.513218,17.186886,16.862366,14.724882,12.5873995,10.449916,8.312433,6.1749506,6.9019485,7.6307597,8.357758,9.084756,9.811753,9.692098,9.572442,9.452786,9.333132,9.211663,8.798307,8.383139,7.9679704,7.552802,7.137634,8.02236,8.907085,9.791811,10.6783495,11.563075,10.827013,10.092763,9.3567,8.62245,7.8882003,7.7757964,7.663393,7.549176,7.4367723,7.324369,5.9392653,4.554162,3.1690586,1.7857682,0.40066472,1.6026589,2.8046532,4.006647,5.2104545,6.412449,7.119504,7.8283725,8.535428,9.242483,9.949538,10.042,10.13446,10.226922,10.319383,10.411844,10.98474,11.557636,12.130532,12.701616,13.274512,14.4420595,15.609608,16.777155,17.944704,19.112251,19.192022,19.271791,19.353376,19.433146,19.512917,16.612177,13.713249,10.812509,7.911769,5.0128417,5.219519,5.42801,5.634688,5.8431783,6.049856,5.600241,5.1506267,4.699199,4.249584,3.7999697,5.2122674,6.624565,8.036863,9.449161,10.863272,9.869768,8.8780775,7.8845744,6.892884,5.89938,5.7779117,5.65463,5.5331616,5.40988,5.2884116,5.812358,6.338117,6.8620634,7.3878226,7.911769,8.912524,9.91328,10.912222,11.912977,12.91192,13.337966,13.762199,14.188245,14.612478,15.036712,12.64904,10.263181,7.8755093,5.487838,3.100166,3.4101827,3.720199,4.0302157,4.3402324,4.650249,4.4526362,4.255023,4.0574102,3.8597972,3.6621845,2.9297476,2.1973107,1.4648738,0.7324369,0.0,0.11059072,0.21936847,0.32995918,0.4405499,0.5493277,0.9481794,1.3452182,1.742257,2.1392958,2.5381477,2.0631514,1.5881553,1.1131591,0.63816285,0.16316663,0.13053331,0.09789998,0.065266654,0.032633327,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.11784257,0.21030366,0.30276474,0.39522585,0.48768693,0.61822027,0.7469406,0.8774739,1.0080072,1.1367276,1.5899682,2.0432088,2.4946365,2.9478772,3.3993049,2.8245957,2.2498865,1.6751775,1.1004683,0.52575916,0.48768693,0.44961473,0.41335547,0.37528324,0.33721104,0.42060733,0.50219065,0.5855869,0.6671702,0.7505665,0.6399758,0.5293851,0.42060733,0.3100166,0.19942589,0.19036107,0.1794833,0.17041849,0.15954071,0.15047589,0.90285534,1.6552348,2.4076142,3.159994,3.9123733,3.5497808,3.1871881,2.8245957,2.4620032,2.0994108,1.8256533,1.550083,1.2745126,1.0007553,0.72518504,0.59283876,0.4604925,0.32814622,0.19579996,0.06164073,0.11421664,0.16679256,0.21936847,0.27194437,0.3245203,0.41335547,0.50037766,0.5873999,0.6744221,0.76325727,0.6979906,0.6327239,0.56745726,0.50219065,0.43692398,1.3977941,2.3568513,3.3177216,4.2767787,5.237649,4.2368937,3.2379513,2.2371957,1.2382535,0.2374981,0.23024625,0.2229944,0.21574254,0.20667773,0.19942589,0.3245203,0.44961473,0.5747091,0.69980353,0.824898,0.774135,0.72518504,0.6744221,0.62547207,0.5747091,0.49675176,0.42060733,0.34264994,0.26469254,0.18673515,0.36259252,0.53663695,0.7124943,0.8883517,1.062396,1.2545701,1.4467441,1.6407311,1.8329052,2.0250793,2.467442,2.909805,3.3521678,3.7945306,4.2368937,4.162562,4.0882306,4.0120864,3.9377546,3.8616104,3.1273603,2.3931105,1.6570477,0.922798,0.18673515,0.2755703,0.36259252,0.44961473,0.53663695,0.62547207,0.7705091,0.9155461,1.0605831,1.2056202,1.3506571,1.1167849,0.88472575,0.6526665,0.42060733,0.18673515,0.17223145,0.15772775,0.14322405,0.12690738,0.11240368,0.16316663,0.21211663,0.26287958,0.31182957,0.36259252,0.53482395,0.7070554,0.8792868,1.0533313,1.2255627,1.0333886,0.83940166,0.64722764,0.4550536,0.26287958,0.5058166,0.7469406,0.9898776,1.2328146,1.4757515,1.1802386,0.88472575,0.58921283,0.2955129,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.034446288,0.07070554,0.10515183,0.13959812,0.17585737,0.70342946,1.2291887,1.7567607,2.2843328,2.811905,3.3757362,3.9377546,4.499773,5.0617914,5.6256227,6.33993,7.0542374,7.7703576,8.484665,9.200785,8.609759,8.020547,7.4295206,6.8403077,6.249282,5.576673,4.9058766,4.233268,3.5606585,2.8880494,3.7147603,4.5432844,5.369995,6.1967063,7.02523,7.3008003,7.574558,7.850128,8.125698,8.399456,8.859948,9.32044,9.77912,10.239613,10.700105,11.920229,13.140353,14.3604765,15.580601,16.800724,17.197763,17.5948,17.99184,18.390692,18.787731,17.859495,16.933071,16.004833,15.07841,14.150173,13.182051,12.215742,11.24762,10.279498,9.313189,9.494485,9.677594,9.860703,10.042,10.225109,12.732436,15.239763,17.747091,20.254417,22.761745,23.729868,24.697989,25.664299,26.63242,27.600542,24.96812,22.333885,19.703278,17.070856,14.436621,15.033086,15.627737,16.22239,16.817041,17.411694,18.075237,18.736969,19.400513,20.062244,20.725788,18.920078,17.114367,15.310469,13.504758,11.700861,10.440851,9.179029,7.9208336,6.6608243,5.4008155,4.9693303,4.539658,4.1099863,3.680314,3.2506418,3.094727,2.9406252,2.7847104,2.6306088,2.474694,3.5171473,4.559601,5.6020546,6.644508,7.686961,6.885632,6.0824895,5.279347,4.478018,3.6748753,3.0747845,2.474694,1.8746033,1.2745126,0.6744221,0.5728962,0.46955732,0.3680314,0.26469254,0.16316663,0.16679256,0.17223145,0.17767033,0.18310922,0.18673515,0.50037766,0.43511102,0.36984438,0.3045777,0.23931105,0.17585737,0.25018883,0.3245203,0.40066472,0.4749962,0.5493277,1.0823387,1.6153497,2.1483607,2.6795588,3.2125697,3.3557937,3.4972048,3.6404288,3.7818398,3.925064,7.0995617,10.274059,13.45037,16.624866,19.799364,16.99471,14.190058,11.385405,8.580752,5.774286,8.423024,11.069949,13.716875,16.365614,19.012539,17.94289,16.873243,15.801782,14.732134,13.662486,16.162561,18.662638,21.162712,23.662788,26.162863,23.447044,20.73304,18.017221,15.303217,12.5873995,13.113158,13.637105,14.162864,14.68681,15.212569,16.004833,16.797098,17.589363,18.381628,19.175705,20.442966,21.710226,22.977488,24.24475,25.512009,26.757515,28.00302,29.246712,30.492218,31.737722,29.527721,27.31772,25.10772,22.897717,20.687716,20.20003,19.712341,19.224655,18.736969,18.24928,19.487535,20.725788,21.962229,23.200481,24.436922,24.614594,24.792263,24.969934,25.147604,25.325274,25.240065,25.154856,25.069647,24.984438,24.89923,22.375584,19.850128,17.32467,14.799213,12.27557,12.400664,12.525759,12.650853,12.774135,12.899229,13.247317,13.595407,13.941682,14.289771,14.63786,13.00438,11.372714,9.739235,8.107569,6.4759026,7.61263,8.749357,9.8878975,11.024626,12.163166,11.1406555,10.118144,9.0956335,8.073122,7.0506115,6.6753283,6.300045,5.924762,5.5494785,5.1741953,6.200332,7.224656,8.2507925,9.275117,10.29944,9.824444,9.349448,8.874452,8.399456,7.9244595,12.674421,17.424383,22.174345,26.924307,31.674269,29.065416,26.45475,23.844084,21.235231,18.624565,19.922646,21.220728,22.516994,23.815077,25.113157,24.050762,22.988365,21.924156,20.861761,19.799364,16.8533,13.905423,10.957546,8.009668,5.0617914,4.2223897,3.3829882,2.5417736,1.7023718,0.8629702,0.7505665,0.63816285,0.52575916,0.41335547,0.2991388,0.2955129,0.29007402,0.28463513,0.27919623,0.2755703,0.32995918,0.38434806,0.4405499,0.4949388,0.5493277,0.9246109,1.2998942,1.6751775,2.0504606,2.4257438,4.0374675,5.6491914,7.262728,8.874452,10.487988,11.347333,12.206677,13.067834,13.927178,14.788336,14.917056,15.047589,15.1781225,15.306843,15.437376,15.995769,16.55235,17.11074,17.66732,18.225714,17.712645,17.199575,16.68832,16.175253,15.662184,13.849221,12.038072,10.225109,8.412147,6.599184,7.3298078,8.0604315,8.789243,9.519867,10.25049,10.13446,10.020245,9.904215,9.789998,9.675781,9.182655,8.689529,8.198216,7.705091,7.211965,7.7322855,8.252605,8.772926,9.293246,9.811753,9.280556,8.747544,8.214534,7.6833353,7.1503243,7.02523,6.9001355,6.775041,6.6499467,6.5248523,5.3554916,4.1843176,3.0149567,1.845596,0.6744221,1.8673514,3.0602808,4.25321,5.4443264,6.637256,6.978093,7.317117,7.6579537,7.996978,8.337815,8.696781,9.057561,9.418341,9.7773075,10.138086,10.894093,11.651911,12.409729,13.167547,13.925365,14.7974,15.6694355,16.543283,17.41532,18.287354,18.434204,18.582867,18.729717,18.87838,19.025229,16.66294,14.300649,11.936545,9.574255,7.211965,7.215591,7.217404,7.219217,7.2228427,7.224656,6.5248523,5.825049,5.125245,4.4254417,3.7256382,4.650249,5.57486,6.4994707,7.4258947,8.350506,7.7776093,7.2047133,6.6318173,6.060734,5.487838,5.217706,4.947575,4.6774435,4.407312,4.137181,4.762653,5.388125,6.011784,6.637256,7.262728,7.750415,8.238102,8.725789,9.211663,9.699349,10.625773,11.5503845,12.474996,13.399607,14.324218,12.562017,10.799818,9.037619,7.2754188,5.5132194,5.1071157,4.702825,4.2967215,3.8924308,3.48814,3.83079,4.171627,4.514277,4.856927,5.199577,4.160749,3.1201086,2.079468,1.0406405,0.0,0.10696479,0.21574254,0.32270733,0.42967212,0.53663695,1.0950294,1.651609,2.2100015,2.7683938,3.3249733,2.6868105,2.0504606,1.4122978,0.774135,0.13778515,0.11059072,0.08339628,0.054388877,0.027194439,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.13415924,0.21936847,0.3045777,0.38978696,0.4749962,0.83577573,1.1947423,1.5555218,1.9144884,2.275268,2.7557032,3.2343252,3.7147603,4.195195,4.6756306,3.925064,3.1744974,2.4257438,1.6751775,0.9246109,0.87566096,0.824898,0.774135,0.72518504,0.6744221,0.678048,0.67986095,0.68167394,0.6852999,0.6871128,0.58014804,0.47318324,0.36440548,0.2574407,0.15047589,0.15410182,0.15954071,0.16497959,0.17041849,0.17585737,0.94274056,1.7096237,2.47832,3.245203,4.0120864,3.5624714,3.1128569,2.663242,2.2118144,1.7621996,1.6624867,1.5627737,1.4630609,1.3633479,1.261822,1.0225109,0.78319985,0.5420758,0.30276474,0.06164073,0.10515183,0.14684997,0.19036107,0.23205921,0.2755703,0.33721104,0.40066472,0.46230546,0.52575916,0.5873999,0.54570174,0.50219065,0.4604925,0.4169814,0.37528324,1.1077201,1.840157,2.572594,3.3050308,4.0374675,3.2869012,2.5381477,1.7875811,1.0370146,0.28826106,0.25925365,0.23205921,0.20486477,0.17767033,0.15047589,0.2755703,0.40066472,0.52575916,0.6508536,0.774135,0.73787576,0.69980353,0.66173136,0.62547207,0.5873999,0.5076295,0.42785916,0.3480888,0.26831847,0.18673515,0.3245203,0.46230546,0.6000906,0.73787576,0.87566096,1.3977941,1.9199274,2.4420607,2.9641938,3.48814,3.9105604,4.3329806,4.7554007,5.177821,5.600241,5.863121,6.1241875,6.3870673,6.6499467,6.9128265,5.580299,4.2477713,2.9152439,1.5827163,0.25018883,0.31182957,0.37528324,0.43692398,0.50037766,0.5620184,0.6526665,0.7433147,0.8321498,0.922798,1.0116332,0.85934424,0.7070554,0.55476654,0.40247768,0.25018883,0.23205921,0.21574254,0.19761293,0.1794833,0.16316663,0.19942589,0.2374981,0.2755703,0.31182957,0.34990177,0.48224804,0.61459434,0.7469406,0.8792868,1.0116332,0.90285534,0.79226464,0.68167394,0.5728962,0.46230546,0.62184614,0.78319985,0.94274056,1.1022812,1.261822,1.0098201,0.75781834,0.5058166,0.2520018,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.045324065,0.09064813,0.13415924,0.1794833,0.22480737,0.7795739,1.3343405,1.8909199,2.4456866,3.000453,3.2869012,3.5751622,3.8616104,4.1498713,4.4381323,4.9802084,5.522284,6.0643597,6.6082487,7.1503243,6.7696023,6.390693,6.009971,5.6292486,5.2503395,4.942136,4.6357455,4.327542,4.019338,3.7129474,4.367427,5.0219064,5.678199,6.3326783,6.987158,7.07418,7.1630154,7.250037,7.3370595,7.4258947,7.9697833,8.515485,9.059374,9.605076,10.150778,11.153346,12.154101,13.15667,14.159238,15.161806,15.531651,15.903308,16.273151,16.642996,17.01284,16.507025,16.003021,15.497204,14.9932,14.487384,13.901797,13.318023,12.732436,12.14685,11.563075,11.176914,10.792566,10.408218,10.022058,9.637709,11.664601,13.693306,15.720199,17.747091,19.775795,20.597069,21.420153,22.243238,23.06451,23.887594,22.06013,20.232662,18.405195,16.57773,14.750263,15.3159075,15.879739,16.445383,17.009214,17.57486,17.638313,17.699953,17.761595,17.825048,17.886688,16.264088,14.641486,13.020698,11.398096,9.775495,8.693155,7.609004,6.526665,5.4443264,4.361988,4.1516843,3.9431937,3.73289,3.5225863,3.3122826,3.1654327,3.0167696,2.8699198,2.72307,2.5744069,3.3231604,4.070101,4.8170414,5.565795,6.3127356,5.620184,4.9276323,4.2350807,3.5425289,2.8499773,2.3876717,1.9253663,1.4630609,1.0007553,0.53663695,0.46955732,0.40247768,0.33539808,0.26831847,0.19942589,0.19761293,0.19579996,0.19217403,0.19036107,0.18673515,0.50037766,0.42785916,0.35534066,0.28282216,0.21030366,0.13778515,0.25018883,0.36259252,0.4749962,0.5873999,0.69980353,1.4431182,2.18462,2.9279346,3.6694362,4.4127507,4.2949085,4.177066,4.059223,3.9431937,3.825351,7.224656,10.625773,14.025079,17.424383,20.8255,17.567608,14.309713,11.05182,7.795739,4.537845,9.327692,14.117539,18.907387,23.697233,28.487082,26.132042,23.777004,21.421967,19.066927,16.71189,18.724277,20.736666,22.750868,24.763256,26.775644,24.377094,21.980358,19.581808,17.185072,14.788336,15.250641,15.712947,16.175253,16.637558,17.099863,17.50778,17.915697,18.3218,18.729717,19.137632,20.531801,21.927782,23.32195,24.717932,26.1121,27.468197,28.82248,30.176762,31.532858,32.887142,30.93458,28.98202,27.029459,25.076899,23.124338,22.038374,20.950596,19.862818,18.77504,17.687263,18.562923,19.436771,20.312433,21.188093,22.061941,22.38465,22.707355,23.030064,23.352772,23.675478,23.760687,23.844084,23.929293,24.014502,24.099712,22.350203,20.600695,18.849373,17.099863,15.350354,15.087475,14.824595,14.561715,14.300649,14.037769,14.090345,14.142921,14.195497,14.248073,14.300649,13.194741,12.090648,10.98474,9.880646,8.774739,9.12464,9.474543,9.824444,10.174346,10.524248,9.659465,8.794682,7.9298983,7.065115,6.200332,6.399758,6.599184,6.8004227,6.9998484,7.1992745,8.549932,9.900589,11.249433,12.60009,13.9507475,13.312584,12.674421,12.038072,11.399909,10.761745,14.474693,18.187641,21.900587,25.611723,29.324669,27.359419,25.394167,23.430729,21.465477,19.500225,20.727602,21.954977,23.182352,24.409729,25.637104,24.737875,23.836832,22.937603,22.038374,21.137331,17.698141,14.257137,10.817947,7.3769445,3.9377546,3.290527,2.6432993,1.9942589,1.3470312,0.69980353,0.6000906,0.50037766,0.40066472,0.2991388,0.19942589,0.21755551,0.23568514,0.2520018,0.27013144,0.28826106,0.3444629,0.40247768,0.4604925,0.5166943,0.5747091,1.0370146,1.49932,1.9616255,2.4257438,2.8880494,4.349297,5.812358,7.2754188,8.736667,10.199727,11.153346,12.105151,13.056956,14.010575,14.96238,15.033086,15.101978,15.172684,15.243389,15.312282,15.841667,16.372866,16.90225,17.431635,17.962833,17.26303,16.563227,15.861609,15.161806,14.462003,12.975373,11.486931,10.000301,8.511859,7.02523,7.757667,8.490104,9.222541,9.954978,10.687414,10.576823,10.468046,10.357455,10.246864,10.138086,9.567003,8.997733,8.42665,7.85738,7.28811,7.4422116,7.5981264,7.752228,7.9081426,8.062244,7.7322855,7.402326,7.072367,6.742408,6.412449,6.2746634,6.1368785,5.999093,5.863121,5.7253356,4.7699046,3.8144734,2.8608549,1.9054236,0.9499924,2.132044,3.3140955,4.49796,5.6800117,6.8620634,6.834869,6.8076744,6.78048,6.7532854,6.7242785,7.3515635,7.9806614,8.607946,9.235231,9.862516,10.805257,11.747997,12.690738,13.631665,14.574407,15.152741,15.729263,16.307598,16.88412,17.462456,17.678198,17.892128,18.10787,18.3218,18.537542,16.71189,14.888049,13.062395,11.236742,9.412902,9.20985,9.006798,8.805559,8.602508,8.399456,7.4494634,6.4994707,5.5494785,4.599486,3.6494937,4.0882306,4.5251546,4.9620786,5.4008155,5.8377395,5.6854506,5.5331616,5.37906,5.2267714,5.0744824,4.6575007,4.2405195,3.8217251,3.4047437,2.9877625,3.7129474,4.4381323,5.163317,5.8866897,6.6118746,6.588306,6.5629244,6.5375433,6.5121617,6.48678,7.911769,9.336758,10.761745,12.186734,13.611723,12.474996,11.338268,10.199727,9.063,7.9244595,6.8058615,5.6854506,4.5650396,3.444629,2.324218,3.207131,4.0900435,4.972956,5.8558693,6.736969,5.389938,4.0429068,2.6958754,1.3470312,0.0,0.10515183,0.21030366,0.3154555,0.42060733,0.52575916,1.2418793,1.9598125,2.6777458,3.395679,4.1117992,3.3122826,2.5127661,1.7132497,0.9119202,0.11240368,0.09064813,0.06707962,0.045324065,0.02175555,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.15228885,0.23024625,0.30820364,0.38434806,0.46230546,1.0533313,1.6425442,2.231757,2.8227828,3.4119956,3.919625,4.4272547,4.934884,5.4425135,5.9501433,5.0255322,4.100921,3.1744974,2.2498865,1.3252757,1.261822,1.2001812,1.1367276,1.0750868,1.0116332,0.9354887,0.8575313,0.7795739,0.7016165,0.62547207,0.52032024,0.41516843,0.3100166,0.20486477,0.099712946,0.11965553,0.13959812,0.15954071,0.1794833,0.19942589,0.9826257,1.7658255,2.5472124,3.3304121,4.1117992,3.5751622,3.0367124,2.5000753,1.9616255,1.4249886,1.49932,1.5754645,1.649796,1.7241274,1.8002719,1.452183,1.1059072,0.75781834,0.40972954,0.06164073,0.09427405,0.12690738,0.15954071,0.19217403,0.22480737,0.26287958,0.2991388,0.33721104,0.37528324,0.41335547,0.39159992,0.37165734,0.35171473,0.33177215,0.31182957,0.81764615,1.3216497,1.8274662,2.333283,2.8372865,2.3369088,1.8383441,1.3379664,0.8375887,0.33721104,0.29007402,0.24293698,0.19579996,0.14684997,0.099712946,0.22480737,0.34990177,0.4749962,0.6000906,0.72518504,0.69980353,0.6744221,0.6508536,0.62547207,0.6000906,0.5166943,0.43511102,0.35171473,0.27013144,0.18673515,0.28826106,0.387974,0.48768693,0.5873999,0.6871128,1.5392052,2.3931105,3.245203,4.0972953,4.949388,5.351866,5.754343,6.156821,6.5592985,6.9617763,7.5618668,8.161958,8.762048,9.362139,9.96223,8.033237,6.1024323,4.171627,2.2426348,0.31182957,0.34990177,0.387974,0.42423326,0.46230546,0.50037766,0.53482395,0.56927025,0.6055295,0.6399758,0.6744221,0.60190356,0.5293851,0.45686656,0.38434806,0.31182957,0.291887,0.27194437,0.2520018,0.23205921,0.21211663,0.2374981,0.26287958,0.28826106,0.31182957,0.33721104,0.42967212,0.52213323,0.61459434,0.7070554,0.7995165,0.77232206,0.7451276,0.7179332,0.69073874,0.66173136,0.73968875,0.81764615,0.89560354,0.97174793,1.0497054,0.83940166,0.629098,0.42060733,0.21030366,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.054388877,0.11059072,0.16497959,0.21936847,0.2755703,0.8575313,1.4394923,2.0232663,2.6052272,3.1871881,3.199879,3.2125697,3.2252605,3.2379513,3.2506418,3.6204863,3.9903307,4.360175,4.7300196,5.0998635,4.9294453,4.76084,4.590421,4.420003,4.249584,4.307599,4.365614,4.421816,4.4798307,4.537845,5.0200934,5.5023413,5.9845896,6.4668374,6.9508986,6.849373,6.7496595,6.6499467,6.550234,6.450521,7.079619,7.71053,8.339628,8.970539,9.599637,10.384649,11.169662,11.954676,12.739688,13.524701,13.867351,14.210001,14.55265,14.895301,15.23795,15.154554,15.072971,14.989574,14.907991,14.824595,14.623356,14.420304,14.217253,14.014201,13.812962,12.859344,11.907538,10.955733,10.002114,9.050309,10.596766,12.145037,13.693306,15.239763,16.788034,17.464268,18.142317,18.820364,19.4966,20.174648,19.152136,18.129625,17.107115,16.084604,15.062093,15.596917,16.13174,16.668379,17.203201,17.738026,17.199575,16.66294,16.124489,15.5878525,15.049402,13.60991,12.170418,10.729113,9.28962,7.850128,6.94546,6.0389786,5.1343102,4.229642,3.3249733,3.3358512,3.3449159,3.3557937,3.3648586,3.3757362,3.2343252,3.094727,2.955129,2.8155308,2.6741197,3.1273603,3.5806012,4.0320287,4.4852695,4.936697,4.3547363,3.7727752,3.1908143,2.6070402,2.0250793,1.7005589,1.3742256,1.0497054,0.72518504,0.40066472,0.3680314,0.33539808,0.30276474,0.27013144,0.2374981,0.22662032,0.21755551,0.20667773,0.19761293,0.18673515,0.50037766,0.42060733,0.34083697,0.25925365,0.1794833,0.099712946,0.25018883,0.40066472,0.5493277,0.69980353,0.85027945,1.8020848,2.7557032,3.7075086,4.6593137,5.612932,5.235836,4.856927,4.4798307,4.102734,3.7256382,7.3497505,10.975676,14.599788,18.225714,21.849825,18.140503,14.429369,10.720048,7.0107265,3.299592,10.232361,17.16513,24.097898,31.030668,37.963436,34.32301,30.682579,27.04215,23.401722,19.763105,21.287807,22.812508,24.33721,25.861912,27.386612,25.307144,23.227676,21.148209,19.066927,16.98746,17.388124,17.786976,18.187641,18.588305,18.987158,19.010725,19.03248,19.054237,19.077805,19.099562,20.62245,22.145338,23.668226,25.189302,26.71219,28.177065,29.64194,31.106812,32.571686,34.038372,32.343254,30.648132,28.953012,27.257893,25.562773,23.874905,22.187037,20.499168,18.813112,17.125244,17.638313,18.149569,18.662638,19.175705,19.68696,20.154705,20.62245,21.090193,21.557938,22.025682,22.279497,22.535126,22.790752,23.044567,23.300196,22.324821,21.349447,20.375887,19.400513,18.425138,17.774284,17.125244,16.474392,15.825351,15.174497,14.9333725,14.690435,14.447499,14.204562,13.961625,13.385102,12.806767,12.230246,11.651911,11.075388,10.636651,10.199727,9.762803,9.325879,8.887142,8.180087,7.473032,6.7641635,6.057108,5.3500524,6.1241875,6.9001355,7.6742706,8.450218,9.224354,10.899531,12.574709,14.249886,15.925063,17.60024,16.800724,15.999394,15.199879,14.400362,13.600845,16.274965,18.949085,21.625017,24.299137,26.97507,25.655233,24.335396,23.01556,21.695723,20.375887,21.532557,22.689226,23.84771,25.00438,26.162863,25.424988,24.68711,23.949236,23.213173,22.475298,18.542982,14.610665,10.676537,6.7442207,2.811905,2.3568513,1.9017978,1.4467441,0.9916905,0.53663695,0.44961473,0.36259252,0.2755703,0.18673515,0.099712946,0.13959812,0.1794833,0.21936847,0.25925365,0.2991388,0.36077955,0.42060733,0.48043507,0.5402629,0.6000906,1.1494182,1.7005589,2.2498865,2.7992141,3.350355,4.6629395,5.975525,7.28811,8.600695,9.91328,10.957546,12.001812,13.047892,14.092158,15.138238,15.147303,15.15818,15.167245,15.1781225,15.187187,15.689378,16.193382,16.695572,17.197763,17.699953,16.813416,15.925063,15.036712,14.150173,13.261822,12.099712,10.937603,9.775495,8.613385,7.4494634,8.185526,8.919776,9.655839,10.390089,11.124338,11.019187,10.915848,10.810696,10.705544,10.600392,9.953164,9.304124,8.656897,8.009668,7.362441,7.1521373,6.9418335,6.733343,6.5230393,6.3127356,6.185828,6.057108,5.9302006,5.803293,5.674573,5.524097,5.375434,5.224958,5.0744824,4.9258194,4.1843176,3.444629,2.70494,1.9652514,1.2255627,2.3967366,3.5697234,4.74271,5.915697,7.0868707,6.6916447,6.298232,5.903006,5.5077806,5.1125546,6.008158,6.9019485,7.797552,8.693155,9.5869465,10.714609,11.842272,12.969934,14.097597,15.22526,15.508082,15.789091,16.071913,16.354736,16.637558,16.92038,17.203201,17.484211,17.767033,18.049856,16.762651,15.475449,14.188245,12.899229,11.612025,11.205922,10.798005,10.390089,9.982172,9.574255,8.375887,7.175706,5.975525,4.7753434,3.5751622,3.5243993,3.4754493,3.4246864,3.3757362,3.3249733,3.5932918,3.8597972,4.1281157,4.3946214,4.6629395,4.0972953,3.531651,2.9678197,2.4021754,1.8383441,2.663242,3.48814,4.313038,5.137936,5.962834,5.424384,4.8877473,4.349297,3.8126602,3.2742105,5.199577,7.124943,9.050309,10.975676,12.899229,12.387974,11.874905,11.361836,10.850581,10.337513,8.502794,6.6680765,4.8315454,2.9968271,1.162109,2.5852847,4.006647,5.429823,6.8529987,8.274362,6.6191263,4.9657044,3.3104696,1.6552348,0.0,0.10333887,0.20486477,0.30820364,0.40972954,0.51306844,1.3905423,2.268016,3.1454902,4.022964,4.900438,3.9377546,2.9750717,2.0123885,1.0497054,0.0870222,0.07070554,0.052575916,0.034446288,0.018129626,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.17041849,0.23931105,0.3100166,0.38072214,0.44961473,1.2708868,2.0903459,2.909805,3.729264,4.550536,5.08536,5.620184,6.155008,6.6898317,7.224656,6.1241875,5.0255322,3.925064,2.8245957,1.7241274,1.649796,1.5754645,1.49932,1.4249886,1.3506571,1.1929294,1.0352017,0.8774739,0.7197462,0.5620184,0.4604925,0.35715362,0.25562772,0.15228885,0.05076295,0.08520924,0.11965553,0.15410182,0.19036107,0.22480737,1.0225109,1.8202144,2.617918,3.4156215,4.213325,3.587853,2.962381,2.3369088,1.7132497,1.0877775,1.3379664,1.5881553,1.8383441,2.08672,2.3369088,1.8818551,1.4268016,0.97174793,0.5166943,0.06164073,0.08520924,0.10696479,0.13053331,0.15228885,0.17585737,0.18673515,0.19942589,0.21211663,0.22480737,0.2374981,0.23931105,0.24293698,0.24474995,0.24837588,0.25018883,0.5275721,0.80495536,1.0823387,1.3597219,1.6371052,1.3869164,1.1367276,0.8883517,0.63816285,0.387974,0.3208944,0.2520018,0.18492219,0.11784257,0.05076295,0.17585737,0.2991388,0.42423326,0.5493277,0.6744221,0.66173136,0.6508536,0.63816285,0.62547207,0.61278135,0.5275721,0.44236287,0.35715362,0.27194437,0.18673515,0.25018883,0.31182957,0.37528324,0.43692398,0.50037766,1.6824293,2.864481,4.0483456,5.230397,6.412449,6.794984,7.177519,7.560054,7.9425893,8.325124,9.262425,10.199727,11.137029,12.07433,13.013446,10.484363,7.957093,5.429823,2.902553,0.37528324,0.387974,0.40066472,0.41335547,0.42423326,0.43692398,0.4169814,0.39703882,0.3770962,0.35715362,0.33721104,0.3444629,0.35171473,0.36077955,0.3680314,0.37528324,0.35171473,0.32995918,0.30820364,0.28463513,0.26287958,0.2755703,0.28826106,0.2991388,0.31182957,0.3245203,0.3770962,0.42967212,0.48224804,0.53482395,0.5873999,0.6417888,0.6979906,0.7523795,0.80676836,0.8629702,0.8575313,0.8520924,0.8466535,0.8430276,0.8375887,0.67079616,0.50219065,0.33539808,0.16679256,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.065266654,0.13053331,0.19579996,0.25925365,0.3245203,0.9354887,1.5446441,2.1556125,2.764768,3.3757362,3.1128569,2.8499773,2.5870976,2.324218,2.0631514,2.2607644,2.4565642,2.6541772,2.8517902,3.049403,3.0892882,3.1291735,3.1708715,3.2107568,3.2506418,3.673062,4.0954823,4.517903,4.940323,5.3627434,5.67276,5.9827766,6.2927933,6.60281,6.9128265,6.624565,6.338117,6.049856,5.763408,5.475147,6.189454,6.9055743,7.6198816,8.334189,9.050309,9.617766,10.185224,10.752681,11.320138,11.887595,12.203052,12.516694,12.8321495,13.147605,13.46306,13.802084,14.142921,14.481945,14.8227825,15.161806,15.343102,15.522586,15.702069,15.883366,16.062849,14.541773,13.022511,11.503247,9.982172,8.46291,9.530745,10.596766,11.664601,12.732436,13.800271,14.333282,14.86448,15.397491,15.930502,16.4617,16.244144,16.026588,15.810846,15.593291,15.375735,15.879739,16.385555,16.889559,17.395376,17.89938,16.762651,15.624111,14.487384,13.3506565,12.212116,10.955733,9.697536,8.439341,7.1829576,5.924762,5.197764,4.4707656,3.7419548,3.0149567,2.2879589,2.518205,2.7466383,2.9768846,3.207131,3.437377,3.3050308,3.1726844,3.0403383,2.907992,2.7756457,2.9333735,3.0892882,3.247016,3.4047437,3.5624714,3.0892882,2.617918,2.1447346,1.6733645,1.2001812,1.0116332,0.824898,0.63816285,0.44961473,0.26287958,0.26469254,0.26831847,0.27013144,0.27194437,0.2755703,0.2574407,0.23931105,0.2229944,0.20486477,0.18673515,0.50037766,0.41335547,0.3245203,0.2374981,0.15047589,0.06164073,0.25018883,0.43692398,0.62547207,0.8122072,1.0007553,2.1628644,3.3249733,4.4870825,5.6491914,6.813113,6.1749506,5.5367875,4.900438,4.262275,3.6241121,7.474845,11.325577,15.174497,19.025229,22.87415,18.7134,14.5508375,10.388275,6.2257137,2.0631514,11.137029,20.212719,29.28841,38.36229,47.43798,42.51216,37.588154,32.662334,27.738327,22.812508,23.849524,24.88835,25.925365,26.96238,27.999393,26.237194,24.474995,22.712795,20.950596,19.188396,19.525606,19.862818,20.20003,20.537241,20.87445,20.511858,20.149265,19.786674,19.425894,19.063301,20.713097,22.362894,24.01269,25.662485,27.31228,28.887745,30.463211,32.03686,33.612328,35.18779,33.75011,32.31243,30.874752,29.437073,27.999393,25.71325,23.42529,21.137331,18.849373,16.563227,16.71189,16.862366,17.01284,17.163317,17.31198,17.92476,18.537542,19.150324,19.763105,20.375887,20.80012,21.224354,21.650398,22.074633,22.500679,22.29944,22.100014,21.900587,21.699348,21.499924,20.462908,19.425894,18.387066,17.350052,16.313038,15.774588,15.23795,14.699501,14.162864,13.6244135,13.575464,13.524701,13.475751,13.424988,13.374225,12.1504755,10.924912,9.699349,8.4756,7.250037,6.70071,6.149569,5.600241,5.049101,4.499773,5.8504305,7.1992745,8.549932,9.900589,11.249433,13.24913,15.250641,17.25034,19.250036,21.249735,20.287052,19.324368,18.361685,17.400814,16.438131,18.075237,19.712341,21.349447,22.988365,24.625471,23.949236,23.274813,22.600391,21.924156,21.249735,22.337511,23.42529,24.513067,25.600845,26.68681,26.1121,25.537392,24.962683,24.387972,23.813263,19.387821,14.96238,10.536939,6.11331,1.6878681,1.4249886,1.162109,0.89922947,0.63816285,0.37528324,0.2991388,0.22480737,0.15047589,0.07433146,0.0,0.06164073,0.12509441,0.18673515,0.25018883,0.31182957,0.37528324,0.43692398,0.50037766,0.5620184,0.62547207,1.261822,1.8999848,2.5381477,3.1744974,3.8126602,4.974769,6.1368785,7.3008003,8.46291,9.625018,10.761745,11.900287,13.037014,14.175554,15.312282,15.263332,15.212569,15.161806,15.112856,15.062093,15.537089,16.012085,16.487082,16.962078,17.437075,16.361988,15.2869005,14.211814,13.136727,12.06164,11.225864,10.388275,9.550687,8.713099,7.8755093,8.613385,9.349448,10.087324,10.825199,11.563075,11.463363,11.361836,11.262123,11.162411,11.062697,10.337513,9.612328,8.887142,8.161958,7.4367723,6.8620634,6.2873545,5.712645,5.137936,4.5632267,4.6375585,4.7118897,4.788034,4.8623657,4.936697,4.7753434,4.612177,4.4508233,4.2876563,4.12449,3.6005437,3.0747845,2.5508385,2.0250793,1.49932,2.663242,3.825351,4.98746,6.149569,7.311678,6.550234,5.7869763,5.0255322,4.262275,3.5008307,4.6629395,5.825049,6.987158,8.149267,9.313189,10.625773,11.938358,13.250943,14.561715,15.8743,15.861609,15.850732,15.838041,15.825351,15.812659,16.162561,16.512463,16.862366,17.212267,17.562168,16.813416,16.062849,15.312282,14.561715,13.812962,13.200181,12.5873995,11.974618,11.361836,10.750868,9.300498,7.850128,6.399758,4.949388,3.5008307,2.962381,2.4257438,1.887294,1.3506571,0.8122072,1.49932,2.1882458,2.8753586,3.5624714,4.249584,3.53709,2.8245957,2.1121013,1.3996071,0.6871128,1.6117238,2.5381477,3.4627585,4.3873696,5.3119802,4.262275,3.2125697,2.1628644,1.1131591,0.06164073,2.4873846,4.9131284,7.3370595,9.762803,12.186734,12.299138,12.413355,12.525759,12.638163,12.750566,10.199727,7.650702,5.0998635,2.5508385,0.0,1.9634385,3.925064,5.8866897,7.850128,9.811753,7.850128,5.8866897,3.925064,1.9616255,0.0,0.099712946,0.19942589,0.2991388,0.40066472,0.50037766,1.5373923,2.5744069,3.6132345,4.650249,5.6872635,4.5632267,3.437377,2.3133402,1.1874905,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.18673515,0.25018883,0.31182957,0.37528324,0.43692398,1.4884423,2.5381477,3.587853,4.6375585,5.6872635,6.249282,6.813113,7.3751316,7.93715,8.499168,7.224656,5.9501433,4.6756306,3.3993049,2.124792,2.03777,1.9507477,1.8619126,1.7748904,1.6878681,1.4503701,1.2128719,0.97537386,0.73787576,0.50037766,0.40066472,0.2991388,0.19942589,0.099712946,0.0,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,1.062396,1.8746033,2.6868105,3.5008307,4.313038,3.6005437,2.8880494,2.175555,1.4630609,0.7505665,1.1747998,1.6008459,2.0250793,2.4493124,2.8753586,2.3133402,1.7495089,1.1874905,0.62547207,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.0870222,0.11240368,0.13778515,0.16316663,0.18673515,0.2374981,0.28826106,0.33721104,0.387974,0.43692398,0.43692398,0.43692398,0.43692398,0.43692398,0.43692398,0.34990177,0.26287958,0.17585737,0.0870222,0.0,0.12509441,0.25018883,0.37528324,0.50037766,0.62547207,0.62547207,0.62547207,0.62547207,0.62547207,0.62547207,0.53663695,0.44961473,0.36259252,0.2755703,0.18673515,0.21211663,0.2374981,0.26287958,0.28826106,0.31182957,1.8256533,3.3376641,4.8496747,6.3616858,7.8755093,8.238102,8.600695,8.963287,9.325879,9.686659,10.962985,12.237497,13.512011,14.788336,16.062849,12.937301,9.811753,6.688019,3.5624714,0.43692398,0.42423326,0.41335547,0.40066472,0.387974,0.37528324,0.2991388,0.22480737,0.15047589,0.07433146,0.0,0.0870222,0.17585737,0.26287958,0.34990177,0.43692398,0.41335547,0.387974,0.36259252,0.33721104,0.31182957,0.31182957,0.31182957,0.31182957,0.31182957,0.31182957,0.3245203,0.33721104,0.34990177,0.36259252,0.37528324,0.51306844,0.6508536,0.7868258,0.9246109,1.062396,0.97537386,0.8883517,0.7995165,0.7124943,0.62547207,0.50037766,0.37528324,0.25018883,0.12509441,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07433146,0.15047589,0.22480737,0.2991388,0.37528324,1.0116332,1.649796,2.2879589,2.9243085,3.5624714,3.0258346,2.4873846,1.9507477,1.4122978,0.87566096,0.89922947,0.9246109,0.9499924,0.97537386,1.0007553,1.2491312,1.49932,1.7495089,1.9996977,2.2498865,3.0367124,3.825351,4.612177,5.4008155,6.187641,6.3254266,6.4632115,6.599184,6.736969,6.874754,6.399758,5.924762,5.4497657,4.974769,4.499773,5.2992897,6.1006193,6.9001355,7.699652,8.499168,8.8508835,9.200785,9.550687,9.900589,10.25049,10.536939,10.825199,11.111648,11.399909,11.6881695,12.449615,13.212872,13.974316,14.737573,15.50083,16.062849,16.624866,17.186886,17.750717,18.312735,16.224201,14.137483,12.050762,9.96223,7.8755093,8.46291,9.050309,9.637709,10.225109,10.812509,11.200482,11.586644,11.974618,12.362592,12.750566,13.337966,13.925365,14.512766,15.100165,15.687565,16.162561,16.637558,17.112555,17.58755,18.062546,16.325727,14.587097,12.850279,11.113461,9.374829,8.299743,7.224656,6.149569,5.0744824,3.9993954,3.4500678,2.9007401,2.3495996,1.8002719,1.2491312,1.7005589,2.1501737,2.5997884,3.049403,3.5008307,3.3757362,3.2506418,3.1255474,3.000453,2.8753586,2.7375734,2.5997884,2.4620032,2.324218,2.1882458,1.8256533,1.4630609,1.1004683,0.73787576,0.37528324,0.3245203,0.2755703,0.22480737,0.17585737,0.12509441,0.16316663,0.19942589,0.2374981,0.2755703,0.31182957,0.28826106,0.26287958,0.2374981,0.21211663,0.18673515,0.40066472,0.33539808,0.27013144,0.20486477,0.13959812,0.07433146,0.23568514,0.39522585,0.55476654,0.71430725,0.87566096,1.8274662,2.7792716,3.73289,4.6846952,5.638314,5.331923,5.027345,4.7227674,4.41819,4.1117992,7.268167,10.422722,13.577277,16.731833,19.888199,17.174194,14.462003,11.74981,9.037619,6.3254266,13.234627,20.14564,27.05484,33.965855,40.875053,37.10772,33.34038,29.573046,25.80571,22.038374,22.529686,23.022812,23.515938,24.00725,24.500376,23.115273,21.73017,20.345066,18.959963,17.57486,17.819609,18.06436,18.310923,18.555672,18.800423,18.637255,18.475903,18.312735,18.149569,17.988214,19.94984,21.913279,23.874905,25.838343,27.799969,29.589363,31.38057,33.169964,34.95936,36.750565,35.731678,34.714607,33.697536,32.68046,31.66158,28.586794,25.512009,22.437225,19.36244,16.287657,16.566853,16.84786,17.127058,17.408066,17.687263,17.995466,18.301857,18.610062,18.918264,19.224655,19.605377,19.984287,20.36501,20.745731,21.12464,20.662334,20.20003,19.737724,19.275417,18.813112,18.252907,17.692701,17.132496,16.57229,16.012085,16.099108,16.187943,16.274965,16.361988,16.450823,16.8533,17.255777,17.658255,18.060734,18.463211,16.630306,14.7974,12.964496,11.13159,9.300498,8.482852,7.665206,6.8475595,6.0299134,5.2122674,6.9055743,8.597069,10.290376,11.98187,13.675177,15.190813,16.704638,18.220274,19.73591,21.249735,20.350506,19.449463,18.550234,17.64919,16.749962,18.055294,19.360628,20.664148,21.96948,23.274813,22.678349,22.08007,21.481794,20.885328,20.287052,20.870825,21.452785,22.034748,22.616709,23.200481,22.408218,21.615953,20.821875,20.02961,19.237347,15.805408,12.373469,8.939718,5.5077806,2.0758421,1.7277533,1.3796645,1.0333886,0.6852999,0.33721104,0.2755703,0.21211663,0.15047589,0.0870222,0.025381476,0.09789998,0.17041849,0.24293698,0.3154555,0.387974,0.49312583,0.5982776,0.7016165,0.80676836,0.9119202,1.649796,2.3876717,3.1255474,3.8616104,4.599486,5.712645,6.825804,7.93715,9.050309,10.161655,11.242181,12.322706,13.403233,14.481945,15.56247,15.54978,15.537089,15.524399,15.511708,15.50083,15.8743,16.249584,16.624866,17.00015,17.375433,16.160748,14.94425,13.729566,12.514881,11.300196,10.674724,10.049252,9.425592,8.80012,8.174648,8.774739,9.374829,9.97492,10.57501,11.175101,11.108022,11.039129,10.97205,10.90497,10.837891,10.424535,10.012992,9.599637,9.188094,8.774739,8.629702,8.484665,8.339628,8.194591,8.049554,7.46578,6.880193,6.294606,5.710832,5.125245,5.527723,5.9302006,6.3326783,6.735156,7.137634,6.399758,5.661882,4.9258194,4.1879435,3.4500678,4.0102735,4.5704784,5.130684,5.6908894,6.249282,6.294606,6.33993,6.3852544,6.430578,6.474089,7.0071006,7.5401115,8.073122,8.604321,9.137331,9.99305,10.846955,11.702674,12.558392,13.412297,13.608097,13.802084,13.997884,14.191871,14.387671,14.922495,15.457319,15.992143,16.526966,17.06179,16.124489,15.187187,14.249886,13.312584,12.375282,11.847711,11.320138,10.792566,10.264994,9.737422,8.859948,7.9824743,7.1050005,6.2275267,5.3500524,4.699199,4.0501585,3.3993049,2.7502642,2.0994108,2.565342,3.0294604,3.4953918,3.9595103,4.4254417,3.7002566,2.9750717,2.2498865,1.5247015,0.7995165,1.550083,2.3006494,3.049403,3.7999697,4.550536,3.7020695,2.855416,2.0069497,1.1602961,0.31182957,2.4402475,4.5668526,6.695271,8.821876,10.950294,10.799818,10.649343,10.500679,10.3502035,10.199727,8.200029,6.200332,4.2006345,2.1991236,0.19942589,1.8202144,3.43919,5.0599785,6.680767,8.299743,6.6571984,5.0146546,3.3721104,1.7295663,0.0870222,0.15410182,0.2229944,0.29007402,0.35715362,0.42423326,1.258196,2.0903459,2.9224956,3.7546456,4.5867953,3.7056956,2.8227828,1.93987,1.0569572,0.17585737,0.14322405,0.11059072,0.07795739,0.045324065,0.012690738,0.09064813,0.16679256,0.24474995,0.32270733,0.40066472,0.39159992,0.38434806,0.3770962,0.36984438,0.36259252,1.3742256,2.3876717,3.3993049,4.4127507,5.424384,5.8359265,6.245656,6.6553855,7.065115,7.474845,6.4178877,5.3609304,4.3021603,3.245203,2.1882458,2.2100015,2.231757,2.2553256,2.277081,2.3006494,1.93987,1.5809034,1.2201238,0.85934424,0.50037766,0.40429065,0.3100166,0.21574254,0.11965553,0.025381476,0.07070554,0.11421664,0.15954071,0.20486477,0.25018883,0.8901646,1.5301404,2.1701162,2.810092,3.4500678,2.8807976,2.3097143,1.7404441,1.1693609,0.6000906,0.94092757,1.2799516,1.6207886,1.9598125,2.3006494,1.8528478,1.405046,0.9572442,0.5094425,0.06164073,0.07070554,0.07795739,0.08520924,0.092461094,0.099712946,0.09064813,0.07977036,0.07070554,0.059827764,0.05076295,0.072518505,0.09427405,0.11784257,0.13959812,0.16316663,0.19942589,0.2374981,0.2755703,0.31182957,0.34990177,0.34990177,0.34990177,0.34990177,0.34990177,0.34990177,0.28282216,0.21574254,0.14684997,0.07977036,0.012690738,0.11421664,0.21755551,0.3208944,0.4224203,0.52575916,0.5293851,0.53482395,0.5402629,0.54570174,0.5493277,0.48043507,0.40972954,0.34083697,0.27013144,0.19942589,0.21755551,0.23568514,0.2520018,0.27013144,0.28826106,1.4956942,2.7031271,3.9105604,5.1179934,6.3254266,6.6155005,6.9055743,7.1956487,7.4857225,7.7757964,9.07569,10.375585,11.675479,12.975373,14.275268,11.490557,8.705847,5.919323,3.1346123,0.34990177,0.73968875,1.1294757,1.5192627,1.9108626,2.3006494,1.8691645,1.4394923,1.0098201,0.58014804,0.15047589,0.19217403,0.23568514,0.27738327,0.3208944,0.36259252,0.37528324,0.387974,0.40066472,0.41335547,0.42423326,0.39522585,0.36440548,0.33539808,0.3045777,0.2755703,0.28282216,0.29007402,0.29732585,0.3045777,0.31182957,0.43511102,0.55839247,0.67986095,0.8031424,0.9246109,0.83940166,0.7541924,0.67079616,0.5855869,0.50037766,0.40066472,0.2991388,0.19942589,0.099712946,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.072518505,0.14503701,0.21755551,0.29007402,0.36259252,0.87022203,1.3778516,1.8854811,2.3931105,2.9007401,2.47832,2.0558996,1.6316663,1.209246,0.7868258,0.7995165,0.8122072,0.824898,0.8375887,0.85027945,1.1403534,1.4304274,1.7205015,2.0105755,2.3006494,3.198066,4.0954823,4.992899,5.8903155,6.787732,6.6898317,6.591932,6.495845,6.397945,6.300045,5.942891,5.5857377,5.2267714,4.8696175,4.512464,5.18326,5.8522434,6.5230393,7.192023,7.8628187,8.205468,8.548119,8.890768,9.231606,9.574255,10.074633,10.57501,11.075388,11.575767,12.07433,12.725184,13.374225,14.025079,14.674119,15.324973,16.109985,16.894999,17.680012,18.465023,19.250036,16.927631,14.6052265,12.282822,9.960417,7.6380115,7.890013,8.1420145,8.39583,8.647832,8.899834,9.63227,10.364707,11.097144,11.829581,12.562017,12.770509,12.977186,13.185677,13.392355,13.600845,14.188245,14.775645,15.363045,15.950445,16.537846,14.927934,13.318023,11.708113,10.098202,8.488291,7.454902,6.4215136,5.389938,4.358362,3.3249733,2.904366,2.4855716,2.0649643,1.6443571,1.2255627,1.5899682,1.9543737,2.3205922,2.6849976,3.049403,2.9224956,2.7955883,2.666868,2.5399606,2.4130533,2.2952106,2.1773682,2.0595255,1.9416829,1.8256533,1.5428312,1.260009,0.97718686,0.69436467,0.41335547,0.36440548,0.31726846,0.27013144,0.2229944,0.17585737,0.19942589,0.22480737,0.25018883,0.2755703,0.2991388,0.3770962,0.4550536,0.533011,0.6091554,0.6871128,0.2991388,0.2574407,0.21574254,0.17223145,0.13053331,0.0870222,0.21936847,0.35171473,0.48587397,0.61822027,0.7505665,1.4920682,2.2353828,2.9768846,3.720199,4.461701,4.4907084,4.517903,4.5450974,4.572292,4.599486,7.059676,9.519867,11.980057,14.440247,16.900436,15.636803,14.37498,13.113158,11.849524,10.587702,15.332225,20.076748,24.823084,29.567606,34.31213,31.703278,29.092611,26.481945,23.87309,21.262424,21.209848,21.157274,21.104698,21.052122,20.999546,19.993351,18.985344,17.977337,16.96933,15.963136,16.115425,16.267714,16.420002,16.57229,16.72458,16.762651,16.800724,16.836983,16.875055,16.913128,19.186583,21.461851,23.73712,26.012386,28.287655,30.292791,32.297928,34.303066,36.3082,38.31334,37.71506,37.116783,36.520317,35.92204,35.325577,31.462152,27.600542,23.73712,19.87551,16.012085,16.421816,16.833357,17.243088,17.652817,18.062546,18.06436,18.067986,18.069798,18.071611,18.075237,18.410635,18.74422,19.079618,19.415016,19.750414,19.025229,18.300045,17.57486,16.849674,16.124489,16.042906,15.95951,15.877926,15.79453,15.712947,16.425442,17.137936,17.85043,18.562923,19.275417,20.129324,20.985043,21.84076,22.694666,23.550385,21.110136,18.66989,16.229641,13.789393,11.349146,10.264994,9.180842,8.094878,7.0107265,5.924762,7.9607186,9.994863,12.03082,14.064963,16.100922,17.130684,18.160446,19.190208,20.219973,21.249735,20.412146,19.574556,18.736969,17.89938,17.06179,18.035353,19.0071,19.980661,20.952408,21.924156,21.40565,20.885328,20.36501,19.844688,19.324368,19.402325,19.480284,19.55824,19.634384,19.712341,18.702522,17.692701,16.682882,15.673061,14.663241,12.222994,9.782746,7.3424983,4.902251,2.4620032,2.030518,1.5972201,1.1657349,0.7324369,0.2991388,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.13234627,0.21574254,0.29732585,0.38072214,0.46230546,0.6091554,0.75781834,0.90466833,1.0533313,1.2001812,2.03777,2.8753586,3.7129474,4.550536,5.388125,6.450521,7.512917,8.575313,9.637709,10.700105,11.722616,12.745127,13.767638,14.790149,15.812659,15.838041,15.861609,15.8869915,15.912373,15.937754,16.213324,16.487082,16.762651,17.038223,17.31198,15.957697,14.603414,13.247317,11.893035,10.536939,10.125396,9.712041,9.300498,8.887142,8.4756,8.937905,9.400211,9.862516,10.324821,10.7871275,10.752681,10.718235,10.681975,10.64753,10.613083,10.51337,10.411844,10.312131,10.212419,10.112705,10.397341,10.681975,10.968424,11.253058,11.537694,10.292189,9.046683,7.802991,6.5574856,5.3119802,6.2801023,7.2482243,8.214534,9.182655,10.150778,9.200785,8.2507925,7.3008003,6.350808,5.4008155,5.3573046,5.315606,5.272095,5.230397,5.186886,6.0407915,6.892884,7.744976,8.597069,9.449161,9.353074,9.255174,9.157274,9.059374,8.963287,9.360326,9.757364,10.154404,10.553255,10.950294,11.352772,11.755249,12.157727,12.5602045,12.962683,13.682428,14.402175,15.121921,15.841667,16.563227,15.437376,14.313339,13.1874895,12.06164,10.937603,10.49524,10.052877,9.610515,9.168152,8.725789,8.419398,8.1148205,7.8102427,7.5056653,7.1992745,6.43783,5.674573,4.9131284,4.1498713,3.386614,3.6295512,3.872488,4.115425,4.358362,4.599486,3.8616104,3.1255474,2.3876717,1.649796,0.9119202,1.4866294,2.0631514,2.6378605,3.2125697,3.787279,3.141864,2.4982624,1.8528478,1.2074331,0.5620184,2.3931105,4.2223897,6.051669,7.8827615,9.712041,9.300498,8.887142,8.4756,8.062244,7.650702,6.200332,4.749962,3.299592,1.8492218,0.40066472,1.6769904,2.955129,4.233268,5.5095935,6.787732,5.464269,4.1426196,2.819157,1.4975071,0.17585737,0.21030366,0.24474995,0.27919623,0.3154555,0.34990177,0.97718686,1.6044719,2.231757,2.8608549,3.48814,2.8481643,2.2081885,1.5682126,0.92823684,0.28826106,0.23568514,0.18310922,0.13053331,0.07795739,0.025381476,0.15591478,0.28463513,0.41516843,0.54570174,0.6744221,0.5982776,0.52032024,0.44236287,0.36440548,0.28826106,1.261822,2.2371957,3.2125697,4.1879435,5.163317,5.4207582,5.678199,5.9356394,6.19308,6.450521,5.6093063,4.7699046,3.930503,3.0892882,2.2498865,2.382233,2.514579,2.6469254,2.7792716,2.911618,2.42937,1.9471219,1.4648738,0.9826257,0.50037766,0.40972954,0.3208944,0.23024625,0.13959812,0.05076295,0.09064813,0.13053331,0.17041849,0.21030366,0.25018883,0.7179332,1.1856775,1.651609,2.1193533,2.5870976,2.1592383,1.7331922,1.305333,0.8774739,0.44961473,0.70524246,0.96087015,1.214685,1.4703126,1.7241274,1.3923552,1.0605831,0.726998,0.39522585,0.06164073,0.065266654,0.06707962,0.07070554,0.072518505,0.07433146,0.06707962,0.059827764,0.052575916,0.045324065,0.038072214,0.058014803,0.07795739,0.09789998,0.11784257,0.13778515,0.16316663,0.18673515,0.21211663,0.2374981,0.26287958,0.26287958,0.26287958,0.26287958,0.26287958,0.26287958,0.21574254,0.16679256,0.11965553,0.072518505,0.025381476,0.10515183,0.18492219,0.26469254,0.3444629,0.42423326,0.43511102,0.44417584,0.4550536,0.46411842,0.4749962,0.4224203,0.36984438,0.31726846,0.26469254,0.21211663,0.2229944,0.23205921,0.24293698,0.2520018,0.26287958,1.1657349,2.0667772,2.9696326,3.872488,4.7753434,4.992899,5.2104545,5.42801,5.6455655,5.863121,7.1883965,8.511859,9.837135,11.162411,12.487686,10.042,7.5981264,5.1524396,2.7067533,0.26287958,1.0551442,1.8474089,2.6396735,3.4319382,4.2242026,3.43919,2.6541772,1.8691645,1.0841516,0.2991388,0.29732585,0.2955129,0.291887,0.29007402,0.28826106,0.33721104,0.387974,0.43692398,0.48768693,0.53663695,0.47680917,0.4169814,0.35715362,0.29732585,0.2374981,0.23931105,0.24293698,0.24474995,0.24837588,0.25018883,0.35715362,0.46411842,0.5728962,0.67986095,0.7868258,0.70524246,0.62184614,0.5402629,0.45686656,0.37528324,0.2991388,0.22480737,0.15047589,0.07433146,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07070554,0.13959812,0.21030366,0.27919623,0.34990177,0.726998,1.1040943,1.4830034,1.8600996,2.2371957,1.9308052,1.6226015,1.3143979,1.0080072,0.69980353,0.69980353,0.69980353,0.69980353,0.69980353,0.69980353,1.0297627,1.3597219,1.6896812,2.0196402,2.3495996,3.3576066,4.365614,5.371808,6.379815,7.3878226,7.0542374,6.722465,6.390693,6.057108,5.7253356,5.484212,5.2449007,5.0055895,4.764466,4.5251546,5.0654173,5.6056805,6.14413,6.684393,7.224656,7.560054,7.895452,8.23085,8.564435,8.899834,9.612328,10.324821,11.037316,11.74981,12.462305,13.000754,13.537392,14.075842,14.612478,15.149116,16.157122,17.16513,18.173138,19.17933,20.187338,17.629248,15.072971,12.514881,9.956791,7.400513,7.317117,7.2355337,7.1521373,7.0705543,6.987158,8.06587,9.142771,10.21967,11.29657,12.375282,12.203052,12.03082,11.856775,11.684544,11.512312,12.212116,12.91192,13.611723,14.313339,15.013144,13.53014,12.047136,10.564133,9.082943,7.5999393,6.6100616,5.620184,4.6303062,3.6404288,2.6505513,2.3604772,2.0704033,1.7803292,1.4902552,1.2001812,1.4793775,1.7603867,2.039583,2.3205922,2.5997884,2.469255,2.3405347,2.2100015,2.079468,1.9507477,1.8528478,1.7549478,1.6570477,1.5591478,1.4630609,1.260009,1.0569572,0.8557183,0.6526665,0.44961473,0.40429065,0.36077955,0.3154555,0.27013144,0.22480737,0.2374981,0.25018883,0.26287958,0.2755703,0.28826106,0.46774435,0.64722764,0.82671094,1.0080072,1.1874905,0.19942589,0.1794833,0.15954071,0.13959812,0.11965553,0.099712946,0.20486477,0.3100166,0.41516843,0.52032024,0.62547207,1.1566701,1.6896812,2.222692,2.7557032,3.2869012,3.6476808,4.006647,4.367427,4.7282066,5.087173,6.8529987,8.617011,10.382836,12.14685,13.912675,14.09941,14.287958,14.474693,14.663241,14.849977,17.429823,20.009668,22.589514,25.16936,27.749205,26.297022,24.84484,23.392656,21.940474,20.48829,19.890013,19.291735,18.69527,18.096992,17.500528,16.869617,16.240519,15.609608,14.98051,14.349599,14.409427,14.4692545,14.529082,14.590723,14.650551,14.888049,15.125546,15.363045,15.600543,15.838041,18.425138,21.012236,23.599335,26.188244,28.775343,30.994408,33.215286,35.434353,37.65523,39.8743,39.69844,39.52077,39.3431,39.165432,38.98776,34.337513,29.687262,25.037014,20.386765,15.738328,16.276777,16.817041,17.357304,17.897566,18.43783,18.135065,17.8323,17.529535,17.22677,16.92582,17.214079,17.504154,17.794228,18.084301,18.374376,17.388124,16.400059,15.411995,14.425743,13.437678,13.832905,14.22813,14.623356,15.016769,15.411995,16.749962,18.087927,19.425894,20.762047,22.100014,23.40716,24.714306,26.023266,27.33041,28.637556,25.589968,22.542377,19.494787,16.447197,13.399607,12.047136,10.694666,9.342196,7.989726,6.637256,9.015862,11.392657,13.769451,16.148058,18.52485,19.070553,19.614443,20.160145,20.705845,21.249735,20.4756,19.699652,18.925516,18.149569,17.375433,18.01541,18.655384,19.29536,19.935337,20.575312,20.13295,19.690586,19.248224,18.80586,18.361685,17.935638,17.50778,17.07992,16.652061,16.224201,14.996826,13.769451,12.542075,11.314699,10.087324,8.640579,7.192023,5.7452784,4.2967215,2.8499773,2.333283,1.8147756,1.2980812,0.7795739,0.26287958,0.22480737,0.18673515,0.15047589,0.11240368,0.07433146,0.16679256,0.25925365,0.35171473,0.44417584,0.53663695,0.726998,0.91735905,1.1077201,1.2980812,1.4866294,2.4257438,3.3630457,4.3003473,5.237649,6.1749506,7.1883965,8.200029,9.211663,10.225109,11.236742,12.203052,13.167547,14.132043,15.098352,16.062849,16.124489,16.187943,16.249584,16.313038,16.374678,16.550535,16.72458,16.900436,17.074482,17.25034,15.754644,14.260764,12.76507,11.269376,9.775495,9.574255,9.374829,9.175404,8.974165,8.774739,9.099259,9.425592,9.750113,10.074633,10.399154,10.397341,10.395528,10.391902,10.390089,10.388275,10.600392,10.812509,11.024626,11.236742,11.450671,12.164979,12.879286,13.595407,14.309713,15.025834,13.12041,11.214987,9.309563,7.404139,5.5005283,7.0324817,8.564435,10.098202,11.630155,13.162108,11.999999,10.837891,9.675781,8.511859,7.3497505,6.7043357,6.060734,5.4153194,4.7699046,4.12449,5.7851634,7.4458375,9.104698,10.765372,12.4242325,11.697234,10.970237,10.243238,9.514427,8.78743,8.727602,8.667774,8.607946,8.548119,8.488291,9.097446,9.706602,10.31757,10.926725,11.537694,12.442362,13.347031,14.2516985,15.15818,16.062849,14.750263,13.437678,12.125093,10.812509,9.499924,9.142771,8.785617,8.42665,8.069496,7.7123427,7.9806614,8.247167,8.515485,8.781991,9.050309,8.174648,7.3008003,6.4251394,5.5494785,4.6756306,4.695573,4.7155156,4.7354584,4.7554007,4.7753434,4.024777,3.2742105,2.525457,1.7748904,1.0243238,1.4249886,1.8256533,2.2245052,2.6251698,3.0258346,2.5816586,2.1392958,1.696933,1.2545701,0.8122072,2.3459735,3.877927,5.40988,6.9418335,8.4756,7.799365,7.124943,6.450521,5.774286,5.0998635,4.2006345,3.299592,2.4003625,1.49932,0.6000906,1.5355793,2.469255,3.4047437,4.3402324,5.275721,4.273153,3.2705846,2.268016,1.2654479,0.26287958,0.26469254,0.26831847,0.27013144,0.27194437,0.2755703,0.6979906,1.1204109,1.5428312,1.9652514,2.3876717,1.9906329,1.5917811,1.1947423,0.79770356,0.40066472,0.32814622,0.25562772,0.18310922,0.11059072,0.038072214,0.21936847,0.40247768,0.5855869,0.7668832,0.9499924,0.8031424,0.6544795,0.5076295,0.36077955,0.21211663,1.1494182,2.08672,3.0258346,3.9631362,4.900438,5.0055895,5.1107416,5.2140803,5.319232,5.424384,4.802538,4.1806917,3.5570326,2.9351864,2.3133402,2.5544643,2.7974012,3.0403383,3.2832751,3.5243993,2.9206827,2.3151531,1.7096237,1.1040943,0.50037766,0.41516843,0.32995918,0.24474995,0.15954071,0.07433146,0.11059072,0.14503701,0.1794833,0.21574254,0.25018883,0.54570174,0.83940166,1.1349145,1.4304274,1.7241274,1.4394923,1.1548572,0.87022203,0.5855869,0.2991388,0.46955732,0.6399758,0.8103943,0.9808127,1.1494182,0.9318628,0.71430725,0.49675176,0.27919623,0.06164073,0.059827764,0.058014803,0.054388877,0.052575916,0.05076295,0.045324065,0.03988518,0.034446288,0.030820364,0.025381476,0.04169814,0.059827764,0.07795739,0.09427405,0.11240368,0.12509441,0.13778515,0.15047589,0.16316663,0.17585737,0.17585737,0.17585737,0.17585737,0.17585737,0.17585737,0.14684997,0.11965553,0.092461094,0.065266654,0.038072214,0.09427405,0.15228885,0.21030366,0.26831847,0.3245203,0.34083697,0.35534066,0.36984438,0.38434806,0.40066472,0.36440548,0.32995918,0.2955129,0.25925365,0.22480737,0.22662032,0.23024625,0.23205921,0.23568514,0.2374981,0.83577573,1.4322405,2.030518,2.6269827,3.2252605,3.3702974,3.5153344,3.6603715,3.8054085,3.9504454,5.2992897,6.6499467,8.000604,9.349448,10.700105,8.595256,6.490406,4.3855567,2.280707,0.17585737,1.3705997,2.565342,3.7600844,4.954827,6.149569,5.009216,3.870675,2.7303216,1.5899682,0.44961473,0.40247768,0.35534066,0.30820364,0.25925365,0.21211663,0.2991388,0.387974,0.4749962,0.5620184,0.6508536,0.56020546,0.46955732,0.38072214,0.29007402,0.19942589,0.19761293,0.19579996,0.19217403,0.19036107,0.18673515,0.27919623,0.37165734,0.46411842,0.55839247,0.6508536,0.56927025,0.4894999,0.40972954,0.32995918,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06707962,0.13415924,0.2030518,0.27013144,0.33721104,0.5855869,0.8321498,1.0805258,1.3270886,1.5754645,1.3832904,1.1893034,0.99712944,0.80495536,0.61278135,0.6000906,0.5873999,0.5747091,0.5620184,0.5493277,0.91917205,1.2908293,1.6606737,2.030518,2.4003625,3.5171473,4.6357455,5.75253,6.869315,7.987913,7.420456,6.8529987,6.285541,5.718084,5.1506267,5.027345,4.9058766,4.782595,4.6593137,4.537845,4.947575,5.3573046,5.767034,6.1767635,6.588306,6.9146395,7.2427855,7.569119,7.897265,8.225411,9.1500225,10.074633,10.999244,11.925668,12.850279,13.274512,13.700559,14.124791,14.5508375,14.975071,16.20426,17.43526,18.66445,19.89545,21.12464,18.332678,15.540715,12.74694,9.954978,7.1630154,6.7442207,6.3272395,5.910258,5.4932766,5.0744824,6.497658,7.9190207,9.342196,10.765372,12.186734,11.635593,11.082641,10.529687,9.976733,9.425592,10.2378,11.050007,11.862214,12.674421,13.486629,12.132345,10.778063,9.421967,8.067683,6.7115874,5.765221,4.8170414,3.870675,2.9224956,1.9743162,1.8147756,1.6552348,1.4956942,1.3343405,1.1747998,1.3705997,1.5645868,1.7603867,1.9543737,2.1501737,2.0178273,1.8854811,1.7531348,1.6207886,1.4866294,1.4104849,1.3325275,1.2545701,1.1766127,1.1004683,0.97718686,0.8557183,0.7324369,0.6091554,0.48768693,0.44417584,0.40247768,0.36077955,0.31726846,0.2755703,0.2755703,0.2755703,0.2755703,0.2755703,0.2755703,0.55839247,0.83940166,1.1222239,1.405046,1.6878681,0.099712946,0.10333887,0.10515183,0.10696479,0.11059072,0.11240368,0.19036107,0.26831847,0.3444629,0.4224203,0.50037766,0.823085,1.1457924,1.4666867,1.789394,2.1121013,2.8046532,3.4972048,4.1897564,4.882308,5.57486,6.644508,7.7141557,8.785617,9.855265,10.924912,12.562017,14.199123,15.838041,17.475147,19.112251,19.52742,19.942589,20.357758,20.772924,21.188093,20.89258,20.597069,20.301556,20.007854,19.712341,18.570175,17.428009,16.284029,15.141864,13.999697,13.747695,13.495693,13.2418785,12.989877,12.737875,12.705242,12.672608,12.639976,12.607342,12.574709,13.011633,13.45037,13.887294,14.324218,14.762955,17.661882,20.562622,23.463362,26.36229,29.26303,31.697838,34.132645,36.567455,39.002266,41.437073,41.680008,41.922947,42.165882,42.40701,42.649944,37.21287,31.775795,26.336908,20.899832,15.462758,16.13174,16.802538,17.473333,18.142317,18.813112,18.20577,17.596615,16.989273,16.38193,15.774588,16.019337,16.264088,16.51065,16.7554,17.00015,15.749206,14.500074,13.24913,11.999999,10.749055,11.622903,12.494938,13.366973,14.240821,15.112856,17.074482,19.03792,20.999546,22.962984,24.92461,26.684996,28.445383,30.20577,31.964344,33.72473,30.069798,26.414865,22.759932,19.105,15.4500675,13.829279,12.210303,10.589515,8.970539,7.3497505,10.069194,12.790451,15.509895,18.22934,20.950596,21.010424,21.070251,21.13008,21.189907,21.249735,20.537241,19.824745,19.112251,18.399757,17.687263,17.995466,18.301857,18.610062,18.918264,19.224655,18.86025,18.495844,18.129625,17.76522,17.400814,16.467138,15.535276,14.601601,13.669738,12.737875,11.292944,9.848013,8.403082,6.9581504,5.5132194,5.0581656,4.603112,4.1480584,3.6930048,3.2379513,2.6342347,2.032331,1.4304274,0.82671094,0.22480737,0.19942589,0.17585737,0.15047589,0.12509441,0.099712946,0.2030518,0.3045777,0.40791658,0.5094425,0.61278135,0.8448406,1.0768998,1.310772,1.5428312,1.7748904,2.811905,3.8507326,4.8877473,5.924762,6.9617763,7.9244595,8.887142,9.849826,10.812509,11.775192,12.681673,13.589968,14.498261,15.404743,16.313038,16.41275,16.512463,16.612177,16.71189,16.813416,16.887747,16.962078,17.038223,17.112555,17.186886,15.553406,13.918114,12.282822,10.64753,9.012237,9.024928,9.037619,9.050309,9.063,9.07569,9.262425,9.449161,9.637709,9.824444,10.012992,10.042,10.07282,10.101828,10.1326475,10.161655,10.687414,11.213174,11.73712,12.262879,12.786825,13.932617,15.076597,16.22239,17.368181,18.512161,15.946819,13.383289,10.817947,8.252605,5.6872635,7.7848616,9.882459,11.980057,14.077655,16.175253,14.799213,13.424988,12.050762,10.674724,9.300498,8.05318,6.8058615,5.5567303,4.309412,3.0620937,5.529536,7.996978,10.46442,12.931862,15.399304,14.043208,12.685299,11.327391,9.969481,8.613385,8.094878,7.5781837,7.059676,6.542982,6.0244746,6.8421206,7.6597667,8.477413,9.295059,10.112705,11.202296,12.291886,13.383289,14.47288,15.56247,14.06315,12.562017,11.062697,9.561564,8.062244,7.7903004,7.518356,7.2445984,6.972654,6.70071,7.5401115,8.379513,9.220728,10.060129,10.899531,9.91328,8.925215,7.93715,6.9508986,5.962834,5.7597823,5.5567303,5.3554916,5.1524396,4.949388,4.1879435,3.4246864,2.663242,1.8999848,1.1367276,1.3633479,1.5881553,1.8129625,2.03777,2.2625773,2.0232663,1.7821422,1.5428312,1.3017071,1.062396,2.2970235,3.531651,4.7680917,6.002719,7.2373466,6.300045,5.3627434,4.4254417,3.48814,2.5508385,2.1991236,1.8492218,1.49932,1.1494182,0.7995165,1.3923552,1.9851941,2.5780327,3.1708715,3.7618973,3.0802233,2.3967366,1.7150626,1.0333886,0.34990177,0.3208944,0.29007402,0.25925365,0.23024625,0.19942589,0.4169814,0.6345369,0.8520924,1.0696479,1.2872034,1.1331016,0.97718686,0.823085,0.6671702,0.51306844,0.42060733,0.32814622,0.23568514,0.14322405,0.05076295,0.28463513,0.52032024,0.7541924,0.9898776,1.2255627,1.0080072,0.7904517,0.5728962,0.35534066,0.13778515,1.0370146,1.938057,2.8372865,3.738329,4.6375585,4.590421,4.5432844,4.494334,4.4471974,4.40006,3.9957695,3.589666,3.1853752,2.7792716,2.374981,2.7266958,3.0802233,3.4319382,3.785466,4.137181,3.4101827,2.6831846,1.9543737,1.2273756,0.50037766,0.42060733,0.34083697,0.25925365,0.1794833,0.099712946,0.13053331,0.15954071,0.19036107,0.21936847,0.25018883,0.37165734,0.4949388,0.61822027,0.73968875,0.8629702,0.7197462,0.57833505,0.43511102,0.291887,0.15047589,0.23568514,0.3208944,0.40429065,0.4894999,0.5747091,0.47318324,0.36984438,0.26831847,0.16497959,0.06164073,0.054388877,0.047137026,0.03988518,0.032633327,0.025381476,0.02175555,0.01994259,0.018129626,0.014503701,0.012690738,0.027194439,0.04169814,0.058014803,0.072518505,0.0870222,0.0870222,0.0870222,0.0870222,0.0870222,0.0870222,0.0870222,0.0870222,0.0870222,0.0870222,0.0870222,0.07977036,0.072518505,0.065266654,0.058014803,0.05076295,0.08520924,0.11965553,0.15410182,0.19036107,0.22480737,0.24474995,0.26469254,0.28463513,0.3045777,0.3245203,0.30820364,0.29007402,0.27194437,0.25562772,0.2374981,0.23205921,0.22662032,0.2229944,0.21755551,0.21211663,0.5058166,0.79770356,1.0895905,1.3832904,1.6751775,1.7476959,1.8202144,1.892733,1.9652514,2.03777,3.4119956,4.788034,6.16226,7.5382986,8.912524,7.1466985,5.382686,3.6168604,1.8528478,0.0870222,1.6842422,3.2832751,4.880495,6.4777155,8.074935,6.5792413,5.08536,3.589666,2.0957847,0.6000906,0.5076295,0.41516843,0.32270733,0.23024625,0.13778515,0.26287958,0.387974,0.51306844,0.63816285,0.76325727,0.6417888,0.52213323,0.40247768,0.28282216,0.16316663,0.15410182,0.14684997,0.13959812,0.13234627,0.12509441,0.2030518,0.27919623,0.35715362,0.43511102,0.51306844,0.43511102,0.35715362,0.27919623,0.2030518,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.065266654,0.13053331,0.19579996,0.25925365,0.3245203,0.44236287,0.56020546,0.678048,0.79589057,0.9119202,0.83577573,0.75781834,0.67986095,0.60190356,0.52575916,0.50037766,0.4749962,0.44961473,0.42423326,0.40066472,0.8103943,1.2201238,1.6298534,2.039583,2.4493124,3.6766882,4.9040637,6.1332526,7.360628,8.588004,7.7848616,6.981719,6.1803894,5.377247,4.574105,4.5704784,4.5650396,4.559601,4.554162,4.550536,4.8297324,5.1107416,5.389938,5.669134,5.9501433,6.2692246,6.590119,6.9092,7.230095,7.549176,8.6877165,9.824444,10.962985,12.099712,13.238253,13.550082,13.861912,14.175554,14.487384,14.799213,16.25321,17.705393,19.157576,20.609758,22.061941,19.034294,16.00846,12.980812,9.953164,6.925517,6.1731377,5.4207582,4.666566,3.9141862,3.1618068,4.9294453,6.697084,8.464723,10.232361,11.999999,11.068136,10.13446,9.202598,8.270736,7.3370595,8.26167,9.188094,10.112705,11.037316,11.961927,10.734551,9.507175,8.2798,7.0524244,5.825049,4.9203806,4.0157123,3.1092308,2.2045624,1.2998942,1.2708868,1.2400664,1.209246,1.1802386,1.1494182,1.260009,1.3705997,1.4793775,1.5899682,1.7005589,1.5645868,1.4304274,1.2944553,1.1602961,1.0243238,0.968122,0.9101072,0.8520924,0.79589057,0.73787576,0.69436467,0.6526665,0.6091554,0.56745726,0.52575916,0.48587397,0.44417584,0.40429065,0.36440548,0.3245203,0.31182957,0.2991388,0.28826106,0.2755703,0.26287958,0.64722764,1.0333886,1.4177368,1.8020848,2.1882458,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.17585737,0.22480737,0.2755703,0.3245203,0.37528324,0.48768693,0.6000906,0.7124943,0.824898,0.93730164,1.9616255,2.9877625,4.0120864,5.038223,6.0625467,6.43783,6.813113,7.1883965,7.5618668,7.93715,11.024626,14.112101,17.199575,20.287052,23.374527,21.625017,19.87551,18.124187,16.374678,14.625169,15.488139,16.349297,17.212267,18.075237,18.938208,17.25034,15.56247,13.874602,12.186734,10.500679,10.625773,10.750868,10.874149,10.999244,11.124338,10.999244,10.874149,10.750868,10.625773,10.500679,11.137029,11.775192,12.413355,13.049705,13.687867,16.900436,20.113007,23.325577,26.538147,29.750715,32.399456,35.050007,37.700558,40.349297,42.999847,43.66339,44.325123,44.986855,45.6504,46.31213,40.08823,33.862514,27.6368,21.4129,15.187187,15.986704,16.788034,17.58755,18.387066,19.188396,18.274662,17.362743,16.450823,15.537089,14.625169,14.824595,15.025834,15.22526,15.4246855,15.624111,14.112101,12.60009,11.088079,9.574255,8.062244,9.412902,10.761745,12.112403,13.46306,14.811904,17.400814,19.987913,22.57501,25.162107,27.749205,29.962833,32.17465,34.388275,36.60009,38.8119,34.54963,30.287354,26.025078,21.762802,17.500528,15.613234,13.72594,11.836833,9.949538,8.062244,11.124338,14.188245,17.25034,20.312433,23.374527,22.950293,22.524246,22.100014,21.675781,21.249735,20.600695,19.94984,19.3008,18.649946,18.000906,17.975525,17.950142,17.92476,17.89938,17.87581,17.58755,17.29929,17.01284,16.72458,16.438131,15.000452,13.562773,12.125093,10.687414,9.249735,7.5872483,5.924762,4.262275,2.5997884,0.93730164,1.4757515,2.0123885,2.5508385,3.0874753,3.6241121,2.9369993,2.2498865,1.5627737,0.87566096,0.18673515,0.17585737,0.16316663,0.15047589,0.13778515,0.12509441,0.2374981,0.34990177,0.46230546,0.5747091,0.6871128,0.96268314,1.2382535,1.5120108,1.7875811,2.0631514,3.199879,4.3366065,5.475147,6.6118746,7.750415,8.662335,9.574255,10.487988,11.399909,12.311829,13.162108,14.012388,14.862667,15.712947,16.563227,16.699198,16.836983,16.97477,17.112555,17.25034,17.224958,17.199575,17.174194,17.150625,17.125244,15.350354,13.575464,11.800573,10.025683,8.2507925,8.4756,8.700407,8.925215,9.1500225,9.374829,9.425592,9.474543,9.525306,9.574255,9.625018,9.686659,9.750113,9.811753,9.875207,9.936848,10.774437,11.612025,12.449615,13.287203,14.124791,15.700256,17.27572,18.849373,20.424837,22.000301,18.77504,15.54978,12.32452,9.099259,5.8758116,8.537241,11.200482,13.861912,16.525154,19.188396,17.60024,16.012085,14.425743,12.837588,11.249433,9.400211,7.549176,5.6999545,3.8507326,1.9996977,5.275721,8.549932,11.825955,15.100165,18.374376,16.38737,14.400362,12.411542,10.424535,8.437528,7.462154,6.48678,5.5132194,4.537845,3.5624714,4.5867953,5.612932,6.637256,7.663393,8.6877165,9.96223,11.236742,12.513068,13.7875805,15.062093,13.374225,11.6881695,10.000301,8.312433,6.624565,6.43783,6.249282,6.0625467,5.8758116,5.6872635,7.0995617,8.511859,9.924157,11.338268,12.750566,11.650098,10.549629,9.449161,8.350506,7.250037,6.825804,6.399758,5.975525,5.5494785,5.125245,4.349297,3.5751622,2.7992141,2.0250793,1.2491312,1.2998942,1.3506571,1.3996071,1.4503701,1.49932,1.4630609,1.4249886,1.3869164,1.3506571,1.3125849,2.2498865,3.1871881,4.12449,5.0617914,6.000906,4.800725,3.6005437,2.4003625,1.2001812,0.0,0.19942589,0.40066472,0.6000906,0.7995165,1.0007553,1.2491312,1.49932,1.7495089,1.9996977,2.2498865,1.887294,1.5247015,1.162109,0.7995165,0.43692398,0.37528324,0.31182957,0.25018883,0.18673515,0.12509441,0.13778515,0.15047589,0.16316663,0.17585737,0.18673515,0.2755703,0.36259252,0.44961473,0.53663695,0.62547207,0.51306844,0.40066472,0.28826106,0.17585737,0.06164073,0.34990177,0.63816285,0.9246109,1.2128719,1.49932,1.2128719,0.9246109,0.63816285,0.34990177,0.06164073,0.9246109,1.7875811,2.6505513,3.5117085,4.3746786,4.175253,3.975827,3.774588,3.5751622,3.3757362,3.1871881,3.000453,2.811905,2.6251698,2.4366217,2.9007401,3.3630457,3.825351,4.2876563,4.749962,3.8996825,3.049403,2.1991236,1.3506571,0.50037766,0.42423326,0.34990177,0.2755703,0.19942589,0.12509441,0.15047589,0.17585737,0.19942589,0.22480737,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.15047589,0.17585737,0.19942589,0.22480737,0.25018883,0.25018883,0.25018883,0.25018883,0.25018883,0.25018883,0.2374981,0.22480737,0.21211663,0.19942589,0.18673515,0.17585737,0.16316663,0.15047589,0.13778515,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,1.5247015,2.9243085,4.325729,5.7253356,7.124943,5.6999545,4.274966,2.8499773,1.4249886,0.0,1.9996977,3.9993954,6.000906,8.000604,10.000301,8.149267,6.300045,4.4508233,2.5997884,0.7505665,0.61278135,0.4749962,0.33721104,0.19942589,0.06164073,0.22480737,0.387974,0.5493277,0.7124943,0.87566096,0.72518504,0.5747091,0.42423326,0.2755703,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.12509441,0.18673515,0.25018883,0.31182957,0.37528324,0.2991388,0.22480737,0.15047589,0.07433146,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06164073,0.12509441,0.18673515,0.25018883,0.31182957,0.2991388,0.28826106,0.2755703,0.26287958,0.25018883,0.28826106,0.3245203,0.36259252,0.40066472,0.43692398,0.40066472,0.36259252,0.3245203,0.28826106,0.25018883,0.69980353,1.1494182,1.6008459,2.0504606,2.5000753,3.8380418,5.1741953,6.5121617,7.850128,9.188094,8.149267,7.112252,6.0752378,5.038223,3.9993954,4.1117992,4.2242026,4.3366065,4.4508233,4.5632267,4.7118897,4.8623657,5.0128417,5.163317,5.3119802,5.6256227,5.9374523,6.249282,6.5629244,6.874754,8.225411,9.574255,10.924912,12.27557,13.6244135,13.825653,14.025079,14.224504,14.425743,14.625169,16.300346,17.975525,19.650702,21.324066,22.999243,19.737724,16.474392,13.212872,9.949538,6.688019,5.600241,4.512464,3.4246864,2.3369088,1.2491312,3.3630457,5.475147,7.5872483,9.699349,11.813264,10.500679,9.188094,7.8755093,6.5629244,5.2503395,6.2873545,7.324369,8.363196,9.400211,10.437225,9.336758,8.238102,7.137634,6.037165,4.936697,4.07554,3.2125697,2.3495996,1.4884423,0.62547207,0.72518504,0.824898,0.9246109,1.0243238,1.1258497,1.1494182,1.1747998,1.2001812,1.2255627,1.2491312,1.1131591,0.97537386,0.8375887,0.69980353,0.5620184,0.52575916,0.48768693,0.44961473,0.41335547,0.37528324,0.41335547,0.44961473,0.48768693,0.52575916,0.5620184,0.52575916,0.48768693,0.44961473,0.41335547,0.37528324,0.34990177,0.3245203,0.2991388,0.2755703,0.25018883,0.73787576,1.2255627,1.7132497,2.1991236,2.6868105,0.06164073,0.08520924,0.10696479,0.13053331,0.15228885,0.17585737,0.31726846,0.4604925,0.60190356,0.7451276,0.8883517,1.067835,1.2473183,1.4268016,1.6080978,1.7875811,2.9206827,4.0519714,5.185073,6.3181744,7.4494634,7.763106,8.074935,8.386765,8.700407,9.012237,11.900287,14.786523,17.674572,20.562622,23.45067,21.880646,20.31062,18.740595,17.170568,15.600543,15.917811,16.23508,16.55235,16.869617,17.186886,15.9431925,14.697688,13.452183,12.206677,10.962985,11.062697,11.162411,11.262123,11.361836,11.463363,11.329204,11.1968565,11.06451,10.932164,10.799818,12.058014,13.314397,14.572594,15.83079,17.087172,20.279799,23.472427,26.665054,29.857681,33.05031,35.369087,37.68968,40.010273,42.330864,44.649643,45.599636,46.549625,47.49962,48.44961,49.399605,43.667015,37.93443,32.201843,26.469254,20.736666,21.697536,22.656593,23.617464,24.57652,25.537392,23.876717,22.217857,20.557182,18.898321,17.237648,17.692701,18.147755,18.60281,19.057863,19.512917,17.870373,16.227829,14.585284,12.9427395,11.300196,11.700861,12.099712,12.500377,12.899229,13.299893,15.140051,16.980207,18.820364,20.660522,22.500679,24.235683,25.97069,27.705694,29.440699,31.175705,29.368181,27.560658,25.753134,23.94561,22.138086,20.939718,19.743162,18.544794,17.34824,16.14987,17.32467,18.49947,19.67427,20.850883,22.025682,22.18341,22.339325,22.497053,22.654781,22.812508,22.49524,22.17797,21.860703,21.541622,21.224354,21.40021,21.574255,21.750113,21.924156,22.100014,20.838192,19.574556,18.312735,17.0491,15.787278,14.512766,13.238253,11.961927,10.687414,9.412902,7.752228,6.093367,4.4326935,2.7720199,1.1131591,2.0649643,3.0167696,3.9703882,4.9221935,5.8758116,4.9294453,3.9848917,3.0403383,2.0957847,1.1494182,0.95180535,0.7541924,0.55839247,0.36077955,0.16316663,0.29732585,0.43329805,0.56745726,0.7016165,0.8375887,1.2273756,1.6171626,2.0069497,2.3967366,2.7883365,3.9341288,5.081734,6.2293396,7.3769445,8.52455,9.599637,10.674724,11.74981,12.824898,13.899984,14.376793,14.855415,15.332225,15.810846,16.287657,16.439945,16.592234,16.744522,16.89681,17.0491,16.900436,16.749962,16.599485,16.450823,16.300346,14.646925,12.995316,11.341894,9.690285,8.036863,8.214534,8.392203,8.569874,8.747544,8.925215,8.985043,9.04487,9.104698,9.164526,9.224354,9.3567,9.490859,9.623205,9.755551,9.8878975,10.547816,11.207735,11.867653,12.527572,13.1874895,14.478319,15.767336,17.058165,18.347181,19.63801,17.786976,15.937754,14.0867195,12.237497,10.388275,12.572895,14.757515,16.942135,19.126755,21.313189,19.337059,17.362743,15.386614,13.412297,11.437981,10.045626,8.653271,7.2591023,5.866747,4.4743915,7.2554765,10.034748,12.815832,15.595104,18.374376,16.084604,13.794832,11.50506,9.215289,6.925517,7.0052876,7.0850577,7.1648283,7.2445984,7.324369,8.178274,9.030367,9.882459,10.734551,11.586644,12.944552,14.302462,15.660371,17.01828,18.374376,15.885179,13.394168,10.90497,8.415772,5.924762,5.6872635,5.4497657,5.2122674,4.974769,4.7372713,5.9900284,7.2427855,8.495543,9.7483,10.999244,10.197914,9.394773,8.59163,7.7903004,6.987158,6.9599633,6.932769,6.9055743,6.87838,6.849373,5.710832,4.5704784,3.4301252,2.2897718,1.1494182,1.1802386,1.209246,1.2400664,1.2708868,1.2998942,1.4268016,1.5555218,1.6824293,1.8093367,1.938057,2.7430124,3.5479677,4.3529234,5.1578784,5.962834,4.8315454,3.7020695,2.572594,1.4431182,0.31182957,0.40972954,0.5076295,0.6055295,0.7016165,0.7995165,1.1403534,1.4793775,1.8202144,2.1592383,2.5000753,2.0722163,1.6443571,1.2183108,0.7904517,0.36259252,0.44780177,0.533011,0.61822027,0.7016165,0.7868258,0.76325727,0.73787576,0.7124943,0.6871128,0.66173136,1.2726997,1.8818551,2.4928236,3.101979,3.7129474,3.147303,2.5816586,2.0178273,1.452183,0.8883517,1.5809034,2.2716422,2.9641938,3.6567454,4.349297,3.5117085,2.6741197,1.8383441,1.0007553,0.16316663,1.5700256,2.9768846,4.3855567,5.7924156,7.1992745,6.7532854,6.305484,5.857682,5.40988,4.9620786,4.836984,4.7118897,4.5867953,4.461701,4.3366065,4.537845,4.7372713,4.936697,5.137936,5.337362,4.4381323,3.53709,2.6378605,1.7368182,0.8375887,0.72518504,0.61278135,0.50037766,0.387974,0.2755703,0.25925365,0.24474995,0.23024625,0.21574254,0.19942589,0.17041849,0.13959812,0.11059072,0.07977036,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.018129626,0.034446288,0.052575916,0.07070554,0.0870222,0.07070554,0.052575916,0.034446288,0.018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.054388877,0.11059072,0.16497959,0.21936847,0.2755703,0.23024625,0.18492219,0.13959812,0.09427405,0.05076295,0.059827764,0.07070554,0.07977036,0.09064813,0.099712946,0.12328146,0.14503701,0.16679256,0.19036107,0.21211663,0.21936847,0.22662032,0.23568514,0.24293698,0.25018883,0.23205921,0.21574254,0.19761293,0.1794833,0.16316663,0.15228885,0.14322405,0.13234627,0.12328146,0.11240368,0.11421664,0.11784257,0.11965553,0.12328146,0.12509441,1.3669738,2.610666,3.8525455,5.0944247,6.338117,5.295664,4.25321,3.2107568,2.1683033,1.1258497,3.7256382,6.3254266,8.925215,11.525003,14.124791,11.419851,8.714911,6.009971,3.3050308,0.6000906,0.4949388,0.38978696,0.28463513,0.1794833,0.07433146,0.20667773,0.34083697,0.47318324,0.6055295,0.73787576,0.61459434,0.49312583,0.36984438,0.24837588,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.11240368,0.16316663,0.21211663,0.26287958,0.31182957,0.2520018,0.19217403,0.13234627,0.072518505,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06164073,0.12509441,0.18673515,0.25018883,0.31182957,0.29007402,0.26831847,0.24474995,0.2229944,0.19942589,0.2574407,0.3154555,0.37165734,0.42967212,0.48768693,0.44417584,0.40247768,0.36077955,0.31726846,0.2755703,0.67079616,1.064209,1.4594349,1.8546607,2.2498865,3.4681973,4.6846952,5.903006,7.119504,8.337815,7.453089,6.5683637,5.6818247,4.797099,3.9123733,4.0519714,4.1933823,4.3329806,4.4725785,4.612177,4.8206677,5.027345,5.235836,5.4425135,5.6491914,5.7072062,5.765221,5.823236,5.8794374,5.9374523,7.137634,8.337815,9.537996,10.738177,11.938358,12.119655,12.302764,12.485873,12.66717,12.850279,14.402175,15.955884,17.50778,19.059675,20.613384,17.6365,14.663241,11.6881695,8.713099,5.7380266,4.9983377,4.256836,3.5171473,2.7774587,2.03777,3.6277382,5.217706,6.8076744,8.397643,9.987611,8.917963,7.846502,6.776854,5.7072062,4.6375585,5.520471,6.4033837,7.2844834,8.167397,9.050309,8.129324,7.210152,6.2891674,5.369995,4.4508233,3.7528327,3.054842,2.3568513,1.6606737,0.96268314,1.0025684,1.0424535,1.0823387,1.1222239,1.162109,1.1602961,1.1566701,1.1548572,1.1530442,1.1494182,1.0497054,0.9499924,0.85027945,0.7505665,0.6508536,0.62184614,0.5946517,0.56745726,0.5402629,0.51306844,0.51306844,0.51306844,0.51306844,0.51306844,0.51306844,0.5293851,0.5475147,0.5656443,0.581961,0.6000906,0.6055295,0.6091554,0.61459434,0.6200332,0.62547207,1.1059072,1.5845293,2.0649643,2.5453994,3.0258346,0.12509441,0.14503701,0.16497959,0.18492219,0.20486477,0.22480737,0.4604925,0.69436467,0.9300498,1.1657349,1.3996071,1.647983,1.8945459,2.1429217,2.3894846,2.6378605,3.877927,5.1179934,6.35806,7.5981264,8.838193,9.088382,9.336758,9.5869465,9.837135,10.087324,12.774135,15.462758,18.149569,20.838192,23.525002,22.13446,20.745731,19.355188,17.964645,16.574104,16.347483,16.120863,15.89243,15.66581,15.437376,14.634234,13.832905,13.029762,12.22662,11.42529,11.499621,11.575767,11.650098,11.724429,11.800573,11.6591625,11.519565,11.379966,11.240368,11.10077,12.977186,14.855415,16.731833,18.610062,20.48829,23.659163,26.831846,30.00453,33.177216,36.3499,38.340534,40.329353,42.319984,44.31062,46.29944,47.537693,48.77413,50.012386,51.25064,52.48708,47.24762,42.008156,36.76688,31.52742,26.287958,27.40837,28.526966,29.647377,30.767788,31.888199,29.480585,27.07297,24.665356,22.257742,19.850128,20.560808,21.269676,21.980358,22.689226,23.399908,21.626831,19.855566,18.082489,16.309412,14.538147,13.987006,13.437678,12.888351,12.337211,11.787883,12.879286,13.972503,15.065719,16.157122,17.25034,18.506721,19.764917,21.023113,22.279497,23.537693,24.184921,24.832148,25.479376,26.128416,26.775644,26.268015,25.760386,25.252756,24.745127,24.237497,23.525002,22.812508,22.100014,21.38752,20.675026,21.414715,22.154404,22.895905,23.635593,24.375282,24.389786,24.40429,24.420607,24.43511,24.449614,24.824896,25.20018,25.575462,25.950747,26.324217,24.08702,21.849825,19.612629,17.375433,15.138238,14.025079,12.91192,11.800573,10.687414,9.574255,7.9172077,6.26016,4.603112,2.9442513,1.2872034,2.6541772,4.022964,5.389938,6.7569118,8.125698,6.921891,5.719897,4.517903,3.3140955,2.1121013,1.7295663,1.3470312,0.9644961,0.581961,0.19942589,0.35715362,0.5148814,0.6726091,0.83033687,0.9880646,1.4920682,1.9978848,2.5018883,3.007705,3.5117085,4.670192,5.826862,6.985345,8.1420145,9.300498,10.536939,11.775192,13.013446,14.249886,15.488139,15.593291,15.6966305,15.801782,15.906934,16.012085,16.18069,16.347483,16.514277,16.682882,16.849674,16.574104,16.300346,16.024776,15.749206,15.475449,13.945308,12.415168,10.885027,9.354887,7.8247466,7.95528,8.0858135,8.214534,8.345067,8.4756,8.544493,8.615198,8.685904,8.754796,8.825501,9.026741,9.229793,9.432844,9.635896,9.837135,10.319383,10.801631,11.285692,11.7679405,12.250188,13.254569,14.260764,15.265145,16.269526,17.27572,16.800724,16.325727,15.850732,15.375735,14.90074,16.606737,18.314548,20.022358,21.73017,23.43798,21.07569,18.7134,16.349297,13.987006,11.624716,10.689227,9.755551,8.820063,7.8845744,6.9508986,9.235231,11.519565,13.80571,16.090042,18.374376,15.781839,13.189302,10.596766,8.00423,5.411693,6.546608,7.6833353,8.81825,9.953164,11.088079,11.7679405,12.447801,13.127662,13.807523,14.487384,15.926876,17.368181,18.807674,20.247166,21.686659,18.394318,15.101978,11.809638,8.517298,5.224958,4.936697,4.650249,4.361988,4.07554,3.787279,4.880495,5.9718986,7.065115,8.158332,9.249735,8.745731,8.239915,7.7340984,7.230095,6.7242785,7.0941224,7.46578,7.835624,8.205468,8.575313,7.0705543,5.565795,4.059223,2.5544643,1.0497054,1.0605831,1.0696479,1.0805258,1.0895905,1.1004683,1.3923552,1.6842422,1.9779422,2.269829,2.561716,3.2343252,3.9069343,4.5795436,5.2521524,5.924762,4.8641787,3.8054085,2.7448254,1.6842422,0.62547207,0.6200332,0.61459434,0.6091554,0.6055295,0.6000906,1.0297627,1.4594349,1.8909199,2.3205922,2.7502642,2.2571385,1.7658255,1.2726997,0.7795739,0.28826106,0.52032024,0.7523795,0.98443866,1.2183108,1.4503701,1.3869164,1.3252757,1.261822,1.2001812,1.1367276,2.269829,3.4029307,4.5342193,5.667321,6.8004227,5.7833505,4.764466,3.7473936,2.7303216,1.7132497,2.810092,3.9069343,5.0055895,6.1024323,7.1992745,5.812358,4.4254417,3.0367124,1.649796,0.26287958,2.2154403,4.168001,6.1205616,8.073122,10.025683,9.329506,8.63514,7.9407763,7.2445984,6.550234,6.48678,6.4251394,6.3616858,6.300045,6.2384043,6.1749506,6.11331,6.049856,5.9882154,5.924762,4.974769,4.024777,3.0747845,2.124792,1.1747998,1.0243238,0.87566096,0.72518504,0.5747091,0.42423326,0.36984438,0.3154555,0.25925365,0.20486477,0.15047589,0.13959812,0.13053331,0.11965553,0.11059072,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0,0.0,0.0,0.0,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.09064813,0.06707962,0.045324065,0.02175555,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.11059072,0.21936847,0.32995918,0.4405499,0.5493277,0.44780177,0.3444629,0.24293698,0.13959812,0.038072214,0.045324065,0.052575916,0.059827764,0.06707962,0.07433146,0.09427405,0.11421664,0.13415924,0.15410182,0.17585737,0.19036107,0.20486477,0.21936847,0.23568514,0.25018883,0.22662032,0.20486477,0.18310922,0.15954071,0.13778515,0.13053331,0.12328146,0.11421664,0.10696479,0.099712946,0.10515183,0.11059072,0.11421664,0.11965553,0.12509441,1.209246,2.2952106,3.3793623,4.465327,5.5494785,4.88956,4.229642,3.5697234,2.909805,2.2498865,5.4497657,8.649645,11.849524,15.049402,18.24928,14.690435,11.129777,7.569119,4.0102735,0.44961473,0.3770962,0.3045777,0.23205921,0.15954071,0.0870222,0.19036107,0.291887,0.39522585,0.49675176,0.6000906,0.5058166,0.40972954,0.3154555,0.21936847,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.099712946,0.13778515,0.17585737,0.21211663,0.25018883,0.20486477,0.15954071,0.11421664,0.07070554,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06164073,0.12509441,0.18673515,0.25018883,0.31182957,0.27919623,0.24837588,0.21574254,0.18310922,0.15047589,0.22662032,0.3045777,0.3825351,0.4604925,0.53663695,0.4894999,0.44236287,0.39522585,0.3480888,0.2991388,0.6399758,0.9808127,1.3198367,1.6606737,1.9996977,3.0983531,4.195195,5.292038,6.390693,7.4875355,6.755099,6.0226617,5.290225,4.557788,3.825351,3.9921436,4.160749,4.327542,4.494334,4.6629395,4.9276323,5.1923246,5.4570174,5.7217097,5.9882154,5.7906027,5.5929894,5.3953767,5.197764,5.0001507,6.049856,7.0995617,8.149267,9.200785,10.25049,10.41547,10.58045,10.745429,10.910409,11.075388,12.5058155,13.93443,15.364858,16.795286,18.225714,15.537089,12.850279,10.161655,7.474845,4.788034,4.3946214,4.0030212,3.6096084,3.2180085,2.8245957,3.8924308,4.9602656,6.0281005,7.0941224,8.161958,7.3352466,6.506723,5.6800117,4.853301,4.024777,4.751775,5.480586,6.207584,6.9345818,7.663393,6.921891,6.1822023,5.4425135,4.702825,3.9631362,3.4301252,2.8971143,2.3641033,1.8329052,1.2998942,1.2799516,1.260009,1.2400664,1.2201238,1.2001812,1.1693609,1.1403534,1.1095331,1.0805258,1.0497054,0.9880646,0.9246109,0.8629702,0.7995165,0.73787576,0.7197462,0.7016165,0.6852999,0.6671702,0.6508536,0.61278135,0.5747091,0.53663695,0.50037766,0.46230546,0.53482395,0.6073425,0.67986095,0.7523795,0.824898,0.85934424,0.89560354,0.9300498,0.9644961,1.0007553,1.4721256,1.9453088,2.4166791,2.8898623,3.3630457,0.18673515,0.20486477,0.2229944,0.23931105,0.2574407,0.2755703,0.60190356,0.9300498,1.258196,1.5845293,1.9126755,2.228131,2.5417736,2.857229,3.1726844,3.48814,4.835171,6.1822023,7.5292335,8.8780775,10.225109,10.411844,10.600392,10.7871275,10.975676,11.162411,13.649796,16.13718,18.624565,21.11195,23.599335,22.390087,21.180841,19.969784,18.760536,17.549479,16.777155,16.004833,15.2325115,14.46019,13.687867,13.327088,12.968122,12.607342,12.248375,11.887595,11.938358,11.9873085,12.038072,12.087022,12.137785,11.989121,11.842272,11.695421,11.546759,11.399909,13.898171,16.39462,18.892883,21.389332,23.887594,27.040337,30.193079,33.34582,36.49675,39.64949,41.310165,42.97084,44.6297,46.290375,47.949234,49.47575,51.00045,52.52515,54.049854,55.574554,50.82822,46.08007,41.33192,36.585587,31.837437,33.117386,34.39734,35.67729,36.95724,38.237194,35.082638,31.928083,28.771717,25.61716,22.462606,23.427103,24.393412,25.357908,26.322403,27.2869,25.385101,23.483305,21.579693,19.677896,17.774284,16.274965,14.775645,13.274512,11.775192,10.274059,10.620335,10.964798,11.30926,11.655537,11.999999,12.779573,13.559147,14.340534,15.120108,15.899682,19.001661,22.105453,25.207432,28.30941,31.413202,31.5945,31.777609,31.960718,32.142014,32.325123,29.725334,27.125546,24.525759,21.924156,19.324368,20.647831,21.96948,23.292944,24.614594,25.938055,26.284332,26.63242,26.980509,27.326784,27.674873,28.249582,28.824291,29.400814,29.975523,30.550232,27.337664,24.125093,20.912523,17.699953,14.487384,13.537392,12.5873995,11.637406,10.687414,9.737422,8.082188,6.4269524,4.7717175,3.1182957,1.4630609,3.245203,5.027345,6.8094873,8.593443,10.375585,8.914337,7.454902,5.995467,4.5342193,3.0747845,2.5073273,1.93987,1.3724127,0.80495536,0.2374981,0.4169814,0.5982776,0.7777609,0.9572442,1.1367276,1.7567607,2.3767939,2.9968271,3.6168604,4.2368937,5.4044414,6.5719895,7.7395372,8.907085,10.074633,11.47424,12.87566,14.275268,15.674874,17.074482,16.807976,16.539658,16.273151,16.004833,15.738328,15.919624,16.102734,16.285843,16.467138,16.650248,16.249584,15.850732,15.4500675,15.049402,14.650551,13.2418785,11.83502,10.428161,9.019489,7.61263,7.6942134,7.7776093,7.859193,7.9425893,8.024173,8.105756,8.185526,8.265296,8.345067,8.424837,8.696781,8.970539,9.242483,9.514427,9.788185,10.092763,10.397341,10.701918,11.008308,11.312886,12.032633,12.752378,13.472125,14.191871,14.911617,15.812659,16.71189,17.612932,18.512161,19.413204,20.642391,21.873394,23.102583,24.33177,25.562773,22.812508,20.062244,17.31198,14.561715,11.813264,11.334642,10.857833,10.37921,9.902402,9.425592,11.214987,13.00438,14.795588,16.584982,18.374376,15.480887,12.585587,9.690285,6.794984,3.8996825,6.089741,8.2798,10.469859,12.659918,14.849977,15.357606,15.865235,16.372866,16.880495,17.388124,18.9092,20.432089,21.954977,23.477865,25.000753,20.905272,16.80979,12.714307,8.620637,4.5251546,4.1879435,3.8507326,3.5117085,3.1744974,2.8372865,3.7691493,4.702825,5.634688,6.5683637,7.500226,7.2917356,7.0850577,6.876567,6.6698895,6.4632115,7.230095,7.996978,8.765674,9.5325575,10.29944,8.430276,6.5592985,4.690134,2.819157,0.9499924,0.93911463,0.9300498,0.91917205,0.9101072,0.89922947,1.357909,1.8147756,2.2716422,2.7303216,3.1871881,3.727451,4.267714,4.8079767,5.3482394,5.8866897,4.896812,3.9069343,2.9170568,1.9271792,0.93730164,0.83033687,0.72337204,0.61459434,0.5076295,0.40066472,0.91917205,1.4394923,1.9598125,2.4801328,3.000453,2.4420607,1.8854811,1.3270886,0.7705091,0.21211663,0.59283876,0.97174793,1.35247,1.7331922,2.1121013,2.0123885,1.9126755,1.8129625,1.7132497,1.6117238,3.2669585,4.9221935,6.5774283,8.232663,9.8878975,8.417585,6.947273,5.47696,4.006647,2.5381477,4.0392804,5.542227,7.0451727,8.548119,10.049252,8.113008,6.1749506,4.2368937,2.3006494,0.36259252,2.8608549,5.3573046,7.855567,10.352016,12.850279,11.907538,10.964798,10.022058,9.079316,8.138389,8.138389,8.138389,8.138389,8.138389,8.138389,7.8120556,7.4875355,7.1630154,6.836682,6.5121617,5.5132194,4.512464,3.5117085,2.5127661,1.5120108,1.3252757,1.1367276,0.9499924,0.76325727,0.5747091,0.48043507,0.38434806,0.29007402,0.19579996,0.099712946,0.11059072,0.11965553,0.13053331,0.13959812,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.0,0.0,0.0,0.0,0.0,0.027194439,0.054388877,0.08339628,0.11059072,0.13778515,0.11059072,0.08339628,0.054388877,0.027194439,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.16497959,0.32995918,0.4949388,0.65991837,0.824898,0.6653573,0.5058166,0.3444629,0.18492219,0.025381476,0.030820364,0.034446288,0.03988518,0.045324065,0.05076295,0.06707962,0.08520924,0.10333887,0.11965553,0.13778515,0.15954071,0.18310922,0.20486477,0.22662032,0.25018883,0.2229944,0.19579996,0.16679256,0.13959812,0.11240368,0.10696479,0.10333887,0.09789998,0.092461094,0.0870222,0.09427405,0.10333887,0.11059072,0.11784257,0.12509441,1.0533313,1.9797552,2.907992,3.834416,4.762653,4.4852695,4.207886,3.930503,3.6531196,3.3757362,7.175706,10.975676,14.775645,18.575615,22.375584,17.959208,13.544643,9.130079,4.7155156,0.2991388,0.25925365,0.21936847,0.1794833,0.13959812,0.099712946,0.17223145,0.24474995,0.31726846,0.38978696,0.46230546,0.39522585,0.32814622,0.25925365,0.19217403,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.0870222,0.11240368,0.13778515,0.16316663,0.18673515,0.15772775,0.12690738,0.09789998,0.06707962,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06164073,0.12509441,0.18673515,0.25018883,0.31182957,0.27013144,0.22662032,0.18492219,0.14322405,0.099712946,0.19761293,0.2955129,0.39159992,0.4894999,0.5873999,0.53482395,0.48224804,0.42967212,0.3770962,0.3245203,0.6091554,0.89560354,1.1802386,1.4648738,1.7495089,2.7266958,3.7056956,4.6828823,5.660069,6.637256,6.057108,5.47696,4.896812,4.3166637,3.738329,3.9323158,4.1281157,4.322103,4.517903,4.7118897,5.034597,5.3573046,5.6800117,6.002719,6.3254266,5.8721857,5.4207582,4.9675174,4.514277,4.062849,4.9620786,5.863121,6.7623506,7.66158,8.562622,8.709473,8.858135,9.004985,9.151835,9.300498,10.607644,11.91479,13.221936,14.529082,15.838041,13.437678,11.037316,8.636953,6.2384043,3.8380418,3.7927177,3.7473936,3.7020695,3.6567454,3.6132345,4.157123,4.702825,5.2467136,5.7924156,6.338117,5.75253,5.1669436,4.5831695,3.9975824,3.4119956,3.9848917,4.557788,5.130684,5.7017674,6.2746634,5.714458,5.1542525,4.59586,4.0356545,3.4754493,3.1074178,2.7393866,2.373168,2.0051367,1.6371052,1.5573349,1.4775645,1.3977941,1.3180238,1.2382535,1.1802386,1.1222239,1.064209,1.0080072,0.9499924,0.9246109,0.89922947,0.87566096,0.85027945,0.824898,0.81764615,0.8103943,0.8031424,0.79589057,0.7868258,0.7124943,0.63816285,0.5620184,0.48768693,0.41335547,0.5402629,0.6671702,0.79589057,0.922798,1.0497054,1.114972,1.1802386,1.2455053,1.310772,1.3742256,1.840157,2.3042755,2.770207,3.2343252,3.7002566,0.25018883,0.26469254,0.27919623,0.2955129,0.3100166,0.3245203,0.7451276,1.1657349,1.5845293,2.0051367,2.4257438,2.808279,3.1908143,3.5733492,3.9558845,4.3384194,5.7924156,7.2482243,8.70222,10.15803,11.612025,11.73712,11.862214,11.9873085,12.112403,12.237497,14.525456,16.811602,19.099562,21.38752,23.675478,22.645716,21.61414,20.584377,19.554615,18.52485,17.206827,15.890617,14.572594,13.254569,11.938358,12.019942,12.103338,12.184921,12.268318,12.349901,12.375282,12.400664,12.4242325,12.449615,12.474996,12.320893,12.164979,12.010877,11.854962,11.700861,14.817343,17.935638,21.052122,24.170418,27.2869,30.419699,33.552498,36.6853,39.818096,42.950897,44.279797,45.61051,46.939415,48.27013,49.60084,51.41199,53.224957,55.037918,56.85088,58.66203,54.407005,50.151985,45.89696,41.641937,37.386913,38.82822,40.26771,41.707203,43.14851,44.588,40.684692,36.7832,32.87989,28.978394,25.075085,26.29521,27.515333,28.735456,29.955582,31.175705,29.143373,27.10923,25.076899,23.044567,21.012236,18.562923,16.1118,13.662486,11.213174,8.762048,8.3595705,7.957093,7.554615,7.1521373,6.7496595,7.0524244,7.3551893,7.6579537,7.9607186,8.26167,13.820213,19.376944,24.935488,30.492218,36.050762,36.922794,37.79483,38.666866,39.540714,40.41275,35.925667,31.438583,26.949688,22.462606,17.975525,19.879135,21.78456,23.689981,25.595406,27.50083,28.18069,28.860552,29.540413,30.220274,30.900135,31.674269,32.45022,33.224354,34.0003,34.774437,30.588305,26.400362,22.212418,18.024473,13.838344,13.049705,12.262879,11.47424,10.687414,9.900589,8.247167,6.5955577,4.942136,3.290527,1.6371052,3.834416,6.0317264,8.23085,10.428161,12.625471,10.906783,9.189907,7.473032,5.754343,4.0374675,3.2850883,2.5327086,1.7803292,1.0279498,0.2755703,0.47680917,0.67986095,0.88291276,1.0841516,1.2872034,2.0232663,2.7575161,3.491766,4.227829,4.9620786,6.1405044,7.317117,8.495543,9.672155,10.850581,12.413355,13.974316,15.537089,17.099863,18.662638,18.022661,17.382685,16.74271,16.102734,15.462758,15.660371,15.857984,16.055597,16.25321,16.450823,15.925063,15.399304,14.875358,14.349599,13.825653,12.540262,11.254871,9.969481,8.684091,7.400513,7.4349594,7.4694057,7.5056653,7.5401115,7.574558,7.665206,7.755854,7.844689,7.935337,8.024173,8.366822,8.709473,9.052122,9.394773,9.737422,9.864329,9.99305,10.119957,10.246864,10.375585,10.810696,11.245807,11.679105,12.114216,12.549327,14.824595,17.099863,19.375132,21.650398,23.925667,24.678047,25.430426,26.182806,26.935184,27.687565,24.549326,21.4129,18.274662,15.138238,11.999999,11.980057,11.9601145,11.940171,11.920229,11.900287,13.194741,14.489197,15.785465,17.07992,18.374376,15.1781225,11.980057,8.781991,5.5857377,2.3876717,5.632875,8.8780775,12.123281,15.368484,18.611874,18.947271,19.282671,19.618069,19.951653,20.287052,21.893335,23.497808,25.10228,26.70675,28.313036,23.414412,18.5176,13.618975,8.722163,3.825351,3.437377,3.049403,2.663242,2.275268,1.887294,2.659616,3.4319382,4.2042603,4.976582,5.750717,5.8395524,5.9302006,6.0208488,6.109684,6.200332,7.364254,8.529989,9.695724,10.859646,12.025381,9.789998,7.554615,5.319232,3.0856624,0.85027945,0.8194591,0.7904517,0.75963134,0.7306239,0.69980353,1.3216497,1.9453088,2.5671551,3.1908143,3.8126602,4.220577,4.6266804,5.034597,5.4425135,5.8504305,4.9294453,4.0102735,3.0892882,2.1701162,1.2491312,1.0406405,0.83033687,0.6200332,0.40972954,0.19942589,0.8103943,1.4195497,2.030518,2.6396735,3.2506418,2.6269827,2.0051367,1.3832904,0.75963134,0.13778515,0.6653573,1.1929294,1.7205015,2.2480736,2.7756457,2.6378605,2.5000753,2.3622901,2.2245052,2.08672,4.265901,6.4432693,8.620637,10.798005,12.975373,11.05182,9.130079,7.208339,5.2847857,3.3630457,5.2702823,7.177519,9.084756,10.991992,12.899229,10.411844,7.9244595,5.4370747,2.94969,0.46230546,3.5044568,6.546608,9.590572,12.632723,15.674874,14.485571,13.294455,12.105151,10.915848,9.724731,9.788185,9.849826,9.91328,9.97492,10.038374,9.449161,8.861761,8.274362,7.686961,7.0995617,6.049856,5.0001507,3.9504454,2.9007401,1.8492218,1.6244144,1.3996071,1.1747998,0.9499924,0.72518504,0.58921283,0.4550536,0.3208944,0.18492219,0.05076295,0.07977036,0.11059072,0.13959812,0.17041849,0.19942589,0.15954071,0.11965553,0.07977036,0.03988518,0.0,0.0,0.0,0.0,0.0,0.0,0.032633327,0.065266654,0.09789998,0.13053331,0.16316663,0.13053331,0.09789998,0.065266654,0.032633327,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.21936847,0.4405499,0.65991837,0.8792868,1.1004683,0.88291276,0.6653573,0.44780177,0.23024625,0.012690738,0.014503701,0.018129626,0.01994259,0.02175555,0.025381476,0.03988518,0.054388877,0.07070554,0.08520924,0.099712946,0.13053331,0.15954071,0.19036107,0.21936847,0.25018883,0.21755551,0.18492219,0.15228885,0.11965553,0.0870222,0.08520924,0.08339628,0.07977036,0.07795739,0.07433146,0.08520924,0.09427405,0.10515183,0.11421664,0.12509441,0.89560354,1.6642996,2.4348087,3.2053177,3.975827,4.079166,4.1843176,4.2894692,4.3946214,4.499773,8.899834,13.299893,17.699953,22.100014,26.500074,21.229792,15.95951,10.689227,5.4207582,0.15047589,0.14322405,0.13415924,0.12690738,0.11965553,0.11240368,0.15410182,0.19761293,0.23931105,0.28282216,0.3245203,0.28463513,0.24474995,0.20486477,0.16497959,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.11059072,0.09427405,0.07977036,0.065266654,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06164073,0.12509441,0.18673515,0.25018883,0.31182957,0.25925365,0.20667773,0.15410182,0.10333887,0.05076295,0.16679256,0.28463513,0.40247768,0.52032024,0.63816285,0.58014804,0.52213323,0.46411842,0.40791658,0.34990177,0.58014804,0.8103943,1.0406405,1.2708868,1.49932,2.3568513,3.2143826,4.071914,4.9294453,5.7869763,5.3591175,4.933071,4.505212,4.077353,3.6494937,3.872488,4.0954823,4.3166637,4.539658,4.762653,5.143375,5.522284,5.903006,6.281915,6.6626377,5.955582,5.2467136,4.539658,3.832603,3.1255474,3.874301,4.6248674,5.375434,6.1241875,6.874754,7.0052876,7.135821,7.264541,7.3950744,7.5256076,8.709473,9.89515,11.080828,12.264692,13.45037,11.336455,9.224354,7.112252,5.0001507,2.8880494,3.1908143,3.491766,3.7945306,4.0972953,4.40006,4.421816,4.445384,4.4671397,4.4907084,4.512464,4.169814,3.827164,3.484514,3.141864,2.7992141,3.2180085,3.63499,4.0519714,4.4707656,4.8877473,4.507025,4.1281157,3.7473936,3.3666716,2.9877625,2.7847104,2.5816586,2.38042,2.1773682,1.9743162,1.8347181,1.69512,1.5555218,1.4141108,1.2745126,1.1893034,1.1040943,1.020698,0.9354887,0.85027945,0.8629702,0.87566096,0.8883517,0.89922947,0.9119202,0.9155461,0.91735905,0.91917205,0.922798,0.9246109,0.8122072,0.69980353,0.5873999,0.4749962,0.36259252,0.54570174,0.726998,0.9101072,1.0932164,1.2745126,1.3705997,1.4648738,1.5591478,1.6552348,1.7495089,2.2081885,2.665055,3.1219215,3.5806012,4.0374675,0.31182957,0.3245203,0.33721104,0.34990177,0.36259252,0.37528324,0.8883517,1.3996071,1.9126755,2.4257438,2.9369993,3.386614,3.8380418,4.2876563,4.7372713,5.186886,6.7496595,8.312433,9.875207,11.437981,13.000754,13.062395,13.125849,13.1874895,13.24913,13.312584,15.399304,17.487837,19.574556,21.66309,23.74981,22.89953,22.049252,21.200785,20.350506,19.500225,17.638313,15.774588,13.912675,12.050762,10.1870365,10.712796,11.236742,11.762501,12.28826,12.812206,12.812206,12.812206,12.812206,12.812206,12.812206,12.650853,12.487686,12.32452,12.163166,11.999999,15.738328,19.474844,23.213173,26.949688,30.688017,33.79906,36.91192,40.024776,43.13763,46.25049,47.24943,48.250187,49.24913,50.249886,51.25064,53.350048,55.44946,57.550686,59.650093,61.749504,57.98761,54.22571,50.462,46.700104,42.938206,44.53724,46.138084,47.737118,49.337963,50.936996,46.286747,41.638313,36.988064,32.337814,27.687565,29.163317,30.637255,32.113007,33.586945,35.062695,32.899834,30.736967,28.574102,26.413052,24.250187,20.850883,17.449764,14.05046,10.649343,7.250037,6.1006193,4.949388,3.7999697,2.6505513,1.49932,1.3252757,1.1494182,0.97537386,0.7995165,0.62547207,8.636953,16.650248,24.663544,32.675026,40.68832,42.24928,43.812054,45.37483,46.937603,48.500374,42.126,35.74981,29.375433,22.999243,16.624866,19.112251,21.599636,24.08702,26.574406,29.06179,30.075235,31.08687,32.100315,33.11195,34.125393,35.10077,36.07433,37.0497,38.025078,39.00045,33.837135,28.675629,23.512312,18.350807,13.1874895,12.562017,11.938358,11.312886,10.687414,10.061942,8.412147,6.7623506,5.1125546,3.4627585,1.8129625,4.4254417,7.037921,9.6504,12.262879,14.875358,12.899229,10.924912,8.950596,6.9744673,5.0001507,4.062849,3.1255474,2.1882458,1.2491312,0.31182957,0.53663695,0.76325727,0.9880646,1.2128719,1.4376793,2.2879589,3.1382382,3.9867048,4.836984,5.6872635,6.874754,8.062244,9.249735,10.437225,11.624716,13.3506565,15.074784,16.800724,18.52485,20.250792,19.237347,18.225714,17.212267,16.200634,15.187187,15.399304,15.613234,15.825351,16.037468,16.249584,15.600543,14.94969,14.300649,13.649796,13.000754,11.836833,10.674724,9.512614,8.350506,7.1883965,7.175706,7.1630154,7.1503243,7.137634,7.124943,7.224656,7.324369,7.4258947,7.5256076,7.6253204,8.036863,8.450218,8.861761,9.275117,9.686659,9.637709,9.5869465,9.537996,9.487233,9.438283,9.5869465,9.737422,9.8878975,10.038374,10.1870365,13.838344,17.487837,21.137331,24.786825,28.438131,28.71189,28.98746,29.26303,29.536787,29.812357,26.287958,22.761745,19.237347,15.712947,12.186734,12.625471,13.062395,13.499319,13.938056,14.37498,15.174497,15.975826,16.775343,17.57486,18.374376,14.875358,11.374527,7.8755093,4.3746786,0.87566096,5.1741953,9.474543,13.77489,18.075237,22.375584,22.536938,22.700104,22.863272,23.024624,23.187792,24.87566,26.561714,28.249582,29.93745,31.625319,25.925365,20.22541,14.525456,8.825501,3.1255474,2.6868105,2.2498865,1.8129625,1.3742256,0.93730164,1.550083,2.1628644,2.7756457,3.386614,3.9993954,4.3873696,4.7753434,5.163317,5.5494785,5.9374523,7.500226,9.063,10.625773,12.186734,13.749508,11.14972,8.549932,5.9501433,3.350355,0.7505665,0.69980353,0.6508536,0.6000906,0.5493277,0.50037766,1.2872034,2.0758421,2.8626678,3.6494937,4.4381323,4.7118897,4.98746,5.2630305,5.5367875,5.812358,4.9620786,4.1117992,3.2633326,2.4130533,1.5627737,1.2491312,0.93730164,0.62547207,0.31182957,0.0,0.69980353,1.3996071,2.0994108,2.7992141,3.5008307,2.811905,2.124792,1.4376793,0.7505665,0.06164073,0.73787576,1.4122978,2.08672,2.762955,3.437377,3.2633326,3.0874753,2.911618,2.7375734,2.561716,5.2630305,7.9625316,10.662033,13.363347,16.062849,13.687867,11.312886,8.937905,6.5629244,4.1879435,6.4994707,8.812811,11.124338,13.437678,15.749206,12.712494,9.675781,6.637256,3.6005437,0.5620184,4.1498713,7.7377243,11.325577,14.91343,18.49947,17.06179,15.625924,14.188245,12.750566,11.312886,11.437981,11.563075,11.6881695,11.813264,11.938358,11.088079,10.2378,9.38752,8.537241,7.686961,6.588306,5.487838,4.3873696,3.2869012,2.1882458,1.9253663,1.6624867,1.3996071,1.1367276,0.87566096,0.69980353,0.52575916,0.34990177,0.17585737,0.0,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.0,0.0,0.0,0.0,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.2755703,0.5493277,0.824898,1.1004683,1.3742256,1.1004683,0.824898,0.5493277,0.2755703,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.099712946,0.13778515,0.17585737,0.21211663,0.25018883,0.21211663,0.17585737,0.13778515,0.099712946,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.73787576,1.3506571,1.9616255,2.5744069,3.1871881,3.6748753,4.162562,4.650249,5.137936,5.6256227,10.625773,15.624111,20.624262,25.624413,30.624563,24.500376,18.374376,12.250188,6.1241875,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.13778515,0.15047589,0.16316663,0.17585737,0.18673515,0.17585737,0.16316663,0.15047589,0.13778515,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06164073,0.12509441,0.18673515,0.25018883,0.31182957,0.25018883,0.18673515,0.12509441,0.06164073,0.0,0.13778515,0.2755703,0.41335547,0.5493277,0.6871128,0.62547207,0.5620184,0.50037766,0.43692398,0.37528324,0.5493277,0.72518504,0.89922947,1.0750868,1.2491312,1.987007,2.7248828,3.4627585,4.2006345,4.936697,4.6629395,4.3873696,4.1117992,3.8380418,3.5624714,3.8126602,4.062849,4.313038,4.5632267,4.8116026,5.2503395,5.6872635,6.1241875,6.5629244,6.9998484,6.037165,5.0744824,4.1117992,3.150929,2.1882458,2.7883365,3.386614,3.9867048,4.5867953,5.186886,5.2992897,5.411693,5.52591,5.638314,5.750717,6.813113,7.8755093,8.937905,10.000301,11.062697,9.237044,7.413204,5.5875506,3.7618973,1.938057,2.5870976,3.2379513,3.8869917,4.537845,5.186886,4.688321,4.1879435,3.6875658,3.1871881,2.6868105,2.5870976,2.4873846,2.3876717,2.2879589,2.1882458,2.4493124,2.712192,2.9750717,3.2379513,3.5008307,3.299592,3.100166,2.9007401,2.6995013,2.5000753,2.4620032,2.4257438,2.3876717,2.3495996,2.3133402,2.1121013,1.9126755,1.7132497,1.5120108,1.3125849,1.2001812,1.0877775,0.97537386,0.8629702,0.7505665,0.7995165,0.85027945,0.89922947,0.9499924,1.0007553,1.0116332,1.0243238,1.0370146,1.0497054,1.062396,0.9119202,0.76325727,0.61278135,0.46230546,0.31182957,0.5493277,0.7868258,1.0243238,1.261822,1.49932,1.6244144,1.7495089,1.8746033,1.9996977,2.124792,2.5744069,3.0258346,3.4754493,3.925064,4.3746786,0.25018883,0.58014804,0.9101072,1.2400664,1.5700256,1.8999848,2.4076142,2.9152439,3.4228733,3.930503,4.4381323,4.646623,4.856927,5.06723,5.277534,5.487838,6.789545,8.093065,9.394773,10.698292,11.999999,12.15954,12.320893,12.480434,12.639976,12.799516,14.277081,15.754644,17.23221,18.709774,20.187338,19.730473,19.271791,18.814926,18.358059,17.89938,16.38193,14.86448,13.347031,11.829581,10.312131,10.852394,11.392657,11.9329195,12.473183,13.011633,12.951805,12.891977,12.8321495,12.772322,12.712494,12.627284,12.542075,12.456866,12.371656,12.28826,15.557032,18.827616,22.098202,25.366972,28.637556,31.630758,34.622147,37.61535,40.606735,43.599937,45.356697,47.115273,48.872032,50.630608,52.387367,54.492218,56.597065,58.701916,60.806767,62.911613,59.03006,55.14851,51.265144,47.38178,43.500225,44.350502,45.200783,46.049248,46.89953,47.74981,43.538296,39.32497,35.111645,30.900135,26.68681,27.975826,29.26303,30.550232,31.837437,33.124638,31.057861,28.989271,26.922495,24.855717,22.787127,20.517298,18.247469,15.977639,13.70781,11.437981,10.455356,9.47273,8.490104,7.507478,6.5248523,5.9718986,5.4207582,4.8678045,4.314851,3.7618973,9.875207,15.986704,22.100014,28.213324,34.32482,35.220425,36.114216,37.00982,37.905422,38.801025,33.76099,28.720953,23.679104,18.64088,13.600845,15.575162,17.549479,19.525606,21.499924,23.47424,24.23931,25.00438,25.76945,26.534521,27.299591,28.080976,28.860552,29.640125,30.419699,31.199272,27.372108,23.544945,19.717781,15.890617,12.06164,11.338268,10.613083,9.8878975,9.162713,8.437528,7.124943,5.812358,4.499773,3.1871881,1.8746033,4.160749,6.445082,8.729415,11.015561,13.299893,11.485118,9.670342,7.855567,6.0407915,4.2242026,3.489953,2.7557032,2.0196402,1.2853905,0.5493277,1.1766127,1.8057107,2.4329958,3.0602808,3.6875658,4.2949085,4.902251,5.5095935,6.1169357,6.7242785,7.574558,8.424837,9.275117,10.125396,10.975676,12.45324,13.930804,15.408369,16.885933,18.361685,17.612932,16.862366,16.1118,15.363045,14.612478,14.795588,14.976884,15.159993,15.343102,15.524399,14.960567,14.394923,13.829279,13.265448,12.699803,11.717177,10.734551,9.751925,8.7693,7.7866745,7.7268467,7.667019,7.607191,7.5473633,7.4875355,7.7141557,7.9425893,8.1692095,8.397643,8.624263,9.11195,9.599637,10.087324,10.57501,11.062697,10.805257,10.547816,10.290376,10.032935,9.775495,10.239613,10.705544,11.169662,11.635593,12.099712,14.969632,17.839552,20.70947,23.579391,26.44931,27.080221,27.70932,28.34023,28.96933,29.60024,26.104849,22.609457,19.114065,15.620485,12.125093,12.420607,12.714307,13.009819,13.305332,13.600845,14.211814,14.824595,15.437376,16.050158,16.66294,14.01964,11.378153,8.734854,6.091554,3.4500678,6.833056,10.2142315,13.597219,16.980207,20.363195,20.580751,20.798307,21.015862,21.233418,21.44916,22.489801,23.530441,24.56927,25.60991,26.65055,21.985798,17.321045,12.654479,7.989726,3.3249733,3.0149567,2.70494,2.3949237,2.084907,1.7748904,2.1229792,2.469255,2.817344,3.1654327,3.5117085,3.8398547,4.168001,4.494334,4.8224807,5.1506267,6.552047,7.95528,9.3567,10.7599325,12.163166,10.2142315,8.267109,6.319988,4.3728657,2.4257438,2.182807,1.93987,1.696933,1.455809,1.2128719,1.84197,2.472881,3.101979,3.73289,4.361988,4.5650396,4.7680917,4.9693303,5.1723824,5.375434,4.550536,3.7256382,2.9007401,2.0758421,1.2491312,1.0823387,0.9155461,0.7469406,0.58014804,0.41335547,0.98443866,1.5573349,2.1302311,2.7031271,3.2742105,2.9351864,2.5943494,2.2553256,1.9144884,1.5754645,2.4094272,3.245203,4.079166,4.914942,5.750717,5.2666564,4.784408,4.3021603,3.8199122,3.3376641,5.2467136,7.157576,9.068439,10.9774885,12.888351,11.6047735,10.323009,9.039432,7.757667,6.474089,7.7177815,8.9596615,10.203354,11.445232,12.687112,10.25049,7.8120556,5.375434,2.9369993,0.50037766,3.3848011,6.2692246,9.155461,12.039885,14.924308,13.800271,12.674421,11.5503845,10.424535,9.300498,9.447348,9.594198,9.742861,9.88971,10.038374,9.333132,8.627889,7.9226465,7.217404,6.5121617,5.560356,4.606738,3.6549325,2.7031271,1.7495089,1.5428312,1.3343405,1.1276628,0.91917205,0.7124943,0.581961,0.45324063,0.32270733,0.19217403,0.06164073,0.09064813,0.11784257,0.14503701,0.17223145,0.19942589,0.15954071,0.11965553,0.07977036,0.03988518,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.03988518,0.06707962,0.09427405,0.12328146,0.15047589,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.045324065,0.065266654,0.08520924,0.10515183,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.2229944,0.44417584,0.6671702,0.8901646,1.1131591,0.90285534,0.69255173,0.48224804,0.27194437,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.07977036,0.11059072,0.13959812,0.17041849,0.19942589,0.17223145,0.14503701,0.11784257,0.09064813,0.06164073,0.059827764,0.058014803,0.054388877,0.052575916,0.05076295,0.059827764,0.07070554,0.07977036,0.09064813,0.099712946,0.59283876,1.0841516,1.5772774,2.0704033,2.561716,3.002266,3.442816,3.8833659,4.322103,4.762653,8.890768,13.017072,17.145187,21.273302,25.399607,20.321497,15.245202,10.167094,5.090799,0.012690738,0.038072214,0.06164073,0.0870222,0.11240368,0.13778515,0.14503701,0.15228885,0.15954071,0.16679256,0.17585737,0.15954071,0.14503701,0.13053331,0.11421664,0.099712946,0.09064813,0.07977036,0.07070554,0.059827764,0.05076295,0.052575916,0.054388877,0.058014803,0.059827764,0.06164073,0.07795739,0.092461094,0.10696479,0.12328146,0.13778515,0.11059072,0.08339628,0.054388877,0.027194439,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.08339628,0.13959812,0.19761293,0.25562772,0.31182957,0.2520018,0.19217403,0.13234627,0.072518505,0.012690738,0.15047589,0.28826106,0.42423326,0.5620184,0.69980353,0.62728506,0.55476654,0.48224804,0.40972954,0.33721104,0.4894999,0.6417888,0.79589057,0.9481794,1.1004683,1.6896812,2.280707,2.8699198,3.4591327,4.0501585,3.966762,3.8851788,3.8017826,3.720199,3.636803,3.9975824,4.358362,4.7173285,5.0781083,5.4370747,5.7779117,6.1169357,6.4577727,6.796797,7.137634,6.1948934,5.2521524,4.309412,3.3666716,2.4257438,2.8427253,3.2597067,3.6766882,4.0954823,4.512464,4.604925,4.6973863,4.7898474,4.882308,4.974769,5.91751,6.8602505,7.802991,8.745731,9.686659,8.149267,6.6118746,5.0744824,3.53709,1.9996977,2.5308957,3.0602808,3.589666,4.120864,4.650249,4.269527,3.8906176,3.5098956,3.1291735,2.7502642,2.665055,2.5798457,2.4946365,2.4094272,2.324218,2.5327086,2.7393866,2.9478772,3.1545548,3.3630457,3.1781235,2.9932013,2.808279,2.6233568,2.4366217,2.4021754,2.3677292,2.333283,2.2970235,2.2625773,2.1048496,1.9471219,1.789394,1.6316663,1.4757515,1.3542831,1.2346275,1.114972,0.99531645,0.87566096,0.922798,0.969935,1.017072,1.064209,1.1131591,1.0605831,1.0080072,0.9554313,0.90285534,0.85027945,0.81583315,0.7795739,0.7451276,0.7106813,0.6744221,0.85027945,1.0243238,1.2001812,1.3742256,1.550083,2.0631514,2.5744069,3.0874753,3.6005437,4.1117992,4.3529234,4.592234,4.8333583,5.0726695,5.3119802,0.18673515,0.83577573,1.4830034,2.1302311,2.7774587,3.4246864,3.926877,4.4308805,4.933071,5.4352617,5.9374523,5.906632,5.8776245,5.846804,5.8177967,5.7869763,6.82943,7.8718834,8.914337,9.956791,10.999244,11.256684,11.514126,11.773379,12.03082,12.28826,13.154857,14.023266,14.889862,15.758271,16.624866,16.5596,16.494333,16.43088,16.365614,16.300346,15.127359,13.954373,12.783199,11.610212,10.437225,10.991992,11.546759,12.103338,12.658105,13.212872,13.093216,12.971747,12.852092,12.732436,12.612781,12.605529,12.598277,12.589212,12.581961,12.574709,15.377548,18.18039,20.983229,23.784256,26.587097,29.460642,32.332375,35.20592,38.077652,40.949387,43.46578,45.98036,48.494938,51.009514,53.525906,55.634384,57.74467,59.85496,61.96525,64.07554,60.072514,56.069492,52.068287,48.065266,44.062244,44.161957,44.26167,44.363194,44.462906,44.562622,40.788033,37.013443,33.23704,29.462456,25.687866,26.788336,27.88699,28.98746,30.087927,31.186583,29.215893,27.24339,25.269072,23.29657,21.325878,20.185526,19.045172,17.904818,16.764465,15.625924,14.810091,13.994258,13.180238,12.364405,11.5503845,10.620335,9.690285,8.760235,7.8301854,6.9001355,11.111648,15.324973,19.538298,23.74981,27.963135,28.189754,28.418188,28.64481,28.873241,29.099863,25.394167,21.690285,17.984589,14.280706,10.57501,12.038072,13.499319,14.96238,16.425442,17.886688,18.405195,18.92189,19.440397,19.957092,20.4756,21.059374,21.64496,22.230547,22.814322,23.399908,20.907085,18.41426,15.92325,13.430427,10.937603,10.112705,9.287807,8.46291,7.6380115,6.813113,5.8377395,4.8623657,3.8869917,2.911618,1.938057,3.8942437,5.8522434,7.8102427,9.768243,11.724429,10.069194,8.415772,6.7605376,5.105303,3.4500678,2.9170568,2.3858588,1.8528478,1.3198367,0.7868258,1.8165885,2.8481643,3.877927,4.9076896,5.9374523,6.301858,6.6680765,7.0324817,7.3968873,7.763106,8.274362,8.78743,9.300498,9.811753,10.324821,11.555823,12.785012,14.014201,15.245202,16.474392,15.986704,15.50083,15.013144,14.525456,14.037769,14.190058,14.342347,14.494636,14.646925,14.799213,14.320591,13.840157,13.359721,12.879286,12.400664,11.597522,10.794379,9.99305,9.189907,8.386765,8.2798,8.172835,8.06587,7.957093,7.850128,8.205468,8.560809,8.914337,9.269678,9.625018,10.1870365,10.750868,11.312886,11.874905,12.436923,11.972805,11.506873,11.042755,10.576823,10.112705,10.89228,11.671853,12.45324,13.232814,14.012388,16.102734,18.193079,20.283426,22.371958,24.462305,25.446743,26.432995,27.417433,28.401873,29.388123,25.92174,22.457167,18.992596,15.528025,12.06164,12.215742,12.368031,12.52032,12.672608,12.824898,13.24913,13.675177,14.09941,14.525456,14.94969,13.165734,11.379966,9.594198,7.8102427,6.0244746,8.490104,10.955733,13.419549,15.885179,18.350807,18.622751,18.894695,19.166641,19.440397,19.712341,20.105755,20.497355,20.890768,21.282368,21.675781,18.044416,14.4148655,10.785315,7.155763,3.5243993,3.343103,3.159994,2.9768846,2.7955883,2.612479,2.6958754,2.7774587,2.8608549,2.9424384,3.0258346,3.29234,3.5606585,3.827164,4.0954823,4.361988,5.6056805,6.8475595,8.089439,9.333132,10.57501,9.280556,7.9842873,6.6898317,5.3953767,4.099108,3.6658103,3.2306993,2.7955883,2.3604772,1.9253663,2.3967366,2.8699198,3.343103,3.8144734,4.2876563,4.41819,4.5469103,4.6774435,4.8079767,4.936697,4.137181,3.3376641,2.5381477,1.7368182,0.93730164,0.9155461,0.8919776,0.87022203,0.8466535,0.824898,1.2708868,1.7150626,2.1592383,2.6052272,3.049403,3.056655,3.0657198,3.0729716,3.0802233,3.0874753,4.082792,5.0781083,6.073425,7.066928,8.062244,7.271793,6.4831543,5.6927023,4.902251,4.1117992,5.23221,6.352621,7.473032,8.59163,9.712041,9.52168,9.333132,9.142771,8.952409,8.762048,8.934279,9.108324,9.280556,9.452786,9.625018,7.7866745,5.9501433,4.1117992,2.275268,0.43692398,2.619731,4.802538,6.985345,9.168152,11.349146,10.536939,9.724731,8.912524,8.100317,7.28811,7.456715,7.6271334,7.797552,7.9679704,8.138389,7.5781837,7.017978,6.4577727,5.8975673,5.337362,4.5324063,3.727451,2.9224956,2.1175404,1.3125849,1.1602961,1.0080072,0.8557183,0.7016165,0.5493277,0.46411842,0.38072214,0.2955129,0.21030366,0.12509441,0.13053331,0.13415924,0.13959812,0.14503701,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.04169814,0.059827764,0.07795739,0.09427405,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.05076295,0.09064813,0.13053331,0.17041849,0.21030366,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.0,0.0,0.0,0.0,0.0,0.17041849,0.34083697,0.5094425,0.67986095,0.85027945,0.70524246,0.56020546,0.41516843,0.27013144,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.059827764,0.08339628,0.10515183,0.12690738,0.15047589,0.13234627,0.11421664,0.09789998,0.07977036,0.06164073,0.058014803,0.052575916,0.047137026,0.04169814,0.038072214,0.045324065,0.052575916,0.059827764,0.06707962,0.07433146,0.44780177,0.8194591,1.1929294,1.5645868,1.938057,2.3296568,2.72307,3.1146698,3.5080826,3.8996825,7.155763,10.410031,13.664299,16.92038,20.174648,16.144432,12.114216,8.084001,4.0555973,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.15047589,0.15228885,0.15410182,0.15772775,0.15954071,0.16316663,0.14503701,0.12690738,0.11059072,0.092461094,0.07433146,0.06707962,0.059827764,0.052575916,0.045324065,0.038072214,0.04169814,0.047137026,0.052575916,0.058014803,0.06164073,0.092461094,0.12328146,0.15228885,0.18310922,0.21211663,0.17041849,0.12690738,0.08520924,0.04169814,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.10333887,0.15410182,0.20667773,0.25925365,0.31182957,0.25562772,0.19761293,0.13959812,0.08339628,0.025381476,0.16316663,0.2991388,0.43692398,0.5747091,0.7124943,0.629098,0.5475147,0.46411842,0.3825351,0.2991388,0.42967212,0.56020546,0.69073874,0.8194591,0.9499924,1.3923552,1.8347181,2.277081,2.7194438,3.1618068,3.2723975,3.3829882,3.491766,3.6023567,3.7129474,4.1825047,4.652062,5.121619,5.5929894,6.0625467,6.305484,6.546608,6.789545,7.0324817,7.2754188,6.352621,5.429823,4.507025,3.584227,2.663242,2.8971143,3.1327994,3.3666716,3.6023567,3.8380418,3.9105604,3.9830787,4.0555973,4.1281157,4.2006345,5.0219064,5.844991,6.6680765,7.4893484,8.312433,7.063302,5.812358,4.5632267,3.3122826,2.0631514,2.472881,2.8826106,3.29234,3.7020695,4.1117992,3.8525455,3.5932918,3.3322253,3.0729716,2.811905,2.7430124,2.6723068,2.6016014,2.5327086,2.4620032,2.6142921,2.7683938,2.9206827,3.0729716,3.2252605,3.054842,2.8844235,2.715818,2.5453994,2.374981,2.3423476,2.3097143,2.277081,2.2444477,2.2118144,2.0975976,1.983381,1.8673514,1.7531348,1.6371052,1.5101979,1.3832904,1.2545701,1.1276628,1.0007553,1.0442665,1.0895905,1.1349145,1.1802386,1.2255627,1.1077201,0.9898776,0.872035,0.7541924,0.63816285,0.7179332,0.79770356,0.8774739,0.9572442,1.0370146,1.1494182,1.261822,1.3742256,1.4866294,1.6008459,2.5000753,3.3993049,4.3003473,5.199577,6.1006193,6.1296263,6.1604466,6.189454,6.2202744,6.249282,0.12509441,1.0895905,2.0540867,3.0203958,3.9848917,4.949388,5.4479527,5.9447045,6.4432693,6.9400206,7.4367723,7.166641,6.8983226,6.628191,6.35806,6.0879283,6.869315,7.652515,8.435715,9.217102,10.000301,10.355642,10.70917,11.06451,11.419851,11.775192,12.032633,12.290073,12.547514,12.804955,13.062395,13.390542,13.716875,14.045021,14.373167,14.699501,13.872789,13.044266,12.217555,11.390844,10.56232,11.13159,11.702674,12.271944,12.843027,13.412297,13.232814,13.05333,12.872034,12.692551,12.513068,12.581961,12.652666,12.7233715,12.792264,12.862969,15.198066,17.533161,19.868258,22.203352,24.536636,27.290525,30.042603,32.79468,35.546757,38.300648,41.573044,44.845444,48.11784,51.390236,54.662636,56.778362,58.892277,61.008003,63.121918,65.23765,61.114967,56.99229,52.869614,48.746937,44.62426,43.97522,43.324368,42.675327,42.02447,41.37543,38.03777,34.700104,31.36244,28.024776,24.68711,25.600845,26.512764,27.424685,28.336605,29.250338,27.372108,25.495693,23.617464,21.739235,19.862818,19.85194,19.842875,19.831997,19.822933,19.812056,19.164827,18.5176,17.870373,17.223145,16.575916,15.266958,13.959812,12.652666,11.34552,10.038374,12.349901,14.663241,16.97477,19.288109,21.599636,21.159086,20.72035,20.279799,19.839249,19.400513,17.029158,14.6596155,12.290073,9.920531,7.549176,8.499168,9.449161,10.399154,11.349146,12.299138,12.569269,12.839401,13.109532,13.379663,13.649796,14.039582,14.429369,14.819156,15.208943,15.600543,14.4420595,13.28539,12.126906,10.970237,9.811753,8.887142,7.9625316,7.037921,6.11331,5.186886,4.550536,3.9123733,3.2742105,2.6378605,1.9996977,3.6295512,5.2594047,6.889258,8.519112,10.150778,8.655084,7.159389,5.6655083,4.169814,2.6741197,2.3441606,2.0142014,1.6842422,1.3542831,1.0243238,2.4583774,3.8906176,5.3228583,6.755099,8.187339,8.31062,8.432089,8.55537,8.676839,8.80012,8.974165,9.1500225,9.325879,9.499924,9.675781,10.656594,11.63922,12.621845,13.604471,14.587097,14.362289,14.137483,13.912675,13.687867,13.46306,13.584529,13.70781,13.829279,13.95256,14.075842,13.680615,13.28539,12.890164,12.494938,12.099712,11.477866,10.854207,10.232361,9.610515,8.9868555,8.832754,8.676839,8.5227375,8.366822,8.212721,8.694968,9.177217,9.659465,10.141713,10.625773,11.262123,11.900287,12.538449,13.174799,13.812962,13.140353,12.467744,11.795135,11.122525,10.449916,11.544946,12.639976,13.735004,14.830034,15.925063,17.235836,18.544794,19.855566,21.164526,22.475298,23.815077,25.154856,26.494635,27.834415,29.174194,25.740442,22.304878,18.869314,15.435563,11.999999,12.010877,12.019942,12.03082,12.039885,12.050762,12.28826,12.525759,12.763257,13.000754,13.238253,12.310016,11.381779,10.455356,9.527119,8.600695,10.147152,11.695421,13.2418785,14.790149,16.336605,16.664753,16.992899,17.319231,17.647377,17.975525,17.719896,17.464268,17.210453,16.954826,16.699198,14.104849,11.510499,8.914337,6.319988,3.7256382,3.6694362,3.6150475,3.5606585,3.5044568,3.4500678,3.2669585,3.0856624,2.902553,2.7194438,2.5381477,2.7448254,2.953316,3.159994,3.3666716,3.5751622,4.6575007,5.7398396,6.8221784,7.9045167,8.9868555,8.345067,7.703278,7.059676,6.4178877,5.774286,5.147001,4.519716,3.8924308,3.2651455,2.6378605,2.953316,3.2669585,3.5824142,3.8978696,4.213325,4.269527,4.327542,4.3855567,4.441758,4.499773,3.7256382,2.94969,2.175555,1.3996071,0.62547207,0.7469406,0.87022203,0.9916905,1.114972,1.2382535,1.5555218,1.8727903,2.1900587,2.5073273,2.8245957,3.1799364,3.5352771,3.8906176,4.2441454,4.599486,5.754343,6.9092,8.06587,9.220728,10.375585,9.27693,8.180087,7.083245,5.9845896,4.8877473,5.217706,5.5476656,5.8776245,6.207584,6.5375433,7.440398,8.343254,9.244296,10.147152,11.050007,10.152591,9.255174,8.357758,7.460341,6.5629244,5.3246713,4.0882306,2.8499773,1.6117238,0.37528324,1.8546607,3.3340383,4.8152285,6.294606,7.7757964,7.2754188,6.775041,6.2746634,5.774286,5.275721,5.467895,5.660069,5.8522434,6.0444174,6.2365913,5.823236,5.408067,4.992899,4.5777307,4.162562,3.5044568,2.8481643,2.1900587,1.5319533,0.87566096,0.7777609,0.67986095,0.581961,0.48587397,0.387974,0.3480888,0.30820364,0.26831847,0.22662032,0.18673515,0.17041849,0.15228885,0.13415924,0.11784257,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.045324065,0.052575916,0.059827764,0.06707962,0.07433146,0.07433146,0.07433146,0.07433146,0.07433146,0.07433146,0.13415924,0.19579996,0.25562772,0.3154555,0.37528324,0.2991388,0.22480737,0.15047589,0.07433146,0.0,0.0,0.0,0.0,0.0,0.0,0.11784257,0.23568514,0.35171473,0.46955732,0.5873999,0.5076295,0.42785916,0.3480888,0.26831847,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.03988518,0.054388877,0.07070554,0.08520924,0.099712946,0.092461094,0.08520924,0.07795739,0.07070554,0.06164073,0.054388877,0.047137026,0.03988518,0.032633327,0.025381476,0.030820364,0.034446288,0.03988518,0.045324065,0.05076295,0.30276474,0.55476654,0.80676836,1.0605831,1.3125849,1.6570477,2.0033236,2.3477864,2.6922495,3.0367124,5.4207582,7.802991,10.185224,12.567456,14.94969,11.967366,8.985043,6.002719,3.0203958,0.038072214,0.06164073,0.0870222,0.11240368,0.13778515,0.16316663,0.15954071,0.15772775,0.15410182,0.15228885,0.15047589,0.13053331,0.11059072,0.09064813,0.07070554,0.05076295,0.045324065,0.03988518,0.034446288,0.030820364,0.025381476,0.032633327,0.03988518,0.047137026,0.054388877,0.06164073,0.10696479,0.15228885,0.19761293,0.24293698,0.28826106,0.23024625,0.17223145,0.11421664,0.058014803,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.12328146,0.17041849,0.21755551,0.26469254,0.31182957,0.2574407,0.2030518,0.14684997,0.092461094,0.038072214,0.17585737,0.31182957,0.44961473,0.5873999,0.72518504,0.6327239,0.5402629,0.44780177,0.35534066,0.26287958,0.36984438,0.47680917,0.5855869,0.69255173,0.7995165,1.0950294,1.3905423,1.6842422,1.9797552,2.275268,2.5780327,2.8807976,3.1817493,3.484514,3.787279,4.367427,4.947575,5.527723,6.107871,6.688019,6.833056,6.978093,7.12313,7.268167,7.413204,6.510349,5.6074934,4.704638,3.8017826,2.9007401,2.953316,3.005892,3.056655,3.1092308,3.1618068,3.2143826,3.2669585,3.3195345,3.3721104,3.4246864,4.1281157,4.8297324,5.5331616,6.2347784,6.9382076,5.975525,5.0128417,4.0501585,3.0874753,2.124792,2.4148662,2.70494,2.9950142,3.2850883,3.5751622,3.435564,3.294153,3.1545548,3.0149567,2.8753586,2.819157,2.764768,2.7103791,2.6541772,2.5997884,2.6976883,2.7955883,2.8916752,2.9895754,3.0874753,2.9333735,2.7774587,2.6233568,2.467442,2.3133402,2.2825198,2.2516994,2.222692,2.1918716,2.1628644,2.0903459,2.0178273,1.9453088,1.8727903,1.8002719,1.6642996,1.5301404,1.3941683,1.260009,1.1258497,1.167548,1.209246,1.2527572,1.2944553,1.3379664,1.1548572,0.97174793,0.7904517,0.6073425,0.42423326,0.6200332,0.81583315,1.0098201,1.2056202,1.3996071,1.4503701,1.49932,1.550083,1.6008459,1.649796,2.9369993,4.2260156,5.5132194,6.8004227,8.087626,7.9081426,7.7268467,7.5473633,7.36788,7.1883965,0.06164073,1.3452182,2.6269827,3.9105604,5.1923246,6.4759026,6.967215,7.460341,7.951654,8.444779,8.937905,8.42665,7.9172077,7.407765,6.8983226,6.3870673,6.9092,7.4331465,7.95528,8.477413,8.999546,9.452786,9.904215,10.357455,10.810696,11.262123,10.910409,10.556881,10.205167,9.851639,9.499924,10.21967,10.939416,11.6591625,12.380721,13.100468,12.618219,12.134158,11.651911,11.169662,10.687414,11.273002,11.856775,12.442362,13.027949,13.611723,13.372412,13.1331005,12.891977,12.652666,12.413355,12.5602045,12.707055,12.855718,13.002567,13.149418,15.016769,16.88412,18.753284,20.620636,22.487988,25.120409,27.75283,30.385252,33.017673,35.650097,39.680313,43.71053,47.740746,51.770958,55.799362,57.92053,60.039883,62.159237,64.2804,66.39976,62.15742,57.91509,53.672756,49.430424,45.18809,43.78667,42.387066,40.987457,39.587852,38.188244,35.287502,32.386765,29.487837,26.587097,23.68817,24.413355,25.136726,25.861912,26.587097,27.31228,25.53014,23.747997,21.96404,20.1819,18.399757,19.520168,20.64058,21.759176,22.879587,23.999998,23.519564,23.040941,22.560507,22.08007,21.599636,19.915394,18.22934,16.545097,14.860854,13.174799,13.588155,13.999697,14.413053,14.824595,15.23795,14.13023,13.022511,11.91479,10.80707,9.699349,8.664148,7.6307597,6.5955577,5.560356,4.5251546,4.9620786,5.4008155,5.8377395,6.2746634,6.7115874,6.735156,6.7569118,6.78048,6.8022356,6.8239913,7.019791,7.215591,7.409578,7.605378,7.799365,7.9770355,8.154706,8.3323765,8.510046,8.6877165,7.663393,6.637256,5.612932,4.5867953,3.5624714,3.2633326,2.962381,2.663242,2.3622901,2.0631514,3.3648586,4.666566,5.9700856,7.271793,8.575313,7.2391596,5.904819,4.5704784,3.2343252,1.8999848,1.7730774,1.6443571,1.5174497,1.3905423,1.261822,3.0983531,4.933071,6.7677894,8.602508,10.437225,10.31757,10.197914,10.078259,9.956791,9.837135,9.675781,9.512614,9.349448,9.188094,9.024928,9.759177,10.49524,11.22949,11.965553,12.699803,12.737875,12.774135,12.812206,12.850279,12.888351,12.980812,13.073273,13.165734,13.258195,13.3506565,13.04064,12.730623,12.420607,12.11059,11.800573,11.358211,10.915848,10.471672,10.029309,9.5869465,9.385707,9.182655,8.979604,8.778365,8.575313,9.184468,9.795437,10.4045925,11.015561,11.624716,12.337211,13.049705,13.762199,14.474693,15.187187,14.3079,13.426801,12.547514,11.668227,10.7871275,12.197612,13.608097,15.016769,16.427254,17.837738,18.367125,18.898321,19.427708,19.957092,20.48829,22.181597,23.876717,25.571836,27.266956,28.962078,25.557333,22.15259,18.747847,15.343102,11.938358,11.804199,11.671853,11.539507,11.407161,11.274815,11.325577,11.374527,11.42529,11.47424,11.525003,11.454298,11.385405,11.314699,11.245807,11.175101,11.804199,12.43511,13.064208,13.695119,14.324218,14.706753,15.089288,15.471823,15.854358,16.236893,15.335851,14.432995,13.53014,12.627284,11.724429,10.165281,8.604321,7.0451727,5.484212,3.925064,3.9975824,4.070101,4.1426196,4.215138,4.2876563,3.8398547,3.392053,2.9442513,2.4982624,2.0504606,2.1973107,2.3441606,2.4928236,2.6396735,2.7883365,3.7093215,4.632119,5.5549173,6.4777155,7.400513,7.409578,7.420456,7.4295206,7.440398,7.4494634,6.630004,5.810545,4.989273,4.169814,3.350355,3.5080826,3.6658103,3.8217251,3.9794528,4.137181,4.122677,4.1081734,4.0918565,4.077353,4.062849,3.3122826,2.561716,1.8129625,1.062396,0.31182957,0.58014804,0.8466535,1.114972,1.3832904,1.649796,1.840157,2.030518,2.220879,2.4094272,2.5997884,3.303218,4.004834,4.708264,5.40988,6.11331,7.4277077,8.7421055,10.058316,11.372714,12.687112,11.282066,9.87702,8.471974,7.066928,5.661882,5.2032027,4.74271,4.2822175,3.8217251,3.3630457,5.3573046,7.3515635,9.347635,11.341894,13.337966,11.369088,9.402024,7.4349594,5.467895,3.5008307,2.8626678,2.2245052,1.5881553,0.9499924,0.31182957,1.0895905,1.8673514,2.6451125,3.4228733,4.2006345,4.0120864,3.825351,3.636803,3.4500678,3.2633326,3.4772623,3.6930048,3.9069343,4.122677,4.3366065,4.068288,3.7981565,3.5280252,3.2578938,2.9877625,2.47832,1.9670644,1.4576219,0.9481794,0.43692398,0.39522585,0.35171473,0.3100166,0.26831847,0.22480737,0.23024625,0.23568514,0.23931105,0.24474995,0.25018883,0.21030366,0.17041849,0.13053331,0.09064813,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.047137026,0.045324065,0.04169814,0.03988518,0.038072214,0.05076295,0.06164073,0.07433146,0.0870222,0.099712946,0.1794833,0.25925365,0.34083697,0.42060733,0.50037766,0.40066472,0.2991388,0.19942589,0.099712946,0.0,0.0,0.0,0.0,0.0,0.0,0.065266654,0.13053331,0.19579996,0.25925365,0.3245203,0.3100166,0.2955129,0.27919623,0.26469254,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.01994259,0.027194439,0.034446288,0.04169814,0.05076295,0.052575916,0.054388877,0.058014803,0.059827764,0.06164073,0.052575916,0.04169814,0.032633327,0.02175555,0.012690738,0.014503701,0.018129626,0.01994259,0.02175555,0.025381476,0.15772775,0.29007402,0.4224203,0.55476654,0.6871128,0.98443866,1.2817645,1.5809034,1.8782293,2.175555,3.6857529,5.1941376,6.7043357,8.214534,9.724731,7.7903004,5.8558693,3.919625,1.9851941,0.05076295,0.07433146,0.099712946,0.12509441,0.15047589,0.17585737,0.16679256,0.15954071,0.15228885,0.14503701,0.13778515,0.11421664,0.092461094,0.07070554,0.047137026,0.025381476,0.02175555,0.01994259,0.018129626,0.014503701,0.012690738,0.02175555,0.032633327,0.04169814,0.052575916,0.06164073,0.12328146,0.18310922,0.24293698,0.30276474,0.36259252,0.29007402,0.21755551,0.14503701,0.072518505,0.0,0.0,0.0,0.0,0.0,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.14322405,0.18492219,0.22662032,0.27013144,0.31182957,0.25925365,0.20667773,0.15410182,0.10333887,0.05076295,0.18673515,0.3245203,0.46230546,0.6000906,0.73787576,0.6345369,0.533011,0.42967212,0.32814622,0.22480737,0.3100166,0.39522585,0.48043507,0.5656443,0.6508536,0.79770356,0.9445535,1.0932164,1.2400664,1.3869164,1.8818551,2.3767939,2.8717327,3.3666716,3.8616104,4.552349,5.243088,5.9320135,6.622752,7.311678,7.360628,7.407765,7.454902,7.502039,7.549176,6.6680765,5.7851634,4.902251,4.019338,3.1382382,3.007705,2.8771715,2.7466383,2.617918,2.4873846,2.520018,2.5526514,2.5852847,2.617918,2.6505513,3.2325122,3.8144734,4.3982472,4.9802084,5.562169,4.8877473,4.213325,3.53709,2.8626678,2.1882458,2.3568513,2.5272698,2.6976883,2.8681068,3.0367124,3.0167696,2.9968271,2.9768846,2.956942,2.9369993,2.8971143,2.857229,2.817344,2.7774587,2.7375734,2.7792716,2.8227828,2.864481,2.907992,2.94969,2.810092,2.6704938,2.5308957,2.3894846,2.2498865,2.222692,2.1954978,2.1683033,2.1392958,2.1121013,2.0830941,2.0522738,2.0232663,1.9924458,1.9616255,1.8202144,1.6769904,1.5355793,1.3923552,1.2491312,1.2908293,1.3307146,1.3705997,1.4104849,1.4503701,1.2019942,0.9554313,0.7070554,0.4604925,0.21211663,0.52213323,0.8321498,1.1421664,1.452183,1.7621996,1.7495089,1.7368182,1.7241274,1.7132497,1.7005589,3.3757362,5.050914,6.7242785,8.399456,10.074633,9.684846,9.295059,8.9052725,8.515485,8.125698,0.0,1.6008459,3.199879,4.800725,6.399758,8.000604,8.488291,8.974165,9.461852,9.949538,10.437225,9.686659,8.937905,8.187339,7.4367723,6.688019,6.9508986,7.211965,7.474845,7.7377243,8.000604,8.549932,9.099259,9.6504,10.199727,10.750868,9.788185,8.825501,7.8628187,6.9001355,5.9374523,7.0506115,8.161958,9.275117,10.388275,11.499621,11.361836,11.225864,11.088079,10.950294,10.812509,11.4126,12.012691,12.612781,13.212872,13.812962,13.512011,13.212872,12.91192,12.612781,12.311829,12.536636,12.763257,12.988064,13.212872,13.437678,14.837286,16.236893,17.638313,19.03792,20.437527,22.950293,25.46306,27.975826,30.486778,32.999546,37.78758,42.575615,47.361835,52.149868,56.937904,59.062695,61.18749,63.31228,65.43707,67.56187,63.199875,58.837887,54.474087,50.1121,45.75011,43.599937,41.449764,39.29959,37.149418,34.99924,32.53724,30.075235,27.613234,25.149418,22.687414,23.225864,23.7625,24.299137,24.837587,25.374224,23.68817,22.000301,20.312433,18.624565,16.936697,19.186583,21.438282,23.68817,25.938055,28.187943,27.8743,27.56247,27.25064,26.936998,26.625168,24.562017,22.500679,20.437527,18.374376,16.313038,14.824595,13.337966,11.849524,10.362894,8.874452,7.0995617,5.3246713,3.5497808,1.7748904,0.0,0.2991388,0.6000906,0.89922947,1.2001812,1.49932,1.4249886,1.3506571,1.2745126,1.2001812,1.1258497,0.89922947,0.6744221,0.44961473,0.22480737,0.0,0.0,0.0,0.0,0.0,0.0,1.5120108,3.0258346,4.537845,6.049856,7.5618668,6.43783,5.3119802,4.1879435,3.0620937,1.938057,1.9743162,2.0123885,2.0504606,2.08672,2.124792,3.100166,4.07554,5.050914,6.0244746,6.9998484,5.825049,4.650249,3.4754493,2.3006494,1.1258497,1.2001812,1.2745126,1.3506571,1.4249886,1.49932,3.738329,5.975525,8.212721,10.449916,12.687112,12.32452,11.961927,11.599335,11.236742,10.874149,10.375585,9.875207,9.374829,8.874452,8.375887,8.861761,9.349448,9.837135,10.324821,10.812509,11.111648,11.4126,11.711739,12.012691,12.311829,12.375282,12.436923,12.500377,12.562017,12.625471,12.400664,12.175857,11.949236,11.724429,11.499621,11.236742,10.975676,10.712796,10.449916,10.1870365,9.936848,9.686659,9.438283,9.188094,8.937905,9.675781,10.411844,11.14972,11.887595,12.625471,13.412297,14.199123,14.9877615,15.774588,16.563227,15.475449,14.387671,13.299893,12.212116,11.124338,12.850279,14.574407,16.300346,18.024473,19.750414,19.500225,19.250036,18.999847,18.749659,18.49947,20.54993,22.600391,24.650852,26.6995,28.74996,25.374224,22.000301,18.624565,15.250641,11.874905,11.599335,11.325577,11.050007,10.774437,10.500679,10.362894,10.225109,10.087324,9.949538,9.811753,10.600392,11.3872175,12.175857,12.962683,13.749508,13.46306,13.174799,12.888351,12.60009,12.311829,12.750566,13.1874895,13.6244135,14.06315,14.500074,12.949992,11.399909,9.849826,8.299743,6.7496595,6.2257137,5.6999545,5.1741953,4.650249,4.12449,4.325729,4.5251546,4.7245803,4.9258194,5.125245,4.4127507,3.7002566,2.9877625,2.275268,1.5627737,1.649796,1.7368182,1.8256533,1.9126755,1.9996977,2.762955,3.5243993,4.2876563,5.050914,5.812358,6.474089,7.137634,7.799365,8.46291,9.12464,8.113008,7.0995617,6.0879283,5.0744824,4.062849,4.062849,4.062849,4.062849,4.062849,4.062849,3.975827,3.8869917,3.7999697,3.7129474,3.6241121,2.9007401,2.175555,1.4503701,0.72518504,0.0,0.41335547,0.824898,1.2382535,1.649796,2.0631514,2.124792,2.1882458,2.2498865,2.3133402,2.374981,3.4246864,4.4743915,5.52591,6.5756154,7.6253204,9.099259,10.57501,12.050762,13.524701,15.000452,13.287203,11.575767,9.862516,8.149267,6.43783,5.186886,3.9377546,2.6868105,1.4376793,0.18673515,3.2760234,6.3616858,9.4509735,12.538449,15.624111,12.5873995,9.550687,6.5121617,3.4754493,0.43692398,0.40066472,0.36259252,0.3245203,0.28826106,0.25018883,0.3245203,0.40066472,0.4749962,0.5493277,0.62547207,0.7505665,0.87566096,1.0007553,1.1258497,1.2491312,1.4866294,1.7241274,1.9616255,2.1991236,2.4366217,2.3133402,2.1882458,2.0631514,1.938057,1.8129625,1.4503701,1.0877775,0.72518504,0.36259252,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.11240368,0.16316663,0.21211663,0.26287958,0.31182957,0.25018883,0.18673515,0.12509441,0.06164073,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.22480737,0.3245203,0.42423326,0.52575916,0.62547207,0.50037766,0.37528324,0.25018883,0.12509441,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.11240368,0.16316663,0.21211663,0.26287958,0.31182957,0.25018883,0.18673515,0.12509441,0.06164073,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.31182957,0.5620184,0.8122072,1.062396,1.3125849,1.9507477,2.5870976,3.2252605,3.8616104,4.499773,3.6132345,2.7248828,1.8383441,0.9499924,0.06164073,0.0870222,0.11240368,0.13778515,0.16316663,0.18673515,0.17585737,0.16316663,0.15047589,0.13778515,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.13778515,0.21211663,0.28826106,0.36259252,0.43692398,0.34990177,0.26287958,0.17585737,0.0870222,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.16316663,0.19942589,0.2374981,0.2755703,0.31182957,0.26287958,0.21211663,0.16316663,0.11240368,0.06164073,0.19942589,0.33721104,0.4749962,0.61278135,0.7505665,0.63816285,0.52575916,0.41335547,0.2991388,0.18673515,0.25018883,0.31182957,0.37528324,0.43692398,0.50037766,0.50037766,0.50037766,0.50037766,0.50037766,0.50037766,1.1874905,1.8746033,2.561716,3.2506418,3.9377546,4.7372713,5.5367875,6.338117,7.137634,7.93715,7.8882003,7.837437,7.7866745,7.7377243,7.686961,6.825804,5.962834,5.0998635,4.2368937,3.3757362,3.0620937,2.7502642,2.4366217,2.124792,1.8129625,1.8256533,1.8383441,1.8492218,1.8619126,1.8746033,2.3369088,2.7992141,3.2633326,3.7256382,4.1879435,3.7999697,3.4119956,3.0258346,2.6378605,2.2498865,2.3006494,2.3495996,2.4003625,2.4493124,2.5000753,2.5997884,2.6995013,2.7992141,2.9007401,3.000453,2.9750717,2.94969,2.9243085,2.9007401,2.8753586,2.8626678,2.8499773,2.8372865,2.8245957,2.811905,2.6868105,2.561716,2.4366217,2.3133402,2.1882458,2.1628644,2.137483,2.1121013,2.08672,2.0631514,2.0758421,2.08672,2.0994108,2.1121013,2.124792,1.9743162,1.8256533,1.6751775,1.5247015,1.3742256,1.4122978,1.4503701,1.4866294,1.5247015,1.5627737,1.2491312,0.93730164,0.62547207,0.31182957,0.0,0.42423326,0.85027945,1.2745126,1.7005589,2.124792,2.0504606,1.9743162,1.8999848,1.8256533,1.7495089,3.8126602,5.8758116,7.93715,10.000301,12.06164,11.463363,10.863272,10.263181,9.663091,9.063,0.43692398,1.7966459,3.1581807,4.517903,5.8776245,7.2373466,7.610817,7.9824743,8.354132,8.727602,9.099259,8.510046,7.9208336,7.3298078,6.740595,6.149569,6.24203,6.3344913,6.4269524,6.5194135,6.6118746,7.135821,7.6579537,8.180087,8.70222,9.224354,8.4756,7.7250338,6.9744673,6.2257137,5.475147,6.78048,8.0858135,9.389333,10.694666,11.999999,11.628342,11.254871,10.883214,10.509744,10.138086,10.857833,11.5775795,12.297325,13.017072,13.736817,13.44493,13.153044,12.859344,12.567456,12.27557,12.456866,12.639976,12.823084,13.00438,13.1874895,14.248073,15.306843,16.367426,17.428009,18.48678,20.437527,22.388275,24.33721,26.287958,28.236893,32.510044,36.7832,41.05454,45.32769,49.60084,52.012085,54.425137,56.83819,59.24943,61.662483,58.187035,54.713398,51.23795,47.7625,44.28705,42.443268,40.59767,38.752075,36.90829,35.062695,31.759478,28.458075,25.154856,21.851639,18.550234,18.97084,19.389635,19.810242,20.23085,20.649643,19.402325,18.155006,16.907688,15.660371,14.413053,16.80979,19.208338,21.605076,24.001812,26.400362,26.347786,26.29521,26.242634,26.190058,26.137482,24.480434,22.823385,21.164526,19.507477,17.85043,15.700256,13.550082,11.399909,9.249735,7.0995617,5.6800117,4.2604623,2.8390994,1.4195497,0.0,0.26287958,0.52575916,0.7868258,1.0497054,1.3125849,1.2473183,1.1820517,1.1167849,1.0533313,0.9880646,0.7904517,0.59283876,0.39522585,0.19761293,0.0,0.0,0.0,0.0,0.0,0.0,1.209246,2.420305,3.6295512,4.84061,6.049856,5.4570174,4.8641787,4.273153,3.680314,3.0874753,3.4555066,3.8217251,4.1897564,4.557788,4.9258194,5.91751,6.9092,7.902704,8.894395,9.8878975,8.225411,6.5629244,4.900438,3.2379513,1.5754645,1.7875811,1.9996977,2.2118144,2.4257438,2.6378605,4.7227674,6.8076744,8.892582,10.9774885,13.062395,12.826711,12.592838,12.357153,12.123281,11.887595,11.651911,11.418038,11.182353,10.946668,10.712796,11.129777,11.546759,11.965553,12.382534,12.799516,12.92461,13.049705,13.174799,13.299893,13.424988,13.3506565,13.274512,13.200181,13.125849,13.049705,12.806767,12.565643,12.322706,12.07977,11.836833,11.615651,11.392657,11.169662,10.946668,10.725487,10.80707,10.890467,10.97205,11.055446,11.137029,11.7679405,12.397038,13.027949,13.657047,14.287958,15.062093,15.838041,16.612177,17.388124,18.16226,17.315605,16.467138,15.620485,14.772019,13.925365,14.819156,15.71476,16.610363,17.504154,18.399757,18.412449,18.425138,18.43783,18.45052,18.463211,19.812056,21.162712,22.513369,23.862213,25.212872,22.266806,19.322556,16.378304,13.43224,10.487988,10.1326475,9.7773075,9.421967,9.066626,8.713099,8.662335,8.613385,8.562622,8.511859,8.46291,9.987611,11.512312,13.037014,14.561715,16.08823,15.000452,13.912675,12.824898,11.73712,10.649343,11.91479,13.180238,14.445685,15.709321,16.97477,14.935185,12.895603,10.854207,8.814624,6.775041,6.35806,5.9392653,5.522284,5.105303,4.688321,4.664753,4.6429973,4.6194286,4.597673,4.574105,4.0918565,3.6096084,3.1273603,2.6451125,2.1628644,2.0957847,2.0268922,1.9598125,1.892733,1.8256533,2.617918,3.4101827,4.2024474,4.994712,5.7869763,6.096993,6.4070096,6.717026,7.027043,7.3370595,6.542982,5.7470913,4.953014,4.157123,3.3630457,3.437377,3.5117085,3.587853,3.6621845,3.738329,3.6041696,3.4718235,3.339477,3.207131,3.0747845,2.4819458,1.8909199,1.2980812,0.70524246,0.11240368,0.48587397,0.8575313,1.2291887,1.6026589,1.9743162,1.9906329,2.0051367,2.0196402,2.034144,2.0504606,3.0675328,4.0846047,5.101677,6.1205616,7.137634,8.99592,10.852394,12.710681,14.567154,16.425442,14.376793,12.329959,10.283124,8.234476,6.187641,5.1596913,4.1317415,3.105605,2.077655,1.0497054,3.3630457,5.674573,7.987913,10.29944,12.612781,10.226922,7.842876,5.4570174,3.0729716,0.6871128,0.8901646,1.0932164,1.2944553,1.4975071,1.7005589,1.7621996,1.8256533,1.887294,1.9507477,2.0123885,2.5798457,3.147303,3.7147603,4.2822175,4.8496747,4.8732433,4.894999,4.9167547,4.940323,4.9620786,4.273153,3.5824142,2.8916752,2.2027495,1.5120108,1.2400664,0.968122,0.69436467,0.4224203,0.15047589,0.13778515,0.12509441,0.11240368,0.099712946,0.0870222,0.12509441,0.16316663,0.19942589,0.2374981,0.2755703,0.21936847,0.16497959,0.11059072,0.054388877,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.19036107,0.26831847,0.3444629,0.4224203,0.50037766,0.40066472,0.2991388,0.19942589,0.099712946,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.09064813,0.13053331,0.17041849,0.21030366,0.25018883,0.23931105,0.23024625,0.21936847,0.21030366,0.19942589,0.15954071,0.11965553,0.07977036,0.03988518,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.42967212,0.8103943,1.1893034,1.5700256,1.9507477,3.9558845,5.959208,7.9643445,9.969481,11.974618,9.684846,7.3950744,5.105303,2.8155308,0.52575916,0.44961473,0.37528324,0.2991388,0.22480737,0.15047589,0.15410182,0.15954071,0.16497959,0.17041849,0.17585737,0.15772775,0.13959812,0.12328146,0.10515183,0.0870222,0.07070554,0.052575916,0.034446288,0.018129626,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.14322405,0.21030366,0.27738327,0.3444629,0.41335547,0.33177215,0.2520018,0.17223145,0.092461094,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.038072214,0.06164073,0.0870222,0.11240368,0.13778515,0.17585737,0.21211663,0.25018883,0.28826106,0.3245203,0.2755703,0.22480737,0.17585737,0.12509441,0.07433146,0.19579996,0.3154555,0.43511102,0.55476654,0.6744221,0.5855869,0.4949388,0.40429065,0.3154555,0.22480737,0.3045777,0.38434806,0.46411842,0.54570174,0.62547207,0.6000906,0.5747091,0.5493277,0.52575916,0.50037766,1.1367276,1.7748904,2.4130533,3.049403,3.6875658,4.3982472,5.1071157,5.8177967,6.526665,7.2373466,7.1883965,7.137634,7.0868707,7.037921,6.987158,6.3671246,5.7470913,5.127058,4.507025,3.8869917,3.4772623,3.0675328,2.657803,2.2480736,1.8383441,1.8147756,1.79302,1.7694515,1.7476959,1.7241274,2.1556125,2.5852847,3.0149567,3.444629,3.874301,3.5443418,3.2143826,2.8844235,2.5544643,2.2245052,2.2933977,2.3604772,2.427557,2.4946365,2.561716,2.659616,2.7575161,2.855416,2.953316,3.049403,3.0222087,2.9950142,2.9678197,2.9406252,2.911618,2.9243085,2.9369993,2.94969,2.962381,2.9750717,2.8517902,2.7303216,2.6070402,2.4855716,2.3622901,2.3042755,2.2480736,2.1900587,2.132044,2.0758421,2.0577126,2.039583,2.0232663,2.0051367,1.987007,1.8582866,1.7277533,1.5972201,1.4666867,1.3379664,1.3270886,1.3180238,1.3071461,1.2980812,1.2872034,1.1349145,0.9826257,0.83033687,0.678048,0.52575916,1.0841516,1.6443571,2.2045624,2.764768,3.3249733,3.141864,2.960568,2.7774587,2.5943494,2.4130533,4.2477713,6.0824895,7.9172077,9.751925,11.586644,10.765372,9.9422865,9.119202,8.29793,7.474845,0.87566096,1.9942589,3.1146698,4.2350807,5.3554916,6.474089,6.733343,6.9907837,7.2482243,7.5056653,7.763106,7.3316207,6.9019485,6.472276,6.0426044,5.612932,5.5349746,5.4570174,5.3808727,5.3029156,5.224958,5.719897,6.2148356,6.7097745,7.2047133,7.699652,7.1630154,6.624565,6.0879283,5.5494785,5.0128417,6.510349,8.007855,9.5053625,11.00287,12.500377,11.893035,11.285692,10.6783495,10.069194,9.461852,10.303066,11.142468,11.98187,12.823084,13.662486,13.377851,13.093216,12.806767,12.522133,12.237497,12.377095,12.516694,12.658105,12.797703,12.937301,13.657047,14.376793,15.098352,15.818098,16.537846,17.92476,19.311678,20.700407,22.087322,23.47424,27.232512,30.98897,34.747242,38.505512,42.26197,44.963284,47.662785,50.36229,53.06179,55.763103,53.174194,50.587093,47.999996,45.4129,42.8258,41.284782,39.74558,38.20456,36.665356,35.124336,30.981718,26.840912,22.696478,18.555672,14.413053,14.715817,15.016769,15.319533,15.622298,15.925063,15.118295,14.309713,13.502945,12.694364,11.887595,14.432995,16.976582,19.52198,22.06738,24.61278,24.819458,25.027948,25.234627,25.443117,25.649796,24.397038,23.14428,21.893335,20.64058,19.387821,16.575916,13.762199,10.950294,8.136576,5.3246713,4.2604623,3.1944401,2.1302311,1.064209,0.0,0.22480737,0.44961473,0.6744221,0.89922947,1.1258497,1.0696479,1.015259,0.96087015,0.90466833,0.85027945,0.67986095,0.5094425,0.34083697,0.17041849,0.0,0.0,0.0,0.0,0.0,0.0,0.90829426,1.8147756,2.72307,3.6295512,4.537845,4.478018,4.41819,4.358362,4.2967215,4.2368937,4.934884,5.632875,6.3308654,7.027043,7.7250338,8.734854,9.744674,10.754494,11.764315,12.774135,10.625773,8.4756,6.3254266,4.175253,2.0250793,2.374981,2.7248828,3.0747845,3.4246864,3.774588,5.7072062,7.6398244,9.572442,11.50506,13.437678,13.330714,13.221936,13.114971,13.008006,12.899229,12.930049,12.96087,12.989877,13.020698,13.049705,13.397794,13.745882,14.092158,14.440247,14.788336,14.737573,14.68681,14.63786,14.587097,14.538147,14.324218,14.112101,13.899984,13.687867,13.475751,13.2146845,12.955431,12.694364,12.43511,12.175857,11.992747,11.809638,11.628342,11.445232,11.262123,11.677292,12.092461,12.507628,12.922797,13.337966,13.860099,14.382232,14.904366,15.428311,15.950445,16.71189,17.475147,18.238403,18.999847,19.763105,19.155762,18.54842,17.939264,17.331923,16.72458,16.789846,16.855114,16.92038,16.985647,17.0491,17.32467,17.60024,17.87581,18.149569,18.425138,19.074179,19.725033,20.375887,21.024927,21.675781,19.15939,16.64481,14.13023,11.615651,9.099259,8.664148,8.23085,7.795739,7.360628,6.925517,6.9617763,6.9998484,7.037921,7.07418,7.112252,9.374829,11.637406,13.899984,16.162561,18.425138,16.537846,14.650551,12.763257,10.874149,8.9868555,11.080828,13.172986,15.265145,17.357304,19.449463,16.92038,14.389484,11.860401,9.329506,6.8004227,6.490406,6.1803894,5.870373,5.560356,5.2503395,5.0055895,4.76084,4.514277,4.269527,4.024777,3.7727752,3.5207734,3.2669585,3.0149567,2.762955,2.5399606,2.3169663,2.0957847,1.8727903,1.649796,2.472881,3.294153,4.117238,4.940323,5.7615952,5.719897,5.678199,5.634688,5.5929894,5.5494785,4.972956,4.3946214,3.8180993,3.2397642,2.663242,2.811905,2.962381,3.1128569,3.2633326,3.4119956,3.2343252,3.056655,2.8807976,2.7031271,2.525457,2.0649643,1.6044719,1.1457924,0.6852999,0.22480737,0.55839247,0.8901646,1.2219368,1.5555218,1.887294,1.8546607,1.8220274,1.789394,1.7567607,1.7241274,2.7103791,3.6948178,4.6792564,5.6655083,6.6499467,8.890768,11.129777,13.370599,15.609608,17.85043,15.468197,13.085964,10.701918,8.319685,5.9374523,5.132497,4.327542,3.5225863,2.7176309,1.9126755,3.4500678,4.98746,6.5248523,8.062244,9.599637,7.8682575,6.1350656,4.401873,2.6704938,0.93730164,1.3796645,1.8220274,2.2643902,2.7067533,3.149116,3.199879,3.2506418,3.299592,3.350355,3.3993049,4.410938,5.4207582,6.430578,7.440398,8.450218,8.258044,8.06587,7.8718834,7.6797094,7.4875355,6.2329655,4.9783955,3.7220123,2.467442,1.2128719,1.0297627,0.8466535,0.6653573,0.48224804,0.2991388,0.26287958,0.22480737,0.18673515,0.15047589,0.11240368,0.13778515,0.16316663,0.18673515,0.21211663,0.2374981,0.19036107,0.14322405,0.09427405,0.047137026,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.15410182,0.21030366,0.26469254,0.3208944,0.37528324,0.2991388,0.22480737,0.15047589,0.07433146,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.06707962,0.09789998,0.12690738,0.15772775,0.18673515,0.23024625,0.27194437,0.3154555,0.35715362,0.40066472,0.3208944,0.23931105,0.15954071,0.07977036,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.5475147,1.0569572,1.5682126,2.077655,2.5870976,5.961021,9.333132,12.705242,16.077353,19.449463,15.756457,12.065266,8.372261,4.6792564,0.9880646,0.8122072,0.63816285,0.46230546,0.28826106,0.11240368,0.13415924,0.15772775,0.1794833,0.2030518,0.22480737,0.21574254,0.20486477,0.19579996,0.18492219,0.17585737,0.13959812,0.10515183,0.07070554,0.034446288,0.0,0.018129626,0.034446288,0.052575916,0.07070554,0.0870222,0.14684997,0.20667773,0.26831847,0.32814622,0.387974,0.3154555,0.24293698,0.17041849,0.09789998,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.15047589,0.18673515,0.22480737,0.26287958,0.2991388,0.33721104,0.28826106,0.2374981,0.18673515,0.13778515,0.0870222,0.19036107,0.291887,0.39522585,0.49675176,0.6000906,0.533011,0.46411842,0.39703882,0.32995918,0.26287958,0.36077955,0.45686656,0.55476654,0.6526665,0.7505665,0.69980353,0.6508536,0.6000906,0.5493277,0.50037766,1.0877775,1.6751775,2.2625773,2.8499773,3.437377,4.0574102,4.6774435,5.297477,5.91751,6.5375433,6.48678,6.43783,6.3870673,6.338117,6.2873545,5.910258,5.5331616,5.1542525,4.7771564,4.40006,3.8924308,3.3848011,2.8771715,2.3695421,1.8619126,1.8057107,1.7476959,1.6896812,1.6316663,1.5754645,1.9725033,2.3695421,2.7683938,3.1654327,3.5624714,3.290527,3.0167696,2.7448254,2.472881,2.1991236,2.2843328,2.3695421,2.4547513,2.5399606,2.6251698,2.7194438,2.8155308,2.909805,3.005892,3.100166,3.0693457,3.0403383,3.009518,2.9805105,2.94969,2.9877625,3.0258346,3.0620937,3.100166,3.1382382,3.0167696,2.8971143,2.7774587,2.657803,2.5381477,2.4474995,2.3568513,2.268016,2.1773682,2.08672,2.039583,1.9924458,1.9453088,1.8981718,1.8492218,1.7404441,1.6298534,1.5192627,1.4104849,1.2998942,1.2418793,1.1856775,1.1276628,1.0696479,1.0116332,1.020698,1.0279498,1.0352017,1.0424535,1.0497054,1.745883,2.4402475,3.1346123,3.83079,4.5251546,4.2350807,3.9450066,3.6549325,3.3648586,3.0747845,4.6828823,6.2909803,7.897265,9.5053625,11.111648,10.067381,9.023115,7.9770355,6.932769,5.8866897,1.3125849,2.1918716,3.0729716,3.9522583,4.8333583,5.712645,5.8558693,5.99728,6.1405044,6.281915,6.4251394,6.155008,5.8848767,5.614745,5.3446136,5.0744824,4.8279195,4.5795436,4.3329806,4.0846047,3.8380418,4.305786,4.7717175,5.239462,5.7072062,6.1749506,5.8504305,5.524097,5.199577,4.8750563,4.550536,6.240217,7.9298983,9.619579,11.30926,13.000754,12.157727,11.314699,10.471672,9.630457,8.78743,9.7483,10.707357,11.668227,12.627284,13.588155,13.310771,13.033388,12.754191,12.476809,12.199425,12.297325,12.395226,12.493125,12.589212,12.687112,13.067834,13.446743,13.827466,14.208188,14.587097,15.411995,16.236893,17.06179,17.886688,18.711586,21.954977,25.196554,28.439943,31.68152,34.92491,37.912674,40.900436,43.8882,46.87415,49.86191,48.163162,46.462605,44.762047,43.0633,41.36274,40.128113,38.891674,37.657047,36.422417,35.18779,30.20577,25.221935,20.239914,15.257894,10.274059,10.4589815,10.645717,10.830639,11.015561,11.200482,10.832452,10.46442,10.098202,9.73017,9.362139,12.054388,14.746637,17.4407,20.13295,22.8252,23.292944,23.760687,24.22662,24.694363,25.162107,24.315454,23.466988,22.620335,21.771868,20.925215,17.449764,13.974316,10.500679,7.02523,3.5497808,2.8390994,2.1302311,1.4195497,0.7106813,0.0,0.18673515,0.37528324,0.5620184,0.7505665,0.93730164,0.8919776,0.8466535,0.8031424,0.75781834,0.7124943,0.56927025,0.42785916,0.28463513,0.14322405,0.0,0.0,0.0,0.0,0.0,0.0,0.6055295,1.209246,1.8147756,2.420305,3.0258346,3.4972048,3.9703882,4.441758,4.914942,5.388125,6.414262,7.4422116,8.470161,9.498111,10.524248,11.552197,12.580148,13.608097,14.634234,15.662184,13.024323,10.388275,7.750415,5.1125546,2.474694,2.962381,3.4500678,3.9377546,4.4254417,4.9131284,6.6916447,8.471974,10.252303,12.032633,13.812962,13.832905,13.852847,13.872789,13.892733,13.912675,14.208188,14.501887,14.7974,15.092914,15.388427,15.66581,15.9431925,16.220575,16.49796,16.775343,16.550535,16.325727,16.100922,15.8743,15.649493,15.299591,14.94969,14.599788,14.249886,13.899984,13.622601,13.345218,13.067834,12.790451,12.513068,12.3698435,12.22662,12.085209,11.941984,11.800573,12.547514,13.294455,14.043208,14.790149,15.537089,15.952258,16.367426,16.782595,17.197763,17.612932,18.361685,19.112251,19.862818,20.613384,21.362139,20.99592,20.627888,20.259857,19.891825,19.525606,18.760536,17.995466,17.230396,16.465326,15.700256,16.236893,16.775343,17.31198,17.85043,18.387066,18.338116,18.287354,18.236591,18.187641,18.136877,16.051971,13.967064,11.882156,9.79725,7.7123427,7.1974616,6.68258,6.167699,5.6528172,5.137936,5.2630305,5.388125,5.5132194,5.638314,5.7615952,8.762048,11.762501,14.762955,17.763407,20.762047,18.075237,15.388427,12.699803,10.012992,7.324369,10.245051,13.165734,16.084604,19.005287,21.92597,18.905573,15.885179,12.864782,9.844387,6.825804,6.622752,6.4197006,6.2166486,6.01541,5.812358,5.3446136,4.876869,4.409125,3.9431937,3.4754493,3.4518807,3.4301252,3.4083695,3.3848011,3.3630457,2.9841363,2.6070402,2.229944,1.8528478,1.4757515,2.327844,3.1799364,4.0320287,4.8841214,5.7380266,5.3428006,4.947575,4.552349,4.157123,3.7618973,3.4029307,3.0421512,2.6831846,2.322405,1.9616255,2.1882458,2.4130533,2.6378605,2.8626678,3.0874753,2.864481,2.6432993,2.420305,2.1973107,1.9743162,1.647983,1.3198367,0.9916905,0.6653573,0.33721104,0.630911,0.922798,1.214685,1.5083848,1.8002719,1.7205015,1.6407311,1.5591478,1.4793775,1.3996071,2.3532255,3.3050308,4.256836,5.2104545,6.16226,8.785617,11.407161,14.030518,16.652061,19.275417,16.557787,13.840157,11.122525,8.404895,5.6872635,5.105303,4.5233417,3.9395678,3.3576066,2.7756457,3.53709,4.3003473,5.0617914,5.825049,6.588306,5.5077806,4.4272547,3.346729,2.268016,1.1874905,1.8691645,2.5526514,3.2343252,3.917812,4.599486,4.6375585,4.6756306,4.7118897,4.749962,4.788034,6.240217,7.6924005,9.144584,10.596766,12.050762,11.642846,11.234929,10.827013,10.420909,10.012992,8.192778,6.3725634,4.552349,2.7321346,0.9119202,0.8194591,0.726998,0.6345369,0.5420758,0.44961473,0.387974,0.3245203,0.26287958,0.19942589,0.13778515,0.15047589,0.16316663,0.17585737,0.18673515,0.19942589,0.15954071,0.11965553,0.07977036,0.03988518,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.018129626,0.034446288,0.052575916,0.07070554,0.0870222,0.11965553,0.15228885,0.18492219,0.21755551,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.045324065,0.065266654,0.08520924,0.10515183,0.12509441,0.21936847,0.3154555,0.40972954,0.5058166,0.6000906,0.48043507,0.36077955,0.23931105,0.11965553,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.6653573,1.305333,1.9453088,2.5852847,3.2252605,7.9661574,12.705242,17.446138,22.185223,26.92612,21.829882,16.735458,11.63922,6.544795,1.4503701,1.1747998,0.89922947,0.62547207,0.34990177,0.07433146,0.11421664,0.15410182,0.19579996,0.23568514,0.2755703,0.27194437,0.27013144,0.26831847,0.26469254,0.26287958,0.21030366,0.15772775,0.10515183,0.052575916,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.15228885,0.20486477,0.2574407,0.3100166,0.36259252,0.29732585,0.23205921,0.16679256,0.10333887,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.06164073,0.0870222,0.11240368,0.13778515,0.16316663,0.19942589,0.2374981,0.2755703,0.31182957,0.34990177,0.2991388,0.25018883,0.19942589,0.15047589,0.099712946,0.18492219,0.27013144,0.35534066,0.4405499,0.52575916,0.48043507,0.43511102,0.38978696,0.3444629,0.2991388,0.41516843,0.5293851,0.64541465,0.75963134,0.87566096,0.7995165,0.72518504,0.6508536,0.5747091,0.50037766,1.0370146,1.5754645,2.1121013,2.6505513,3.1871881,3.7183862,4.2477713,4.7771564,5.3083544,5.8377395,5.7869763,5.7380266,5.6872635,5.638314,5.5875506,5.4515786,5.317419,5.18326,5.047288,4.9131284,4.307599,3.7020695,3.0983531,2.4928236,1.887294,1.794833,1.7023718,1.6099107,1.5174497,1.4249886,1.789394,2.1556125,2.520018,2.8844235,3.2506418,3.0348995,2.819157,2.6052272,2.3894846,2.175555,2.277081,2.38042,2.4819458,2.5852847,2.6868105,2.7792716,2.8717327,2.9641938,3.056655,3.149116,3.1182957,3.0856624,3.053029,3.0203958,2.9877625,3.049403,3.1128569,3.1744974,3.2379513,3.299592,3.1817493,3.0657198,2.9478772,2.8300345,2.712192,2.5907235,2.467442,2.3441606,2.222692,2.0994108,2.0232663,1.9453088,1.8673514,1.789394,1.7132497,1.6226015,1.5319533,1.4431182,1.35247,1.261822,1.1566701,1.0533313,0.9481794,0.8430276,0.73787576,0.90466833,1.0732739,1.2400664,1.4068589,1.5754645,2.4058013,3.2343252,4.064662,4.894999,5.7253356,5.328297,4.9294453,4.5324063,4.135368,3.738329,5.1179934,6.497658,7.877322,9.256987,10.636651,9.3693905,8.10213,6.834869,5.567608,4.3003473,1.7495089,2.3894846,3.0294604,3.6694362,4.309412,4.949388,4.976582,5.0055895,5.032784,5.0599785,5.087173,4.976582,4.8678045,4.7572136,4.646623,4.537845,4.120864,3.7020695,3.2850883,2.8681068,2.4493124,2.8898623,3.3304121,3.7691493,4.209699,4.650249,4.537845,4.4254417,4.313038,4.2006345,4.0882306,5.9700856,7.851941,9.735609,11.617464,13.499319,12.42242,11.34552,10.266808,9.189907,8.113008,9.19172,10.272246,11.352772,12.433297,13.512011,13.2418785,12.971747,12.701616,12.433297,12.163166,12.217555,12.271944,12.328146,12.382534,12.436923,12.476809,12.516694,12.556579,12.598277,12.638163,12.899229,13.162108,13.424988,13.687867,13.9507475,16.677443,19.404139,22.132647,24.859343,27.587852,30.862062,34.138084,37.412296,40.68832,43.96253,43.150322,42.338116,41.524094,40.711887,39.89968,38.96963,38.03958,37.10953,36.17948,35.24943,29.428009,23.604773,17.781536,11.9601145,6.1368785,6.205771,6.2728505,6.33993,6.4070096,6.474089,6.546608,6.6191263,6.6916447,6.7641635,6.836682,9.677594,12.516694,15.357606,18.196705,21.037619,21.764616,22.491613,23.220425,23.947422,24.674421,24.232058,23.789696,23.347332,22.90497,22.462606,18.325426,14.188245,10.049252,5.9120708,1.7748904,1.4195497,1.064209,0.7106813,0.35534066,0.0,0.15047589,0.2991388,0.44961473,0.6000906,0.7505665,0.71430725,0.67986095,0.64541465,0.6091554,0.5747091,0.4604925,0.3444629,0.23024625,0.11421664,0.0,0.0,0.0,0.0,0.0,0.0,0.30276474,0.6055295,0.90829426,1.209246,1.5120108,2.518205,3.5225863,4.5269675,5.5331616,6.5375433,7.895452,9.253361,10.609457,11.967366,13.325275,14.369541,15.415621,16.459887,17.505966,18.550234,15.4246855,12.300951,9.175404,6.049856,2.9243085,3.5497808,4.175253,4.800725,5.424384,6.049856,7.6778965,9.304124,10.932164,12.5602045,14.188245,14.335095,14.481945,14.630608,14.777458,14.924308,15.484513,16.04472,16.604925,17.16513,17.725336,17.932013,18.140503,18.347181,18.555672,18.76235,18.361685,17.962833,17.562168,17.163317,16.762651,16.274965,15.787278,15.299591,14.811904,14.324218,14.030518,13.735004,13.439491,13.145792,12.850279,12.74694,12.645414,12.542075,12.440549,12.337211,13.417736,14.498261,15.576975,16.6575,17.738026,18.044416,18.352621,18.660824,18.967215,19.275417,20.013294,20.749357,21.487232,22.22511,22.962984,22.834263,22.707355,22.580448,22.451729,22.324821,20.729414,19.13582,17.540413,15.945006,14.349599,15.149116,15.950445,16.749962,17.549479,18.350807,17.60024,16.849674,16.099108,15.350354,14.599788,12.944552,11.289318,9.634083,7.9806614,6.3254266,5.730775,5.1343102,4.539658,3.9450066,3.350355,3.5624714,3.774588,3.9867048,4.2006345,4.4127507,8.149267,11.887595,15.625924,19.36244,23.100769,19.612629,16.124489,12.638163,9.1500225,5.661882,9.409276,13.15667,16.905876,20.653269,24.400663,20.890768,17.380873,13.8691635,10.359268,6.849373,6.755099,6.6608243,6.5647373,6.4704633,6.3743763,5.6854506,4.994712,4.305786,3.6150475,2.9243085,3.1327994,3.339477,3.5479677,3.7546456,3.9631362,3.4301252,2.8971143,2.3641033,1.8329052,1.2998942,2.182807,3.0657198,3.9468195,4.8297324,5.712645,4.9657044,4.216951,3.4700103,2.72307,1.9743162,1.8329052,1.6896812,1.54827,1.405046,1.261822,1.5627737,1.8619126,2.1628644,2.4620032,2.762955,2.4946365,2.228131,1.9598125,1.693307,1.4249886,1.2291887,1.0352017,0.83940166,0.64541465,0.44961473,0.7016165,0.9554313,1.2074331,1.4594349,1.7132497,1.5845293,1.4576219,1.3307146,1.2019942,1.0750868,1.9942589,2.9152439,3.834416,4.7554007,5.674573,8.680465,11.684544,14.690435,17.694515,20.700407,17.647377,14.594349,11.543133,8.490104,5.4370747,5.0781083,4.7173285,4.358362,3.9975824,3.636803,3.6241121,3.6132345,3.6005437,3.587853,3.5751622,3.147303,2.7194438,2.2915847,1.8655385,1.4376793,2.3604772,3.2832751,4.2042603,5.127058,6.049856,6.0752378,6.1006193,6.1241875,6.149569,6.1749506,8.069496,9.965856,11.860401,13.754947,15.649493,15.027647,14.405801,13.782142,13.1602955,12.536636,10.152591,7.7667317,5.382686,2.9968271,0.61278135,0.6091554,0.6073425,0.6055295,0.60190356,0.6000906,0.51306844,0.42423326,0.33721104,0.25018883,0.16316663,0.16316663,0.16316663,0.16316663,0.16316663,0.16316663,0.13053331,0.09789998,0.065266654,0.032633327,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.08520924,0.09427405,0.10515183,0.11421664,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.02175555,0.032633327,0.04169814,0.052575916,0.06164073,0.21030366,0.35715362,0.5058166,0.6526665,0.7995165,0.6399758,0.48043507,0.3208944,0.15954071,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.78319985,1.551896,2.322405,3.092914,3.8616104,9.971294,16.077353,22.185223,28.293095,34.400967,27.901495,21.40565,14.907991,8.410334,1.9126755,1.5373923,1.162109,0.7868258,0.41335547,0.038072214,0.09427405,0.15228885,0.21030366,0.26831847,0.3245203,0.32995918,0.33539808,0.34083697,0.3444629,0.34990177,0.27919623,0.21030366,0.13959812,0.07070554,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.15772775,0.2030518,0.24837588,0.291887,0.33721104,0.27919623,0.2229944,0.16497959,0.10696479,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.07433146,0.099712946,0.12509441,0.15047589,0.17585737,0.21211663,0.25018883,0.28826106,0.3245203,0.36259252,0.31182957,0.26287958,0.21211663,0.16316663,0.11240368,0.1794833,0.24837588,0.3154555,0.3825351,0.44961473,0.42785916,0.40429065,0.3825351,0.36077955,0.33721104,0.46955732,0.60190356,0.73424983,0.8665961,1.0007553,0.89922947,0.7995165,0.69980353,0.6000906,0.50037766,0.9880646,1.4757515,1.9616255,2.4493124,2.9369993,3.3775494,3.8180993,4.256836,4.6973863,5.137936,5.087173,5.038223,4.98746,4.936697,4.8877473,4.994712,5.101677,5.2104545,5.317419,5.424384,4.7227674,4.019338,3.3177216,2.6142921,1.9126755,1.7857682,1.6570477,1.5301404,1.403233,1.2745126,1.6080978,1.93987,2.2716422,2.6052272,2.9369993,2.7792716,2.6233568,2.465629,2.3079014,2.1501737,2.269829,2.3894846,2.5091403,2.6306088,2.7502642,2.8409123,2.9297476,3.0203958,3.1092308,3.199879,3.1654327,3.1291735,3.094727,3.0602808,3.0258346,3.1128569,3.199879,3.2869012,3.3757362,3.4627585,3.346729,3.2325122,3.1182957,3.002266,2.8880494,2.7321346,2.5780327,2.422118,2.268016,2.1121013,2.0051367,1.8981718,1.789394,1.6824293,1.5754645,1.504759,1.4358664,1.3651608,1.2944553,1.2255627,1.0732739,0.91917205,0.7668832,0.61459434,0.46230546,0.7904517,1.1167849,1.4449311,1.7730774,2.0994108,3.0657198,4.0302157,4.994712,5.959208,6.925517,6.4197006,5.915697,5.40988,4.9058766,4.40006,5.5531044,6.7043357,7.85738,9.010424,10.161655,8.673213,7.1829576,5.6927023,4.2024474,2.712192,2.1882458,2.5870976,2.9877625,3.386614,3.787279,4.1879435,4.099108,4.0120864,3.925064,3.8380418,3.7492065,3.7999697,3.8507326,3.8996825,3.9504454,3.9993954,3.4119956,2.8245957,2.2371957,1.649796,1.062396,1.4757515,1.887294,2.3006494,2.712192,3.1255474,3.2252605,3.3249733,3.4246864,3.5243993,3.6241121,5.6999545,7.7757964,9.849826,11.925668,13.999697,12.687112,11.374527,10.061942,8.749357,7.4367723,8.636953,9.837135,11.037316,12.237497,13.437678,13.174799,12.91192,12.650853,12.387974,12.125093,12.137785,12.1504755,12.163166,12.175857,12.186734,11.887595,11.586644,11.287505,10.988366,10.687414,10.388275,10.087324,9.788185,9.487233,9.188094,11.399909,13.611723,15.825351,18.037165,20.250792,23.813263,27.375734,30.938206,34.50068,38.06315,38.13748,38.21181,38.287956,38.36229,38.43662,37.81296,37.18749,36.562016,35.93836,35.312885,28.650248,21.98761,15.324973,8.662335,1.9996977,1.9507477,1.8999848,1.8492218,1.8002719,1.7495089,2.2625773,2.7756457,3.2869012,3.7999697,4.313038,7.3008003,10.28675,13.274512,16.262274,19.250036,20.238102,21.224354,22.212418,23.200481,24.186733,24.150475,24.112402,24.07433,24.03807,23.999998,19.199274,14.400362,9.599637,4.800725,0.0,0.0,0.0,0.0,0.0,0.0,0.11240368,0.22480737,0.33721104,0.44961473,0.5620184,0.53663695,0.51306844,0.48768693,0.46230546,0.43692398,0.34990177,0.26287958,0.17585737,0.0870222,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.5373923,3.0747845,4.612177,6.149569,7.686961,9.374829,11.062697,12.750566,14.436621,16.124489,17.186886,18.24928,19.311678,20.375887,21.438282,17.825048,14.211814,10.600392,6.987158,3.3757362,4.137181,4.900438,5.661882,6.4251394,7.1883965,8.662335,10.138086,11.612025,13.087777,14.561715,14.837286,15.112856,15.386614,15.662184,15.937754,16.762651,17.58755,18.412449,19.237347,20.062244,20.20003,20.337814,20.4756,20.613384,20.749357,20.174648,19.59994,19.025229,18.45052,17.87581,17.25034,16.624866,15.999394,15.375735,14.750263,14.436621,14.124791,13.812962,13.499319,13.1874895,13.125849,13.062395,13.000754,12.937301,12.87566,14.287958,15.700256,17.112555,18.52485,19.93715,20.138388,20.337814,20.537241,20.736666,20.937904,21.66309,22.388275,23.111647,23.836832,24.562017,24.674421,24.786825,24.89923,25.011631,25.125849,22.700104,20.27436,17.85043,15.4246855,13.000754,14.06315,15.125546,16.187943,17.25034,18.312735,16.862366,15.411995,13.961625,12.513068,11.062697,9.837135,8.613385,7.3878226,6.16226,4.936697,4.262275,3.587853,2.911618,2.2371957,1.5627737,1.8619126,2.1628644,2.4620032,2.762955,3.0620937,7.5382986,12.012691,16.487082,20.963285,25.437677,21.15002,16.862366,12.574709,8.287052,3.9993954,8.575313,13.149418,17.725336,22.29944,26.875357,22.875961,18.874754,14.875358,10.874149,6.874754,6.887445,6.9001355,6.9128265,6.925517,6.9382076,6.0244746,5.1125546,4.2006345,3.2869012,2.374981,2.811905,3.2506418,3.6875658,4.12449,4.5632267,3.874301,3.1871881,2.5000753,1.8129625,1.1258497,2.03777,2.94969,3.8634233,4.7753434,5.6872635,4.5867953,3.48814,2.3876717,1.2872034,0.18673515,0.26287958,0.33721104,0.41335547,0.48768693,0.5620184,0.93730164,1.3125849,1.6878681,2.0631514,2.4366217,2.124792,1.8129625,1.49932,1.1874905,0.87566096,0.8122072,0.7505665,0.6871128,0.62547207,0.5620184,0.774135,0.9880646,1.2001812,1.4122978,1.6244144,1.4503701,1.2745126,1.1004683,0.9246109,0.7505665,1.6371052,2.525457,3.4119956,4.3003473,5.186886,8.575313,11.961927,15.350354,18.736969,22.125395,18.736969,15.350354,11.961927,8.575313,5.186886,5.049101,4.9131284,4.7753434,4.6375585,4.499773,3.7129474,2.9243085,2.137483,1.3506571,0.5620184,0.7868258,1.0116332,1.2382535,1.4630609,1.6878681,2.8499773,4.0120864,5.1741953,6.338117,7.500226,7.512917,7.5256076,7.5382986,7.549176,7.5618668,9.900589,12.237497,14.574407,16.913128,19.250036,18.412449,17.57486,16.73727,15.899682,15.062093,12.112403,9.162713,6.2130227,3.2633326,0.31182957,0.40066472,0.48768693,0.5747091,0.66173136,0.7505665,0.63816285,0.52575916,0.41335547,0.2991388,0.18673515,0.17585737,0.16316663,0.15047589,0.13778515,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.19942589,0.40066472,0.6000906,0.7995165,1.0007553,0.7995165,0.6000906,0.40066472,0.19942589,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.89922947,1.8002719,2.6995013,3.6005437,4.499773,11.974618,19.449463,26.92612,34.400967,41.87581,33.97492,26.07584,18.17495,10.274059,2.374981,1.8999848,1.4249886,0.9499924,0.4749962,0.0,0.07433146,0.15047589,0.22480737,0.2991388,0.37528324,0.387974,0.40066472,0.41335547,0.42423326,0.43692398,0.34990177,0.26287958,0.17585737,0.0870222,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.16316663,0.19942589,0.2374981,0.2755703,0.31182957,0.26287958,0.21211663,0.16316663,0.11240368,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.0870222,0.11240368,0.13778515,0.16316663,0.18673515,0.22480737,0.26287958,0.2991388,0.33721104,0.37528324,0.3245203,0.2755703,0.22480737,0.17585737,0.12509441,0.17585737,0.22480737,0.2755703,0.3245203,0.37528324,0.37528324,0.37528324,0.37528324,0.37528324,0.37528324,0.52575916,0.6744221,0.824898,0.97537386,1.1258497,1.0007553,0.87566096,0.7505665,0.62547207,0.50037766,0.93730164,1.3742256,1.8129625,2.2498865,2.6868105,3.0367124,3.386614,3.738329,4.0882306,4.4381323,4.3873696,4.3366065,4.2876563,4.2368937,4.1879435,4.537845,4.8877473,5.237649,5.5875506,5.9374523,5.137936,4.3384194,3.53709,2.7375734,1.938057,1.7748904,1.6117238,1.4503701,1.2872034,1.1258497,1.4249886,1.7241274,2.0250793,2.324218,2.6251698,2.525457,2.4257438,2.324218,2.2245052,2.124792,2.2625773,2.4003625,2.5381477,2.6741197,2.811905,2.9007401,2.9877625,3.0747845,3.1618068,3.2506418,3.2125697,3.1744974,3.1382382,3.100166,3.0620937,3.1744974,3.2869012,3.3993049,3.5117085,3.6241121,3.5117085,3.3993049,3.2869012,3.1744974,3.0620937,2.8753586,2.6868105,2.5000753,2.3133402,2.124792,1.987007,1.8492218,1.7132497,1.5754645,1.4376793,1.3869164,1.3379664,1.2872034,1.2382535,1.1874905,0.9880646,0.7868258,0.5873999,0.387974,0.18673515,0.6744221,1.162109,1.649796,2.137483,2.6251698,3.7256382,4.8242936,5.924762,7.02523,8.125698,7.512917,6.9001355,6.2873545,5.674573,5.0617914,5.9882154,6.9128265,7.837437,8.762048,9.686659,7.9752226,6.261973,4.550536,2.8372865,1.1258497,2.2118144,2.5979755,2.9823234,3.3666716,3.7528327,4.137181,3.9867048,3.8380418,3.6875658,3.53709,3.386614,3.39024,3.392053,3.395679,3.397492,3.3993049,2.8971143,2.3949237,1.892733,1.3905423,0.8883517,1.2328146,1.5772774,1.9217403,2.268016,2.612479,2.8282216,3.0421512,3.2578938,3.4718235,3.6875658,5.866747,8.047741,10.226922,12.407916,14.587097,13.049705,11.512312,9.97492,8.437528,6.9001355,8.107569,9.3150015,10.522435,11.729868,12.937301,12.634536,12.331772,12.03082,11.728055,11.42529,11.612025,11.800573,11.9873085,12.175857,12.362592,13.366973,14.373167,15.377548,16.38193,17.388124,19.53286,21.677593,23.822329,25.967064,28.111797,27.571535,27.033085,26.492823,25.952559,25.412296,27.696629,29.982775,32.26711,34.553253,36.837585,38.501884,40.168,41.8323,43.496597,45.162712,42.724277,40.287655,37.84922,35.412598,32.974163,26.71219,20.450218,14.186432,7.9244595,1.6624867,1.6207886,1.5772774,1.5355793,1.4920682,1.4503701,1.8492218,2.2498865,2.6505513,3.049403,3.4500678,5.8866897,8.325124,10.761745,13.200181,15.636803,16.797098,17.957394,19.117691,20.277987,21.438282,21.010424,20.582563,20.154705,19.726847,19.3008,15.441002,11.579392,7.7195945,3.8597972,0.0,0.0,0.0,0.0,0.0,0.0,0.09427405,0.19036107,0.28463513,0.38072214,0.4749962,0.44961473,0.42423326,0.40066472,0.37528324,0.34990177,0.27919623,0.21030366,0.13959812,0.07070554,0.0,0.0,0.0,0.0,0.0,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,1.4376793,2.762955,4.0882306,5.411693,6.736969,8.375887,10.012992,11.650098,13.287203,14.924308,16.557787,18.189453,19.822933,21.4546,23.088078,19.469404,15.852545,12.235684,8.617011,5.0001507,5.527723,6.055295,6.582867,7.1104393,7.6380115,8.727602,9.817192,10.906783,11.998186,13.087777,13.664299,14.242634,14.819156,15.397491,15.975826,16.59042,17.205015,17.819609,18.434204,19.050611,19.38057,19.71053,20.04049,20.370447,20.700407,20.624262,20.54993,20.4756,20.399454,20.325123,20.142014,19.960718,19.777609,19.5945,19.413204,19.291735,19.17208,19.052423,18.932768,18.813112,18.684393,18.557486,18.430578,18.301857,18.17495,19.112251,20.049553,20.986855,21.924156,22.863272,22.130835,21.398397,20.664148,19.931711,19.199274,19.485722,19.770357,20.054993,20.339626,20.624262,20.542679,20.459282,20.377699,20.294304,20.212719,18.390692,16.566853,14.744824,12.922797,11.10077,12.279196,13.4594345,14.639673,15.819912,17.00015,15.509895,14.01964,12.529385,11.039129,9.550687,8.792869,8.03505,7.2772317,6.5194135,5.7615952,5.1179934,4.4725785,3.827164,3.1817493,2.5381477,2.7430124,2.9478772,3.152742,3.3576066,3.5624714,7.572745,11.583018,15.593291,19.601751,23.612024,19.618069,15.622298,11.626529,7.6325727,3.636803,8.323311,13.008006,17.692701,22.377398,27.062092,23.129776,19.19746,15.265145,11.332829,7.400513,7.066928,6.735156,6.4033837,6.069799,5.7380266,5.0617914,4.3873696,3.7129474,3.0367124,2.3622901,2.666868,2.9732587,3.2778363,3.5824142,3.8869917,3.3304121,2.7720199,2.2154403,1.6570477,1.1004683,1.8202144,2.5399606,3.2597067,3.9794528,4.699199,3.8416677,2.9841363,2.126605,1.2708868,0.41335547,0.43329805,0.45324063,0.47318324,0.49312583,0.51306844,0.9354887,1.357909,1.7803292,2.2027495,2.6251698,2.3931105,2.1592383,1.9271792,1.69512,1.4630609,1.2726997,1.0823387,0.8919776,0.7016165,0.51306844,0.69980353,0.8883517,1.0750868,1.261822,1.4503701,1.305333,1.1602961,1.015259,0.87022203,0.72518504,1.4195497,2.1157274,2.810092,3.5044568,4.2006345,7.309865,10.419096,13.53014,16.63937,19.750414,16.63937,13.53014,10.419096,7.309865,4.2006345,4.1933823,4.1843176,4.177066,4.169814,4.162562,3.5552197,2.9478772,2.3405347,1.7331922,1.1258497,1.2001812,1.2745126,1.3506571,1.4249886,1.49932,2.5997884,3.7002566,4.800725,5.89938,6.9998484,7.083245,7.1648283,7.2482243,7.3298078,7.413204,9.117389,10.821573,12.527572,14.231756,15.937754,15.867048,15.798156,15.72745,15.656745,15.5878525,12.549327,9.512614,6.474089,3.437377,0.40066472,0.57833505,0.7541924,0.9318628,1.1095331,1.2872034,1.0950294,0.90285534,0.7106813,0.5166943,0.3245203,0.27919623,0.23568514,0.19036107,0.14503701,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.15954071,0.3208944,0.48043507,0.6399758,0.7995165,0.6399758,0.48043507,0.3208944,0.15954071,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.7197462,1.4394923,2.1592383,2.8807976,3.6005437,9.579695,15.5606575,21.539808,27.520773,33.499924,27.218008,20.936092,14.652364,8.370448,2.08672,1.6697385,1.2527572,0.83577573,0.4169814,0.0,0.065266654,0.13053331,0.19579996,0.25925365,0.3245203,0.3770962,0.42967212,0.48224804,0.53482395,0.5873999,0.46955732,0.35171473,0.23568514,0.11784257,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.15228885,0.1794833,0.20667773,0.23568514,0.26287958,0.21936847,0.17767033,0.13415924,0.092461094,0.05076295,0.12690738,0.20486477,0.28282216,0.36077955,0.43692398,0.3825351,0.32814622,0.27194437,0.21755551,0.16316663,0.20667773,0.2520018,0.29732585,0.34264994,0.387974,0.33539808,0.28282216,0.23024625,0.17767033,0.12509441,0.17041849,0.21574254,0.25925365,0.3045777,0.34990177,0.36259252,0.37528324,0.387974,0.40066472,0.41335547,0.5493277,0.6871128,0.824898,0.96268314,1.1004683,0.99712944,0.89560354,0.79226464,0.69073874,0.5873999,1.0043813,1.4231756,1.840157,2.2571385,2.6741197,2.907992,3.1400511,3.3721104,3.6041696,3.8380418,3.919625,4.0030212,4.0846047,4.168001,4.249584,4.4925213,4.7354584,4.9783955,5.219519,5.462456,4.764466,4.068288,3.3702974,2.6723068,1.9743162,1.8220274,1.6697385,1.5174497,1.3651608,1.2128719,1.4721256,1.7331922,1.9924458,2.2516994,2.5127661,2.3931105,2.2716422,2.1519866,2.032331,1.9126755,2.030518,2.1483607,2.2643902,2.382233,2.5000753,2.6922495,2.8844235,3.0784104,3.2705846,3.4627585,3.397492,3.3322253,3.2669585,3.2016919,3.1382382,3.2216346,3.3068438,3.392053,3.4772623,3.5624714,3.4029307,3.2415771,3.0820365,2.9224956,2.762955,2.5979755,2.4329958,2.268016,2.1030366,1.938057,1.7966459,1.6570477,1.5174497,1.3778516,1.2382535,1.1802386,1.1222239,1.064209,1.0080072,0.9499924,0.81764615,0.6852999,0.5529536,0.42060733,0.28826106,0.6852999,1.0823387,1.4793775,1.8782293,2.275268,3.2397642,4.2042603,5.1705694,6.1350656,7.0995617,6.5556726,6.009971,5.464269,4.9203806,4.3746786,5.235836,6.09518,6.9545245,7.8156815,8.675026,7.155763,5.634688,4.115425,2.5943494,1.0750868,2.2371957,2.6070402,2.9768846,3.346729,3.7183862,4.0882306,3.874301,3.6621845,3.4500678,3.2379513,3.0258346,2.9805105,2.9351864,2.8898623,2.8445382,2.7992141,2.382233,1.9652514,1.54827,1.1294757,0.7124943,0.9898776,1.2672608,1.5446441,1.8220274,2.0994108,2.42937,2.759329,3.0892882,3.4192474,3.7492065,6.035352,8.319685,10.605831,12.890164,15.174497,13.412297,11.650098,9.8878975,8.125698,6.3616858,7.5781837,8.792869,10.007553,11.222239,12.436923,12.094274,11.751623,11.410787,11.068136,10.725487,11.088079,11.450671,11.813264,12.175857,12.536636,14.848164,17.157877,19.467592,21.777306,24.08702,28.677443,33.267864,37.858284,42.44689,47.037315,43.744976,40.452633,37.160294,33.867954,30.575613,31.581808,32.589817,33.597824,34.60583,35.612022,38.868103,42.12237,45.378452,48.63272,51.88699,47.637405,43.38782,39.138237,34.88684,30.637255,24.775948,18.912827,13.049705,7.1865835,1.3252757,1.2908293,1.2545701,1.2201238,1.1856775,1.1494182,1.4376793,1.7241274,2.0123885,2.3006494,2.5870976,4.4743915,6.3616858,8.2507925,10.138086,12.025381,13.357908,14.690435,16.022963,17.355492,18.688019,17.870373,17.052727,16.23508,15.417434,14.599788,11.680918,8.760235,5.8395524,2.9206827,0.0,0.0,0.0,0.0,0.0,0.0,0.07795739,0.15410182,0.23205921,0.3100166,0.387974,0.36259252,0.33721104,0.31182957,0.28826106,0.26287958,0.21030366,0.15772775,0.10515183,0.052575916,0.0,0.0,0.0,0.0,0.0,0.0,0.045324065,0.09064813,0.13415924,0.1794833,0.22480737,1.3379664,2.4493124,3.5624714,4.6756306,5.7869763,7.3751316,8.963287,10.549629,12.137785,13.724127,15.926876,18.129625,20.332375,22.535126,24.737875,21.115576,17.493277,13.8691635,10.246864,6.624565,6.9182653,7.210152,7.502039,7.795739,8.087626,8.792869,9.498111,10.203354,10.906783,11.612025,12.493125,13.372412,14.2516985,15.132799,16.012085,16.41819,16.82248,17.22677,17.632874,18.037165,18.559298,19.083244,19.605377,20.12751,20.649643,21.07569,21.499924,21.924156,22.350203,22.774435,23.035503,23.294756,23.555822,23.815077,24.07433,24.146849,24.219368,24.291885,24.364405,24.436922,24.24475,24.052574,23.860401,23.668226,23.47424,23.938358,24.400663,24.862968,25.325274,25.78758,24.12328,22.457167,20.792868,19.126755,17.462456,17.308353,17.15244,16.998337,16.842422,16.68832,16.409124,16.13174,15.854358,15.576975,15.299591,14.079468,12.859344,11.63922,10.419096,9.200785,10.497053,11.795135,13.093216,14.389484,15.687565,14.157425,12.627284,11.097144,9.567003,8.036863,7.746789,7.456715,7.166641,6.87838,6.588306,5.9718986,5.3573046,4.74271,4.1281157,3.5117085,3.6222992,3.73289,3.8416677,3.9522583,4.062849,7.607191,11.151533,14.697688,18.24203,21.788185,18.084301,14.382232,10.680162,6.978093,3.2742105,8.069496,12.864782,17.660069,22.455355,27.25064,23.385405,19.520168,15.654932,11.789696,7.9244595,7.2482243,6.5701766,5.8921285,5.2140803,4.537845,4.099108,3.6621845,3.2252605,2.7883365,2.3495996,2.521831,2.6958754,2.8681068,3.0403383,3.2125697,2.7847104,2.3568513,1.9308052,1.502946,1.0750868,1.6026589,2.1302311,2.657803,3.1853752,3.7129474,3.0983531,2.4819458,1.8673514,1.2527572,0.63816285,0.60190356,0.56745726,0.533011,0.49675176,0.46230546,0.9318628,1.403233,1.8727903,2.3423476,2.811905,2.659616,2.5073273,2.3550384,2.2027495,2.0504606,1.7331922,1.4141108,1.0968424,0.7795739,0.46230546,0.62547207,0.7868258,0.9499924,1.1131591,1.2745126,1.1602961,1.0442665,0.9300498,0.81583315,0.69980353,1.2019942,1.7041848,2.2081885,2.7103791,3.2125697,6.0444174,8.8780775,11.709926,14.541773,17.375433,14.541773,11.709926,8.8780775,6.0444174,3.2125697,3.3358512,3.4573197,3.5806012,3.7020695,3.825351,3.397492,2.9696326,2.5417736,2.1157274,1.6878681,1.6117238,1.5373923,1.4630609,1.3869164,1.3125849,2.3495996,3.386614,4.4254417,5.462456,6.4994707,6.6517596,6.8058615,6.9581504,7.1104393,7.262728,8.334189,9.407463,10.480737,11.552197,12.625471,13.321649,14.01964,14.71763,15.415621,16.1118,12.988064,9.862516,6.736969,3.6132345,0.48768693,0.7541924,1.0225109,1.2908293,1.5573349,1.8256533,1.551896,1.2799516,1.0080072,0.73424983,0.46230546,0.38434806,0.30820364,0.23024625,0.15228885,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.11965553,0.23931105,0.36077955,0.48043507,0.6000906,0.48043507,0.36077955,0.23931105,0.11965553,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.5402629,1.0805258,1.6207886,2.1592383,2.6995013,7.1847706,11.67004,16.15531,20.64058,25.124035,20.459282,15.79453,11.129777,6.4650245,1.8002719,1.4394923,1.0805258,0.7197462,0.36077955,0.0,0.054388877,0.11059072,0.16497959,0.21936847,0.2755703,0.3680314,0.4604925,0.5529536,0.64541465,0.73787576,0.58921283,0.44236287,0.2955129,0.14684997,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.14322405,0.15954071,0.17767033,0.19579996,0.21211663,0.17767033,0.14322405,0.10696479,0.072518505,0.038072214,0.19217403,0.3480888,0.50219065,0.65810543,0.8122072,0.678048,0.5420758,0.40791658,0.27194437,0.13778515,0.19036107,0.24293698,0.2955129,0.3480888,0.40066472,0.3444629,0.29007402,0.23568514,0.1794833,0.12509441,0.16497959,0.20486477,0.24474995,0.28463513,0.3245203,0.34990177,0.37528324,0.40066472,0.42423326,0.44961473,0.5747091,0.69980353,0.824898,0.9499924,1.0750868,0.99531645,0.9155461,0.83577573,0.7541924,0.6744221,1.0732739,1.4703126,1.8673514,2.2643902,2.663242,2.7774587,2.8916752,3.007705,3.1219215,3.2379513,3.4518807,3.6676233,3.8833659,4.0972953,4.313038,4.4471974,4.5831695,4.7173285,4.853301,4.98746,4.3928084,3.7981565,3.2016919,2.6070402,2.0123885,1.8691645,1.7277533,1.5845293,1.4431182,1.2998942,1.5192627,1.7404441,1.9598125,2.179181,2.4003625,2.2607644,2.1193533,1.9797552,1.840157,1.7005589,1.7966459,1.8945459,1.9924458,2.0903459,2.1882458,2.4855716,2.7828975,3.0802233,3.3775494,3.6748753,3.5824142,3.489953,3.397492,3.3050308,3.2125697,3.2705846,3.3267863,3.3848011,3.442816,3.5008307,3.29234,3.0856624,2.8771715,2.6704938,2.4620032,2.3205922,2.1773682,2.034144,1.892733,1.7495089,1.6080978,1.4648738,1.3216497,1.1802386,1.0370146,0.97174793,0.90829426,0.8430276,0.7777609,0.7124943,0.64722764,0.581961,0.5166943,0.45324063,0.387974,0.69436467,1.0025684,1.310772,1.6171626,1.9253663,2.7557032,3.584227,4.4145637,5.2449007,6.0752378,5.5966153,5.1198063,4.6429973,4.164375,3.6875658,4.4816437,5.277534,6.071612,6.867502,7.663393,6.3344913,5.0074024,3.680314,2.3532255,1.0243238,2.2625773,2.617918,2.9732587,3.3267863,3.682127,4.0374675,3.7618973,3.48814,3.2125697,2.9369993,2.663242,2.570781,2.47832,2.3858588,2.2915847,2.1991236,1.8673514,1.5355793,1.2019942,0.87022203,0.53663695,0.7469406,0.9572442,1.167548,1.3778516,1.5881553,2.032331,2.47832,2.9224956,3.3666716,3.8126602,6.202145,8.59163,10.982927,13.372412,15.761897,13.77489,11.787883,9.799063,7.8120556,5.825049,7.0469856,8.270736,9.492672,10.714609,11.938358,11.555823,11.173288,10.790753,10.408218,10.025683,10.56232,11.10077,11.637406,12.175857,12.712494,16.327541,19.942589,23.557636,27.172684,30.787731,37.822025,44.85813,51.89243,58.928535,65.96283,59.918415,53.873997,47.827766,41.783348,35.737118,35.466988,35.196857,34.926723,34.656593,34.388275,39.23251,44.076748,48.922794,53.767033,58.61308,52.550533,46.487988,40.425438,34.362892,28.300346,22.837889,17.375433,11.912977,6.450521,0.9880646,0.96087015,0.9318628,0.90466833,0.8774739,0.85027945,1.0243238,1.2001812,1.3742256,1.550083,1.7241274,3.0620937,4.40006,5.7380266,7.07418,8.412147,9.916905,11.421664,12.928236,14.432995,15.937754,14.730321,13.522888,12.3154545,11.108022,9.900589,7.9190207,5.9392653,3.9595103,1.9797552,0.0,0.0,0.0,0.0,0.0,0.0,0.059827764,0.11965553,0.1794833,0.23931105,0.2991388,0.2755703,0.25018883,0.22480737,0.19942589,0.17585737,0.13959812,0.10515183,0.07070554,0.034446288,0.0,0.0,0.0,0.0,0.0,0.0,0.06707962,0.13415924,0.2030518,0.27013144,0.33721104,1.2382535,2.137483,3.0367124,3.9377546,4.836984,6.3743763,7.911769,9.449161,10.988366,12.525759,15.297778,18.069798,20.841818,23.61565,26.38767,22.759932,19.132195,15.504456,11.876718,8.2507925,8.306994,8.365009,8.423024,8.479226,8.537241,8.858135,9.177217,9.498111,9.817192,10.138086,11.320138,12.50219,13.684241,14.868106,16.050158,16.244144,16.439945,16.635744,16.829731,17.025532,17.73984,18.454145,19.170267,19.884573,20.600695,21.525305,22.449915,23.374527,24.300951,25.225561,25.927177,26.630608,27.332224,28.035654,28.73727,29.001963,29.268469,29.533161,29.797853,30.062546,29.805105,29.547665,29.290224,29.032784,28.775343,28.762651,28.74996,28.73727,28.724579,28.71189,26.115726,23.51775,20.919775,18.3218,15.725637,15.129172,14.534521,13.939869,13.345218,12.750566,12.277383,11.804199,11.332829,10.859646,10.386462,9.770056,9.151835,8.535428,7.9172077,7.3008003,8.714911,10.129022,11.544946,12.96087,14.37498,12.804955,11.234929,9.664904,8.094878,6.5248523,6.7025228,6.880193,7.057863,7.2355337,7.413204,6.827617,6.24203,5.658256,5.0726695,4.4870825,4.503399,4.517903,4.5324063,4.5469103,4.5632267,7.6416373,10.721861,13.802084,16.882307,19.96253,16.55235,13.142166,9.731983,6.3218007,2.911618,7.817495,12.721559,17.627436,22.533312,27.437376,23.63922,19.842875,16.04472,12.246562,8.450218,7.4277077,6.4051967,5.382686,4.360175,3.3376641,3.1382382,2.9369993,2.7375734,2.5381477,2.3369088,2.3767939,2.4166791,2.4583774,2.4982624,2.5381477,2.2408218,1.9416829,1.6443571,1.3470312,1.0497054,1.3851035,1.7205015,2.0540867,2.3894846,2.7248828,2.3532255,1.9797552,1.6080978,1.2346275,0.8629702,0.77232206,0.68167394,0.59283876,0.50219065,0.41335547,0.9300498,1.4467441,1.9652514,2.4819458,3.000453,2.9279346,2.855416,2.7828975,2.7103791,2.6378605,2.1918716,1.7476959,1.3017071,0.8575313,0.41335547,0.5493277,0.6871128,0.824898,0.96268314,1.1004683,1.015259,0.9300498,0.8448406,0.75963134,0.6744221,0.98443866,1.2944553,1.6044719,1.9144884,2.2245052,4.780782,7.3352466,9.88971,12.444175,15.000452,12.444175,9.88971,7.3352466,4.780782,2.2245052,2.47832,2.7303216,2.9823234,3.2343252,3.48814,3.2397642,2.9932013,2.7448254,2.4982624,2.2498865,2.0250793,1.8002719,1.5754645,1.3506571,1.1258497,2.0994108,3.0747845,4.0501585,5.0255322,5.999093,6.2220874,6.445082,6.6680765,6.889258,7.112252,7.552802,7.991539,8.432089,8.872639,9.313189,10.778063,12.242936,13.70781,15.172684,16.637558,13.424988,10.212419,6.9998484,3.787279,0.5747091,0.9318628,1.2908293,1.647983,2.0051367,2.3622901,2.0105755,1.6570477,1.305333,0.95180535,0.6000906,0.4894999,0.38072214,0.27013144,0.15954071,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07977036,0.15954071,0.23931105,0.3208944,0.40066472,0.3208944,0.23931105,0.15954071,0.07977036,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.36077955,0.7197462,1.0805258,1.4394923,1.8002719,4.7898474,7.7794223,10.770811,13.760386,16.749962,13.702372,10.654781,7.607191,4.559601,1.5120108,1.209246,0.90829426,0.6055295,0.30276474,0.0,0.045324065,0.09064813,0.13415924,0.1794833,0.22480737,0.35715362,0.4894999,0.62184614,0.7541924,0.8883517,0.7106813,0.533011,0.35534066,0.17767033,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.13234627,0.13959812,0.14684997,0.15410182,0.16316663,0.13415924,0.10696479,0.07977036,0.052575916,0.025381476,0.2574407,0.4894999,0.72337204,0.9554313,1.1874905,0.97174793,0.75781834,0.5420758,0.32814622,0.11240368,0.17223145,0.23205921,0.291887,0.35171473,0.41335547,0.35534066,0.29732585,0.23931105,0.18310922,0.12509441,0.15954071,0.19579996,0.23024625,0.26469254,0.2991388,0.33721104,0.37528324,0.41335547,0.44961473,0.48768693,0.6000906,0.7124943,0.824898,0.93730164,1.0497054,0.9916905,0.9354887,0.8774739,0.8194591,0.76325727,1.1403534,1.5174497,1.8945459,2.2716422,2.6505513,2.6469254,2.6451125,2.6432993,2.6396735,2.6378605,2.9841363,3.3322253,3.680314,4.02659,4.3746786,4.401873,4.4308805,4.458075,4.4852695,4.512464,4.019338,3.5280252,3.0348995,2.5417736,2.0504606,1.9181144,1.7857682,1.651609,1.5192627,1.3869164,1.5682126,1.7476959,1.9271792,2.1066625,2.2879589,2.126605,1.9670644,1.8075237,1.647983,1.4866294,1.5645868,1.6425442,1.7205015,1.7966459,1.8746033,2.277081,2.6795588,3.0820365,3.484514,3.8869917,3.7673361,3.6476808,3.5280252,3.4083695,3.2869012,3.3177216,3.346729,3.3775494,3.4083695,3.437377,3.1817493,2.9279346,2.6723068,2.4166791,2.1628644,2.0432088,1.9217403,1.8020848,1.6824293,1.5627737,1.4177368,1.2726997,1.1276628,0.9826257,0.8375887,0.7650702,0.69255173,0.6200332,0.5475147,0.4749962,0.47680917,0.48043507,0.48224804,0.48587397,0.48768693,0.70524246,0.922798,1.1403534,1.357909,1.5754645,2.269829,2.9641938,3.6603715,4.3547363,5.049101,4.6393714,4.229642,3.8199122,3.4101827,3.000453,3.729264,4.459888,5.1905117,5.919323,6.6499467,5.5150323,4.3801174,3.245203,2.1102884,0.97537386,2.2879589,2.6269827,2.9678197,3.3068438,3.6476808,3.9867048,3.6494937,3.3122826,2.9750717,2.6378605,2.3006494,2.1592383,2.0196402,1.8800422,1.7404441,1.6008459,1.35247,1.1059072,0.8575313,0.6091554,0.36259252,0.5058166,0.64722764,0.7904517,0.9318628,1.0750868,1.6352923,2.1954978,2.7557032,3.3159087,3.874301,6.3707504,8.865387,11.3600235,13.85466,16.349297,14.137483,11.925668,9.712041,7.500226,5.2865987,6.5176005,7.746789,8.977791,10.20698,11.437981,11.015561,10.593141,10.17072,9.7483,9.325879,10.038374,10.750868,11.463363,12.175857,12.888351,17.80692,22.727299,27.64768,32.568058,37.48844,46.96661,56.44659,65.92838,75.40836,84.88834,76.09004,67.29355,58.49524,49.69693,40.900436,39.352165,37.80571,36.25744,34.709167,33.162712,39.596916,46.032932,52.467136,58.903152,65.33736,57.46185,49.588154,41.712643,33.837135,25.961624,20.899832,15.838041,10.774437,5.712645,0.6508536,0.629098,0.6091554,0.58921283,0.56927025,0.5493277,0.61278135,0.6744221,0.73787576,0.7995165,0.8629702,1.649796,2.4366217,3.2252605,4.0120864,4.800725,6.4777155,8.154706,9.8316965,11.510499,13.1874895,11.59027,9.99305,8.394017,6.796797,5.199577,4.160749,3.1201086,2.079468,1.0406405,0.0,0.0,0.0,0.0,0.0,0.0,0.04169814,0.08520924,0.12690738,0.17041849,0.21211663,0.18673515,0.16316663,0.13778515,0.11240368,0.0870222,0.07070554,0.052575916,0.034446288,0.018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.09064813,0.1794833,0.27013144,0.36077955,0.44961473,1.1367276,1.8256533,2.5127661,3.199879,3.8869917,5.375434,6.8620634,8.350506,9.837135,11.325577,14.666867,18.00997,21.353073,24.694363,28.037466,24.40429,20.772924,17.139748,13.506571,9.875207,9.697536,9.519867,9.342196,9.164526,8.9868555,8.923402,8.858135,8.792869,8.727602,8.662335,10.147152,11.631968,13.116784,14.603414,16.08823,16.071913,16.05741,16.042906,16.026588,16.012085,16.92038,17.82686,18.735155,19.641636,20.54993,21.97492,23.399908,24.824896,26.249886,27.674873,28.820665,29.964645,31.110437,32.254417,33.40021,33.857075,34.315754,34.77262,35.22949,35.688168,35.36546,35.042755,34.720047,34.39734,34.07463,33.586945,33.09926,32.613384,32.125698,31.63801,28.108171,24.578333,21.046682,17.516844,13.987006,12.951805,11.916603,10.883214,9.848013,8.812811,8.145641,7.476658,6.8094873,6.1423173,5.475147,5.4606433,5.4443264,5.429823,5.4153194,5.4008155,6.932769,8.464723,9.9966755,11.530442,13.062395,11.452485,9.842574,8.232663,6.622752,5.0128417,5.658256,6.301858,6.947273,7.592687,8.238102,7.6833353,7.1267557,6.5719895,6.017223,5.462456,5.382686,5.3029156,5.223145,5.143375,5.0617914,7.6778965,10.292189,12.908294,15.522586,18.136877,15.020395,11.9021,8.785617,5.667321,2.5508385,7.5654926,12.580148,17.5948,22.609457,27.624111,23.894846,20.165583,16.434505,12.705242,8.974165,7.607191,6.240217,4.8732433,3.5044568,2.137483,2.175555,2.2118144,2.2498865,2.2879589,2.324218,2.231757,2.1392958,2.0468347,1.9543737,1.8619126,1.69512,1.5283275,1.3597219,1.1929294,1.0243238,1.167548,1.310772,1.452183,1.5954071,1.7368182,1.6080978,1.4775645,1.3470312,1.2183108,1.0877775,0.94274056,0.79770356,0.6526665,0.5076295,0.36259252,0.92823684,1.4920682,2.0577126,2.6233568,3.1871881,3.1944401,3.2016919,3.2107568,3.2180085,3.2252605,2.6523643,2.079468,1.5083848,0.9354887,0.36259252,0.4749962,0.5873999,0.69980353,0.8122072,0.9246109,0.87022203,0.81583315,0.75963134,0.70524246,0.6508536,0.7668832,0.88472575,1.0025684,1.1204109,1.2382535,3.5153344,5.7924156,8.069496,10.348391,12.625471,10.346578,8.069496,5.7924156,3.5153344,1.2382535,1.6207886,2.0033236,2.3858588,2.7683938,3.149116,3.0820365,3.0149567,2.9478772,2.8807976,2.811905,2.4366217,2.0631514,1.6878681,1.3125849,0.93730164,1.8492218,2.762955,3.6748753,4.5867953,5.5005283,5.7924156,6.0843024,6.378002,6.6698895,6.9617763,6.7696023,6.5774283,6.3852544,6.19308,5.999093,8.232663,10.46442,12.697989,14.929747,17.163317,13.861912,10.56232,7.262728,3.9631362,0.66173136,1.1095331,1.5573349,2.0051367,2.4529383,2.9007401,2.467442,2.034144,1.6026589,1.1693609,0.73787576,0.5946517,0.45324063,0.3100166,0.16679256,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03988518,0.07977036,0.11965553,0.15954071,0.19942589,0.15954071,0.11965553,0.07977036,0.03988518,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1794833,0.36077955,0.5402629,0.7197462,0.89922947,2.3949237,3.8906176,5.384499,6.880193,8.374074,6.94546,5.5150323,4.0846047,2.6541772,1.2255627,0.9808127,0.73424983,0.4894999,0.24474995,0.0,0.034446288,0.07070554,0.10515183,0.13959812,0.17585737,0.3480888,0.52032024,0.69255173,0.86478317,1.0370146,0.83033687,0.62184614,0.41516843,0.20667773,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.12328146,0.11965553,0.11784257,0.11421664,0.11240368,0.092461094,0.072518505,0.052575916,0.032633327,0.012690738,0.32270733,0.6327239,0.94274056,1.2527572,1.5627737,1.2672608,0.97174793,0.678048,0.3825351,0.0870222,0.15410182,0.2229944,0.29007402,0.35715362,0.42423326,0.36440548,0.3045777,0.24474995,0.18492219,0.12509441,0.15410182,0.18492219,0.21574254,0.24474995,0.2755703,0.3245203,0.37528324,0.42423326,0.4749962,0.52575916,0.62547207,0.72518504,0.824898,0.9246109,1.0243238,0.9898776,0.9554313,0.91917205,0.88472575,0.85027945,1.2074331,1.5645868,1.9217403,2.280707,2.6378605,2.518205,2.3967366,2.277081,2.1574254,2.03777,2.518205,2.9968271,3.4772623,3.9576974,4.4381323,4.358362,4.2767787,4.1970086,4.117238,4.0374675,3.6476808,3.2578938,2.8681068,2.47832,2.08672,1.9652514,1.84197,1.7205015,1.5972201,1.4757515,1.6153497,1.7549478,1.8945459,2.034144,2.175555,1.9942589,1.8147756,1.6352923,1.455809,1.2745126,1.3325275,1.3905423,1.4467441,1.504759,1.5627737,2.0704033,2.5780327,3.0856624,3.5932918,4.099108,3.9522583,3.8054085,3.6567454,3.5098956,3.3630457,3.3648586,3.3666716,3.3702974,3.3721104,3.3757362,3.0729716,2.770207,2.467442,2.1646774,1.8619126,1.7658255,1.6679256,1.5700256,1.4721256,1.3742256,1.2273756,1.0805258,0.9318628,0.7850128,0.63816285,0.55839247,0.47680917,0.39703882,0.31726846,0.2374981,0.30820364,0.3770962,0.44780177,0.5166943,0.5873999,0.71430725,0.8430276,0.969935,1.0968424,1.2255627,1.7857682,2.3441606,2.904366,3.4645715,4.024777,3.682127,3.339477,2.9968271,2.6541772,2.3133402,2.9768846,3.6422417,4.307599,4.972956,5.638314,4.695573,3.7528327,2.810092,1.8673514,0.9246109,2.3133402,2.6378605,2.962381,3.2869012,3.6132345,3.9377546,3.53709,3.1382382,2.7375734,2.3369088,1.938057,1.7495089,1.5627737,1.3742256,1.1874905,1.0007553,0.8375887,0.6744221,0.51306844,0.34990177,0.18673515,0.26287958,0.33721104,0.41335547,0.48768693,0.5620184,1.2382535,1.9126755,2.5870976,3.2633326,3.9377546,6.5375433,9.137331,11.73712,14.336908,16.936697,14.500074,12.063453,9.625018,7.1865835,4.749962,5.9882154,7.224656,8.46291,9.699349,10.937603,10.475298,10.012992,9.550687,9.088382,8.624263,9.512614,10.399154,11.287505,12.175857,13.062395,19.288109,25.512009,31.737722,37.963436,44.187336,56.113007,68.03686,79.962524,91.8882,103.81205,92.26348,80.7131,69.16271,57.612324,46.06194,43.237343,40.41275,37.588154,34.761745,31.93715,39.963135,47.987305,56.01329,64.03747,72.06164,62.374977,52.68832,42.999847,33.313187,23.624716,18.961775,14.300649,9.637709,4.974769,0.31182957,0.2991388,0.28826106,0.2755703,0.26287958,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.2374981,0.4749962,0.7124943,0.9499924,1.1874905,3.0367124,4.8877473,6.736969,8.588004,10.437225,8.450218,6.4632115,4.4743915,2.4873846,0.50037766,0.40066472,0.2991388,0.19942589,0.099712946,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.11240368,0.22480737,0.33721104,0.44961473,0.5620184,1.0370146,1.5120108,1.987007,2.4620032,2.9369993,4.3746786,5.812358,7.250037,8.6877165,10.125396,14.037769,17.950142,21.862516,25.774889,29.687262,26.050459,22.411844,18.77504,15.138238,11.499621,11.088079,10.674724,10.263181,9.849826,9.438283,8.9868555,8.537241,8.087626,7.6380115,7.1883965,8.974165,10.761745,12.549327,14.336908,16.124489,15.899682,15.674874,15.4500675,15.22526,15.000452,16.099108,17.199575,18.300045,19.400513,20.499168,22.424534,24.349901,26.275267,28.200632,30.124186,31.712341,33.300495,34.88684,36.474995,38.06315,38.71219,39.363045,40.012085,40.662937,41.311977,40.925816,40.53784,40.149868,39.761894,39.375732,38.41305,37.450367,36.487686,35.525,34.562317,30.100618,25.637104,21.175404,16.71189,12.250188,10.774437,9.300498,7.8247466,6.350808,4.8750563,4.0120864,3.150929,2.2879589,1.4249886,0.5620184,1.1494182,1.7368182,2.324218,2.911618,3.5008307,5.1506267,6.8004227,8.450218,10.100015,11.74981,10.100015,8.450218,6.8004227,5.1506267,3.5008307,4.612177,5.7253356,6.836682,7.949841,9.063,8.537241,8.013294,7.4875355,6.9617763,6.43783,6.261973,6.0879283,5.9120708,5.7380266,5.562169,7.7123427,9.862516,12.012691,14.162864,16.313038,13.488441,10.662033,7.837437,5.0128417,2.1882458,7.311678,12.436923,17.562168,22.687414,27.812658,24.150475,20.48829,16.824293,13.162108,9.499924,7.7866745,6.0752378,4.361988,2.6505513,0.93730164,1.2128719,1.4866294,1.7621996,2.03777,2.3133402,2.08672,1.8619126,1.6371052,1.4122978,1.1874905,1.1494182,1.1131591,1.0750868,1.0370146,1.0007553,0.9499924,0.89922947,0.85027945,0.7995165,0.7505665,0.8629702,0.97537386,1.0877775,1.2001812,1.3125849,1.1131591,0.9119202,0.7124943,0.51306844,0.31182957,0.9246109,1.5373923,2.1501737,2.762955,3.3757362,3.4627585,3.5497808,3.636803,3.7256382,3.8126602,3.1128569,2.4130533,1.7132497,1.0116332,0.31182957,0.40066472,0.48768693,0.5747091,0.66173136,0.7505665,0.72518504,0.69980353,0.6744221,0.6508536,0.62547207,0.5493277,0.4749962,0.40066472,0.3245203,0.25018883,2.2498865,4.249584,6.249282,8.2507925,10.25049,8.24898,6.249282,4.249584,2.2498865,0.25018883,0.76325727,1.2745126,1.7875811,2.3006494,2.811905,2.9243085,3.0367124,3.149116,3.2633326,3.3757362,2.8499773,2.324218,1.8002719,1.2745126,0.7505665,1.6008459,2.4493124,3.299592,4.1498713,5.0001507,5.3627434,5.7253356,6.0879283,6.450521,6.813113,5.9882154,5.163317,4.3366065,3.5117085,2.6868105,5.6872635,8.6877165,11.6881695,14.68681,17.687263,14.300649,10.912222,7.5256076,4.137181,0.7505665,1.2872034,1.8256533,2.3622901,2.9007401,3.437377,2.9243085,2.4130533,1.8999848,1.3869164,0.87566096,0.69980353,0.52575916,0.34990177,0.17585737,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.18673515,0.37528324,0.5620184,0.7505665,0.93730164,0.7505665,0.5620184,0.37528324,0.18673515,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.33721104,0.5493277,0.76325727,0.97537386,1.1874905,0.9499924,0.7124943,0.4749962,0.2374981,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.387974,0.774135,1.162109,1.550083,1.938057,1.5627737,1.1874905,0.8122072,0.43692398,0.06164073,0.13778515,0.21211663,0.28826106,0.36259252,0.43692398,0.37528324,0.31182957,0.25018883,0.18673515,0.12509441,0.15047589,0.17585737,0.19942589,0.22480737,0.25018883,0.31182957,0.37528324,0.43692398,0.50037766,0.5620184,0.6508536,0.73787576,0.824898,0.9119202,1.0007553,0.9880646,0.97537386,0.96268314,0.9499924,0.93730164,1.2745126,1.6117238,1.9507477,2.2879589,2.6251698,2.3876717,2.1501737,1.9126755,1.6751775,1.4376793,2.0504606,2.663242,3.2742105,3.8869917,4.499773,4.313038,4.12449,3.9377546,3.7492065,3.5624714,3.2742105,2.9877625,2.6995013,2.4130533,2.124792,2.0123885,1.8999848,1.7875811,1.6751775,1.5627737,1.6624867,1.7621996,1.8619126,1.9616255,2.0631514,1.8619126,1.6624867,1.4630609,1.261822,1.062396,1.1004683,1.1367276,1.1747998,1.2128719,1.2491312,1.8619126,2.474694,3.0874753,3.7002566,4.313038,4.137181,3.9631362,3.787279,3.6132345,3.437377,3.4119956,3.386614,3.3630457,3.3376641,3.3122826,2.962381,2.612479,2.2625773,1.9126755,1.5627737,1.4866294,1.4122978,1.3379664,1.261822,1.1874905,1.0370146,0.8883517,0.73787576,0.5873999,0.43692398,0.34990177,0.26287958,0.17585737,0.0870222,0.0,0.13778515,0.2755703,0.41335547,0.5493277,0.6871128,0.72518504,0.76325727,0.7995165,0.8375887,0.87566096,1.2998942,1.7259403,2.1501737,2.5744069,3.000453,2.7248828,2.4493124,2.175555,1.8999848,1.6244144,2.2245052,2.8245957,3.4246864,4.024777,4.6248674,3.874301,3.1255474,2.374981,1.6244144,0.87566096,2.9369993,2.9877625,3.0367124,3.0874753,3.1382382,3.1871881,2.8971143,2.6070402,2.3169663,2.0268922,1.7368182,1.5627737,1.3869164,1.2128719,1.0370146,0.8629702,0.7505665,0.63816285,0.52575916,0.41335547,0.2991388,0.35715362,0.41516843,0.47318324,0.5293851,0.5873999,1.4775645,2.3677292,3.2578938,4.1480584,5.038223,6.9490857,8.861761,10.774437,12.687112,14.599788,12.964496,11.329204,9.695724,8.0604315,6.4251394,7.3298078,8.234476,9.139144,10.045626,10.950294,10.874149,10.799818,10.725487,10.649343,10.57501,12.099712,13.6244135,15.149116,16.67563,18.20033,25.20018,32.200027,39.19988,46.199726,53.199574,62.170113,71.13884,80.109375,89.07992,98.05045,87.07478,76.100914,65.125244,54.149567,43.175705,41.237648,39.29959,37.363346,35.42529,33.487232,38.795586,44.102127,49.41048,54.717022,60.02538,52.49977,44.975975,37.450367,29.92476,22.399153,17.970085,13.541018,9.110137,4.6792564,0.25018883,0.24837588,0.24474995,0.24293698,0.23931105,0.2374981,0.21574254,0.19217403,0.17041849,0.14684997,0.12509441,0.3045777,0.48587397,0.6653573,0.8448406,1.0243238,2.4928236,3.9595103,5.42801,6.8946967,8.363196,6.773228,5.18326,3.5932918,2.0033236,0.41335547,0.34083697,0.26831847,0.19579996,0.12328146,0.05076295,0.06707962,0.08520924,0.10333887,0.11965553,0.13778515,0.13053331,0.12328146,0.11421664,0.10696479,0.099712946,0.11421664,0.13053331,0.14503701,0.15954071,0.17585737,0.40429065,0.6345369,0.86478317,1.0950294,1.3252757,1.3379664,1.3506571,1.3633479,1.3742256,1.3869164,1.2745126,1.162109,1.0497054,0.93730164,0.824898,1.5428312,2.2607644,2.9768846,3.6948178,4.4127507,5.6999545,6.987158,8.274362,9.563377,10.850581,13.878228,16.904062,19.933523,22.959358,25.987005,23.704485,21.421967,19.139446,16.856926,14.574407,13.809336,13.044266,12.279196,11.514126,10.750868,10.627586,10.504305,10.382836,10.259555,10.138086,11.757062,13.377851,14.996826,16.617615,18.236591,17.932013,17.627436,17.322857,17.01828,16.71189,17.669134,18.628191,19.585434,20.542679,21.499924,22.089136,22.680162,23.269375,23.860401,24.449614,26.24082,28.030214,29.819609,31.610815,33.40021,33.434654,33.470917,33.50536,33.539806,33.574253,33.731983,33.88971,34.047436,34.205166,34.362892,33.15002,31.93715,30.724277,29.513218,28.300346,24.792263,21.285994,17.77791,14.269829,10.761745,9.510801,8.258044,7.0052876,5.75253,4.499773,3.785466,3.0693457,2.3550384,1.6407311,0.9246109,3.0820365,5.239462,7.3968873,9.554313,11.711739,11.617464,11.5231905,11.427103,11.332829,11.236742,10.729113,10.223296,9.715667,9.208037,8.700407,9.104698,9.510801,9.915092,10.319383,10.725487,10.587702,10.449916,10.312131,10.174346,10.036561,9.481794,8.927028,8.372261,7.817495,7.262728,9.19172,11.122525,13.05333,14.982323,16.913128,14.144734,11.378153,8.609759,5.8431783,3.0747845,7.137634,11.200482,15.263332,19.324368,23.387217,20.263483,17.137936,14.012388,10.88684,7.763106,6.6100616,5.4570174,4.305786,3.152742,1.9996977,2.1556125,2.3097143,2.465629,2.619731,2.7756457,2.4493124,2.124792,1.8002719,1.4757515,1.1494182,1.1059072,1.0605831,1.015259,0.969935,0.9246109,0.87566096,0.824898,0.774135,0.72518504,0.6744221,1.1566701,1.6407311,2.1229792,2.6052272,3.0874753,2.764768,2.4420607,2.1193533,1.7966459,1.4757515,1.7223145,1.9706904,2.2172532,2.465629,2.712192,2.8844235,3.056655,3.2306993,3.4029307,3.5751622,2.9224956,2.269829,1.6171626,0.9644961,0.31182957,0.40429065,0.49675176,0.58921283,0.68167394,0.774135,0.7324369,0.69073874,0.64722764,0.6055295,0.5620184,0.5166943,0.47318324,0.42785916,0.3825351,0.33721104,2.1429217,3.9468195,5.75253,7.558241,9.362139,7.552802,5.7434654,3.9323158,2.1229792,0.31182957,0.7324369,1.1530442,1.5718386,1.9924458,2.4130533,2.4928236,2.572594,2.6523643,2.7321346,2.811905,2.3949237,1.9779422,1.5591478,1.1421664,0.72518504,1.4249886,2.124792,2.8245957,3.5243993,4.2242026,4.539658,4.855114,5.1705694,5.484212,5.7996674,5.1923246,4.5849824,3.97764,3.3702974,2.762955,5.0599785,7.3570023,9.655839,11.952863,14.249886,12.018129,9.784559,7.552802,5.319232,3.0874753,3.0820365,3.0765975,3.0729716,3.0675328,3.0620937,2.7828975,2.5018883,2.222692,1.9416829,1.6624867,1.3325275,1.0025684,0.6726091,0.34264994,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.07070554,0.07795739,0.08520924,0.092461094,0.099712946,0.08520924,0.07070554,0.054388877,0.03988518,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.15047589,0.2991388,0.44961473,0.6000906,0.7505665,0.6000906,0.44961473,0.2991388,0.15047589,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.2955129,0.47680917,0.65991837,0.8430276,1.0243238,0.83940166,0.6544795,0.46955732,0.28463513,0.099712946,0.10696479,0.11421664,0.12328146,0.13053331,0.13778515,0.13234627,0.12690738,0.12328146,0.11784257,0.11240368,0.09064813,0.06707962,0.045324065,0.02175555,0.0,0.33177215,0.6653573,0.99712944,1.3307146,1.6624867,1.357909,1.0533313,0.7469406,0.44236287,0.13778515,0.19942589,0.26287958,0.3245203,0.387974,0.44961473,0.3825351,0.3154555,0.24837588,0.1794833,0.11240368,0.13415924,0.15772775,0.1794833,0.2030518,0.22480737,0.28826106,0.34990177,0.41335547,0.4749962,0.53663695,0.6091554,0.68167394,0.7541924,0.82671094,0.89922947,0.8901646,0.8792868,0.87022203,0.85934424,0.85027945,1.1276628,1.405046,1.6824293,1.9598125,2.2371957,2.0722163,1.9072367,1.742257,1.5772774,1.4122978,1.9326181,2.4529383,2.9732587,3.491766,4.0120864,3.8942437,3.778214,3.6603715,3.5425289,3.4246864,3.1944401,2.9641938,2.7357605,2.5055144,2.275268,2.2081885,2.1392958,2.0722163,2.0051367,1.938057,1.9471219,1.9579996,1.9670644,1.9779422,1.987007,1.7676386,1.54827,1.3270886,1.1077201,0.8883517,0.9119202,0.93730164,0.96268314,0.9880646,1.0116332,1.5881553,2.1628644,2.7375734,3.3122826,3.8869917,3.7002566,3.5117085,3.3249733,3.1382382,2.94969,2.907992,2.864481,2.8227828,2.7792716,2.7375734,2.4529383,2.1683033,1.8818551,1.5972201,1.3125849,1.2491312,1.1874905,1.1258497,1.062396,1.0007553,0.8919776,0.7850128,0.678048,0.56927025,0.46230546,0.387974,0.31182957,0.2374981,0.16316663,0.0870222,0.18310922,0.27738327,0.37165734,0.46774435,0.5620184,0.6327239,0.7016165,0.77232206,0.8430276,0.9119202,1.2473183,1.5827163,1.9181144,2.2516994,2.5870976,2.4402475,2.2915847,2.1447346,1.9978848,1.8492218,2.4420607,3.0348995,3.6277382,4.220577,4.8116026,4.0157123,3.2180085,2.420305,1.6226015,0.824898,3.5624714,3.3376641,3.1128569,2.8880494,2.663242,2.4366217,2.2571385,2.077655,1.8981718,1.7168756,1.5373923,1.3742256,1.2128719,1.0497054,0.8883517,0.72518504,0.66173136,0.6000906,0.53663695,0.4749962,0.41335547,0.45324063,0.49312583,0.533011,0.5728962,0.61278135,1.7168756,2.8227828,3.926877,5.032784,6.1368785,7.362441,8.588004,9.811753,11.037316,12.262879,11.430729,10.596766,9.764616,8.9324665,8.100317,8.673213,9.244296,9.817192,10.390089,10.962985,11.274815,11.586644,11.900287,12.212116,12.525759,14.68681,16.849674,19.012539,21.175404,23.338266,31.112251,38.888046,46.66203,54.437828,62.21181,68.22722,74.24263,80.25804,86.27345,92.28705,81.88789,71.48693,61.087772,50.68681,40.287655,39.23795,38.188244,37.136726,36.08702,35.037315,37.628036,40.21695,42.80767,45.396584,47.987305,42.624565,37.26182,31.899076,26.538147,21.175404,16.978395,12.779573,8.582565,4.3855567,0.18673515,0.19579996,0.2030518,0.21030366,0.21755551,0.22480737,0.23024625,0.23568514,0.23931105,0.24474995,0.25018883,0.37165734,0.4949388,0.61822027,0.73968875,0.8629702,1.9471219,3.0330863,4.117238,5.2032027,6.2873545,5.0944247,3.9033084,2.7103791,1.5174497,0.3245203,0.27919623,0.23568514,0.19036107,0.14503701,0.099712946,0.13415924,0.17041849,0.20486477,0.23931105,0.2755703,0.23568514,0.19579996,0.15410182,0.11421664,0.07433146,0.13053331,0.18492219,0.23931105,0.2955129,0.34990177,0.8103943,1.2708868,1.7295663,2.1900587,2.6505513,2.6741197,2.6995013,2.7248828,2.7502642,2.7756457,2.4366217,2.0994108,1.7621996,1.4249886,1.0877775,2.0468347,3.007705,3.966762,4.9276323,5.8866897,7.02523,8.161958,9.300498,10.437225,11.575767,13.716875,15.859797,18.002718,20.14564,22.286749,21.360325,20.432089,19.505665,18.577427,17.64919,16.532406,15.415621,14.297023,13.180238,12.06164,12.268318,12.473183,12.678047,12.882912,13.087777,14.53996,15.992143,17.444326,18.898321,20.350506,19.964344,19.579996,19.195648,18.809486,18.425138,19.239159,20.054993,20.870825,21.684845,22.500679,21.75555,21.010424,20.265295,19.520168,18.77504,20.767487,22.759932,24.752378,26.744823,28.73727,28.157122,27.576973,26.996826,26.416677,25.838343,26.539959,27.241575,27.945005,28.646622,29.350052,27.88699,26.425743,24.962683,23.49962,22.03656,19.485722,16.933071,14.380419,11.827768,9.275117,8.245354,7.215591,6.185828,5.1542525,4.12449,3.5570326,2.9895754,2.422118,1.8546607,1.2872034,5.0146546,8.7421055,12.469557,16.197008,19.92446,18.084301,16.245958,14.405801,12.565643,10.725487,11.3600235,11.99456,12.63091,13.265448,13.899984,13.597219,13.294455,12.99169,12.690738,12.387974,12.638163,12.888351,13.136727,13.386916,13.637105,12.703429,11.7679405,10.832452,9.896963,8.963287,10.672911,12.382534,14.092158,15.801782,17.513218,14.802839,12.092461,9.382081,6.6717024,3.9631362,6.9617763,9.96223,12.962683,15.963136,18.961775,16.374678,13.7875805,11.200482,8.611572,6.0244746,5.431636,4.84061,4.2477713,3.6549325,3.0620937,3.0983531,3.1327994,3.1672456,3.2016919,3.2379513,2.811905,2.3876717,1.9616255,1.5373923,1.1131591,1.0605831,1.0080072,0.9554313,0.90285534,0.85027945,0.7995165,0.7505665,0.69980353,0.6508536,0.6000906,1.452183,2.3042755,3.1581807,4.0102735,4.8623657,4.41819,3.972201,3.5280252,3.0820365,2.6378605,2.520018,2.4021754,2.2843328,2.1683033,2.0504606,2.3079014,2.565342,2.8227828,3.0802233,3.3376641,2.7321346,2.128418,1.5228885,0.91735905,0.31182957,0.40972954,0.5076295,0.6055295,0.7016165,0.7995165,0.73968875,0.67986095,0.6200332,0.56020546,0.50037766,0.48587397,0.46955732,0.4550536,0.4405499,0.42423326,2.035957,3.644055,5.2557783,6.8656893,8.4756,6.8548117,5.235836,3.6150475,1.9942589,0.37528324,0.7016165,1.0297627,1.357909,1.6842422,2.0123885,2.0595255,2.1066625,2.1556125,2.2027495,2.2498865,1.93987,1.6298534,1.3198367,1.0098201,0.69980353,1.2491312,1.8002719,2.3495996,2.9007401,3.4500678,3.7183862,3.9848917,4.25321,4.519716,4.788034,4.3982472,4.006647,3.6168604,3.2270734,2.8372865,4.4326935,6.0281005,7.6216946,9.217102,10.812509,9.735609,8.656897,7.5799966,6.5030966,5.424384,4.876869,4.329355,3.7818398,3.2343252,2.6868105,2.6396735,2.5925364,2.5453994,2.4982624,2.4493124,1.9652514,1.4793775,0.99531645,0.5094425,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.09064813,0.11784257,0.14503701,0.17223145,0.19942589,0.17041849,0.13959812,0.11059072,0.07977036,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.11240368,0.22480737,0.33721104,0.44961473,0.5620184,0.44961473,0.33721104,0.22480737,0.11240368,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.2520018,0.40429065,0.55839247,0.7106813,0.8629702,0.7306239,0.5982776,0.46411842,0.33177215,0.19942589,0.19036107,0.1794833,0.17041849,0.15954071,0.15047589,0.15228885,0.15410182,0.15772775,0.15954071,0.16316663,0.13053331,0.09789998,0.065266654,0.032633327,0.0,0.27738327,0.55476654,0.8321498,1.1095331,1.3869164,1.1530442,0.91735905,0.68167394,0.44780177,0.21211663,0.26287958,0.31182957,0.36259252,0.41335547,0.46230546,0.38978696,0.31726846,0.24474995,0.17223145,0.099712946,0.11965553,0.13959812,0.15954071,0.1794833,0.19942589,0.26287958,0.3245203,0.387974,0.44961473,0.51306844,0.56927025,0.62728506,0.6852999,0.7433147,0.7995165,0.79226464,0.7850128,0.7777609,0.7705091,0.76325727,0.9808127,1.1983683,1.4141108,1.6316663,1.8492218,1.7567607,1.6642996,1.5718386,1.4793775,1.3869164,1.8147756,2.2426348,2.6704938,3.0983531,3.5243993,3.4772623,3.4301252,3.3829882,3.3358512,3.2869012,3.1146698,2.9424384,2.770207,2.5979755,2.4257438,2.4021754,2.38042,2.3568513,2.335096,2.3133402,2.231757,2.1519866,2.0722163,1.9924458,1.9126755,1.6733645,1.4322405,1.1929294,0.95180535,0.7124943,0.72518504,0.73787576,0.7505665,0.76325727,0.774135,1.3125849,1.8492218,2.3876717,2.9243085,3.4627585,3.2633326,3.0620937,2.8626678,2.663242,2.4620032,2.4021754,2.3423476,2.2825198,2.222692,2.1628644,1.9416829,1.7223145,1.502946,1.2817645,1.062396,1.0116332,0.96268314,0.9119202,0.8629702,0.8122072,0.7469406,0.68167394,0.61822027,0.5529536,0.48768693,0.42423326,0.36259252,0.2991388,0.2374981,0.17585737,0.22662032,0.27919623,0.33177215,0.38434806,0.43692398,0.5402629,0.6417888,0.7451276,0.8466535,0.9499924,1.1947423,1.4394923,1.6842422,1.9308052,2.175555,2.1556125,2.13567,2.1157274,2.0957847,2.0758421,2.659616,3.245203,3.83079,4.4145637,5.0001507,4.15531,3.3104696,2.465629,1.6207886,0.774135,4.1879435,3.6875658,3.1871881,2.6868105,2.1882458,1.6878681,1.6171626,1.54827,1.4775645,1.4068589,1.3379664,1.1874905,1.0370146,0.8883517,0.73787576,0.5873999,0.5747091,0.5620184,0.5493277,0.53663695,0.52575916,0.5475147,0.56927025,0.59283876,0.61459434,0.63816285,1.9579996,3.2778363,4.597673,5.91751,7.2373466,7.7757964,8.312433,8.8508835,9.38752,9.924157,9.89515,9.864329,9.835322,9.804502,9.775495,10.014805,10.255929,10.49524,10.734551,10.975676,11.675479,12.375282,13.075087,13.77489,14.474693,17.27572,20.074934,22.875961,25.675177,28.47439,37.024323,45.574253,54.126,62.67593,71.22586,74.28433,77.34461,80.40489,83.46517,86.52545,76.699196,66.87475,57.05031,47.22405,37.399605,37.23825,37.075085,36.91192,36.750565,36.5874,36.46049,36.33177,36.204865,36.077957,35.949234,32.749355,29.549477,26.349598,23.14972,19.94984,15.984891,12.019942,8.054993,4.0900435,0.12509441,0.14322405,0.15954071,0.17767033,0.19579996,0.21211663,0.24474995,0.27738327,0.3100166,0.34264994,0.37528324,0.4405499,0.5058166,0.56927025,0.6345369,0.69980353,1.403233,2.1048496,2.808279,3.5098956,4.213325,3.4174345,2.6233568,1.8274662,1.0315757,0.2374981,0.21936847,0.2030518,0.18492219,0.16679256,0.15047589,0.2030518,0.25562772,0.30820364,0.36077955,0.41335547,0.34083697,0.26831847,0.19579996,0.12328146,0.05076295,0.14503701,0.23931105,0.33539808,0.42967212,0.52575916,1.214685,1.9054236,2.5943494,3.2850883,3.975827,4.0120864,4.0501585,4.0882306,4.12449,4.162562,3.6005437,3.0367124,2.474694,1.9126755,1.3506571,2.5526514,3.7546456,4.9584527,6.1604466,7.362441,8.350506,9.336758,10.324821,11.312886,12.299138,13.557334,14.81553,16.071913,17.330109,18.586493,19.01435,19.442211,19.87007,20.29793,20.725788,19.255476,17.785164,16.31485,14.844538,13.374225,13.907236,14.440247,14.973258,15.504456,16.037468,17.322857,18.608248,19.891825,21.177216,22.462606,21.996675,21.532557,21.068438,20.602507,20.138388,20.809185,21.481794,22.154404,22.827011,23.49962,21.420153,19.340685,17.259403,15.179935,13.100468,15.294152,17.48965,19.685148,21.880646,24.07433,22.879587,21.684845,20.490103,19.29536,18.100618,19.347937,20.595255,21.842573,23.089891,24.33721,22.625772,20.912523,19.199274,17.487837,15.774588,14.177367,12.580148,10.982927,9.385707,7.7866745,6.979906,6.1731377,5.3645563,4.557788,3.7492065,3.3304121,2.909805,2.4891977,2.0704033,1.649796,6.947273,12.244749,17.542227,22.839703,28.137178,24.552952,20.966911,17.382685,13.796645,10.212419,11.989121,13.767638,15.544341,17.322857,19.099562,18.08974,17.07992,16.0701,15.06028,14.05046,14.68681,15.324973,15.963136,16.599485,17.237648,15.92325,14.607039,13.292642,11.978244,10.662033,12.152288,13.642544,15.132799,16.623055,18.11331,15.460945,12.806767,10.154404,7.502039,4.8496747,6.787732,8.725789,10.662033,12.60009,14.538147,12.487686,10.437225,8.386765,6.338117,4.2876563,4.255023,4.2223897,4.1897564,4.157123,4.12449,4.0392804,3.9558845,3.870675,3.785466,3.7002566,3.1744974,2.6505513,2.124792,1.6008459,1.0750868,1.015259,0.9554313,0.89560354,0.83577573,0.774135,0.72518504,0.6744221,0.62547207,0.5747091,0.52575916,1.7476959,2.9696326,4.1933823,5.4153194,6.637256,6.069799,5.5023413,4.934884,4.367427,3.7999697,3.3177216,2.8354735,2.3532255,1.8691645,1.3869164,1.7295663,2.0722163,2.4148662,2.7575161,3.100166,2.5417736,1.9851941,1.4268016,0.87022203,0.31182957,0.41516843,0.5166943,0.6200332,0.72337204,0.824898,0.7469406,0.67079616,0.59283876,0.5148814,0.43692398,0.45324063,0.46774435,0.48224804,0.49675176,0.51306844,1.9271792,3.343103,4.7572136,6.1731377,7.5872483,6.156821,4.7282066,3.2977788,1.8673514,0.43692398,0.6726091,0.90829426,1.1421664,1.3778516,1.6117238,1.6280404,1.6425442,1.6570477,1.6733645,1.6878681,1.4848163,1.2817645,1.0805258,0.8774739,0.6744221,1.0750868,1.4757515,1.8746033,2.275268,2.6741197,2.8953013,3.1146698,3.3358512,3.5552197,3.774588,3.6023567,3.4301252,3.2578938,3.0856624,2.911618,3.8054085,4.6973863,5.5893636,6.4831543,7.3751316,7.453089,7.5292335,7.607191,7.6851482,7.763106,6.6717024,5.582112,4.4925213,3.4029307,2.3133402,2.4982624,2.6831846,2.8681068,3.053029,3.2379513,2.5979755,1.9579996,1.3180238,0.678048,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.11059072,0.15772775,0.20486477,0.2520018,0.2991388,0.25562772,0.21030366,0.16497959,0.11965553,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07433146,0.15047589,0.22480737,0.2991388,0.37528324,0.2991388,0.22480737,0.15047589,0.07433146,0.0,0.018129626,0.034446288,0.052575916,0.07070554,0.0870222,0.21030366,0.33177215,0.4550536,0.57833505,0.69980353,0.6200332,0.5402629,0.4604925,0.38072214,0.2991388,0.27194437,0.24474995,0.21755551,0.19036107,0.16316663,0.17223145,0.18310922,0.19217403,0.2030518,0.21211663,0.17041849,0.12690738,0.08520924,0.04169814,0.0,0.2229944,0.44417584,0.6671702,0.8901646,1.1131591,0.9481794,0.78319985,0.61822027,0.45324063,0.28826106,0.3245203,0.36259252,0.40066472,0.43692398,0.4749962,0.39703882,0.3208944,0.24293698,0.16497959,0.0870222,0.10515183,0.12328146,0.13959812,0.15772775,0.17585737,0.2374981,0.2991388,0.36259252,0.42423326,0.48768693,0.5293851,0.5728962,0.61459434,0.65810543,0.69980353,0.69436467,0.69073874,0.6852999,0.67986095,0.6744221,0.8321498,0.9898776,1.1476053,1.305333,1.4630609,1.4431182,1.4231756,1.403233,1.3832904,1.3633479,1.696933,2.032331,2.3677292,2.7031271,3.0367124,3.0602808,3.0820365,3.105605,3.1273603,3.149116,3.0348995,2.9206827,2.8046532,2.6904364,2.5744069,2.5979755,2.619731,2.6432993,2.665055,2.6868105,2.518205,2.3477864,2.1773682,2.0069497,1.8383441,1.5772774,1.3180238,1.0569572,0.79770356,0.53663695,0.53663695,0.53663695,0.53663695,0.53663695,0.53663695,1.0370146,1.5373923,2.03777,2.5381477,3.0367124,2.8245957,2.612479,2.4003625,2.1882458,1.9743162,1.8981718,1.8202144,1.742257,1.6642996,1.5881553,1.4322405,1.2781386,1.1222239,0.968122,0.8122072,0.774135,0.73787576,0.69980353,0.66173136,0.62547207,0.60190356,0.58014804,0.55839247,0.53482395,0.51306844,0.46230546,0.41335547,0.36259252,0.31182957,0.26287958,0.27194437,0.28282216,0.291887,0.30276474,0.31182957,0.44780177,0.581961,0.7179332,0.8520924,0.9880646,1.1421664,1.2980812,1.452183,1.6080978,1.7621996,1.8691645,1.9779422,2.084907,2.1918716,2.3006494,2.8771715,3.4555066,4.0320287,4.610364,5.186886,4.2949085,3.4029307,2.5091403,1.6171626,0.72518504,4.8134155,4.0374675,3.2633326,2.4873846,1.7132497,0.93730164,0.97718686,1.017072,1.0569572,1.0968424,1.1367276,1.0007553,0.8629702,0.72518504,0.5873999,0.44961473,0.48768693,0.52575916,0.5620184,0.6000906,0.63816285,0.6417888,0.64722764,0.6526665,0.65810543,0.66173136,2.1973107,3.73289,5.2666564,6.8022356,8.337815,8.187339,8.036863,7.8882003,7.7377243,7.5872483,8.3595705,9.131892,9.904215,10.6783495,11.450671,11.358211,11.26575,11.173288,11.080828,10.988366,12.07433,13.162108,14.249886,15.337664,16.425442,19.862818,23.300196,26.737572,30.17495,33.612328,42.938206,52.26227,61.58815,70.91222,80.2381,80.34325,80.4484,80.55174,80.65689,80.76205,71.51231,62.262573,53.01284,43.763103,34.511555,35.23674,35.961926,36.68711,37.412296,38.13748,35.292942,32.448402,29.602053,26.757515,23.912977,22.87415,21.837133,20.80012,19.763105,18.724277,14.9932,11.26031,7.5274205,3.7945306,0.06164073,0.09064813,0.11784257,0.14503701,0.17223145,0.19942589,0.25925365,0.3208944,0.38072214,0.4405499,0.50037766,0.5076295,0.5148814,0.52213323,0.5293851,0.53663695,0.8575313,1.1766127,1.4975071,1.8165885,2.137483,1.7404441,1.3415923,0.9445535,0.5475147,0.15047589,0.15954071,0.17041849,0.1794833,0.19036107,0.19942589,0.27013144,0.34083697,0.40972954,0.48043507,0.5493277,0.44417584,0.34083697,0.23568514,0.13053331,0.025381476,0.15954071,0.2955129,0.42967212,0.5656443,0.69980353,1.6207886,2.5399606,3.4609456,4.3801174,5.2992897,5.3500524,5.4008155,5.4497657,5.5005283,5.5494785,4.762653,3.975827,3.1871881,2.4003625,1.6117238,3.056655,4.501586,5.9483304,7.3932614,8.838193,9.675781,10.51337,11.349146,12.186734,13.024323,13.397794,13.769451,14.142921,14.514579,14.888049,16.67019,18.452333,20.234476,22.01843,23.800573,21.976732,20.154705,18.332678,16.51065,14.68681,15.547967,16.40731,17.266655,18.127813,18.987158,20.105755,21.22254,22.339325,23.457922,24.574707,24.030819,23.485117,22.939415,22.395527,21.849825,22.37921,22.910408,23.439793,23.96918,24.500376,21.084755,17.670946,14.255324,10.839704,7.424082,9.822631,12.219368,14.617917,17.014654,19.413204,17.602055,15.792717,13.981567,12.172231,10.362894,12.154101,13.947122,15.740141,17.533161,19.324368,17.362743,15.399304,13.437678,11.47424,9.512614,8.870826,8.227224,7.5854354,6.9418335,6.300045,5.714458,5.130684,4.5450974,3.9595103,3.3757362,3.101979,2.8300345,2.5580902,2.2843328,2.0123885,8.87989,15.747393,22.614895,29.482397,36.3499,31.01979,25.68968,20.35957,15.02946,9.699349,12.620032,15.540715,18.459585,21.380268,24.300951,22.582262,20.865387,19.146698,17.429823,15.712947,16.73727,17.763407,18.787731,19.812056,20.838192,19.143072,17.447952,15.752831,14.057712,12.362592,13.631665,14.902553,16.173439,17.442513,18.7134,16.117237,13.522888,10.926725,8.3323765,5.7380266,6.6118746,7.4875355,8.363196,9.237044,10.112705,8.600695,7.0868707,5.57486,4.062849,2.5508385,3.0765975,3.6041696,4.1317415,4.6593137,5.186886,4.9820213,4.7771564,4.572292,4.367427,4.162562,3.53709,2.911618,2.2879589,1.6624867,1.0370146,0.969935,0.90285534,0.83577573,0.7668832,0.69980353,0.6508536,0.6000906,0.5493277,0.50037766,0.44961473,2.0432088,3.63499,5.2267714,6.8203654,8.412147,7.723221,7.0324817,6.341743,5.6528172,4.9620786,4.115425,3.2669585,2.420305,1.5718386,0.72518504,1.1530442,1.5790904,2.0069497,2.4348087,2.8626678,2.3532255,1.84197,1.3325275,0.823085,0.31182957,0.42060733,0.5275721,0.6345369,0.7433147,0.85027945,0.7541924,0.65991837,0.5656443,0.46955732,0.37528324,0.42060733,0.46411842,0.5094425,0.55476654,0.6000906,1.8202144,3.0403383,4.2604623,5.480586,6.70071,5.4606433,4.220577,2.9805105,1.7404441,0.50037766,0.6417888,0.7850128,0.92823684,1.0696479,1.2128719,1.1947423,1.1766127,1.1602961,1.1421664,1.1258497,1.0297627,0.9354887,0.83940166,0.7451276,0.6508536,0.89922947,1.1494182,1.3996071,1.649796,1.8999848,2.0722163,2.2444477,2.4166791,2.5907235,2.762955,2.808279,2.8517902,2.8971143,2.9424384,2.9877625,3.1781235,3.3666716,3.5570326,3.7473936,3.9377546,5.1705694,6.401571,7.6343856,8.8672,10.100015,8.466536,6.834869,5.2032027,3.5697234,1.938057,2.3550384,2.7720199,3.1908143,3.6077955,4.024777,3.2306993,2.4348087,1.6407311,0.8448406,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.13053331,0.19761293,0.26469254,0.33177215,0.40066472,0.34083697,0.27919623,0.21936847,0.15954071,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.16679256,0.25925365,0.35171473,0.44417584,0.53663695,0.5094425,0.48224804,0.4550536,0.42785916,0.40066472,0.35534066,0.3100166,0.26469254,0.21936847,0.17585737,0.19217403,0.21030366,0.22662032,0.24474995,0.26287958,0.21030366,0.15772775,0.10515183,0.052575916,0.0,0.16679256,0.33539808,0.50219065,0.67079616,0.8375887,0.7433147,0.64722764,0.5529536,0.45686656,0.36259252,0.387974,0.41335547,0.43692398,0.46230546,0.48768693,0.40429065,0.32270733,0.23931105,0.15772775,0.07433146,0.09064813,0.10515183,0.11965553,0.13415924,0.15047589,0.21211663,0.2755703,0.33721104,0.40066472,0.46230546,0.4894999,0.5166943,0.54570174,0.5728962,0.6000906,0.5982776,0.5946517,0.59283876,0.58921283,0.5873999,0.6852999,0.78319985,0.8792868,0.97718686,1.0750868,1.1276628,1.1802386,1.2328146,1.2853905,1.3379664,1.5809034,1.8220274,2.0649643,2.3079014,2.5508385,2.6432993,2.7357605,2.8282216,2.9206827,3.0131438,2.955129,2.8971143,2.8390994,2.7828975,2.7248828,2.7919624,2.8608549,2.9279346,2.9950142,3.0620937,2.8028402,2.5417736,2.2825198,2.0232663,1.7621996,1.4830034,1.2019942,0.922798,0.6417888,0.36259252,0.34990177,0.33721104,0.3245203,0.31182957,0.2991388,0.76325727,1.2255627,1.6878681,2.1501737,2.612479,2.3876717,2.1628644,1.938057,1.7132497,1.4866294,1.3923552,1.2980812,1.2019942,1.1077201,1.0116332,0.922798,0.8321498,0.7433147,0.6526665,0.5620184,0.53663695,0.51306844,0.48768693,0.46230546,0.43692398,0.45686656,0.47680917,0.49675176,0.5166943,0.53663695,0.50037766,0.46230546,0.42423326,0.387974,0.34990177,0.31726846,0.28463513,0.2520018,0.21936847,0.18673515,0.35534066,0.52213323,0.69073874,0.8575313,1.0243238,1.0895905,1.1548572,1.2201238,1.2853905,1.3506571,1.5845293,1.8202144,2.0558996,2.2897718,2.525457,3.094727,3.6658103,4.2350807,4.804351,5.375434,4.4345064,3.4953918,2.5544643,1.6153497,0.6744221,5.4370747,4.3873696,3.3376641,2.2879589,1.2382535,0.18673515,0.33721104,0.48768693,0.63816285,0.7868258,0.93730164,0.8122072,0.6871128,0.5620184,0.43692398,0.31182957,0.40066472,0.48768693,0.5747091,0.66173136,0.7505665,0.73787576,0.72518504,0.7124943,0.69980353,0.6871128,2.4366217,4.1879435,5.9374523,7.686961,9.438283,8.600695,7.763106,6.925517,6.0879283,5.2503395,6.825804,8.399456,9.97492,11.5503845,13.125849,12.699803,12.27557,11.849524,11.42529,10.999244,12.474996,13.9507475,15.4246855,16.900436,18.374376,22.449915,26.525455,30.600996,34.67472,38.750263,48.850277,58.95029,69.05031,79.15032,89.250336,86.40036,83.55038,80.7004,77.850426,75.00045,66.325424,57.6504,48.975372,40.300346,31.625319,33.23704,34.85058,36.462303,38.07584,39.687565,34.125393,28.563225,22.999243,17.437075,11.874905,13.000754,14.124791,15.250641,16.374678,17.500528,13.999697,10.500679,6.9998484,3.5008307,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.2755703,0.36259252,0.44961473,0.53663695,0.62547207,0.5747091,0.52575916,0.4749962,0.42423326,0.37528324,0.31182957,0.25018883,0.18673515,0.12509441,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.099712946,0.13778515,0.17585737,0.21211663,0.25018883,0.33721104,0.42423326,0.51306844,0.6000906,0.6871128,0.5493277,0.41335547,0.2755703,0.13778515,0.0,0.17585737,0.34990177,0.52575916,0.69980353,0.87566096,2.0250793,3.1744974,4.325729,5.475147,6.624565,6.688019,6.7496595,6.813113,6.874754,6.9382076,5.924762,4.9131284,3.8996825,2.8880494,1.8746033,3.5624714,5.2503395,6.9382076,8.624263,10.312131,10.999244,11.6881695,12.375282,13.062395,13.749508,13.238253,12.725184,12.212116,11.700861,11.187792,14.324218,17.462456,20.600695,23.73712,26.875357,24.699802,22.524246,20.350506,18.17495,15.999394,17.186886,18.374376,19.561867,20.749357,21.936848,22.886839,23.836832,24.786825,25.736816,26.68681,26.06315,25.437677,24.812206,24.186733,23.563074,23.949236,24.33721,24.725183,25.113157,25.49932,20.749357,15.999394,11.249433,6.4994707,1.7495089,4.349297,6.9490857,9.550687,12.1504755,14.750263,12.32452,9.900589,7.474845,5.049101,2.6251698,4.9620786,7.3008003,9.637709,11.974618,14.313339,12.099712,9.8878975,7.6742706,5.462456,3.2506418,3.5624714,3.874301,4.1879435,4.499773,4.8116026,4.4508233,4.0882306,3.7256382,3.3630457,3.000453,2.8753586,2.7502642,2.6251698,2.5000753,2.374981,10.812509,19.250036,27.687565,36.12509,44.562622,37.48844,30.412447,23.336454,16.262274,9.188094,13.24913,17.31198,21.374828,25.437677,29.500526,27.074783,24.650852,22.22511,19.799364,17.375433,18.787731,20.20003,21.612328,23.024624,24.436922,22.362894,20.287052,18.213022,16.13718,14.06315,15.112856,16.162561,17.212267,18.261972,19.311678,16.775343,14.237195,11.699047,9.162713,6.624565,6.43783,6.249282,6.0625467,5.8758116,5.6872635,4.7118897,3.738329,2.762955,1.7875811,0.8122072,1.8999848,2.9877625,4.07554,5.163317,6.249282,5.924762,5.600241,5.275721,4.949388,4.6248674,3.8996825,3.1744974,2.4493124,1.7241274,1.0007553,0.9246109,0.85027945,0.774135,0.69980353,0.62547207,0.5747091,0.52575916,0.4749962,0.42423326,0.37528324,2.3369088,4.3003473,6.261973,8.225411,10.1870365,9.374829,8.562622,7.750415,6.9382076,6.1241875,4.9131284,3.7002566,2.4873846,1.2745126,0.06164073,0.5747091,1.0877775,1.6008459,2.1121013,2.6251698,2.1628644,1.7005589,1.2382535,0.774135,0.31182957,0.42423326,0.53663695,0.6508536,0.76325727,0.87566096,0.76325727,0.6508536,0.53663695,0.42423326,0.31182957,0.387974,0.46230546,0.53663695,0.61278135,0.6871128,1.7132497,2.7375734,3.7618973,4.788034,5.812358,4.762653,3.7129474,2.663242,1.6117238,0.5620184,0.61278135,0.66173136,0.7124943,0.76325727,0.8122072,0.76325727,0.7124943,0.66173136,0.61278135,0.5620184,0.5747091,0.5873999,0.6000906,0.61278135,0.62547207,0.72518504,0.824898,0.9246109,1.0243238,1.1258497,1.2491312,1.3742256,1.49932,1.6244144,1.7495089,2.0123885,2.275268,2.5381477,2.7992141,3.0620937,2.5508385,2.03777,1.5247015,1.0116332,0.50037766,2.8880494,5.275721,7.663393,10.049252,12.436923,10.263181,8.087626,5.9120708,3.738329,1.5627737,2.2118144,2.8626678,3.5117085,4.162562,4.8116026,3.8616104,2.913431,1.9616255,1.0116332,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.15047589,0.2374981,0.3245203,0.41335547,0.50037766,0.42423326,0.34990177,0.2755703,0.19942589,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.12509441,0.18673515,0.25018883,0.31182957,0.37528324,0.40066472,0.42423326,0.44961473,0.4749962,0.50037766,0.43692398,0.37528324,0.31182957,0.25018883,0.18673515,0.21211663,0.2374981,0.26287958,0.28826106,0.31182957,0.25018883,0.18673515,0.12509441,0.06164073,0.0,0.11240368,0.22480737,0.33721104,0.44961473,0.5620184,0.53663695,0.51306844,0.48768693,0.46230546,0.43692398,0.44961473,0.46230546,0.4749962,0.48768693,0.50037766,0.41335547,0.3245203,0.2374981,0.15047589,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.18673515,0.25018883,0.31182957,0.37528324,0.43692398,0.44961473,0.46230546,0.4749962,0.48768693,0.50037766,0.50037766,0.50037766,0.50037766,0.50037766,0.50037766,0.53663695,0.5747091,0.61278135,0.6508536,0.6871128,0.8122072,0.93730164,1.062396,1.1874905,1.3125849,1.4630609,1.6117238,1.7621996,1.9126755,2.0631514,2.2245052,2.3876717,2.5508385,2.712192,2.8753586,2.8753586,2.8753586,2.8753586,2.8753586,2.8753586,2.9877625,3.100166,3.2125697,3.3249733,3.437377,3.0874753,2.7375734,2.3876717,2.03777,1.6878681,1.3869164,1.0877775,0.7868258,0.48768693,0.18673515,0.16316663,0.13778515,0.11240368,0.0870222,0.06164073,0.48768693,0.9119202,1.3379664,1.7621996,2.1882458,1.9507477,1.7132497,1.4757515,1.2382535,1.0007553,0.8883517,0.774135,0.66173136,0.5493277,0.43692398,0.41335547,0.387974,0.36259252,0.33721104,0.31182957,0.2991388,0.28826106,0.2755703,0.26287958,0.25018883,0.31182957,0.37528324,0.43692398,0.50037766,0.5620184,0.53663695,0.51306844,0.48768693,0.46230546,0.43692398,0.36259252,0.28826106,0.21211663,0.13778515,0.06164073,0.26287958,0.46230546,0.66173136,0.8629702,1.062396,1.0370146,1.0116332,0.9880646,0.96268314,0.93730164,1.2998942,1.6624867,2.0250793,2.3876717,2.7502642,3.3122826,3.874301,4.4381323,5.0001507,5.562169,4.574105,3.587853,2.5997884,1.6117238,0.62547207,4.461701,3.6458678,2.8282216,2.0105755,1.1929294,0.37528324,0.46411842,0.55476654,0.64541465,0.73424983,0.824898,0.73787576,0.6508536,0.5620184,0.4749962,0.387974,0.50219065,0.61822027,0.7324369,0.8466535,0.96268314,0.96087015,0.9572442,0.9554313,0.95180535,0.9499924,2.4130533,3.874301,5.337362,6.8004227,8.26167,7.8827615,7.502039,7.12313,6.742408,6.3616858,7.6307597,8.898021,10.165281,11.432542,12.699803,12.371656,12.045323,11.717177,11.390844,11.062697,12.692551,14.322405,15.952258,17.582111,19.211964,22.388275,25.562773,28.73727,31.911768,35.088078,42.802235,50.518204,58.232357,65.948326,73.66248,70.972046,68.283424,65.59299,62.90255,60.212112,53.42982,46.647526,39.865234,33.082943,26.300648,28.349297,30.399757,32.45022,34.50068,36.549324,31.862818,27.174496,22.487988,17.799667,13.113158,13.611723,14.112101,14.612478,15.112856,15.613234,12.513068,9.412902,6.3127356,3.2125697,0.11240368,0.25018883,0.387974,0.52575916,0.66173136,0.7995165,0.7469406,0.69436467,0.6417888,0.58921283,0.53663695,0.50037766,0.46230546,0.42423326,0.387974,0.34990177,0.32814622,0.3045777,0.28282216,0.25925365,0.2374981,0.32995918,0.4224203,0.5148814,0.6073425,0.69980353,0.6091554,0.52032024,0.42967212,0.34083697,0.25018883,0.3245203,0.40066472,0.4749962,0.5493277,0.62547207,0.52575916,0.42423326,0.3245203,0.22480737,0.12509441,0.75963134,1.3941683,2.030518,2.665055,3.299592,4.077353,4.855114,5.632875,6.4106355,7.1883965,6.9545245,6.722465,6.490406,6.258347,6.0244746,5.1198063,4.215138,3.3104696,2.4058013,1.49932,3.045777,4.590421,6.1350656,7.6797094,9.224354,10.127209,11.030065,11.9329195,12.835775,13.736817,13.399607,13.062395,12.725184,12.387974,12.050762,14.9932,17.935638,20.878077,23.820515,26.762953,25.08415,23.40716,21.73017,20.053179,18.374376,19.304426,20.234476,21.164526,22.094576,23.024624,23.747997,24.469557,25.192928,25.914488,26.63786,26.24082,25.841969,25.44493,25.047892,24.650852,24.806767,24.964495,25.122223,25.279951,25.437677,22.295815,19.152136,16.010273,12.866595,9.724731,11.427103,13.129475,14.831847,16.534218,18.236591,15.760084,13.281764,10.805257,8.326937,5.8504305,8.357758,10.865085,13.372412,15.879739,18.387066,16.682882,14.976884,13.272699,11.566701,9.862516,10.067381,10.272246,10.477111,10.681975,10.88684,9.295059,7.703278,6.109684,4.517903,2.9243085,2.9968271,3.0693457,3.141864,3.2143826,3.2869012,9.871581,16.458075,23.042755,29.627434,36.212116,31.489347,26.768393,22.045626,17.322857,12.60009,17.527721,22.455355,27.382986,32.31062,37.23825,32.8672,28.49796,24.126905,19.757666,15.388427,17.81417,20.241728,22.669285,25.096842,27.524399,26.184618,24.84484,23.50506,22.165281,20.8255,20.290678,19.755854,19.219215,18.684393,18.149569,16.389181,14.630608,12.870221,11.109835,9.349448,9.461852,9.574255,9.686659,9.799063,9.91328,8.1148205,6.3181744,4.519716,2.72307,0.9246109,1.9217403,2.9206827,3.917812,4.914942,5.9120708,5.634688,5.3573046,5.0799212,4.802538,4.5251546,4.099108,3.6748753,3.2506418,2.8245957,2.4003625,2.0504606,1.7005589,1.3506571,1.0007553,0.6508536,1.0116332,1.3742256,1.7368182,2.0994108,2.4620032,3.7600844,5.0581656,6.354434,7.652515,8.950596,8.140202,7.3298078,6.5194135,5.710832,4.900438,4.3819304,3.8652363,3.346729,2.8300345,2.3133402,2.3931105,2.472881,2.5526514,2.6324217,2.712192,2.2353828,1.7567607,1.2799516,0.8031424,0.3245203,0.4224203,0.52032024,0.61822027,0.71430725,0.8122072,0.7433147,0.6726091,0.60190356,0.533011,0.46230546,0.50037766,0.53663695,0.5747091,0.61278135,0.6508536,1.502946,2.3550384,3.207131,4.059223,4.9131284,4.077353,3.24339,2.4076142,1.5718386,0.73787576,0.7668832,0.79770356,0.82671094,0.8575313,0.8883517,0.85027945,0.8122072,0.774135,0.73787576,0.69980353,0.7124943,0.72518504,0.73787576,0.7505665,0.76325727,0.82671094,0.8919776,0.9572442,1.0225109,1.0877775,1.167548,1.2473183,1.3270886,1.4068589,1.4866294,1.7767034,2.0667772,2.3568513,2.6469254,2.9369993,2.4583774,1.9779422,1.4975071,1.017072,0.53663695,2.4946365,4.4526362,6.4106355,8.366822,10.324821,8.557183,6.789545,5.0219064,3.254268,1.4866294,1.9598125,2.4329958,2.904366,3.3775494,3.8507326,3.0892882,2.3296568,1.5700256,0.8103943,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.01994259,0.027194439,0.034446288,0.04169814,0.05076295,0.13959812,0.23024625,0.3208944,0.40972954,0.50037766,0.44961473,0.40066472,0.34990177,0.2991388,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.027194439,0.04169814,0.058014803,0.072518505,0.0870222,0.15047589,0.21211663,0.2755703,0.33721104,0.40066472,0.40791658,0.41516843,0.4224203,0.42967212,0.43692398,0.387974,0.33721104,0.28826106,0.2374981,0.18673515,0.21574254,0.24293698,0.27013144,0.29732585,0.3245203,0.25925365,0.19579996,0.13053331,0.065266654,0.0,0.092461094,0.18492219,0.27738327,0.36984438,0.46230546,0.47318324,0.48224804,0.49312583,0.50219065,0.51306844,0.52032024,0.5275721,0.53482395,0.5420758,0.5493277,0.44961473,0.34990177,0.25018883,0.15047589,0.05076295,0.065266654,0.07977036,0.09427405,0.11059072,0.12509441,0.17223145,0.21936847,0.26831847,0.3154555,0.36259252,0.40791658,0.45324063,0.49675176,0.5420758,0.5873999,0.5656443,0.5420758,0.52032024,0.49675176,0.4749962,0.5094425,0.54570174,0.58014804,0.61459434,0.6508536,0.7451276,0.83940166,0.9354887,1.0297627,1.1258497,1.2382535,1.3506571,1.4630609,1.5754645,1.6878681,1.8691645,2.0522738,2.2353828,2.4166791,2.5997884,2.6052272,2.610666,2.6142921,2.619731,2.6251698,2.712192,2.7992141,2.8880494,2.9750717,3.0620937,2.811905,2.561716,2.3133402,2.0631514,1.8129625,1.4848163,1.1566701,0.83033687,0.50219065,0.17585737,0.15410182,0.13415924,0.11421664,0.09427405,0.07433146,0.41335547,0.7505665,1.0877775,1.4249886,1.7621996,1.5790904,1.3977941,1.214685,1.0333886,0.85027945,0.7668832,0.6852999,0.60190356,0.52032024,0.43692398,0.4405499,0.44236287,0.44417584,0.44780177,0.44961473,0.43329805,0.41516843,0.39703882,0.38072214,0.36259252,0.3825351,0.40247768,0.4224203,0.44236287,0.46230546,0.4405499,0.4169814,0.39522585,0.37165734,0.34990177,0.29007402,0.23024625,0.17041849,0.11059072,0.05076295,0.21211663,0.37528324,0.53663695,0.69980353,0.8629702,1.1131591,1.3633479,1.6117238,1.8619126,2.1121013,3.0167696,3.923251,4.8279195,5.732588,6.637256,6.2257137,5.812358,5.4008155,4.98746,4.5759177,3.7691493,2.9641938,2.1592383,1.3542831,0.5493277,3.48814,2.902553,2.3169663,1.7331922,1.1476053,0.5620184,0.59283876,0.62184614,0.6526665,0.68167394,0.7124943,0.66173136,0.61278135,0.5620184,0.51306844,0.46230546,0.6055295,0.7469406,0.8901646,1.0333886,1.1747998,1.1820517,1.1893034,1.1983683,1.2056202,1.2128719,2.3876717,3.5624714,4.7372713,5.9120708,7.0868707,7.1648283,7.2427855,7.320743,7.3968873,7.474845,8.435715,9.394773,10.355642,11.314699,12.27557,12.045323,11.815077,11.584831,11.354585,11.124338,12.910107,14.694061,16.47983,18.265598,20.049553,22.324821,24.60009,26.875357,29.150625,31.42408,36.75419,42.0843,47.41441,52.744522,58.07463,55.545547,53.014652,50.48557,47.954674,45.42559,40.534218,35.644657,30.755096,25.865538,20.974165,23.461548,25.950747,28.438131,30.925516,33.4129,29.60024,25.78758,21.97492,18.16226,14.349599,14.224504,14.09941,13.974316,13.849221,13.724127,11.024626,8.325124,5.6256227,2.9243085,0.22480737,0.46230546,0.69980353,0.93730164,1.1747998,1.4122978,1.2201238,1.0279498,0.83577573,0.6417888,0.44961473,0.42423326,0.40066472,0.37528324,0.34990177,0.3245203,0.34264994,0.36077955,0.3770962,0.39522585,0.41335547,0.5982776,0.78319985,0.968122,1.1530442,1.3379664,1.1204109,0.90285534,0.6852999,0.46774435,0.25018883,0.31182957,0.37528324,0.43692398,0.50037766,0.5620184,0.50037766,0.43692398,0.37528324,0.31182957,0.25018883,1.3452182,2.4402475,3.5352771,4.6303062,5.7253356,6.1296263,6.53573,6.9400206,7.344311,7.750415,7.2228427,6.695271,6.167699,5.6401267,5.1125546,4.314851,3.5171473,2.7194438,1.9217403,1.1258497,2.5272698,3.930503,5.331923,6.735156,8.138389,9.255174,10.371959,11.490557,12.607342,13.724127,13.562773,13.399607,13.238253,13.075087,12.91192,15.660371,18.40701,21.15546,23.9021,26.65055,25.470312,24.290073,23.109835,21.929596,20.749357,21.421967,22.094576,22.767183,23.439793,24.112402,24.607342,25.10228,25.59722,26.092157,26.587097,26.416677,26.248072,26.077654,25.907236,25.736816,25.664299,25.59178,25.51926,25.446743,25.374224,23.840458,22.304878,20.769299,19.235533,17.699953,18.50491,19.309864,20.11482,20.919775,21.724731,19.195648,16.664753,14.13567,11.6047735,9.07569,11.751623,14.429369,17.107115,19.78486,22.462606,21.264238,20.067682,18.869314,17.67276,16.474392,16.57229,16.67019,16.768091,16.864178,16.962078,14.139296,11.318325,8.495543,5.67276,2.8499773,3.1201086,3.39024,3.6603715,3.930503,4.2006345,8.9324665,13.664299,18.397943,23.129776,27.861609,25.492067,23.122524,20.752983,18.381628,16.012085,21.8045,27.596916,33.38933,39.181747,44.974163,38.659615,32.345066,26.030518,19.714155,13.399607,16.842422,20.285238,23.728054,27.17087,30.611874,30.008156,29.402628,28.797098,28.19338,27.587852,25.466686,23.347332,21.22798,19.106813,16.98746,16.004833,15.022208,14.039582,13.056956,12.07433,12.487686,12.899229,13.312584,13.72594,14.137483,11.517752,8.898021,6.2782893,3.6567454,1.0370146,1.9453088,2.8517902,3.7600844,4.668379,5.57486,5.3446136,5.1143675,4.8841214,4.655688,4.4254417,4.3003473,4.175253,4.0501585,3.925064,3.7999697,3.1744974,2.5508385,1.9253663,1.2998942,0.6744221,1.4503701,2.2245052,3.000453,3.774588,4.550536,5.18326,5.814171,6.446895,7.079619,7.7123427,6.9055743,6.096993,5.290225,4.4816437,3.6748753,3.8525455,4.0302157,4.207886,4.3855567,4.5632267,4.209699,3.8579843,3.5044568,3.152742,2.7992141,2.3079014,1.8147756,1.3216497,0.83033687,0.33721104,0.42060733,0.50219065,0.5855869,0.6671702,0.7505665,0.72337204,0.69436467,0.6671702,0.6399758,0.61278135,0.61278135,0.61278135,0.61278135,0.61278135,0.61278135,1.2926424,1.9725033,2.6523643,3.3322253,4.0120864,3.392053,2.7720199,2.1519866,1.5319533,0.9119202,0.922798,0.9318628,0.94274056,0.95180535,0.96268314,0.93730164,0.9119202,0.8883517,0.8629702,0.8375887,0.85027945,0.8629702,0.87566096,0.8883517,0.89922947,0.9300498,0.96087015,0.9898776,1.020698,1.0497054,1.0841516,1.1204109,1.1548572,1.1893034,1.2255627,1.5428312,1.8600996,2.1773682,2.4946365,2.811905,2.3641033,1.9181144,1.4703126,1.0225109,0.5747091,2.1030366,3.6295512,5.1578784,6.684393,8.212721,6.8529987,5.4932766,4.1317415,2.7720199,1.4122978,1.7078108,2.0033236,2.2970235,2.5925364,2.8880494,2.3169663,1.7476959,1.1766127,0.6073425,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.027194439,0.030820364,0.032633327,0.034446288,0.038072214,0.13053331,0.2229944,0.3154555,0.40791658,0.50037766,0.4749962,0.44961473,0.42423326,0.40066472,0.37528324,0.2991388,0.22480737,0.15047589,0.07433146,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.04169814,0.059827764,0.07795739,0.09427405,0.11240368,0.17585737,0.2374981,0.2991388,0.36259252,0.42423326,0.41516843,0.40429065,0.39522585,0.38434806,0.37528324,0.33721104,0.2991388,0.26287958,0.22480737,0.18673515,0.21755551,0.24837588,0.27738327,0.30820364,0.33721104,0.27013144,0.2030518,0.13415924,0.06707962,0.0,0.072518505,0.14503701,0.21755551,0.29007402,0.36259252,0.40791658,0.45324063,0.49675176,0.5420758,0.5873999,0.58921283,0.59283876,0.5946517,0.5982776,0.6000906,0.48768693,0.37528324,0.26287958,0.15047589,0.038072214,0.054388877,0.072518505,0.09064813,0.10696479,0.12509441,0.15772775,0.19036107,0.2229944,0.25562772,0.28826106,0.36440548,0.44236287,0.52032024,0.5982776,0.6744221,0.629098,0.5855869,0.5402629,0.4949388,0.44961473,0.48224804,0.5148814,0.5475147,0.58014804,0.61278135,0.678048,0.7433147,0.80676836,0.872035,0.93730164,1.0116332,1.0877775,1.162109,1.2382535,1.3125849,1.5156367,1.7168756,1.9199274,2.1229792,2.324218,2.335096,2.3441606,2.3550384,2.3641033,2.374981,2.4366217,2.5000753,2.561716,2.6251698,2.6868105,2.5381477,2.3876717,2.2371957,2.08672,1.938057,1.5827163,1.2273756,0.872035,0.5166943,0.16316663,0.14684997,0.13234627,0.11784257,0.10333887,0.0870222,0.33721104,0.5873999,0.8375887,1.0877775,1.3379664,1.209246,1.0823387,0.9554313,0.82671094,0.69980353,0.64722764,0.5946517,0.5420758,0.4894999,0.43692398,0.46774435,0.49675176,0.5275721,0.55839247,0.5873999,0.5656443,0.5420758,0.52032024,0.49675176,0.4749962,0.45324063,0.42967212,0.40791658,0.38434806,0.36259252,0.34264994,0.32270733,0.30276474,0.28282216,0.26287958,0.21755551,0.17223145,0.12690738,0.08339628,0.038072214,0.16316663,0.28826106,0.41335547,0.53663695,0.66173136,1.1874905,1.7132497,2.2371957,2.762955,3.2869012,4.7354584,6.1822023,7.6307597,9.077503,10.524248,9.137331,7.750415,6.3616858,4.974769,3.587853,2.9641938,2.3423476,1.7205015,1.0968424,0.4749962,2.5127661,2.1592383,1.8075237,1.455809,1.1022812,0.7505665,0.7197462,0.69073874,0.65991837,0.629098,0.6000906,0.5873999,0.5747091,0.5620184,0.5493277,0.53663695,0.7070554,0.8774739,1.0478923,1.2183108,1.3869164,1.405046,1.4231756,1.4394923,1.4576219,1.4757515,2.3622901,3.2506418,4.137181,5.0255322,5.9120708,6.446895,6.981719,7.518356,8.05318,8.588004,9.24067,9.893337,10.54419,11.1968565,11.849524,11.717177,11.584831,11.452485,11.320138,11.187792,13.127662,15.067532,17.007402,18.947271,20.887142,22.26318,23.637405,25.011631,26.38767,27.761896,30.70796,33.65221,36.596462,39.542526,42.48678,40.117237,37.747692,35.37634,33.006798,30.637255,27.640427,24.641787,21.64496,18.648132,15.649493,18.575615,21.499924,24.424232,27.350353,30.274662,27.337664,24.400663,21.461851,18.52485,15.5878525,14.837286,14.0867195,13.337966,12.5873995,11.836833,9.537996,7.2373466,4.936697,2.6378605,0.33721104,0.6744221,1.0116332,1.3506571,1.6878681,2.0250793,1.693307,1.3597219,1.0279498,0.69436467,0.36259252,0.34990177,0.33721104,0.3245203,0.31182957,0.2991388,0.35715362,0.41516843,0.47318324,0.5293851,0.5873999,0.86478317,1.1421664,1.4195497,1.696933,1.9743162,1.6298534,1.2853905,0.93911463,0.5946517,0.25018883,0.2991388,0.34990177,0.40066472,0.44961473,0.50037766,0.4749962,0.44961473,0.42423326,0.40066472,0.37528324,1.9308052,3.484514,5.040036,6.5955577,8.149267,8.1819,8.214534,8.247167,8.2798,8.312433,7.4893484,6.6680765,5.844991,5.0219064,4.2006345,3.5098956,2.819157,2.1302311,1.4394923,0.7505665,2.0105755,3.2705846,4.5305934,5.7906027,7.0506115,8.383139,9.715667,11.048194,12.380721,13.713249,13.724127,13.736817,13.749508,13.762199,13.77489,16.327541,18.880192,21.432844,23.985495,26.538147,25.85466,25.172985,24.489498,23.807825,23.124338,23.539507,23.954674,24.369843,24.785011,25.20018,25.466686,25.735004,26.003323,26.269827,26.538147,26.594349,26.652363,26.710379,26.768393,26.824594,26.52183,26.220879,25.918114,25.615349,25.312584,25.385101,25.45762,25.53014,25.602657,25.675177,25.582714,25.490253,25.397793,25.305332,25.212872,22.629398,20.04774,17.464268,14.882609,12.300951,15.147303,17.995466,20.841818,23.689981,26.538147,25.847408,25.158482,24.467743,23.777004,23.088078,23.0772,23.068136,23.057259,23.048193,23.037315,18.985344,14.9333725,10.879588,6.827617,2.7756457,3.24339,3.7093215,4.177066,4.64481,5.1125546,7.991539,10.872336,13.753134,16.632118,19.512917,19.494787,19.476658,19.46034,19.442211,19.425894,26.083092,32.74029,39.39749,46.054688,52.711887,44.45203,36.192173,27.932314,19.672457,11.4126,15.870674,20.326937,24.785011,29.243086,33.69935,33.829884,33.960415,34.09095,34.21967,34.3502,30.644506,26.940624,23.234928,19.529232,15.825351,15.620485,15.415621,15.210756,15.005891,14.799213,15.511708,16.224201,16.938509,17.651003,18.363499,14.920682,11.477866,8.03505,4.592234,1.1494182,1.9670644,2.7847104,3.6023567,4.420003,5.237649,5.0545397,4.8732433,4.690134,4.507025,4.325729,4.499773,4.6756306,4.8496747,5.0255322,5.199577,4.3003473,3.3993049,2.5000753,1.6008459,0.69980353,1.887294,3.0747845,4.262275,5.4497657,6.637256,6.604623,6.5719895,6.539356,6.506723,6.474089,5.669134,4.8641787,4.059223,3.254268,2.4493124,3.3231604,4.195195,5.06723,5.9392653,6.813113,6.0281005,5.243088,4.458075,3.673062,2.8880494,2.38042,1.8727903,1.3651608,0.8575313,0.34990177,0.4169814,0.48587397,0.5529536,0.6200332,0.6871128,0.7016165,0.7179332,0.7324369,0.7469406,0.76325727,0.72518504,0.6871128,0.6508536,0.61278135,0.5747091,1.0823387,1.5899682,2.0975976,2.6052272,3.1128569,2.7067533,2.3024626,1.8981718,1.4920682,1.0877775,1.0768998,1.067835,1.0569572,1.0478923,1.0370146,1.0243238,1.0116332,1.0007553,0.9880646,0.97537386,0.9880646,1.0007553,1.0116332,1.0243238,1.0370146,1.0333886,1.0279498,1.0225109,1.017072,1.0116332,1.0025684,0.9916905,0.9826257,0.97174793,0.96268314,1.3071461,1.651609,1.9978848,2.3423476,2.6868105,2.2716422,1.8582866,1.4431182,1.0279498,0.61278135,1.7096237,2.808279,3.9051213,5.0019636,6.1006193,5.147001,4.195195,3.2415771,2.2897718,1.3379664,1.455809,1.5718386,1.6896812,1.8075237,1.9253663,1.5446441,1.1657349,0.7850128,0.40429065,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.034446288,0.032633327,0.030820364,0.027194439,0.025381476,0.11965553,0.21574254,0.3100166,0.40429065,0.50037766,0.50037766,0.50037766,0.50037766,0.50037766,0.50037766,0.40066472,0.2991388,0.19942589,0.099712946,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.058014803,0.07795739,0.09789998,0.11784257,0.13778515,0.19942589,0.26287958,0.3245203,0.387974,0.44961473,0.4224203,0.39522585,0.3680314,0.34083697,0.31182957,0.28826106,0.26287958,0.2374981,0.21211663,0.18673515,0.21936847,0.2520018,0.28463513,0.31726846,0.34990177,0.27919623,0.21030366,0.13959812,0.07070554,0.0,0.052575916,0.10515183,0.15772775,0.21030366,0.26287958,0.34264994,0.4224203,0.50219065,0.581961,0.66173136,0.65991837,0.65810543,0.6544795,0.6526665,0.6508536,0.52575916,0.40066472,0.2755703,0.15047589,0.025381476,0.045324065,0.065266654,0.08520924,0.10515183,0.12509441,0.14322405,0.15954071,0.17767033,0.19579996,0.21211663,0.32270733,0.43329805,0.5420758,0.6526665,0.76325727,0.69436467,0.62728506,0.56020546,0.49312583,0.42423326,0.4550536,0.48587397,0.5148814,0.54570174,0.5747091,0.6091554,0.64541465,0.67986095,0.71430725,0.7505665,0.7868258,0.824898,0.8629702,0.89922947,0.93730164,1.1602961,1.3832904,1.6044719,1.8274662,2.0504606,2.0649643,2.079468,2.0957847,2.1102884,2.124792,2.1628644,2.1991236,2.2371957,2.275268,2.3133402,2.2625773,2.2118144,2.1628644,2.1121013,2.0631514,1.6806163,1.2980812,0.9155461,0.533011,0.15047589,0.13959812,0.13053331,0.11965553,0.11059072,0.099712946,0.26287958,0.42423326,0.5873999,0.7505665,0.9119202,0.83940166,0.7668832,0.69436467,0.62184614,0.5493277,0.5275721,0.5058166,0.48224804,0.4604925,0.43692398,0.4949388,0.5529536,0.6091554,0.6671702,0.72518504,0.6979906,0.67079616,0.6417888,0.61459434,0.5873999,0.52213323,0.45686656,0.39159992,0.32814622,0.26287958,0.24474995,0.22662032,0.21030366,0.19217403,0.17585737,0.14503701,0.11421664,0.08520924,0.054388877,0.025381476,0.11240368,0.19942589,0.28826106,0.37528324,0.46230546,1.261822,2.0631514,2.8626678,3.6621845,4.461701,6.452334,8.442966,10.431787,12.42242,14.413053,12.050762,9.686659,7.324369,4.9620786,2.5997884,2.1592383,1.7205015,1.2799516,0.83940166,0.40066472,1.5373923,1.4177368,1.2980812,1.1766127,1.0569572,0.93730164,0.8466535,0.75781834,0.6671702,0.57833505,0.48768693,0.51306844,0.53663695,0.5620184,0.5873999,0.61278135,0.8103943,1.0080072,1.2056202,1.403233,1.6008459,1.6280404,1.6552348,1.6824293,1.7096237,1.7368182,2.3369088,2.9369993,3.53709,4.137181,4.7372713,5.730775,6.722465,7.7141557,8.70766,9.699349,10.045626,10.390089,10.734551,11.080828,11.42529,11.390844,11.354585,11.320138,11.285692,11.249433,13.345218,15.439189,17.534973,19.630758,21.724731,22.199726,22.674723,23.14972,23.624716,24.099712,24.659918,25.220123,25.780329,26.340534,26.898926,24.688925,22.480736,20.26892,18.05892,15.848919,14.744824,13.640731,12.534823,11.430729,10.324821,13.687867,17.0491,20.412146,23.77519,27.138237,25.075085,23.011934,20.950596,18.887444,16.824293,15.4500675,14.075842,12.699803,11.325577,9.949538,8.049554,6.149569,4.249584,2.3495996,0.44961473,0.8883517,1.3252757,1.7621996,2.1991236,2.6378605,2.1646774,1.693307,1.2201238,0.7469406,0.2755703,0.2755703,0.2755703,0.2755703,0.2755703,0.2755703,0.37165734,0.46955732,0.56745726,0.6653573,0.76325727,1.1331016,1.502946,1.8727903,2.2426348,2.612479,2.1392958,1.6679256,1.1947423,0.72337204,0.25018883,0.28826106,0.3245203,0.36259252,0.40066472,0.43692398,0.44961473,0.46230546,0.4749962,0.48768693,0.50037766,2.514579,4.5305934,6.544795,8.560809,10.57501,10.234174,9.89515,9.554313,9.215289,8.874452,7.757667,6.640882,5.522284,4.405499,3.2869012,2.70494,2.1229792,1.5392052,0.9572442,0.37528324,1.4920682,2.610666,3.727451,4.844236,5.962834,7.509291,9.057561,10.605831,12.152288,13.700559,13.887294,14.075842,14.262577,14.449312,14.63786,16.99471,19.351562,21.710226,24.067078,26.425743,26.24082,26.055899,25.869164,25.68424,25.49932,25.657047,25.814774,25.972502,26.13023,26.287958,26.327843,26.367727,26.407614,26.447498,26.487383,26.772018,27.056654,27.343102,27.627737,27.912373,27.37936,26.848164,26.315151,25.78214,25.24913,26.929747,28.610363,30.29098,31.969782,33.6504,32.660522,31.670643,30.680765,29.690887,28.699198,26.064962,23.430729,20.794682,18.160446,15.524399,18.542982,21.559752,24.578333,27.595104,30.611874,30.430576,30.247467,30.064358,29.883062,29.699953,29.582111,29.464268,29.348238,29.230396,29.112553,23.82958,18.54842,13.265448,7.9824743,2.6995013,3.3648586,4.0302157,4.695573,5.3591175,6.0244746,7.0524244,8.080374,9.108324,10.13446,11.162411,13.497506,15.8326025,18.167698,20.502794,22.837889,30.35987,37.881855,45.405647,52.92763,60.44961,50.244446,40.041092,29.834112,19.628946,9.425592,14.897114,20.370447,25.841969,31.315302,36.786823,37.65342,38.518204,39.382988,40.24777,41.112553,35.822327,30.532103,25.241879,19.951653,14.663241,15.234324,15.80722,16.380117,16.953012,17.52591,18.537542,19.549175,20.562622,21.574255,22.5877,18.3218,14.057712,9.791811,5.527723,1.261822,1.9906329,2.7176309,3.444629,4.171627,4.900438,4.764466,4.6303062,4.494334,4.360175,4.2242026,4.699199,5.1741953,5.6491914,6.1241875,6.599184,5.424384,4.249584,3.0747845,1.8999848,0.72518504,2.324218,3.925064,5.52591,7.124943,8.725789,8.027799,7.3298078,6.6318173,5.9356394,5.237649,4.4345064,3.633177,2.8300345,2.0268922,1.2255627,2.7919624,4.360175,5.9283876,7.494787,9.063,7.844689,6.628191,5.40988,4.1933823,2.9750717,2.4529383,1.9308052,1.4068589,0.88472575,0.36259252,0.41516843,0.46774435,0.52032024,0.5728962,0.62547207,0.68167394,0.73968875,0.79770356,0.8557183,0.9119202,0.8375887,0.76325727,0.6871128,0.61278135,0.53663695,0.872035,1.2074331,1.5428312,1.8782293,2.2118144,2.0232663,1.8329052,1.6425442,1.452183,1.261822,1.2328146,1.2019942,1.1729867,1.1421664,1.1131591,1.1131591,1.1131591,1.1131591,1.1131591,1.1131591,1.1258497,1.1367276,1.1494182,1.162109,1.1747998,1.1349145,1.0950294,1.0551442,1.015259,0.97537386,0.91917205,0.86478317,0.8103943,0.7541924,0.69980353,1.0732739,1.4449311,1.8184015,2.1900587,2.561716,2.179181,1.7966459,1.4141108,1.0333886,0.6508536,1.3180238,1.9851941,2.6523643,3.3195345,3.9867048,3.442816,2.8971143,2.3532255,1.8075237,1.261822,1.2019942,1.1421664,1.0823387,1.0225109,0.96268314,0.77232206,0.581961,0.39159992,0.2030518,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.04169814,0.034446288,0.027194439,0.01994259,0.012690738,0.11059072,0.20667773,0.3045777,0.40247768,0.50037766,0.52575916,0.5493277,0.5747091,0.6000906,0.62547207,0.50037766,0.37528324,0.25018883,0.12509441,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.072518505,0.09427405,0.11784257,0.13959812,0.16316663,0.22480737,0.28826106,0.34990177,0.41335547,0.4749962,0.42967212,0.38434806,0.34083697,0.2955129,0.25018883,0.2374981,0.22480737,0.21211663,0.19942589,0.18673515,0.2229944,0.2574407,0.291887,0.32814622,0.36259252,0.29007402,0.21755551,0.14503701,0.072518505,0.0,0.032633327,0.065266654,0.09789998,0.13053331,0.16316663,0.27738327,0.39159992,0.5076295,0.62184614,0.73787576,0.7306239,0.72337204,0.71430725,0.7070554,0.69980353,0.5620184,0.42423326,0.28826106,0.15047589,0.012690738,0.034446288,0.058014803,0.07977036,0.10333887,0.12509441,0.12690738,0.13053331,0.13234627,0.13415924,0.13778515,0.27919623,0.4224203,0.5656443,0.7070554,0.85027945,0.75963134,0.67079616,0.58014804,0.4894999,0.40066472,0.42785916,0.4550536,0.48224804,0.5094425,0.53663695,0.5420758,0.5475147,0.5529536,0.55839247,0.5620184,0.5620184,0.5620184,0.5620184,0.5620184,0.5620184,0.80495536,1.0478923,1.2908293,1.5319533,1.7748904,1.794833,1.8147756,1.8347181,1.8546607,1.8746033,1.887294,1.8999848,1.9126755,1.9253663,1.938057,1.987007,2.03777,2.08672,2.137483,2.1882458,1.7767034,1.3669738,0.9572442,0.5475147,0.13778515,0.13234627,0.12690738,0.12328146,0.11784257,0.11240368,0.18673515,0.26287958,0.33721104,0.41335547,0.48768693,0.46955732,0.45324063,0.43511102,0.4169814,0.40066472,0.40791658,0.41516843,0.4224203,0.42967212,0.43692398,0.52213323,0.6073425,0.69255173,0.7777609,0.8629702,0.83033687,0.79770356,0.7650702,0.7324369,0.69980353,0.59283876,0.48587397,0.3770962,0.27013144,0.16316663,0.14684997,0.13234627,0.11784257,0.10333887,0.0870222,0.072518505,0.058014803,0.04169814,0.027194439,0.012690738,0.06164073,0.11240368,0.16316663,0.21211663,0.26287958,1.3379664,2.4130533,3.48814,4.5632267,5.638314,8.171022,10.703732,13.234627,15.767336,18.300045,14.96238,11.624716,8.287052,4.949388,1.6117238,1.3542831,1.0968424,0.83940166,0.581961,0.3245203,0.5620184,0.6744221,0.7868258,0.89922947,1.0116332,1.1258497,0.97537386,0.824898,0.6744221,0.52575916,0.37528324,0.43692398,0.50037766,0.5620184,0.62547207,0.6871128,0.9119202,1.1367276,1.3633479,1.5881553,1.8129625,1.8492218,1.887294,1.9253663,1.9616255,1.9996977,2.3133402,2.6251698,2.9369993,3.2506418,3.5624714,5.0128417,6.4632115,7.911769,9.362139,10.812509,10.850581,10.88684,10.924912,10.962985,10.999244,11.062697,11.124338,11.187792,11.249433,11.312886,13.562773,15.812659,18.062546,20.312433,22.562319,22.138086,21.71204,21.287807,20.861761,20.437527,18.611874,16.788034,14.96238,13.136727,11.312886,9.262425,7.211965,5.163317,3.1128569,1.062396,1.8492218,2.6378605,3.4246864,4.213325,5.0001507,8.80012,12.60009,16.400059,20.20003,23.999998,22.812508,21.625017,20.437527,19.250036,18.062546,16.062849,14.06315,12.06164,10.061942,8.062244,6.5629244,5.0617914,3.5624714,2.0631514,0.5620184,1.1004683,1.6371052,2.175555,2.712192,3.2506418,2.6378605,2.0250793,1.4122978,0.7995165,0.18673515,0.19942589,0.21211663,0.22480737,0.2374981,0.25018883,0.387974,0.52575916,0.66173136,0.7995165,0.93730164,1.3996071,1.8619126,2.324218,2.7883365,3.2506418,2.6505513,2.0504606,1.4503701,0.85027945,0.25018883,0.2755703,0.2991388,0.3245203,0.34990177,0.37528324,0.42423326,0.4749962,0.52575916,0.5747091,0.62547207,3.100166,5.57486,8.049554,10.524248,13.000754,12.28826,11.575767,10.863272,10.150778,9.438283,8.024173,6.6118746,5.199577,3.787279,2.374981,1.8999848,1.4249886,0.9499924,0.4749962,0.0,0.97537386,1.9507477,2.9243085,3.8996825,4.8750563,6.637256,8.399456,10.161655,11.925668,13.687867,14.05046,14.413053,14.775645,15.138238,15.50083,17.661882,19.824745,21.98761,24.150475,26.31334,26.625168,26.936998,27.25064,27.56247,27.8743,27.774588,27.674873,27.575161,27.475449,27.375734,27.187187,27.000452,26.811903,26.625168,26.43662,26.949688,27.462757,27.975826,28.487082,29.000149,28.236893,27.475449,26.71219,25.950747,25.187489,28.47439,31.763105,35.050007,38.336906,41.62562,39.738327,37.84922,35.961926,34.07463,32.187336,29.500526,26.811903,24.125093,21.438282,18.749659,21.936848,25.124035,28.313036,31.500225,34.687412,35.011932,35.33827,35.66279,35.98731,36.31183,36.08702,35.862213,35.637405,35.412598,35.18779,28.675629,22.163467,15.649493,9.137331,2.6251698,3.48814,4.349297,5.2122674,6.0752378,6.9382076,6.11331,5.2884116,4.461701,3.636803,2.811905,7.500226,12.186734,16.875055,21.563377,26.249886,34.63665,43.025227,51.41199,59.80057,68.18733,56.03686,43.8882,31.737722,19.587248,7.4367723,13.925365,20.412146,26.90074,33.38752,39.8743,41.475143,43.074177,44.675022,46.27587,47.874905,41.00015,34.125393,27.25064,20.374073,13.499319,14.849977,16.200634,17.549479,18.900135,20.250792,21.563377,22.87415,24.186733,25.49932,26.811903,21.724731,16.637558,11.5503845,6.4632115,1.3742256,2.0123885,2.6505513,3.2869012,3.925064,4.5632267,4.4743915,4.3873696,4.3003473,4.213325,4.12449,4.900438,5.674573,6.450521,7.224656,8.000604,6.550234,5.0998635,3.6494937,2.1991236,0.7505665,2.762955,4.7753434,6.787732,8.80012,10.812509,9.449161,8.087626,6.7242785,5.3627434,3.9993954,3.199879,2.4003625,1.6008459,0.7995165,0.0,2.2625773,4.5251546,6.787732,9.050309,11.312886,9.663091,8.013294,6.3616858,4.7118897,3.0620937,2.525457,1.987007,1.4503701,0.9119202,0.37528324,0.41335547,0.44961473,0.48768693,0.52575916,0.5620184,0.66173136,0.76325727,0.8629702,0.96268314,1.062396,0.9499924,0.8375887,0.72518504,0.61278135,0.50037766,0.66173136,0.824898,0.9880646,1.1494182,1.3125849,1.3379664,1.3633479,1.3869164,1.4122978,1.4376793,1.3869164,1.3379664,1.2872034,1.2382535,1.1874905,1.2001812,1.2128719,1.2255627,1.2382535,1.2491312,1.261822,1.2745126,1.2872034,1.2998942,1.3125849,1.2382535,1.162109,1.0877775,1.0116332,0.93730164,0.8375887,0.73787576,0.63816285,0.53663695,0.43692398,0.8375887,1.2382535,1.6371052,2.03777,2.4366217,2.08672,1.7368182,1.3869164,1.0370146,0.6871128,0.9246109,1.162109,1.3996071,1.6371052,1.8746033,1.7368182,1.6008459,1.4630609,1.3252757,1.1874905,0.9499924,0.7124943,0.4749962,0.2374981,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.099712946,0.19942589,0.2991388,0.40066472,0.50037766,0.5493277,0.6000906,0.6508536,0.69980353,0.7505665,0.6000906,0.44961473,0.2991388,0.15047589,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.0870222,0.11240368,0.13778515,0.16316663,0.18673515,0.25018883,0.31182957,0.37528324,0.43692398,0.50037766,0.43692398,0.37528324,0.31182957,0.25018883,0.18673515,0.18673515,0.18673515,0.18673515,0.18673515,0.18673515,0.22480737,0.26287958,0.2991388,0.33721104,0.37528324,0.2991388,0.22480737,0.15047589,0.07433146,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.21211663,0.36259252,0.51306844,0.66173136,0.8122072,0.7995165,0.7868258,0.774135,0.76325727,0.7505665,0.6000906,0.44961473,0.2991388,0.15047589,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.2374981,0.41335547,0.5873999,0.76325727,0.93730164,0.824898,0.7124943,0.6000906,0.48768693,0.37528324,0.40066472,0.42423326,0.44961473,0.4749962,0.50037766,0.4749962,0.44961473,0.42423326,0.40066472,0.37528324,0.33721104,0.2991388,0.26287958,0.22480737,0.18673515,0.44961473,0.7124943,0.97537386,1.2382535,1.49932,1.5247015,1.550083,1.5754645,1.6008459,1.6244144,1.6117238,1.6008459,1.5881553,1.5754645,1.5627737,1.7132497,1.8619126,2.0123885,2.1628644,2.3133402,1.8746033,1.4376793,1.0007553,0.5620184,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.099712946,0.13778515,0.17585737,0.21211663,0.25018883,0.28826106,0.3245203,0.36259252,0.40066472,0.43692398,0.5493277,0.66173136,0.774135,0.8883517,1.0007553,0.96268314,0.9246109,0.8883517,0.85027945,0.8122072,0.66173136,0.51306844,0.36259252,0.21211663,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,1.4122978,2.762955,4.1117992,5.462456,6.813113,9.8878975,12.962683,16.037468,19.112251,22.187037,17.873999,13.562773,9.249735,4.93851,0.62547207,0.5493277,0.4749962,0.40066472,0.3245203,0.25018883,0.61278135,0.7016165,0.79226464,0.88291276,0.97174793,1.062396,0.969935,0.8774739,0.7850128,0.69255173,0.6000906,0.7197462,0.83940166,0.96087015,1.0805258,1.2001812,1.3669738,1.5355793,1.7023718,1.8691645,2.03777,2.0033236,1.9670644,1.9326181,1.8981718,1.8619126,2.0903459,2.3169663,2.5453994,2.7720199,3.000453,4.3347936,5.669134,7.0052876,8.339628,9.675781,10.022058,10.370146,10.718235,11.06451,11.4126,11.844085,12.277383,12.710681,13.142166,13.575464,14.824595,16.075539,17.32467,18.575615,19.824745,19.665205,19.505665,19.34431,19.18477,19.025229,17.26303,15.50083,13.736817,11.974618,10.212419,8.415772,6.6173134,4.8206677,3.0222087,1.2255627,1.9471219,2.6704938,3.392053,4.115425,4.836984,8.319685,11.802386,15.285088,18.767788,22.25049,21.197159,20.14564,19.092308,18.04079,16.98746,14.989574,12.99169,10.995618,8.997733,6.9998484,5.922949,4.844236,3.7673361,2.6904364,1.6117238,1.9598125,2.3079014,2.6541772,3.002266,3.350355,2.762955,2.175555,1.5881553,1.0007553,0.41335547,0.6055295,0.79770356,0.9898776,1.1820517,1.3742256,2.1556125,2.9351864,3.7147603,4.494334,5.275721,5.4570174,5.6401267,5.823236,6.004532,6.187641,4.989273,3.7927177,2.5943494,1.3977941,0.19942589,0.26469254,0.32995918,0.39522585,0.4604925,0.52575916,0.83033687,1.1349145,1.4394923,1.745883,2.0504606,4.360175,6.6698895,8.979604,11.289318,13.600845,12.685299,11.769753,10.854207,9.940474,9.024928,7.605378,6.185828,4.764466,3.3449159,1.9253663,1.5428312,1.1602961,0.7777609,0.39522585,0.012690738,0.83577573,1.6570477,2.4801328,3.303218,4.12449,5.569421,7.0143523,8.459284,9.904215,11.349146,11.635593,11.920229,12.2048645,12.489499,12.775948,14.626982,16.47983,18.332678,20.185526,22.038374,22.239613,22.442663,22.645716,22.846954,23.050007,23.644657,24.23931,24.835773,25.430426,26.025078,27.062092,28.099108,29.137934,30.17495,31.211964,32.568058,33.922344,35.276627,36.63272,37.987003,36.645412,35.302006,33.960415,32.61701,31.275417,33.313187,35.349144,37.386913,39.424683,41.462456,40.3076,39.15274,37.997883,36.843025,35.688168,33.059372,30.43239,27.805407,25.17661,22.54963,24.63816,26.724882,28.813414,30.900135,32.986855,32.95966,32.932465,32.90527,32.878075,32.850883,34.243237,35.635593,37.027946,38.420303,39.812656,33.771866,27.73289,21.692097,15.653119,9.612328,10.435412,11.256684,12.07977,12.902855,13.724127,12.284635,10.845142,9.40565,7.9643445,6.5248523,10.346578,14.170115,17.99184,21.815378,25.637104,32.622448,39.60779,46.59314,53.578484,60.562016,49.680614,38.797398,27.914185,17.032784,6.149569,12.154101,18.160446,24.164978,30.16951,36.175854,38.0704,39.964947,41.859493,43.75585,45.6504,39.19081,32.729412,26.269827,19.810242,13.3506565,14.811904,16.274965,17.738026,19.199274,20.662334,21.655838,22.647528,23.63922,24.632723,25.624413,21.095633,16.565039,12.034446,7.5056653,2.9750717,3.1273603,3.2796493,3.4319382,3.584227,3.738329,3.825351,3.9123733,3.9993954,4.0882306,4.175253,5.224958,6.2746634,7.324369,8.375887,9.425592,8.127511,6.82943,5.5331616,4.2350807,2.9369993,4.256836,5.576673,6.8983226,8.21816,9.537996,8.406708,7.2772317,6.147756,5.0182805,3.8869917,3.1182957,2.3477864,1.5772774,0.80676836,0.038072214,1.840157,3.6422417,5.4443264,7.2482243,9.050309,7.744976,6.439643,5.1343102,3.83079,2.525457,2.1175404,1.7096237,1.3017071,0.89560354,0.48768693,0.5855869,0.68167394,0.7795739,0.8774739,0.97537386,0.9572442,0.93911463,0.922798,0.90466833,0.8883517,0.8103943,0.7324369,0.6544795,0.57833505,0.50037766,0.65810543,0.81583315,0.97174793,1.1294757,1.2872034,1.2908293,1.2926424,1.2944553,1.2980812,1.2998942,1.2726997,1.2455053,1.2183108,1.1893034,1.162109,1.1747998,1.1874905,1.2001812,1.2128719,1.2255627,1.2183108,1.209246,1.2019942,1.1947423,1.1874905,1.1131591,1.0370146,0.96268314,0.8883517,0.8122072,0.7197462,0.62728506,0.53482395,0.44236287,0.34990177,0.68167394,1.015259,1.3470312,1.6806163,2.0123885,1.7350051,1.4576219,1.1802386,0.90285534,0.62547207,0.7995165,0.97537386,1.1494182,1.3252757,1.49932,1.3996071,1.2998942,1.2001812,1.1004683,1.0007553,0.7995165,0.6000906,0.40066472,0.19942589,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.065266654,0.13053331,0.19579996,0.25925365,0.3245203,0.25925365,0.19579996,0.13053331,0.065266654,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.07977036,0.15954071,0.23931105,0.3208944,0.40066472,0.4405499,0.48043507,0.52032024,0.56020546,0.6000906,0.48043507,0.36077955,0.23931105,0.11965553,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.07795739,0.10515183,0.13234627,0.15954071,0.18673515,0.24837588,0.30820364,0.3680314,0.42785916,0.48768693,0.4405499,0.39159992,0.3444629,0.29732585,0.25018883,0.23205921,0.21574254,0.19761293,0.1794833,0.16316663,0.20667773,0.2520018,0.29732585,0.34264994,0.387974,0.31726846,0.24837588,0.17767033,0.10696479,0.038072214,0.03988518,0.04169814,0.045324065,0.047137026,0.05076295,0.18492219,0.3208944,0.4550536,0.58921283,0.72518504,0.726998,0.7306239,0.7324369,0.73424983,0.73787576,0.59283876,0.44780177,0.30276474,0.15772775,0.012690738,0.030820364,0.047137026,0.065266654,0.08339628,0.099712946,0.09427405,0.09064813,0.08520924,0.07977036,0.07433146,0.21211663,0.34990177,0.48768693,0.62547207,0.76325727,0.6871128,0.61278135,0.53663695,0.46230546,0.387974,0.40791658,0.42785916,0.44780177,0.46774435,0.48768693,0.47680917,0.46774435,0.45686656,0.44780177,0.43692398,0.38978696,0.34264994,0.2955129,0.24837588,0.19942589,0.40247768,0.6055295,0.80676836,1.0098201,1.2128719,1.2382535,1.261822,1.2872034,1.3125849,1.3379664,1.3506571,1.3633479,1.3742256,1.3869164,1.3996071,1.5718386,1.745883,1.9181144,2.0903459,2.2625773,1.845596,1.4268016,1.0098201,0.59283876,0.17585737,0.17223145,0.17041849,0.16679256,0.16497959,0.16316663,0.15954071,0.15772775,0.15410182,0.15228885,0.15047589,0.17041849,0.19036107,0.21030366,0.23024625,0.25018883,0.3245203,0.40066472,0.4749962,0.5493277,0.62547207,0.7850128,0.9445535,1.1040943,1.2654479,1.4249886,1.2745126,1.1258497,0.97537386,0.824898,0.6744221,0.5493277,0.42423326,0.2991388,0.17585737,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.02175555,0.032633327,0.04169814,0.052575916,0.06164073,1.4703126,2.8771715,4.2858434,5.6927023,7.0995617,9.336758,11.575767,13.812962,16.050158,18.287354,14.762955,11.236742,7.7123427,4.1879435,0.66173136,0.6055295,0.5475147,0.4894999,0.43329805,0.37528324,0.66173136,0.7306239,0.79770356,0.86478317,0.9318628,1.0007553,0.9644961,0.9300498,0.89560354,0.85934424,0.824898,1.0025684,1.1802386,1.357909,1.5355793,1.7132497,1.8220274,1.9326181,2.0432088,2.1519866,2.2625773,2.1556125,2.0468347,1.93987,1.8329052,1.7241274,1.8673514,2.0105755,2.1519866,2.2952106,2.4366217,3.6567454,4.876869,6.096993,7.317117,8.537241,9.195346,9.851639,10.509744,11.16785,11.8241415,12.627284,13.430427,14.231756,15.034899,15.838041,16.08823,16.336605,16.586794,16.836983,17.087172,17.192324,17.297476,17.402628,17.50778,17.612932,15.912373,14.211814,12.513068,10.812509,9.11195,7.567306,6.0226617,4.478018,2.9333735,1.3869164,2.0450218,2.7031271,3.3594196,4.017525,4.6756306,7.83925,11.004683,14.170115,17.335548,20.499168,19.581808,18.66445,17.747091,16.829731,15.912373,13.918114,11.922042,9.927783,7.931711,5.9374523,5.282973,4.6266804,3.972201,3.3177216,2.663242,2.819157,2.9768846,3.1346123,3.29234,3.4500678,2.8880494,2.324218,1.7621996,1.2001812,0.63816285,1.0098201,1.3832904,1.7549478,2.128418,2.5000753,3.923251,5.3446136,6.7677894,8.189152,9.612328,9.514427,9.418341,9.32044,9.222541,9.12464,7.3298078,5.5349746,3.7401419,1.9453088,0.15047589,0.25562772,0.36077955,0.46411842,0.56927025,0.6744221,1.2346275,1.794833,2.3550384,2.9152439,3.4754493,5.620184,7.764919,9.909654,12.054388,14.199123,13.082338,11.965553,10.846955,9.73017,8.613385,7.1847706,5.7579694,4.329355,2.902553,1.4757515,1.1856775,0.89560354,0.6055295,0.3154555,0.025381476,0.69436467,1.3651608,2.034144,2.70494,3.3757362,4.501586,5.6292486,6.7569118,7.8845744,9.012237,9.220728,9.427405,9.634083,9.842574,10.049252,11.592083,13.134913,14.677745,16.220575,17.761595,17.85587,17.94833,18.04079,18.133251,18.225714,19.514729,20.80556,22.094576,23.385405,24.674421,26.936998,29.199575,31.462152,33.72473,35.98731,38.184616,40.381927,42.57924,44.778362,46.975674,45.05212,43.13038,41.206825,39.285088,37.363346,38.150173,38.936996,39.725636,40.512463,41.299286,40.87687,40.45445,40.03203,39.609608,39.187187,36.62003,34.052876,31.485722,28.916754,26.349598,27.337664,28.325727,29.31198,30.300043,31.288109,30.907387,30.526665,30.147755,29.767033,29.388123,32.39764,35.407158,38.41849,41.42801,44.437527,38.86992,33.30231,27.734701,22.167093,16.599485,17.382685,18.165886,18.947271,19.730473,20.511858,18.457771,16.401873,14.347786,12.291886,10.2378,13.194741,16.151684,19.11044,22.06738,25.024323,30.608248,36.190357,41.772472,47.354584,52.936695,43.322556,33.708412,24.09246,14.476506,4.8623657,10.384649,15.906934,21.43103,26.953314,32.475597,34.665657,36.855717,39.045776,41.235832,43.42408,37.37966,31.335245,25.289015,19.244598,13.200181,14.775645,16.349297,17.92476,19.500225,21.07569,21.748299,22.419096,23.091705,23.764313,24.436922,20.464722,16.492521,12.52032,8.548119,4.5759177,4.2423325,3.9105604,3.576975,3.245203,2.911618,3.1744974,3.437377,3.7002566,3.9631362,4.2242026,5.5494785,6.874754,8.200029,9.525306,10.850581,9.704789,8.560809,7.415017,6.2692246,5.125245,5.75253,6.379815,7.0071006,7.6343856,8.26167,7.364254,6.4668374,5.569421,4.6720047,3.774588,3.0348995,2.2952106,1.5555218,0.81583315,0.07433146,1.4177368,2.759329,4.102734,5.4443264,6.787732,5.826862,4.8678045,3.9069343,2.9478772,1.987007,1.7096237,1.4322405,1.1548572,0.8774739,0.6000906,0.75781834,0.9155461,1.0732739,1.2291887,1.3869164,1.2527572,1.1167849,0.9826257,0.8466535,0.7124943,0.67079616,0.62728506,0.5855869,0.5420758,0.50037766,0.6526665,0.80495536,0.9572442,1.1095331,1.261822,1.2418793,1.2219368,1.2019942,1.1820517,1.162109,1.1566701,1.1530442,1.1476053,1.1421664,1.1367276,1.1494182,1.162109,1.1747998,1.1874905,1.2001812,1.1729867,1.1457924,1.1167849,1.0895905,1.062396,0.9880646,0.9119202,0.8375887,0.76325727,0.6871128,0.60190356,0.5166943,0.43329805,0.3480888,0.26287958,0.5275721,0.79226464,1.0569572,1.3216497,1.5881553,1.3832904,1.1766127,0.97174793,0.7668832,0.5620184,0.6744221,0.7868258,0.89922947,1.0116332,1.1258497,1.062396,1.0007553,0.93730164,0.87566096,0.8122072,0.6508536,0.48768693,0.3245203,0.16316663,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.10515183,0.21030366,0.3154555,0.42060733,0.52575916,0.42060733,0.3154555,0.21030366,0.10515183,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.059827764,0.11965553,0.1794833,0.23931105,0.2991388,0.32995918,0.36077955,0.38978696,0.42060733,0.44961473,0.36077955,0.27013144,0.1794833,0.09064813,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.06707962,0.09789998,0.12690738,0.15772775,0.18673515,0.24474995,0.30276474,0.36077955,0.4169814,0.4749962,0.44236287,0.40972954,0.3770962,0.3444629,0.31182957,0.27738327,0.24293698,0.20667773,0.17223145,0.13778515,0.19036107,0.24293698,0.2955129,0.3480888,0.40066472,0.33539808,0.27013144,0.20486477,0.13959812,0.07433146,0.06707962,0.059827764,0.052575916,0.045324065,0.038072214,0.15772775,0.27738327,0.39703882,0.5166943,0.63816285,0.6544795,0.6726091,0.69073874,0.7070554,0.72518504,0.5855869,0.44417584,0.3045777,0.16497959,0.025381476,0.034446288,0.045324065,0.054388877,0.065266654,0.07433146,0.07795739,0.07977036,0.08339628,0.08520924,0.0870222,0.18673515,0.28826106,0.387974,0.48768693,0.5873999,0.5493277,0.51306844,0.4749962,0.43692398,0.40066472,0.41516843,0.42967212,0.44417584,0.4604925,0.4749962,0.48043507,0.48587397,0.4894999,0.4949388,0.50037766,0.44236287,0.38434806,0.32814622,0.27013144,0.21211663,0.35534066,0.49675176,0.6399758,0.78319985,0.9246109,0.9499924,0.97537386,1.0007553,1.0243238,1.0497054,1.0877775,1.1258497,1.162109,1.2001812,1.2382535,1.4322405,1.6280404,1.8220274,2.0178273,2.2118144,1.8147756,1.4177368,1.020698,0.62184614,0.22480737,0.21936847,0.21574254,0.21030366,0.20486477,0.19942589,0.20667773,0.21574254,0.2229944,0.23024625,0.2374981,0.23931105,0.24293698,0.24474995,0.24837588,0.25018883,0.36259252,0.4749962,0.5873999,0.69980353,0.8122072,1.020698,1.2273756,1.4358664,1.6425442,1.8492218,1.5881553,1.3252757,1.062396,0.7995165,0.53663695,0.43692398,0.33721104,0.2374981,0.13778515,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.032633327,0.03988518,0.047137026,0.054388877,0.06164073,1.5283275,2.9932013,4.458075,5.922949,7.3878226,8.78743,10.1870365,11.586644,12.988064,14.387671,11.650098,8.912524,6.1749506,3.437377,0.69980353,0.65991837,0.6200332,0.58014804,0.5402629,0.50037766,0.7124943,0.75781834,0.8031424,0.8466535,0.8919776,0.93730164,0.96087015,0.9826257,1.0043813,1.0279498,1.0497054,1.2853905,1.5192627,1.7549478,1.9906329,2.2245052,2.277081,2.3296568,2.382233,2.4348087,2.4873846,2.3079014,2.126605,1.9471219,1.7676386,1.5881553,1.6443571,1.7023718,1.7603867,1.8165885,1.8746033,2.9805105,4.0846047,5.1905117,6.294606,7.400513,8.366822,9.334945,10.303066,11.269376,12.237497,13.410484,14.581658,15.754644,16.927631,18.100618,17.350052,16.599485,15.850732,15.100165,14.349599,14.719443,15.089288,15.459132,15.83079,16.200634,14.561715,12.92461,11.287505,9.6504,8.013294,6.720652,5.42801,4.135368,2.8427253,1.550083,2.1429217,2.7357605,3.3267863,3.919625,4.512464,7.360628,10.20698,13.055143,15.903308,18.749659,17.968271,17.185072,16.401873,15.620485,14.837286,12.84484,10.852394,8.859948,6.867502,4.8750563,4.6429973,4.409125,4.177066,3.9450066,3.7129474,3.680314,3.6476808,3.6150475,3.5824142,3.5497808,3.0131438,2.474694,1.938057,1.3996071,0.8629702,1.4141108,1.9670644,2.520018,3.0729716,3.625925,5.6908894,7.755854,9.820818,11.885782,13.9507475,13.571837,13.194741,12.817645,12.440549,12.063453,9.670342,7.2772317,4.8841214,2.4928236,0.099712946,0.24474995,0.38978696,0.53482395,0.67986095,0.824898,1.6407311,2.4547513,3.2705846,4.0846047,4.900438,6.880193,8.859948,10.839704,12.819458,14.799213,13.479377,12.15954,10.839704,9.519867,8.200029,6.7641635,5.33011,3.8942437,2.4601903,1.0243238,0.82671094,0.629098,0.43329805,0.23568514,0.038072214,0.55476654,1.0732739,1.5899682,2.1066625,2.6251698,3.435564,4.2441454,5.0545397,5.864934,6.6753283,6.8040485,6.9345818,7.065115,7.1956487,7.324369,8.557183,9.789998,11.022813,12.255627,13.486629,13.470312,13.452183,13.434052,13.417736,13.399607,15.384801,17.369995,19.355188,21.340382,23.325577,26.811903,30.300043,33.788185,37.27451,40.76265,43.80299,46.843327,49.883667,52.92219,55.96253,53.46064,50.95694,48.45505,45.953163,43.449463,42.987156,42.52485,42.062546,41.60024,41.137936,41.447952,41.75797,42.067986,42.378002,42.68802,40.18069,37.673363,35.164223,32.656895,30.149569,30.037165,29.92476,29.812357,29.699953,29.58755,28.855112,28.122675,27.390238,26.657803,25.925365,30.552046,35.18054,39.80722,44.435715,49.062393,43.967968,38.873543,33.777306,28.68288,23.588457,24.329958,25.073273,25.814774,26.558088,27.299591,24.630909,21.960415,19.289923,16.619429,13.9507475,16.042906,18.135065,20.227224,22.319382,24.413355,28.592234,32.772926,36.951805,41.132496,45.311375,36.964493,28.617615,20.26892,11.922042,3.5751622,8.615198,13.655234,18.69527,23.735306,28.775343,31.2591,33.74467,36.230244,38.715816,41.199574,35.570328,29.939264,24.310015,18.680767,13.049705,14.737573,16.425442,18.11331,19.799364,21.487232,21.84076,22.192474,22.54419,22.897717,23.249432,19.835623,16.420002,13.00438,9.590572,6.1749506,5.3573046,4.539658,3.7220123,2.904366,2.08672,2.525457,2.962381,3.3993049,3.8380418,4.274966,5.8758116,7.474845,9.07569,10.674724,12.27557,11.282066,10.290376,9.296872,8.3051815,7.311678,7.2482243,7.1829576,7.117691,7.0524244,6.987158,6.3218007,5.658256,4.992899,4.327542,3.6621845,2.953316,2.2426348,1.5319533,0.823085,0.11240368,0.99531645,1.8782293,2.759329,3.6422417,4.5251546,3.9105604,3.294153,2.6795588,2.0649643,1.4503701,1.3017071,1.1548572,1.0080072,0.85934424,0.7124943,0.9300498,1.1476053,1.3651608,1.5827163,1.8002719,1.54827,1.2944553,1.0424535,0.7904517,0.53663695,0.5293851,0.52213323,0.5148814,0.5076295,0.50037766,0.64722764,0.79589057,0.94274056,1.0895905,1.2382535,1.1947423,1.1530442,1.1095331,1.067835,1.0243238,1.0424535,1.0605831,1.0768998,1.0950294,1.1131591,1.1258497,1.1367276,1.1494182,1.162109,1.1747998,1.1276628,1.0805258,1.0333886,0.98443866,0.93730164,0.8629702,0.7868258,0.7124943,0.63816285,0.5620184,0.48587397,0.40791658,0.32995918,0.2520018,0.17585737,0.37165734,0.56927025,0.7668832,0.9644961,1.162109,1.0297627,0.8974165,0.7650702,0.6327239,0.50037766,0.5493277,0.6000906,0.6508536,0.69980353,0.7505665,0.72518504,0.69980353,0.6744221,0.6508536,0.62547207,0.50037766,0.37528324,0.25018883,0.12509441,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14503701,0.29007402,0.43511102,0.58014804,0.72518504,0.58014804,0.43511102,0.29007402,0.14503701,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.03988518,0.07977036,0.11965553,0.15954071,0.19942589,0.21936847,0.23931105,0.25925365,0.27919623,0.2991388,0.23931105,0.1794833,0.11965553,0.059827764,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.058014803,0.09064813,0.12328146,0.15410182,0.18673515,0.24293698,0.29732585,0.35171473,0.40791658,0.46230546,0.44417584,0.42785916,0.40972954,0.39159992,0.37528324,0.32270733,0.27013144,0.21755551,0.16497959,0.11240368,0.17223145,0.23205921,0.291887,0.35171473,0.41335547,0.35171473,0.291887,0.23205921,0.17223145,0.11240368,0.09427405,0.07795739,0.059827764,0.04169814,0.025381476,0.13053331,0.23568514,0.34083697,0.44417584,0.5493277,0.581961,0.61459434,0.64722764,0.67986095,0.7124943,0.57833505,0.44236287,0.30820364,0.17223145,0.038072214,0.03988518,0.04169814,0.045324065,0.047137026,0.05076295,0.059827764,0.07070554,0.07977036,0.09064813,0.099712946,0.16316663,0.22480737,0.28826106,0.34990177,0.41335547,0.41335547,0.41335547,0.41335547,0.41335547,0.41335547,0.4224203,0.43329805,0.44236287,0.45324063,0.46230546,0.48224804,0.50219065,0.52213323,0.5420758,0.5620184,0.4949388,0.42785916,0.36077955,0.291887,0.22480737,0.30820364,0.38978696,0.47318324,0.55476654,0.63816285,0.66173136,0.6871128,0.7124943,0.73787576,0.76325727,0.824898,0.8883517,0.9499924,1.0116332,1.0750868,1.2926424,1.5101979,1.7277533,1.9453088,2.1628644,1.7857682,1.4068589,1.0297627,0.6526665,0.2755703,0.26831847,0.25925365,0.2520018,0.24474995,0.2374981,0.25562772,0.27194437,0.29007402,0.30820364,0.3245203,0.3100166,0.2955129,0.27919623,0.26469254,0.25018883,0.40066472,0.5493277,0.69980353,0.85027945,1.0007553,1.2545701,1.5101979,1.7658255,2.0196402,2.275268,1.8999848,1.5247015,1.1494182,0.774135,0.40066472,0.3245203,0.25018883,0.17585737,0.099712946,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.04169814,0.047137026,0.052575916,0.058014803,0.06164073,1.5845293,3.1074178,4.6303062,6.153195,7.6742706,8.238102,8.80012,9.362139,9.924157,10.487988,8.537241,6.586493,4.6375585,2.6868105,0.73787576,0.71430725,0.69255173,0.67079616,0.64722764,0.62547207,0.76325727,0.7850128,0.80676836,0.83033687,0.8520924,0.87566096,0.9554313,1.0352017,1.114972,1.1947423,1.2745126,1.5682126,1.8600996,2.1519866,2.4456866,2.7375734,2.7321346,2.7266958,2.72307,2.7176309,2.712192,2.4601903,2.2081885,1.9543737,1.7023718,1.4503701,1.4231756,1.3941683,1.3669738,1.3397794,1.3125849,2.3024626,3.29234,4.2822175,5.272095,6.261973,7.5401115,8.81825,10.094576,11.372714,12.650853,14.191871,15.734702,17.277533,18.820364,20.363195,18.611874,16.862366,15.112856,13.363347,11.612025,12.246562,12.882912,13.517449,14.151986,14.788336,13.212872,11.637406,10.061942,8.488291,6.9128265,5.8721857,4.8333583,3.7927177,2.752077,1.7132497,2.2408218,2.7665808,3.294153,3.8217251,4.349297,6.880193,9.409276,11.940171,14.4692545,17.00015,16.352922,15.705695,15.056654,14.409427,13.762199,11.773379,9.782746,7.7921133,5.803293,3.8126602,4.0030212,4.1933823,4.3819304,4.572292,4.762653,4.539658,4.3166637,4.0954823,3.872488,3.6494937,3.1382382,2.6251698,2.1121013,1.6008459,1.0877775,1.8202144,2.5526514,3.2850883,4.017525,4.749962,7.456715,10.165281,12.872034,15.580601,18.287354,17.629248,16.972956,16.31485,15.656745,15.000452,12.010877,9.019489,6.0299134,3.0403383,0.05076295,0.23568514,0.42060733,0.6055295,0.7904517,0.97537386,2.0450218,3.1146698,4.1843176,5.2557783,6.3254266,8.140202,9.954978,11.769753,13.584529,15.399304,13.878228,12.35534,10.832452,9.309563,7.7866745,6.345369,4.902251,3.4591327,2.0178273,0.5747091,0.46955732,0.36440548,0.25925365,0.15410182,0.05076295,0.41516843,0.7795739,1.1457924,1.5101979,1.8746033,2.3677292,2.8608549,3.3521678,3.8452935,4.3366065,4.3891826,4.441758,4.494334,4.5469103,4.599486,5.522284,6.445082,7.36788,8.290678,9.211663,9.084756,8.957849,8.829127,8.70222,8.575313,11.254871,13.93443,16.615803,19.29536,21.97492,26.68681,31.400513,36.1124,40.82429,45.537994,49.419548,53.302914,57.184467,61.067833,64.94939,61.867348,58.785313,55.703274,52.619427,49.537388,47.825954,46.1127,44.399452,42.68802,40.974766,42.01722,43.059673,44.102127,45.14458,46.187035,43.739536,41.292034,38.844536,36.397038,33.94954,32.736664,31.525606,30.312735,29.099863,27.88699,26.80284,25.716875,24.632723,23.546759,22.462606,28.708263,34.952106,41.19776,47.443417,53.68726,49.06602,44.442966,39.819912,35.196857,30.575613,31.277231,31.98066,32.682278,33.385708,34.087322,30.802235,27.517145,24.232058,20.94697,17.661882,18.889257,20.116632,21.345821,22.573196,23.800573,26.578032,29.35549,32.13295,34.910408,37.687866,30.608248,23.526815,16.447197,9.367578,2.2879589,6.8457465,11.401722,15.95951,20.517298,25.075085,27.854357,30.63544,33.414715,36.195797,38.97507,33.759174,28.545095,23.329203,18.115122,12.899229,14.699501,16.499773,18.300045,20.100317,21.900587,21.933222,21.965855,21.996675,22.029308,22.061941,19.204712,16.347483,13.490254,10.633025,7.7757964,6.472276,5.1705694,3.8670492,2.565342,1.261822,1.8746033,2.4873846,3.100166,3.7129474,4.325729,6.200332,8.074935,9.949538,11.8241415,13.700559,12.859344,12.019942,11.18054,10.339326,9.499924,8.7421055,7.9842873,7.228282,6.4704633,5.712645,5.279347,4.847862,4.4145637,3.9830787,3.5497808,2.8699198,2.1900587,1.5101979,0.83033687,0.15047589,0.5728962,0.99531645,1.4177368,1.840157,2.2625773,1.9924458,1.7223145,1.452183,1.1820517,0.9119202,0.89560354,0.8774739,0.85934424,0.8430276,0.824898,1.1022812,1.3796645,1.6570477,1.9344311,2.2118144,1.84197,1.4721256,1.1022812,0.7324369,0.36259252,0.38978696,0.4169814,0.44417584,0.47318324,0.50037766,0.6417888,0.7850128,0.92823684,1.0696479,1.2128719,1.1476053,1.0823387,1.017072,0.95180535,0.8883517,0.92823684,0.968122,1.0080072,1.0478923,1.0877775,1.1004683,1.1131591,1.1258497,1.1367276,1.1494182,1.0823387,1.015259,0.9481794,0.8792868,0.8122072,0.73787576,0.66173136,0.5873999,0.51306844,0.43692398,0.3680314,0.29732585,0.22662032,0.15772775,0.0870222,0.21755551,0.3480888,0.47680917,0.6073425,0.73787576,0.678048,0.61822027,0.55839247,0.49675176,0.43692398,0.42423326,0.41335547,0.40066472,0.387974,0.37528324,0.387974,0.40066472,0.41335547,0.42423326,0.43692398,0.34990177,0.26287958,0.17585737,0.0870222,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.18492219,0.36984438,0.55476654,0.73968875,0.9246109,0.73968875,0.55476654,0.36984438,0.18492219,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.11059072,0.11965553,0.13053331,0.13959812,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.047137026,0.08339628,0.11784257,0.15228885,0.18673515,0.23931105,0.291887,0.3444629,0.39703882,0.44961473,0.44780177,0.44417584,0.44236287,0.4405499,0.43692398,0.3680314,0.29732585,0.22662032,0.15772775,0.0870222,0.15410182,0.2229944,0.29007402,0.35715362,0.42423326,0.36984438,0.3154555,0.25925365,0.20486477,0.15047589,0.12328146,0.09427405,0.06707962,0.03988518,0.012690738,0.10333887,0.19217403,0.28282216,0.37165734,0.46230546,0.5094425,0.55839247,0.6055295,0.6526665,0.69980353,0.56927025,0.4405499,0.3100166,0.1794833,0.05076295,0.045324065,0.03988518,0.034446288,0.030820364,0.025381476,0.04169814,0.059827764,0.07795739,0.09427405,0.11240368,0.13778515,0.16316663,0.18673515,0.21211663,0.2374981,0.2755703,0.31182957,0.34990177,0.387974,0.42423326,0.42967212,0.43511102,0.4405499,0.44417584,0.44961473,0.48587397,0.52032024,0.55476654,0.58921283,0.62547207,0.5475147,0.46955732,0.39159992,0.3154555,0.2374981,0.25925365,0.28282216,0.3045777,0.32814622,0.34990177,0.37528324,0.40066472,0.42423326,0.44961473,0.4749962,0.5620184,0.6508536,0.73787576,0.824898,0.9119202,1.1530442,1.3923552,1.6316663,1.8727903,2.1121013,1.7549478,1.3977941,1.0406405,0.68167394,0.3245203,0.3154555,0.3045777,0.2955129,0.28463513,0.2755703,0.30276474,0.32995918,0.35715362,0.38434806,0.41335547,0.38072214,0.3480888,0.3154555,0.28282216,0.25018883,0.43692398,0.62547207,0.8122072,1.0007553,1.1874905,1.4902552,1.79302,2.0957847,2.3967366,2.6995013,2.2118144,1.7241274,1.2382535,0.7505665,0.26287958,0.21211663,0.16316663,0.11240368,0.06164073,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.052575916,0.054388877,0.058014803,0.059827764,0.06164073,1.6425442,3.2234476,4.802538,6.3816285,7.9625316,7.686961,7.413204,7.137634,6.8620634,6.588306,5.424384,4.262275,3.100166,1.938057,0.774135,0.7705091,0.7650702,0.75963134,0.7541924,0.7505665,0.8122072,0.8122072,0.8122072,0.8122072,0.8122072,0.8122072,0.9499924,1.0877775,1.2255627,1.3633479,1.49932,1.8492218,2.1991236,2.5508385,2.9007401,3.2506418,3.1871881,3.1255474,3.0620937,3.000453,2.9369993,2.612479,2.2879589,1.9616255,1.6371052,1.3125849,1.2001812,1.0877775,0.97537386,0.8629702,0.7505665,1.6244144,2.5000753,3.3757362,4.249584,5.125245,6.7115874,8.299743,9.8878975,11.47424,13.062395,14.975071,16.887747,18.800423,20.713097,22.625772,19.87551,17.125244,14.37498,11.624716,8.874452,9.775495,10.674724,11.575767,12.474996,13.374225,11.862214,10.3502035,8.838193,7.324369,5.812358,5.0255322,4.2368937,3.4500678,2.663242,1.8746033,2.3369088,2.7992141,3.2633326,3.7256382,4.1879435,6.399758,8.611572,10.825199,13.037014,15.250641,14.737573,14.224504,13.713249,13.200181,12.687112,10.700105,8.713099,6.7242785,4.7372713,2.7502642,3.3630457,3.975827,4.5867953,5.199577,5.812358,5.4008155,4.98746,4.574105,4.162562,3.7492065,3.2633326,2.7756457,2.2879589,1.8002719,1.3125849,2.2245052,3.1382382,4.0501585,4.9620786,5.8758116,9.224354,12.574709,15.925063,19.275417,22.625772,21.686659,20.749357,19.812056,18.874754,17.937452,14.349599,10.761745,7.175706,3.587853,0.0,0.22480737,0.44961473,0.6744221,0.89922947,1.1258497,2.4493124,3.774588,5.0998635,6.4251394,7.750415,9.400211,11.050007,12.699803,14.349599,15.999394,14.275268,12.549327,10.825199,9.099259,7.3751316,5.924762,4.4743915,3.0258346,1.5754645,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.2755703,0.48768693,0.69980353,0.9119202,1.1258497,1.2998942,1.4757515,1.649796,1.8256533,1.9996977,1.9743162,1.9507477,1.9253663,1.8999848,1.8746033,2.4873846,3.100166,3.7129474,4.325729,4.936697,4.699199,4.461701,4.2242026,3.9867048,3.7492065,7.124943,10.500679,13.874602,17.25034,20.624262,26.561714,32.49917,38.43843,44.375885,50.31334,55.037918,59.762497,64.487076,69.21347,73.93805,70.27587,66.61187,62.949688,59.287502,55.625317,52.662937,49.700558,46.738174,43.775795,40.8116,42.588303,44.363194,46.138084,47.912975,49.687866,47.300194,44.91252,42.52485,40.13718,37.749508,35.43798,33.124638,30.813112,28.499771,26.188244,24.750565,23.312885,21.875206,20.437527,18.999847,26.862667,34.725487,42.588303,50.44931,58.31213,54.16226,50.012386,45.862514,41.712643,37.56277,38.224503,38.888046,39.549778,40.21332,40.875053,36.975372,33.07569,29.174194,25.274511,21.374828,21.737421,22.100014,22.462606,22.8252,23.187792,24.562017,25.938055,27.31228,28.68832,30.062546,24.250187,18.43783,12.625471,6.813113,1.0007553,5.0744824,9.1500225,13.225562,17.29929,21.374828,24.449614,27.524399,30.600996,33.67578,36.750565,31.949839,27.150928,22.350203,17.549479,12.750566,14.663241,16.574104,18.48678,20.399454,22.31213,22.025682,21.737421,21.44916,21.162712,20.87445,18.575615,16.274965,13.974316,11.675479,9.374829,7.5872483,5.7996674,4.0120864,2.2245052,0.43692398,1.2255627,2.0123885,2.7992141,3.587853,4.3746786,6.5248523,8.675026,10.825199,12.975373,15.125546,14.436621,13.749508,13.062395,12.375282,11.6881695,10.2378,8.78743,7.3370595,5.8866897,4.4381323,4.2368937,4.0374675,3.8380418,3.636803,3.437377,2.7883365,2.137483,1.4866294,0.8375887,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.07433146,0.15047589,0.22480737,0.2991388,0.37528324,0.48768693,0.6000906,0.7124943,0.824898,0.93730164,1.2745126,1.6117238,1.9507477,2.2879589,2.6251698,2.137483,1.649796,1.162109,0.6744221,0.18673515,0.25018883,0.31182957,0.37528324,0.43692398,0.50037766,0.63816285,0.774135,0.9119202,1.0497054,1.1874905,1.1004683,1.0116332,0.9246109,0.8375887,0.7505665,0.8122072,0.87566096,0.93730164,1.0007553,1.062396,1.0750868,1.0877775,1.1004683,1.1131591,1.1258497,1.0370146,0.9499924,0.8629702,0.774135,0.6871128,0.61278135,0.53663695,0.46230546,0.387974,0.31182957,0.25018883,0.18673515,0.12509441,0.06164073,0.0,0.06164073,0.12509441,0.18673515,0.25018883,0.31182957,0.3245203,0.33721104,0.34990177,0.36259252,0.37528324,0.2991388,0.22480737,0.15047589,0.07433146,0.0,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.22480737,0.44961473,0.6744221,0.89922947,1.1258497,0.89922947,0.6744221,0.44961473,0.22480737,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.2374981,0.28826106,0.33721104,0.387974,0.43692398,0.44961473,0.46230546,0.4749962,0.48768693,0.50037766,0.41335547,0.3245203,0.2374981,0.15047589,0.06164073,0.13778515,0.21211663,0.28826106,0.36259252,0.43692398,0.387974,0.33721104,0.28826106,0.2374981,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.07433146,0.15047589,0.22480737,0.2991388,0.37528324,0.43692398,0.50037766,0.5620184,0.62547207,0.6871128,0.5620184,0.43692398,0.31182957,0.18673515,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.13778515,0.21211663,0.28826106,0.36259252,0.43692398,0.43692398,0.43692398,0.43692398,0.43692398,0.43692398,0.48768693,0.53663695,0.5873999,0.63816285,0.6871128,0.6000906,0.51306844,0.42423326,0.33721104,0.25018883,0.21211663,0.17585737,0.13778515,0.099712946,0.06164073,0.0870222,0.11240368,0.13778515,0.16316663,0.18673515,0.2991388,0.41335547,0.52575916,0.63816285,0.7505665,1.0116332,1.2745126,1.5373923,1.8002719,2.0631514,1.7241274,1.3869164,1.0497054,0.7124943,0.37528324,0.36259252,0.34990177,0.33721104,0.3245203,0.31182957,0.34990177,0.387974,0.42423326,0.46230546,0.50037766,0.44961473,0.40066472,0.34990177,0.2991388,0.25018883,0.4749962,0.69980353,0.9246109,1.1494182,1.3742256,1.7241274,2.0758421,2.4257438,2.7756457,3.1255474,2.525457,1.9253663,1.3252757,0.72518504,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,1.7005589,3.3376641,4.974769,6.6118746,8.2507925,7.137634,6.0244746,4.9131284,3.7999697,2.6868105,2.3133402,1.938057,1.5627737,1.1874905,0.8122072,0.824898,0.8375887,0.85027945,0.8629702,0.87566096,1.0877775,1.0007553,0.9119202,0.824898,0.73787576,0.6508536,0.83033687,1.0098201,1.1893034,1.3705997,1.550083,1.8528478,2.1556125,2.4583774,2.759329,3.0620937,2.9243085,2.7883365,2.6505513,2.5127661,2.374981,2.1592383,1.9453088,1.7295663,1.5156367,1.2998942,1.4195497,1.5392052,1.6606737,1.7803292,1.8999848,2.7448254,3.589666,4.4345064,5.279347,6.1241875,7.494787,8.865387,10.234174,11.6047735,12.975373,14.382232,15.789091,17.197763,18.604622,20.013294,17.797853,15.582414,13.366973,11.153346,8.937905,9.739235,10.542377,11.34552,12.14685,12.949992,11.49237,10.034748,8.577126,7.119504,5.661882,5.143375,4.6230545,4.102734,3.5824142,3.0620937,3.9649491,4.8678045,5.77066,6.6717024,7.574558,9.137331,10.700105,12.262879,13.825653,15.386614,14.663241,13.938056,13.212872,12.487686,11.762501,9.987611,8.212721,6.43783,4.6629395,2.8880494,3.3576066,3.827164,4.2967215,4.7680917,5.237649,4.9657044,4.691947,4.420003,4.1480584,3.874301,3.3122826,2.7502642,2.1882458,1.6244144,1.062396,1.9507477,2.8372865,3.7256382,4.612177,5.5005283,9.2044115,12.910107,16.615803,20.319685,24.025381,22.620335,21.215288,19.810242,18.405195,17.00015,13.742256,10.484363,7.228282,3.9703882,0.7124943,0.88472575,1.0569572,1.2291887,1.403233,1.5754645,3.1219215,4.670192,6.2166486,7.764919,9.313189,10.741803,12.172231,13.602658,15.033086,16.4617,14.860854,13.258195,11.655537,10.052877,8.450218,7.0451727,5.6401267,4.2350807,2.8300345,1.4249886,1.1494182,0.87566096,0.6000906,0.3245203,0.05076295,0.21936847,0.38978696,0.56020546,0.7306239,0.89922947,1.0406405,1.1802386,1.3198367,1.4594349,1.6008459,2.0595255,2.520018,2.9805105,3.43919,3.8996825,5.3391747,6.78048,8.219973,9.659465,11.10077,10.725487,10.3502035,9.97492,9.599637,9.224354,11.992747,14.759329,17.527721,20.294304,23.062696,26.684996,30.307295,33.929596,37.551895,41.176006,44.898018,48.62003,52.34204,56.06587,59.78788,58.509743,57.233418,55.955276,54.67714,53.400814,50.35322,47.305634,44.25804,41.210453,38.16286,39.32497,40.48708,41.651,42.81311,43.97522,41.83955,39.705692,37.570023,35.434353,33.300495,31.757666,30.214834,28.672003,27.129171,25.588154,23.793322,21.996675,20.201841,18.40701,16.612177,23.249432,29.886688,36.525757,43.163013,49.80027,46.49524,43.19021,39.885178,36.580147,33.275116,33.590572,33.904213,34.21967,34.535126,34.85058,32.239914,29.629248,27.020395,24.409729,21.800875,22.950293,24.099712,25.24913,26.400362,27.54978,27.653118,27.754644,27.857983,27.959509,28.062847,23.069948,18.07705,13.084151,8.093065,3.100166,7.0868707,11.075388,15.062093,19.050611,23.037315,25.589968,28.142618,30.695269,33.24792,35.80057,33.46729,31.135818,28.802536,26.469254,24.137783,23.167849,22.197914,21.22798,20.258043,19.288109,20.653269,22.016617,23.381779,24.746939,26.1121,22.81976,19.52742,16.23508,12.9427395,9.6504,8.113008,6.5756154,5.038223,3.5008307,1.9616255,2.5780327,3.1926272,3.8072214,4.421816,5.038223,6.4577727,7.877322,9.296872,10.718235,12.137785,11.691795,11.24762,10.801631,10.357455,9.91328,10.00574,10.098202,10.190662,10.283124,10.375585,8.854509,7.3352466,5.814171,4.2949085,2.7756457,2.3441606,1.9144884,1.4848163,1.0551442,0.62547207,2.0649643,3.5044568,4.945762,6.3852544,7.8247466,6.7242785,5.6256227,4.5251546,3.4246864,2.324218,2.0105755,1.69512,1.3796645,1.064209,0.7505665,1.7857682,2.819157,3.8543584,4.88956,5.924762,4.954827,3.9848917,3.0149567,2.0450218,1.0750868,0.94274056,0.8103943,0.678048,0.54570174,0.41335547,0.52032024,0.62728506,0.73424983,0.8430276,0.9499924,0.88472575,0.8194591,0.7541924,0.69073874,0.62547207,0.69073874,0.7541924,0.8194591,0.88472575,0.9499924,0.9499924,0.9499924,0.9499924,0.9499924,0.9499924,0.90829426,0.86478317,0.823085,0.7795739,0.73787576,0.64722764,0.55839247,0.46774435,0.3770962,0.28826106,0.23205921,0.17767033,0.12328146,0.06707962,0.012690738,0.06164073,0.11240368,0.16316663,0.21211663,0.26287958,0.27194437,0.28282216,0.291887,0.30276474,0.31182957,0.25018883,0.18673515,0.12509441,0.06164073,0.0,0.03988518,0.07977036,0.11965553,0.15954071,0.19942589,0.15954071,0.11965553,0.07977036,0.03988518,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1794833,0.36077955,0.5402629,0.7197462,0.89922947,0.7197462,0.5402629,0.36077955,0.1794833,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.19942589,0.25018883,0.2991388,0.34990177,0.40066472,0.42060733,0.4405499,0.4604925,0.48043507,0.50037766,0.41516843,0.32995918,0.24474995,0.15954071,0.07433146,0.13959812,0.20486477,0.27013144,0.33539808,0.40066472,0.36259252,0.3245203,0.28826106,0.25018883,0.21211663,0.17585737,0.13778515,0.099712946,0.06164073,0.025381476,0.07977036,0.13415924,0.19036107,0.24474995,0.2991388,0.3680314,0.43511102,0.50219065,0.56927025,0.63816285,0.5275721,0.4169814,0.30820364,0.19761293,0.0870222,0.07070554,0.052575916,0.034446288,0.018129626,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.099712946,0.099712946,0.099712946,0.099712946,0.099712946,0.15047589,0.19942589,0.25018883,0.2991388,0.34990177,0.36077955,0.36984438,0.38072214,0.38978696,0.40066472,0.46774435,0.53482395,0.60190356,0.67079616,0.73787576,0.64541465,0.5529536,0.4604925,0.3680314,0.2755703,0.23205921,0.19036107,0.14684997,0.10515183,0.06164073,0.092461094,0.12328146,0.15228885,0.18310922,0.21211663,0.2955129,0.3770962,0.4604925,0.5420758,0.62547207,0.83577573,1.0442665,1.2545701,1.4648738,1.6751775,1.405046,1.1349145,0.86478317,0.5946517,0.3245203,0.31726846,0.3100166,0.30276474,0.2955129,0.28826106,0.33177215,0.3770962,0.4224203,0.46774435,0.51306844,0.46230546,0.41335547,0.36259252,0.31182957,0.26287958,0.46955732,0.678048,0.88472575,1.0932164,1.2998942,1.5700256,1.840157,2.1102884,2.38042,2.6505513,2.1392958,1.6298534,1.1204109,0.6091554,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.03988518,0.06707962,0.09427405,0.12328146,0.15047589,0.16679256,0.18492219,0.2030518,0.21936847,0.2374981,1.7621996,3.2869012,4.8134155,6.338117,7.8628187,6.7242785,5.5875506,4.4508233,3.3122826,2.175555,1.889107,1.6044719,1.3198367,1.0352017,0.7505665,0.7505665,0.7505665,0.7505665,0.7505665,0.7505665,1.3633479,1.1874905,1.0116332,0.8375887,0.66173136,0.48768693,0.7106813,0.9318628,1.1548572,1.3778516,1.6008459,1.8546607,2.1102884,2.3641033,2.619731,2.8753586,2.663242,2.4493124,2.2371957,2.0250793,1.8129625,1.7078108,1.6026589,1.4975071,1.3923552,1.2872034,1.6407311,1.9924458,2.3441606,2.6976883,3.049403,3.8652363,4.6792564,5.4950895,6.3109226,7.124943,8.2779875,9.429218,10.582263,11.735307,12.888351,13.789393,14.692248,15.595104,16.49796,17.400814,15.720199,14.039582,12.360779,10.680162,8.999546,9.704789,10.410031,11.115273,11.820516,12.525759,11.122525,9.719293,8.317872,6.9146395,5.5132194,5.2594047,5.0074024,4.7554007,4.503399,4.249584,5.5929894,6.9345818,8.2779875,9.619579,10.962985,11.874905,12.786825,13.700559,14.612478,15.524399,14.587097,13.649796,12.712494,11.775192,10.837891,9.275117,7.7123427,6.149569,4.5867953,3.0258346,3.3521678,3.680314,4.006647,4.3347936,4.6629395,4.5305934,4.3982472,4.265901,4.1317415,3.9993954,3.3630457,2.7248828,2.08672,1.4503701,0.8122072,1.6751775,2.5381477,3.3993049,4.262275,5.125245,9.184468,13.245504,17.304728,21.365765,25.424988,23.552197,21.679407,19.806616,17.935638,16.062849,13.134913,10.20698,7.2790446,4.3529234,1.4249886,1.5446441,1.6642996,1.7857682,1.9054236,2.0250793,3.7945306,5.565795,7.3352466,9.104698,10.874149,12.085209,13.294455,14.505513,15.71476,16.92582,15.444629,13.965251,12.48406,11.004683,9.525306,8.165584,6.8058615,5.4443264,4.0846047,2.7248828,2.1882458,1.649796,1.1131591,0.5747091,0.038072214,0.16497959,0.291887,0.42060733,0.5475147,0.6744221,0.7795739,0.88472575,0.9898776,1.0950294,1.2001812,2.1447346,3.0892882,4.0356545,4.9802084,5.924762,8.192778,10.460794,12.726997,14.995013,17.26303,16.749962,16.236893,15.725637,15.212569,14.699501,16.860552,19.01979,21.180841,23.34008,25.49932,26.808277,28.115423,29.42257,30.729715,32.03686,34.758118,37.477562,40.197006,42.918262,45.637707,46.745426,47.853146,48.96087,50.066776,51.174496,48.041695,44.91071,41.77791,38.64511,35.51231,36.061638,36.612778,37.162106,37.71325,38.262577,36.380722,34.49705,32.615196,30.733341,28.849674,28.07735,27.305029,26.532707,25.760386,24.988064,22.834263,20.682278,18.53029,16.378304,14.224504,19.63801,25.049704,30.463211,35.874905,41.2866,38.82822,36.36803,33.90784,31.447649,28.98746,28.954826,28.922192,28.889559,28.856926,28.824291,27.504456,26.184618,24.864782,23.544945,22.22511,24.163166,26.09941,28.037466,29.975523,31.911768,30.742407,29.573046,28.401873,27.232512,26.06315,21.88971,17.718082,13.544643,9.373016,5.199577,9.099259,13.000754,16.900436,20.80012,24.699802,26.73032,28.760838,30.789543,32.82006,34.85058,34.984737,35.120712,35.25487,35.390842,35.525,31.672457,27.81991,23.967365,20.11482,16.262274,19.279043,22.297626,25.314396,28.33298,31.349749,27.065718,22.779875,18.494032,14.210001,9.924157,8.636953,7.3497505,6.0625467,4.7753434,3.48814,3.930503,4.3728657,4.8152285,5.2575917,5.6999545,6.390693,7.079619,7.7703576,8.459284,9.1500225,8.94697,8.745731,8.54268,8.339628,8.138389,9.771869,11.407161,13.042453,14.677745,16.313038,13.472125,10.633025,7.7921133,4.953014,2.1121013,1.9017978,1.693307,1.4830034,1.2726997,1.062396,3.9794528,6.8983226,9.815379,12.732436,15.649493,13.374225,11.10077,8.825501,6.550234,4.274966,3.531651,2.7901495,2.0468347,1.305333,0.5620184,2.2952106,4.02659,5.7597823,7.4929743,9.224354,7.7721705,6.319988,4.8678045,3.4156215,1.9616255,1.6352923,1.3071461,0.9808127,0.6526665,0.3245203,0.40247768,0.48043507,0.55839247,0.6345369,0.7124943,0.67079616,0.62728506,0.5855869,0.5420758,0.50037766,0.56745726,0.6345369,0.7016165,0.7705091,0.8375887,0.824898,0.8122072,0.7995165,0.7868258,0.774135,0.7777609,0.7795739,0.78319985,0.7850128,0.7868258,0.68167394,0.57833505,0.47318324,0.3680314,0.26287958,0.21574254,0.16679256,0.11965553,0.072518505,0.025381476,0.06164073,0.099712946,0.13778515,0.17585737,0.21211663,0.21936847,0.22662032,0.23568514,0.24293698,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13415924,0.27013144,0.40429065,0.5402629,0.6744221,0.5402629,0.40429065,0.27013144,0.13415924,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.16316663,0.21211663,0.26287958,0.31182957,0.36259252,0.38978696,0.4169814,0.44417584,0.47318324,0.50037766,0.4169814,0.33539808,0.2520018,0.17041849,0.0870222,0.14322405,0.19761293,0.2520018,0.30820364,0.36259252,0.33721104,0.31182957,0.28826106,0.26287958,0.2374981,0.19942589,0.16316663,0.12509441,0.0870222,0.05076295,0.08520924,0.11965553,0.15410182,0.19036107,0.22480737,0.29732585,0.36984438,0.44236287,0.5148814,0.5873999,0.49312583,0.39703882,0.30276474,0.20667773,0.11240368,0.09064813,0.06707962,0.045324065,0.02175555,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.13778515,0.16316663,0.18673515,0.21211663,0.2374981,0.26287958,0.28282216,0.30276474,0.32270733,0.34264994,0.36259252,0.44780177,0.533011,0.61822027,0.7016165,0.7868258,0.69073874,0.59283876,0.4949388,0.39703882,0.2991388,0.2520018,0.20486477,0.15772775,0.11059072,0.06164073,0.09789998,0.13234627,0.16679256,0.2030518,0.2374981,0.29007402,0.34264994,0.39522585,0.44780177,0.50037766,0.65810543,0.81583315,0.97174793,1.1294757,1.2872034,1.0841516,0.88291276,0.67986095,0.47680917,0.2755703,0.27194437,0.27013144,0.26831847,0.26469254,0.26287958,0.3154555,0.3680314,0.42060733,0.47318324,0.52575916,0.4749962,0.42423326,0.37528324,0.3245203,0.2755703,0.46411842,0.6544795,0.8448406,1.0352017,1.2255627,1.4141108,1.6044719,1.794833,1.9851941,2.175555,1.7549478,1.3343405,0.9155461,0.4949388,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.06707962,0.11059072,0.15228885,0.19579996,0.2374981,0.27194437,0.30820364,0.34264994,0.3770962,0.41335547,1.8256533,3.2379513,4.650249,6.0625467,7.474845,6.3127356,5.1506267,3.9867048,2.8245957,1.6624867,1.4666867,1.2726997,1.0768998,0.88291276,0.6871128,0.6744221,0.66173136,0.6508536,0.63816285,0.62547207,1.6371052,1.3742256,1.1131591,0.85027945,0.5873999,0.3245203,0.58921283,0.8557183,1.1204109,1.3851035,1.649796,1.8582866,2.0649643,2.2716422,2.4801328,2.6868105,2.4003625,2.1121013,1.8256533,1.5373923,1.2491312,1.2545701,1.260009,1.2654479,1.2708868,1.2745126,1.8600996,2.4456866,3.0294604,3.6150475,4.2006345,4.985647,5.77066,6.5556726,7.3406854,8.125698,9.059374,9.994863,10.930351,11.86584,12.799516,13.198368,13.595407,13.992445,14.389484,14.786523,13.642544,12.496751,11.352772,10.20698,9.063,9.670342,10.277685,10.885027,11.49237,12.099712,10.752681,9.40565,8.056806,6.7097745,5.3627434,5.377247,5.391751,5.408067,5.422571,5.4370747,7.219217,9.003172,10.785315,12.567456,14.349599,14.612478,14.875358,15.138238,15.399304,15.662184,14.512766,13.363347,12.212116,11.062697,9.91328,8.562622,7.211965,5.863121,4.512464,3.1618068,3.346729,3.531651,3.7183862,3.9033084,4.0882306,4.0954823,4.102734,4.1099863,4.117238,4.12449,3.4119956,2.6995013,1.987007,1.2745126,0.5620184,1.3996071,2.2371957,3.0747845,3.9123733,4.749962,9.164526,13.57909,17.995466,22.41003,26.824594,24.485872,22.145338,19.804804,17.464268,15.125546,12.527572,9.929596,7.3316207,4.7354584,2.137483,2.2045624,2.2716422,2.3405347,2.4076142,2.474694,4.4671397,6.4595857,8.452031,10.444477,12.436923,13.426801,14.416678,15.408369,16.398247,17.388124,16.030214,14.672306,13.314397,11.958302,10.600392,9.284182,7.9697833,6.6553855,5.3391747,4.024777,3.2252605,2.4257438,1.6244144,0.824898,0.025381476,0.11059072,0.19579996,0.27919623,0.36440548,0.44961473,0.52032024,0.58921283,0.65991837,0.7306239,0.7995165,2.229944,3.6603715,5.090799,6.5194135,7.949841,11.044568,14.139296,17.235836,20.330563,23.42529,22.774435,22.125395,21.474543,20.8255,20.174648,21.728357,23.280252,24.832148,26.385857,27.937754,26.929747,25.92174,24.915545,23.907537,22.89953,24.616405,26.335094,28.05197,29.768847,31.487534,34.9793,38.472878,41.964645,45.458225,48.94999,45.73198,42.515785,39.297775,36.07977,32.86176,32.800117,32.736664,32.675026,32.611572,32.54993,30.920076,29.290224,27.66037,26.030518,24.400663,24.397038,24.395224,24.391598,24.389786,24.387972,21.87702,19.36788,16.856926,14.347786,11.836833,16.024776,20.212719,24.400663,28.586794,32.77474,31.159388,29.544039,27.930502,26.315151,24.699802,24.31908,23.94017,23.559448,23.18054,22.799818,22.768997,22.73999,22.70917,22.680162,22.649342,25.374224,28.099108,30.825802,33.550686,36.27557,33.833508,31.389635,28.947573,26.505512,24.06164,20.70947,17.357304,14.005136,10.652968,7.3008003,11.111648,14.924308,18.736969,22.54963,26.36229,27.870674,29.377245,30.88563,32.392204,33.90059,36.50219,39.105602,41.707203,44.31062,46.91222,40.177063,33.44372,26.70675,19.971596,13.238253,17.906631,22.576822,27.247015,31.917206,36.5874,31.309864,26.03233,20.754795,15.477262,10.199727,9.162713,8.125698,7.0868707,6.049856,5.0128417,5.282973,5.5531044,5.823236,6.093367,6.3616858,6.3218007,6.281915,6.24203,6.202145,6.16226,6.202145,6.24203,6.281915,6.3218007,6.3616858,9.539809,12.717933,15.896056,19.072367,22.25049,18.08974,13.930804,9.770056,5.6093063,1.4503701,1.4594349,1.4703126,1.4793775,1.4902552,1.49932,5.8957543,10.290376,14.684997,19.079618,23.476053,20.024172,16.575916,13.125849,9.675781,6.2257137,5.0545397,3.8851788,2.715818,1.5446441,0.37528324,2.8046532,5.235836,7.665206,10.094576,12.525759,10.589515,8.655084,6.720652,4.784408,2.8499773,2.327844,1.8057107,1.2817645,0.75963134,0.2374981,0.28463513,0.33177215,0.38072214,0.42785916,0.4749962,0.4550536,0.43511102,0.41516843,0.39522585,0.37528324,0.44417584,0.5148814,0.5855869,0.6544795,0.72518504,0.69980353,0.6744221,0.6508536,0.62547207,0.6000906,0.64722764,0.69436467,0.7433147,0.7904517,0.8375887,0.7179332,0.5982776,0.47680917,0.35715362,0.2374981,0.19761293,0.15772775,0.11784257,0.07795739,0.038072214,0.06164073,0.0870222,0.11240368,0.13778515,0.16316663,0.16679256,0.17223145,0.17767033,0.18310922,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.09064813,0.1794833,0.27013144,0.36077955,0.44961473,0.36077955,0.27013144,0.1794833,0.09064813,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.12509441,0.17585737,0.22480737,0.2755703,0.3245203,0.36077955,0.39522585,0.42967212,0.46411842,0.50037766,0.42060733,0.34083697,0.25925365,0.1794833,0.099712946,0.14503701,0.19036107,0.23568514,0.27919623,0.3245203,0.31182957,0.2991388,0.28826106,0.2755703,0.26287958,0.22480737,0.18673515,0.15047589,0.11240368,0.07433146,0.09064813,0.10515183,0.11965553,0.13415924,0.15047589,0.22662032,0.3045777,0.3825351,0.4604925,0.53663695,0.45686656,0.3770962,0.29732585,0.21755551,0.13778515,0.11059072,0.08339628,0.054388877,0.027194439,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.07433146,0.099712946,0.12509441,0.15047589,0.17585737,0.17585737,0.17585737,0.17585737,0.17585737,0.17585737,0.20486477,0.23568514,0.26469254,0.2955129,0.3245203,0.42785916,0.5293851,0.6327239,0.73424983,0.8375887,0.73424983,0.6327239,0.5293851,0.42785916,0.3245203,0.27194437,0.21936847,0.16679256,0.11421664,0.06164073,0.10333887,0.14322405,0.18310922,0.2229944,0.26287958,0.28463513,0.30820364,0.32995918,0.35171473,0.37528324,0.48043507,0.5855869,0.69073874,0.79407763,0.89922947,0.7650702,0.629098,0.4949388,0.36077955,0.22480737,0.22662032,0.23024625,0.23205921,0.23568514,0.2374981,0.29732585,0.35715362,0.4169814,0.47680917,0.53663695,0.48768693,0.43692398,0.387974,0.33721104,0.28826106,0.4604925,0.6327239,0.80495536,0.97718686,1.1494182,1.260009,1.3705997,1.4793775,1.5899682,1.7005589,1.3705997,1.0406405,0.7106813,0.38072214,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.09427405,0.15228885,0.21030366,0.26831847,0.3245203,0.3770962,0.42967212,0.48224804,0.53482395,0.5873999,1.887294,3.1871881,4.4870825,5.7869763,7.0868707,5.89938,4.7118897,3.5243993,2.3369088,1.1494182,1.0442665,0.93911463,0.83577573,0.7306239,0.62547207,0.6000906,0.5747091,0.5493277,0.52575916,0.50037766,1.9126755,1.5627737,1.2128719,0.8629702,0.51306844,0.16316663,0.46955732,0.7777609,1.0841516,1.3923552,1.7005589,1.8600996,2.0196402,2.179181,2.3405347,2.5000753,2.137483,1.7748904,1.4122978,1.0497054,0.6871128,0.8031424,0.91735905,1.0333886,1.1476053,1.261822,2.079468,2.8971143,3.7147603,4.5324063,5.3500524,6.104245,6.8602505,7.614443,8.370448,9.12464,9.842574,10.560507,11.276628,11.99456,12.712494,12.605529,12.496751,12.389787,12.282822,12.175857,11.564888,10.955733,10.344765,9.735609,9.12464,9.635896,10.145339,10.654781,11.164224,11.675479,10.382836,9.090195,7.797552,6.5049095,5.2122674,5.4950895,5.7779117,6.060734,6.341743,6.624565,8.847258,11.069949,13.292642,15.515334,17.738026,17.350052,16.962078,16.575916,16.187943,15.799969,14.436621,13.075087,11.711739,10.3502035,8.9868555,7.850128,6.7134004,5.57486,4.4381323,3.299592,3.343103,3.3848011,3.4283123,3.4700103,3.5117085,3.6603715,3.8072214,3.9558845,4.102734,4.249584,3.4627585,2.6741197,1.887294,1.1004683,0.31182957,1.1258497,1.938057,2.7502642,3.5624714,4.3746786,9.144584,13.914488,18.684393,23.454296,28.224201,25.417736,22.609457,19.80299,16.99471,14.188245,11.920229,9.652213,7.3841968,5.1179934,2.8499773,2.864481,2.8807976,2.8953013,2.909805,2.9243085,5.139749,7.3551893,9.570629,11.784257,13.999697,14.770206,15.540715,16.309412,17.07992,17.85043,16.615803,15.379361,14.144734,12.910107,11.675479,10.4045925,9.135518,7.8646317,6.5955577,5.3246713,4.262275,3.199879,2.137483,1.0750868,0.012690738,0.054388877,0.09789998,0.13959812,0.18310922,0.22480737,0.25925365,0.2955129,0.32995918,0.36440548,0.40066472,2.3151531,4.229642,6.145943,8.0604315,9.97492,13.898171,17.819609,21.74286,25.664299,29.58755,28.800724,28.012085,27.22526,26.438433,25.649796,26.594349,27.540714,28.485268,29.429821,30.374374,27.053028,23.729868,20.406708,17.08536,13.762199,14.476506,15.192626,15.906934,16.623055,17.33736,23.214987,29.092611,34.970234,40.84786,46.725483,43.422268,40.12086,36.817646,33.514427,30.213022,29.536787,28.862364,28.187943,27.511707,26.837286,25.459433,24.081581,22.705544,21.327692,19.94984,20.716722,21.48542,22.252302,23.019186,23.787882,20.919775,18.051668,15.185374,12.317267,9.449161,12.411542,15.375735,18.338116,21.300497,24.262878,23.492369,22.72186,21.953163,21.182655,20.412146,19.685148,18.958149,18.22934,17.50234,16.775343,18.035353,19.29536,20.55537,21.815378,23.075388,26.587097,30.100618,33.612328,37.125847,40.637558,36.922794,33.208035,29.493275,25.776703,22.061941,19.529232,16.998337,14.465629,11.9329195,9.400211,13.125849,16.849674,20.575312,24.300951,28.024776,29.009214,29.995466,30.979904,31.964344,32.950596,38.019638,43.090496,48.15954,53.230396,58.29944,48.683483,39.06572,29.44795,19.830185,10.212419,16.534218,22.857832,29.179632,35.503246,41.825047,35.55582,29.284784,23.01556,16.744522,10.475298,9.686659,8.899834,8.113008,7.324369,6.5375433,6.635443,6.733343,6.82943,6.92733,7.02523,6.2547207,5.484212,4.7155156,3.9450066,3.1744974,3.4573197,3.7401419,4.022964,4.305786,4.5867953,9.30775,14.026892,18.747847,23.466988,28.187943,22.707355,17.228584,11.747997,6.2674117,0.7868258,1.017072,1.2473183,1.4775645,1.7078108,1.938057,7.8102427,13.682428,19.554615,25.4268,31.300798,26.674118,22.051064,17.424383,12.799516,8.174648,6.5774283,4.9802084,3.3829882,1.7857682,0.18673515,3.3159087,6.4432693,9.570629,12.697989,15.825351,13.406858,10.990179,8.571687,6.155008,3.738329,3.0203958,2.3024626,1.5845293,0.8665961,0.15047589,0.16679256,0.18492219,0.2030518,0.21936847,0.2374981,0.23931105,0.24293698,0.24474995,0.24837588,0.25018883,0.32270733,0.39522585,0.46774435,0.5402629,0.61278135,0.5747091,0.53663695,0.50037766,0.46230546,0.42423326,0.5166943,0.6091554,0.7016165,0.79589057,0.8883517,0.7523795,0.61822027,0.48224804,0.3480888,0.21211663,0.1794833,0.14684997,0.11421664,0.08339628,0.05076295,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.11421664,0.11784257,0.11965553,0.12328146,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.045324065,0.09064813,0.13415924,0.1794833,0.22480737,0.1794833,0.13415924,0.09064813,0.045324065,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.0870222,0.13778515,0.18673515,0.2374981,0.28826106,0.32995918,0.37165734,0.41516843,0.45686656,0.50037766,0.4224203,0.3444629,0.26831847,0.19036107,0.11240368,0.14684997,0.18310922,0.21755551,0.2520018,0.28826106,0.28826106,0.28826106,0.28826106,0.28826106,0.28826106,0.25018883,0.21211663,0.17585737,0.13778515,0.099712946,0.09427405,0.09064813,0.08520924,0.07977036,0.07433146,0.15772775,0.23931105,0.32270733,0.40429065,0.48768693,0.4224203,0.35715362,0.291887,0.22662032,0.16316663,0.13053331,0.09789998,0.065266654,0.032633327,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.06164073,0.099712946,0.13778515,0.17585737,0.21211663,0.18673515,0.16316663,0.13778515,0.11240368,0.0870222,0.12690738,0.16679256,0.20667773,0.24837588,0.28826106,0.40791658,0.5275721,0.64722764,0.7668832,0.8883517,0.7795739,0.6726091,0.5656443,0.45686656,0.34990177,0.291887,0.23568514,0.17767033,0.11965553,0.06164073,0.10696479,0.15228885,0.19761293,0.24293698,0.28826106,0.27919623,0.27194437,0.26469254,0.2574407,0.25018883,0.30276474,0.35534066,0.40791658,0.4604925,0.51306844,0.44417584,0.3770962,0.3100166,0.24293698,0.17585737,0.18310922,0.19036107,0.19761293,0.20486477,0.21211663,0.27919623,0.3480888,0.41516843,0.48224804,0.5493277,0.50037766,0.44961473,0.40066472,0.34990177,0.2991388,0.4550536,0.6091554,0.7650702,0.91917205,1.0750868,1.1040943,1.1349145,1.1657349,1.1947423,1.2255627,0.98443866,0.7451276,0.5058166,0.26469254,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.12328146,0.19579996,0.26831847,0.34083697,0.41335547,0.48224804,0.5529536,0.62184614,0.69255173,0.76325727,1.9507477,3.1382382,4.325729,5.5132194,6.70071,5.487838,4.274966,3.0620937,1.8492218,0.63816285,0.62184614,0.6073425,0.59283876,0.57833505,0.5620184,0.52575916,0.48768693,0.44961473,0.41335547,0.37528324,2.1882458,1.7495089,1.3125849,0.87566096,0.43692398,0.0,0.34990177,0.69980353,1.0497054,1.3996071,1.7495089,1.8619126,1.9743162,2.08672,2.1991236,2.3133402,1.8746033,1.4376793,1.0007553,0.5620184,0.12509441,0.34990177,0.5747091,0.7995165,1.0243238,1.2491312,2.3006494,3.350355,4.40006,5.4497657,6.4994707,7.224656,7.949841,8.675026,9.400211,10.125396,10.625773,11.124338,11.624716,12.125093,12.625471,12.012691,11.399909,10.7871275,10.174346,9.563377,9.487233,9.412902,9.336758,9.262425,9.188094,9.599637,10.012992,10.424535,10.837891,11.249433,10.012992,8.774739,7.5382986,6.300045,5.0617914,5.612932,6.16226,6.7134004,7.262728,7.8120556,10.475298,13.136727,15.799969,18.463211,21.12464,20.087626,19.050611,18.011784,16.97477,15.937754,14.362289,12.786825,11.213174,9.637709,8.062244,7.137634,6.2130227,5.2865987,4.361988,3.437377,3.3376641,3.2379513,3.1382382,3.0367124,2.9369993,3.2252605,3.5117085,3.7999697,4.0882306,4.3746786,3.5117085,2.6505513,1.7875811,0.9246109,0.06164073,0.85027945,1.6371052,2.4257438,3.2125697,3.9993954,9.12464,14.249886,19.375132,24.500376,29.625622,26.349598,23.075388,19.799364,16.525154,13.24913,11.312886,9.374829,7.4367723,5.5005283,3.5624714,3.5243993,3.48814,3.4500678,3.4119956,3.3757362,5.812358,8.2507925,10.687414,13.125849,15.56247,16.1118,16.66294,17.212267,17.763407,18.312735,17.199575,16.08823,14.975071,13.861912,12.750566,11.525003,10.29944,9.07569,7.850128,6.624565,5.2992897,3.975827,2.6505513,1.3252757,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.4003625,4.800725,7.1992745,9.599637,11.999999,16.749962,21.499924,26.249886,30.999847,35.74981,34.8252,33.90059,32.974163,32.049553,31.12494,31.462152,31.799364,32.13839,32.475597,32.81281,27.174496,21.537996,15.899682,10.263181,4.6248674,4.3366065,4.0501585,3.7618973,3.4754493,3.1871881,11.450671,19.712341,27.975826,36.237495,44.49917,41.112553,37.725937,34.337513,30.949083,27.56247,26.275267,24.988064,23.70086,22.411844,21.12464,20.000603,18.874754,17.750717,16.624866,15.50083,17.038223,18.575615,20.113007,21.650398,23.187792,19.96253,16.73727,13.512011,10.28675,7.063302,8.80012,10.536939,12.27557,14.012388,15.749206,15.825351,15.899682,15.975826,16.050158,16.124489,15.049402,13.974316,12.899229,11.8241415,10.750868,13.299893,15.850732,18.399757,20.950596,23.49962,27.799969,32.100315,36.40066,40.699196,44.999546,40.012085,35.024624,30.037165,25.049704,20.062244,18.350807,16.637558,14.924308,13.212872,11.499621,15.138238,18.77504,22.411844,26.050459,29.687262,30.149569,30.611874,31.074179,31.538298,32.000603,39.537086,47.075386,54.611874,62.15017,69.68665,57.18809,44.687714,32.187336,19.68696,7.1883965,15.161806,23.137028,31.112251,39.087475,47.062695,39.79997,32.53724,25.274511,18.011784,10.750868,10.212419,9.675781,9.137331,8.600695,8.062244,7.987913,7.911769,7.837437,7.763106,7.686961,6.187641,4.688321,3.1871881,1.6878681,0.18673515,0.7124943,1.2382535,1.7621996,2.2879589,2.811905,9.07569,15.337664,21.599636,27.863422,34.125393,27.324972,20.52455,13.724127,6.925517,0.12509441,0.5747091,1.0243238,1.4757515,1.9253663,2.374981,9.724731,17.074482,24.426044,31.775795,39.125546,33.324066,27.524399,21.724731,15.925063,10.125396,8.100317,6.0752378,4.0501585,2.0250793,0.0,3.825351,7.650702,11.47424,15.299591,19.124943,16.224201,13.325275,10.424535,7.5256076,4.6248674,3.7129474,2.7992141,1.887294,0.97537386,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.19942589,0.2755703,0.34990177,0.42423326,0.50037766,0.44961473,0.40066472,0.34990177,0.2991388,0.25018883,0.387974,0.52575916,0.66173136,0.7995165,0.93730164,0.7868258,0.63816285,0.48768693,0.33721104,0.18673515,0.16316663,0.13778515,0.11240368,0.0870222,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06164073,0.12509441,0.18673515,0.25018883,0.31182957,0.25018883,0.18673515,0.12509441,0.06164073,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,0.2991388,0.34990177,0.40066472,0.44961473,0.50037766,0.42423326,0.34990177,0.2755703,0.19942589,0.12509441,0.15047589,0.17585737,0.19942589,0.22480737,0.25018883,0.26287958,0.2755703,0.28826106,0.2991388,0.31182957,0.2755703,0.2374981,0.19942589,0.16316663,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0870222,0.17585737,0.26287958,0.34990177,0.43692398,0.387974,0.33721104,0.28826106,0.2374981,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.0,0.0,0.0,0.0,0.0,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,0.387974,0.52575916,0.66173136,0.7995165,0.93730164,0.824898,0.7124943,0.6000906,0.48768693,0.37528324,0.31182957,0.25018883,0.18673515,0.12509441,0.06164073,0.11240368,0.16316663,0.21211663,0.26287958,0.31182957,0.2755703,0.2374981,0.19942589,0.16316663,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.13778515,0.15047589,0.16316663,0.17585737,0.18673515,0.26287958,0.33721104,0.41335547,0.48768693,0.5620184,0.51306844,0.46230546,0.41335547,0.36259252,0.31182957,0.44961473,0.5873999,0.72518504,0.8629702,1.0007553,0.9499924,0.89922947,0.85027945,0.7995165,0.7505665,0.6000906,0.44961473,0.2991388,0.15047589,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.15047589,0.2374981,0.3245203,0.41335547,0.50037766,0.5873999,0.6744221,0.76325727,0.85027945,0.93730164,2.0123885,3.0874753,4.162562,5.237649,6.3127356,5.0744824,3.8380418,2.5997884,1.3633479,0.12509441,0.19942589,0.2755703,0.34990177,0.42423326,0.50037766,0.44961473,0.40066472,0.34990177,0.2991388,0.25018883,2.3876717,1.9199274,1.452183,0.98443866,0.5166943,0.05076295,0.32814622,0.6055295,0.88291276,1.1602961,1.4376793,1.6026589,1.7676386,1.9326181,2.0975976,2.2625773,1.9181144,1.5718386,1.2273756,0.88291276,0.53663695,0.8629702,1.1874905,1.5120108,1.8383441,2.1628644,3.1944401,4.227829,5.2594047,6.2927933,7.324369,7.7757964,8.225411,8.675026,9.12464,9.574255,9.835322,10.094576,10.355642,10.614896,10.874149,10.431787,9.989424,9.547061,9.104698,8.662335,9.046683,9.432844,9.817192,10.203354,10.587702,11.082641,11.5775795,12.072517,12.567456,13.062395,11.307447,9.5525,7.797552,6.0426044,4.2876563,4.9276323,5.567608,6.207584,6.8475595,7.4875355,9.610515,11.731681,13.85466,15.977639,18.100618,17.308353,16.514277,15.722012,14.929747,14.137483,12.92461,11.711739,10.500679,9.287807,8.074935,7.115878,6.155008,5.1941376,4.2350807,3.2742105,3.1327994,2.9895754,2.8481643,2.70494,2.561716,3.1128569,3.6621845,4.213325,4.762653,5.3119802,4.4526362,3.5932918,2.7321346,1.8727903,1.0116332,1.5083848,2.0033236,2.4982624,2.9932013,3.48814,7.8483152,12.206677,16.566853,20.927027,25.287203,22.460793,19.632572,16.80435,13.9779415,11.14972,9.527119,7.9045167,6.281915,4.6593137,3.0367124,3.0330863,3.0276475,3.0222087,3.0167696,3.0131438,5.0599785,7.1068134,9.155461,11.202296,13.24913,13.667925,14.084907,14.501887,14.920682,15.337664,14.68681,14.037769,13.386916,12.737875,12.087022,11.024626,9.96223,8.899834,7.837437,6.775041,6.6118746,6.450521,6.2873545,6.1241875,5.962834,6.9980354,8.033237,9.066626,10.101828,11.137029,10.05469,8.972352,7.890013,6.8076744,5.7253356,6.7569118,7.7903004,8.821876,9.855265,10.88684,14.4692545,18.051668,21.635895,25.21831,28.800724,28.762651,28.724579,28.68832,28.650248,28.612175,29.310165,30.008156,30.704334,31.402325,32.100315,26.420303,20.740292,15.06028,9.380268,3.7002566,3.8652363,4.0302157,4.195195,4.360175,4.5251546,10.852394,17.179634,23.506872,29.835926,36.163166,33.465477,30.767788,28.070099,25.372412,22.674723,21.626831,20.580751,19.53286,18.484966,17.437075,17.355492,17.272095,17.190512,17.107115,17.025532,17.533161,18.04079,18.54842,19.054237,19.561867,17.322857,15.082036,12.843027,10.602205,8.363196,9.313189,10.263181,11.213174,12.163166,13.113158,13.1602955,13.207433,13.254569,13.301706,13.3506565,15.105604,16.860552,18.6155,20.370447,22.125395,25.047892,27.970387,30.892883,33.815376,36.737873,37.056953,37.37785,37.69693,38.017826,38.336906,34.660217,30.98353,27.305029,23.628342,19.94984,19.244598,18.539356,17.834112,17.130684,16.425442,18.94002,21.4546,23.96918,26.48557,29.000149,28.717327,28.434505,28.151684,27.870674,27.587852,34.30488,41.021904,47.740746,54.45777,61.174797,50.53452,39.896053,29.253963,18.6155,7.9752226,13.999697,20.024172,26.050459,32.074936,38.099407,32.627888,27.154554,21.683033,16.209698,10.738177,9.924157,9.11195,8.299743,7.4875355,6.6753283,6.5701766,6.4650245,6.359873,6.2547207,6.149569,5.081734,4.0157123,2.9478772,1.8800422,0.8122072,1.6824293,2.5526514,3.4228733,4.2930956,5.163317,9.7773075,14.39311,19.0071,23.622902,28.236893,22.8252,17.413506,11.999999,6.588306,1.1747998,1.3270886,1.4793775,1.6316663,1.7857682,1.938057,8.049554,14.162864,20.27436,26.38767,32.50098,27.634989,22.77081,17.904818,13.04064,8.174648,7.95528,7.7340984,7.51473,7.2953615,7.07418,8.9596615,10.845142,12.730623,14.614291,16.499773,14.895301,13.290829,11.684544,10.080072,8.4756,7.2971745,6.1205616,4.942136,3.7655232,2.5870976,2.077655,1.5682126,1.0569572,0.5475147,0.038072214,0.059827764,0.08339628,0.10515183,0.12690738,0.15047589,0.20667773,0.26469254,0.32270733,0.38072214,0.43692398,0.42423326,0.41335547,0.40066472,0.387974,0.37528324,0.46955732,0.5656443,0.65991837,0.7541924,0.85027945,0.7179332,0.5855869,0.45324063,0.3208944,0.18673515,0.16679256,0.14684997,0.12690738,0.10696479,0.0870222,0.08520924,0.08339628,0.07977036,0.07795739,0.07433146,0.07795739,0.07977036,0.08339628,0.08520924,0.0870222,0.07070554,0.052575916,0.034446288,0.018129626,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.059827764,0.10696479,0.15410182,0.2030518,0.25018883,0.23931105,0.23024625,0.21936847,0.21030366,0.19942589,0.15954071,0.11965553,0.07977036,0.03988518,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.030820364,0.047137026,0.065266654,0.08339628,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.04169814,0.08520924,0.12690738,0.17041849,0.21211663,0.25925365,0.30820364,0.35534066,0.40247768,0.44961473,0.38978696,0.32995918,0.27013144,0.21030366,0.15047589,0.17041849,0.19036107,0.21030366,0.23024625,0.25018883,0.2520018,0.25562772,0.2574407,0.25925365,0.26287958,0.23024625,0.19761293,0.16497959,0.13234627,0.099712946,0.08339628,0.065266654,0.047137026,0.030820364,0.012690738,0.0870222,0.16316663,0.2374981,0.31182957,0.387974,0.3680314,0.3480888,0.32814622,0.30820364,0.28826106,0.23024625,0.17223145,0.11421664,0.058014803,0.0,0.0,0.0,0.0,0.0,0.0,0.03988518,0.07977036,0.11965553,0.15954071,0.19942589,0.16316663,0.12509441,0.0870222,0.05076295,0.012690738,0.058014803,0.10333887,0.14684997,0.19217403,0.2374981,0.3934129,0.5475147,0.7016165,0.8575313,1.0116332,0.88291276,0.7523795,0.62184614,0.49312583,0.36259252,0.3100166,0.2574407,0.20486477,0.15228885,0.099712946,0.13959812,0.1794833,0.21936847,0.25925365,0.2991388,0.35171473,0.40429065,0.45686656,0.5094425,0.5620184,0.47318324,0.3825351,0.291887,0.2030518,0.11240368,0.11240368,0.11240368,0.11240368,0.11240368,0.11240368,0.11965553,0.12690738,0.13415924,0.14322405,0.15047589,0.21030366,0.27013144,0.32995918,0.38978696,0.44961473,0.4169814,0.38434806,0.35171473,0.3208944,0.28826106,0.40791658,0.5275721,0.64722764,0.7668832,0.8883517,0.8321498,0.7777609,0.72337204,0.6671702,0.61278135,0.49312583,0.37165734,0.2520018,0.13234627,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.02175555,0.032633327,0.04169814,0.052575916,0.06164073,0.13234627,0.2030518,0.27194437,0.34264994,0.41335547,0.5058166,0.5982776,0.69073874,0.78319985,0.87566096,1.7857682,2.6958754,3.6041696,4.514277,5.424384,4.3783045,3.3304121,2.2825198,1.2346275,0.18673515,0.23024625,0.27194437,0.3154555,0.35715362,0.40066472,0.36440548,0.32995918,0.2955129,0.25925365,0.22480737,2.5870976,2.0903459,1.5917811,1.0950294,0.5982776,0.099712946,0.3045777,0.5094425,0.71430725,0.91917205,1.1258497,1.3415923,1.5591478,1.7767034,1.9942589,2.2118144,1.9598125,1.7078108,1.455809,1.2019942,0.9499924,1.3742256,1.8002719,2.2245052,2.6505513,3.0747845,4.0900435,5.105303,6.1205616,7.135821,8.149267,8.325124,8.499168,8.675026,8.8508835,9.024928,9.04487,9.064813,9.084756,9.104698,9.12464,8.852696,8.580752,8.306994,8.03505,7.763106,8.607946,9.452786,10.297627,11.142468,11.9873085,12.565643,13.142166,13.720501,14.297023,14.875358,12.601903,10.330261,8.056806,5.7851634,3.5117085,4.2423325,4.972956,5.7017674,6.432391,7.1630154,8.745731,10.326634,11.909351,13.492067,15.074784,14.527269,13.979754,13.43224,12.884725,12.337211,11.486931,10.636651,9.788185,8.937905,8.087626,7.0923095,6.096993,5.101677,4.1081734,3.1128569,2.9279346,2.7430124,2.5580902,2.373168,2.1882458,3.000453,3.8126602,4.6248674,5.4370747,6.249282,5.391751,4.5342193,3.6766882,2.819157,1.9616255,2.1646774,2.3677292,2.570781,2.7720199,2.9750717,6.5701766,10.165281,13.760386,17.355492,20.950596,18.570175,16.189756,13.809336,11.430729,9.050309,7.743163,6.434204,5.127058,3.8199122,2.5127661,2.5399606,2.5671551,2.5943494,2.6233568,2.6505513,4.307599,5.964647,7.6216946,9.280556,10.937603,11.222239,11.506873,11.793322,12.077957,12.362592,12.175857,11.9873085,11.800573,11.612025,11.42529,10.524248,9.625018,8.725789,7.8247466,6.925517,7.9244595,8.925215,9.924157,10.924912,11.925668,13.994258,16.064661,18.135065,20.205467,22.275871,20.10938,17.944704,15.780026,13.615349,11.450671,11.115273,10.779876,10.444477,10.110892,9.775495,12.19036,14.6052265,17.020092,19.43496,21.849825,22.700104,23.550385,24.400663,25.24913,26.09941,27.15818,28.215137,29.272095,30.330864,31.387821,25.664299,19.942589,14.219066,8.497355,2.7756457,3.392053,4.0102735,4.6266804,5.2449007,5.863121,10.254116,14.646925,19.039734,23.43254,27.82535,25.816587,23.809637,21.802689,19.795738,17.786976,16.980207,16.171627,15.364858,14.558089,13.749508,14.710379,15.6694355,16.630306,17.589363,18.550234,18.0281,17.504154,16.982021,16.459887,15.937754,14.683184,13.426801,12.172231,10.917661,9.663091,9.824444,9.987611,10.150778,10.312131,10.475298,10.49524,10.515183,10.535126,10.555068,10.57501,15.159993,19.744976,24.329958,28.91494,33.499924,36.795887,40.090042,43.38601,46.68016,49.97431,46.315754,42.655384,38.99501,35.33464,31.674269,29.308353,26.940624,24.572895,22.205166,19.837437,20.140202,20.442966,20.745731,21.046682,21.349447,22.741802,24.134157,25.528326,26.920681,28.313036,27.285088,26.257137,25.229187,24.20305,23.1751,29.072668,34.970234,40.8678,46.76537,52.662937,43.88276,35.10258,26.322403,17.542227,8.762048,12.837588,16.913128,20.986855,25.062395,29.137934,25.455807,21.771868,18.08974,14.407614,10.725487,9.637709,8.549932,7.462154,6.3743763,5.2865987,5.1524396,5.0182805,4.882308,4.748149,4.612177,3.97764,3.343103,2.7067533,2.0722163,1.4376793,2.6523643,3.8670492,5.081734,6.298232,7.512917,10.480737,13.446743,16.414564,19.382383,22.350203,18.325426,14.300649,10.274059,6.249282,2.2245052,2.079468,1.9344311,1.789394,1.6443571,1.49932,6.376189,11.249433,16.124489,20.999546,25.874601,21.9441,18.01541,14.084907,10.154404,6.2257137,7.8102427,9.394773,10.979301,12.565643,14.150173,14.095784,14.039582,13.985193,13.930804,13.874602,13.564586,13.254569,12.944552,12.634536,12.32452,10.883214,9.440096,7.996978,6.5556726,5.1125546,4.1045475,3.0983531,2.0903459,1.0823387,0.07433146,0.09427405,0.11421664,0.13415924,0.15410182,0.17585737,0.21574254,0.25562772,0.2955129,0.33539808,0.37528324,0.40066472,0.42423326,0.44961473,0.4749962,0.50037766,0.5529536,0.6055295,0.65810543,0.7106813,0.76325727,0.64722764,0.533011,0.4169814,0.30276474,0.18673515,0.17223145,0.15772775,0.14322405,0.12690738,0.11240368,0.10696479,0.10333887,0.09789998,0.092461094,0.0870222,0.092461094,0.09789998,0.10333887,0.10696479,0.11240368,0.09064813,0.06707962,0.045324065,0.02175555,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.058014803,0.09064813,0.12328146,0.15410182,0.18673515,0.23024625,0.27194437,0.3154555,0.35715362,0.40066472,0.3208944,0.23931105,0.15954071,0.07977036,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.059827764,0.09427405,0.13053331,0.16497959,0.19942589,0.15954071,0.11965553,0.07977036,0.03988518,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.034446288,0.07070554,0.10515183,0.13959812,0.17585737,0.21936847,0.26469254,0.3100166,0.35534066,0.40066472,0.35534066,0.3100166,0.26469254,0.21936847,0.17585737,0.19036107,0.20486477,0.21936847,0.23568514,0.25018883,0.24293698,0.23568514,0.22662032,0.21936847,0.21211663,0.18492219,0.15772775,0.13053331,0.10333887,0.07433146,0.065266654,0.054388877,0.045324065,0.034446288,0.025381476,0.0870222,0.15047589,0.21211663,0.2755703,0.33721104,0.3480888,0.35715362,0.3680314,0.3770962,0.387974,0.3100166,0.23205921,0.15410182,0.07795739,0.0,0.0,0.0,0.0,0.0,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.065266654,0.10515183,0.14503701,0.18492219,0.22480737,0.39703882,0.56927025,0.7433147,0.9155461,1.0877775,0.93911463,0.79226464,0.64541465,0.49675176,0.34990177,0.30820364,0.26469254,0.2229944,0.1794833,0.13778515,0.16679256,0.19761293,0.22662032,0.2574407,0.28826106,0.42967212,0.5728962,0.71430725,0.8575313,1.0007553,0.8194591,0.6399758,0.4604925,0.27919623,0.099712946,0.099712946,0.099712946,0.099712946,0.099712946,0.099712946,0.10333887,0.10515183,0.10696479,0.11059072,0.11240368,0.15772775,0.2030518,0.24837588,0.291887,0.33721104,0.32270733,0.30820364,0.291887,0.27738327,0.26287958,0.36440548,0.46774435,0.56927025,0.6726091,0.774135,0.71430725,0.6544795,0.5946517,0.53482395,0.4749962,0.38434806,0.2955129,0.20486477,0.11421664,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.032633327,0.03988518,0.047137026,0.054388877,0.06164073,0.11421664,0.16679256,0.21936847,0.27194437,0.3245203,0.4224203,0.52032024,0.61822027,0.71430725,0.8122072,1.5573349,2.3024626,3.04759,3.7927177,4.537845,3.680314,2.8227828,1.9652514,1.1077201,0.25018883,0.25925365,0.27013144,0.27919623,0.29007402,0.2991388,0.27919623,0.25925365,0.23931105,0.21936847,0.19942589,2.7883365,2.2607644,1.7331922,1.2056202,0.678048,0.15047589,0.28282216,0.41516843,0.5475147,0.67986095,0.8122072,1.0823387,1.35247,1.6226015,1.892733,2.1628644,2.0033236,1.84197,1.6824293,1.5228885,1.3633479,1.887294,2.4130533,2.9369993,3.4627585,3.9867048,4.985647,5.9827766,6.979906,7.9770355,8.974165,8.874452,8.774739,8.675026,8.575313,8.4756,8.254418,8.03505,7.8156815,7.5945,7.3751316,7.271793,7.170267,7.066928,6.965402,6.8620634,8.167397,9.47273,10.778063,12.083396,13.386916,14.046834,14.706753,15.366671,16.028402,16.68832,13.898171,11.108022,8.317872,5.527723,2.7375734,3.5570326,4.3783045,5.197764,6.017223,6.836682,7.8791356,8.921589,9.965856,11.008308,12.050762,11.747997,11.445232,11.142468,10.839704,10.536939,10.049252,9.563377,9.07569,8.588004,8.100317,7.0705543,6.0407915,5.009216,3.9794528,2.94969,2.72307,2.4946365,2.268016,2.039583,1.8129625,2.8880494,3.9631362,5.038223,6.11331,7.1883965,6.3326783,5.47696,4.6230545,3.7673361,2.913431,2.8227828,2.7321346,2.6432993,2.5526514,2.4620032,5.292038,8.122072,10.952107,13.782142,16.612177,14.679558,12.74694,10.8143215,8.881703,6.9490857,5.957395,4.9657044,3.972201,2.9805105,1.987007,2.0468347,2.1066625,2.1683033,2.228131,2.2879589,3.5552197,4.8224807,6.089741,7.3570023,8.624263,8.776552,8.930654,9.082943,9.235231,9.38752,9.663091,9.936848,10.212419,10.487988,10.761745,10.025683,9.287807,8.549932,7.8120556,7.07418,9.237044,11.399909,13.562773,15.725637,17.888502,20.992294,24.097898,27.203503,30.307295,33.4129,30.165884,26.917055,23.67004,20.423023,17.176008,15.471823,13.769451,12.067079,10.364707,8.662335,9.909654,11.156972,12.40429,13.651608,14.898927,16.637558,18.374376,20.113007,21.849825,23.586643,25.00438,26.422117,27.839853,29.25759,30.675327,24.910107,19.144884,13.379663,7.614443,1.8492218,2.9206827,3.9903307,5.0599785,6.1296263,7.1992745,9.657652,12.114216,14.572594,17.029158,19.487535,18.169512,16.851488,15.535276,14.217253,12.899229,12.331772,11.764315,11.1968565,10.629399,10.061942,12.065266,14.066776,16.0701,18.073423,20.074934,18.523039,16.96933,15.417434,13.865538,12.311829,12.0416975,11.771566,11.503247,11.233116,10.962985,10.337513,9.712041,9.086569,8.46291,7.837437,7.8301854,7.8229337,7.8156815,7.806617,7.799365,15.214382,22.629398,30.046228,37.461246,44.87445,48.542072,52.209698,55.87732,59.544945,63.212566,55.572742,47.93292,40.293095,32.651455,25.011631,23.954674,22.897717,21.84076,20.78199,19.725033,21.035805,22.344765,23.655537,24.964495,26.275267,26.545399,26.815529,27.08566,27.355793,27.624111,25.852846,24.07977,22.306692,20.535427,18.76235,23.840458,28.916754,33.99486,39.07297,44.149265,37.229187,30.31092,23.38903,16.470764,9.550687,11.675479,13.800271,15.925063,18.049856,20.174648,18.281914,16.389181,14.4964485,12.605529,10.712796,9.349448,7.987913,6.624565,5.2630305,3.8996825,3.7347028,3.5697234,3.4047437,3.2397642,3.0747845,2.8717327,2.6704938,2.467442,2.2643902,2.0631514,3.6222992,5.18326,6.742408,8.303369,9.862516,11.182353,12.50219,13.822026,15.141864,16.4617,13.825653,11.187792,8.549932,5.9120708,3.2742105,2.8318477,2.3894846,1.9471219,1.504759,1.062396,4.701012,8.337815,11.974618,15.613234,19.250036,16.255022,13.260008,10.264994,7.26998,4.274966,7.665206,11.055446,14.445685,17.835926,21.224354,19.230095,17.235836,15.239763,13.245504,11.249433,12.235684,13.220123,14.204562,15.190813,16.175253,14.467442,12.75963,11.05182,9.345822,7.6380115,6.1332526,4.6284933,3.1219215,1.6171626,0.11240368,0.13053331,0.14684997,0.16497959,0.18310922,0.19942589,0.2229944,0.24474995,0.26831847,0.29007402,0.31182957,0.37528324,0.43692398,0.50037766,0.5620184,0.62547207,0.6345369,0.64541465,0.6544795,0.6653573,0.6744221,0.57833505,0.48043507,0.3825351,0.28463513,0.18673515,0.17767033,0.16679256,0.15772775,0.14684997,0.13778515,0.13053331,0.12328146,0.11421664,0.10696479,0.099712946,0.10696479,0.11421664,0.12328146,0.13053331,0.13778515,0.11059072,0.08339628,0.054388877,0.027194439,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.054388877,0.072518505,0.09064813,0.10696479,0.12509441,0.21936847,0.3154555,0.40972954,0.5058166,0.6000906,0.48043507,0.36077955,0.23931105,0.11965553,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.09064813,0.14322405,0.19579996,0.24837588,0.2991388,0.23931105,0.1794833,0.11965553,0.059827764,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.09064813,0.06707962,0.045324065,0.02175555,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.027194439,0.054388877,0.08339628,0.11059072,0.13778515,0.1794833,0.2229944,0.26469254,0.30820364,0.34990177,0.3208944,0.29007402,0.25925365,0.23024625,0.19942589,0.21030366,0.21936847,0.23024625,0.23931105,0.25018883,0.23205921,0.21574254,0.19761293,0.1794833,0.16316663,0.13959812,0.11784257,0.09427405,0.072518505,0.05076295,0.047137026,0.045324065,0.04169814,0.03988518,0.038072214,0.0870222,0.13778515,0.18673515,0.2374981,0.28826106,0.32814622,0.3680314,0.40791658,0.44780177,0.48768693,0.38978696,0.291887,0.19579996,0.09789998,0.0,0.0,0.0,0.0,0.0,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.0870222,0.07433146,0.06164073,0.05076295,0.038072214,0.072518505,0.10696479,0.14322405,0.17767033,0.21211663,0.40247768,0.59283876,0.78319985,0.97174793,1.162109,0.99712944,0.8321498,0.6671702,0.50219065,0.33721104,0.3045777,0.27194437,0.23931105,0.20667773,0.17585737,0.19579996,0.21574254,0.23568514,0.25562772,0.2755703,0.5076295,0.73968875,0.97174793,1.2056202,1.4376793,1.167548,0.8974165,0.62728506,0.35715362,0.0870222,0.0870222,0.0870222,0.0870222,0.0870222,0.0870222,0.08520924,0.08339628,0.07977036,0.07795739,0.07433146,0.10515183,0.13415924,0.16497959,0.19579996,0.22480737,0.22662032,0.23024625,0.23205921,0.23568514,0.2374981,0.32270733,0.40791658,0.49312583,0.57833505,0.66173136,0.5982776,0.533011,0.46774435,0.40247768,0.33721104,0.27738327,0.21755551,0.15772775,0.09789998,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.04169814,0.047137026,0.052575916,0.058014803,0.06164073,0.09789998,0.13234627,0.16679256,0.2030518,0.2374981,0.34083697,0.44236287,0.54570174,0.64722764,0.7505665,1.3307146,1.9108626,2.4891977,3.0693457,3.6494937,2.9823234,2.3151531,1.647983,0.9808127,0.31182957,0.29007402,0.26831847,0.24474995,0.2229944,0.19942589,0.19579996,0.19036107,0.18492219,0.1794833,0.17585737,2.9877625,2.42937,1.8727903,1.3143979,0.75781834,0.19942589,0.25925365,0.3208944,0.38072214,0.4405499,0.50037766,0.823085,1.1457924,1.4666867,1.789394,2.1121013,2.0450218,1.9779422,1.9108626,1.84197,1.7748904,2.4003625,3.0258346,3.6494937,4.274966,4.900438,5.8794374,6.8602505,7.83925,8.820063,9.800876,9.425592,9.050309,8.675026,8.299743,7.9244595,7.46578,7.0052876,6.544795,6.0843024,5.6256227,5.6927023,5.7597823,5.826862,5.8957543,5.962834,7.7268467,9.492672,11.256684,13.022511,14.788336,15.529838,16.273151,17.014654,17.757969,18.49947,15.192626,11.885782,8.577126,5.2702823,1.9616255,2.8717327,3.7818398,4.691947,5.6020546,6.5121617,7.0143523,7.518356,8.020547,8.5227375,9.024928,8.966913,8.910711,8.852696,8.794682,8.736667,8.613385,8.488291,8.363196,8.238102,8.113008,7.0469856,5.9827766,4.9167547,3.8525455,2.7883365,2.518205,2.2480736,1.9779422,1.7078108,1.4376793,2.7756457,4.1117992,5.4497657,6.787732,8.125698,7.271793,6.4197006,5.567608,4.7155156,3.8616104,3.4808881,3.0983531,2.715818,2.333283,1.9507477,4.0157123,6.0806766,8.145641,10.210606,12.27557,10.790753,9.304124,7.819308,6.3344913,4.8496747,4.171627,3.4953918,2.817344,2.1392958,1.4630609,1.5555218,1.647983,1.7404441,1.8329052,1.9253663,2.8028402,3.680314,4.557788,5.4352617,6.3127356,6.3326783,6.352621,6.3725634,6.392506,6.412449,7.1503243,7.8882003,8.624263,9.362139,10.100015,9.525306,8.950596,8.374074,7.799365,7.224656,10.549629,13.874602,17.199575,20.52455,23.849524,27.99033,32.129322,36.27013,40.410934,44.54993,40.220573,35.88941,31.560053,27.230698,22.89953,19.830185,16.76084,13.68968,10.620335,7.549176,7.6307597,7.71053,7.7903004,7.8700705,7.949841,10.57501,13.200181,15.825351,18.45052,21.07569,22.852394,24.629097,26.407614,28.184317,29.962833,24.155914,18.347181,12.540262,6.73153,0.9246109,2.4474995,3.9703882,5.4932766,7.0143523,8.537241,9.059374,9.583321,10.1054535,10.627586,11.14972,10.522435,9.89515,9.267865,8.640579,8.013294,7.6851482,7.3570023,7.0306687,6.7025228,6.3743763,9.420154,12.464118,15.509895,18.555672,21.599636,19.017977,16.434505,13.852847,11.269376,8.6877165,9.402024,10.118144,10.832452,11.546759,12.262879,10.850581,9.438283,8.024173,6.6118746,5.199577,5.1651306,5.130684,5.0944247,5.0599785,5.0255322,15.270584,25.515635,35.76069,46.005737,56.25079,60.29007,64.32935,68.370445,72.40973,76.45082,64.82973,53.210453,41.589363,29.970085,18.348995,18.60281,18.85481,19.106813,19.360628,19.612629,21.929596,24.246561,26.56534,28.882307,31.199272,30.347181,29.495089,28.642996,27.789091,26.936998,24.420607,21.902401,19.384195,16.867804,14.349599,18.608248,22.865084,27.12192,31.38057,35.637405,30.577427,25.517448,20.45747,15.397491,10.337513,10.51337,10.687414,10.863272,11.037316,11.213174,11.109835,11.008308,10.90497,10.801631,10.700105,9.063,7.4258947,5.7869763,4.1498713,2.5127661,2.3169663,2.1229792,1.9271792,1.7331922,1.5373923,1.7676386,1.9978848,2.228131,2.4583774,2.6868105,4.592234,6.497658,8.403082,10.306692,12.212116,11.885782,11.557636,11.22949,10.903157,10.57501,9.324066,8.074935,6.825804,5.57486,4.325729,3.584227,2.8445382,2.1048496,1.3651608,0.62547207,3.0258346,5.424384,7.8247466,10.225109,12.625471,10.564133,8.504607,6.445082,4.3855567,2.324218,7.520169,12.714307,17.910257,23.104395,28.300346,24.364405,20.430275,16.494333,12.5602045,8.624263,10.90497,13.185677,15.464571,17.745277,20.024172,18.051668,16.080978,14.106662,12.134158,10.161655,8.160145,6.156821,4.15531,2.1519866,0.15047589,0.16497959,0.1794833,0.19579996,0.21030366,0.22480737,0.23024625,0.23568514,0.23931105,0.24474995,0.25018883,0.34990177,0.44961473,0.5493277,0.6508536,0.7505665,0.7179332,0.6852999,0.6526665,0.6200332,0.5873999,0.5076295,0.42785916,0.3480888,0.26831847,0.18673515,0.18310922,0.17767033,0.17223145,0.16679256,0.16316663,0.15228885,0.14322405,0.13234627,0.12328146,0.11240368,0.12328146,0.13234627,0.14322405,0.15228885,0.16316663,0.13053331,0.09789998,0.065266654,0.032633327,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.052575916,0.054388877,0.058014803,0.059827764,0.06164073,0.21030366,0.35715362,0.5058166,0.6526665,0.7995165,0.6399758,0.48043507,0.3208944,0.15954071,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.11965553,0.19036107,0.25925365,0.32995918,0.40066472,0.3208944,0.23931105,0.15954071,0.07977036,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.13959812,0.1794833,0.21936847,0.25925365,0.2991388,0.28463513,0.27013144,0.25562772,0.23931105,0.22480737,0.23024625,0.23568514,0.23931105,0.24474995,0.25018883,0.2229944,0.19579996,0.16679256,0.13959812,0.11240368,0.09427405,0.07795739,0.059827764,0.04169814,0.025381476,0.030820364,0.034446288,0.03988518,0.045324065,0.05076295,0.0870222,0.12509441,0.16316663,0.19942589,0.2374981,0.30820364,0.3770962,0.44780177,0.5166943,0.5873999,0.46955732,0.35171473,0.23568514,0.11784257,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.07977036,0.11059072,0.13959812,0.17041849,0.19942589,0.40791658,0.61459434,0.823085,1.0297627,1.2382535,1.0551442,0.872035,0.69073874,0.5076295,0.3245203,0.30276474,0.27919623,0.2574407,0.23568514,0.21211663,0.2229944,0.23205921,0.24293698,0.2520018,0.26287958,0.5855869,0.90829426,1.2291887,1.551896,1.8746033,1.5156367,1.1548572,0.79589057,0.43511102,0.07433146,0.07433146,0.07433146,0.07433146,0.07433146,0.07433146,0.06707962,0.059827764,0.052575916,0.045324065,0.038072214,0.052575916,0.06707962,0.08339628,0.09789998,0.11240368,0.13234627,0.15228885,0.17223145,0.19217403,0.21211663,0.27919623,0.3480888,0.41516843,0.48224804,0.5493277,0.48043507,0.40972954,0.34083697,0.27013144,0.19942589,0.17041849,0.13959812,0.11059072,0.07977036,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.052575916,0.054388877,0.058014803,0.059827764,0.06164073,0.07977036,0.09789998,0.11421664,0.13234627,0.15047589,0.2574407,0.36440548,0.47318324,0.58014804,0.6871128,1.1022812,1.5174497,1.9326181,2.3477864,2.762955,2.2843328,1.8075237,1.3307146,0.8520924,0.37528324,0.3208944,0.26469254,0.21030366,0.15410182,0.099712946,0.11059072,0.11965553,0.13053331,0.13959812,0.15047589,3.1871881,2.5997884,2.0123885,1.4249886,0.8375887,0.25018883,0.2374981,0.22480737,0.21211663,0.19942589,0.18673515,0.5620184,0.93730164,1.3125849,1.6878681,2.0631514,2.08672,2.1121013,2.137483,2.1628644,2.1882458,2.911618,3.636803,4.361988,5.087173,5.812358,6.775041,7.7377243,8.700407,9.663091,10.625773,9.97492,9.325879,8.675026,8.024173,7.3751316,6.6753283,5.975525,5.275721,4.574105,3.874301,4.1117992,4.349297,4.5867953,4.8242936,5.0617914,7.28811,9.512614,11.73712,13.963438,16.187943,17.01284,17.837738,18.662638,19.487535,20.312433,16.487082,12.661731,8.838193,5.0128417,1.1874905,2.1882458,3.1871881,4.1879435,5.186886,6.187641,6.149569,6.11331,6.0752378,6.037165,6.000906,6.187641,6.3743763,6.5629244,6.7496595,6.9382076,7.175706,7.413204,7.650702,7.8882003,8.125698,7.02523,5.924762,4.8242936,3.7256382,2.6251698,2.3133402,1.9996977,1.6878681,1.3742256,1.062396,2.663242,4.262275,5.863121,7.462154,9.063,8.212721,7.362441,6.5121617,5.661882,4.8116026,4.137181,3.4627585,2.7883365,2.1121013,1.4376793,2.7375734,4.0374675,5.337362,6.637256,7.93715,6.9001355,5.863121,4.8242936,3.787279,2.7502642,2.3876717,2.0250793,1.6624867,1.2998942,0.93730164,1.062396,1.1874905,1.3125849,1.4376793,1.5627737,2.0504606,2.5381477,3.0258346,3.5117085,3.9993954,3.8869917,3.774588,3.6621845,3.5497808,3.437377,4.6375585,5.8377395,7.037921,8.238102,9.438283,9.024928,8.613385,8.200029,7.7866745,7.3751316,11.862214,16.349297,20.838192,25.325274,29.812357,34.986553,40.16256,45.336754,50.512764,55.68696,50.275265,44.86176,39.450066,34.03656,28.624866,24.186733,19.750414,15.312282,10.874149,6.43783,5.3500524,4.262275,3.1744974,2.08672,1.0007553,4.512464,8.024173,11.537694,15.049402,18.562923,20.700407,22.837889,24.975372,27.112856,29.250338,23.399908,17.549479,11.699047,5.8504305,0.0,1.9743162,3.9504454,5.924762,7.900891,9.875207,8.46291,7.0506115,5.638314,4.2242026,2.811905,2.8753586,2.9369993,3.000453,3.0620937,3.1255474,3.0367124,2.94969,2.8626678,2.7756457,2.6868105,6.775041,10.863272,14.94969,19.03792,23.124338,19.512917,15.899682,12.28826,8.675026,5.0617914,6.7623506,8.46291,10.161655,11.862214,13.562773,11.361836,9.162713,6.9617763,4.762653,2.561716,2.5000753,2.4366217,2.374981,2.3133402,2.2498865,15.324973,28.400059,41.475143,54.550232,67.62532,72.03807,76.449005,80.861755,85.274506,89.687256,74.08853,58.487988,42.887444,27.2869,11.6881695,13.24913,14.811904,16.374678,17.937452,19.500225,22.8252,26.150173,29.475145,32.800117,36.12509,34.150776,32.17465,30.20033,28.224201,26.249886,22.988365,19.725033,16.4617,13.200181,9.936848,13.374225,16.811602,20.250792,23.68817,27.125546,23.925667,20.725788,17.524096,14.324218,11.124338,9.349448,7.574558,5.7996674,4.024777,2.2498865,3.9377546,5.6256227,7.311678,8.999546,10.687414,8.774739,6.8620634,4.949388,3.0367124,1.1258497,0.89922947,0.6744221,0.44961473,0.22480737,0.0,0.66173136,1.3252757,1.987007,2.6505513,3.3122826,5.562169,7.8120556,10.061942,12.311829,14.561715,12.5873995,10.613083,8.636953,6.6626377,4.688321,4.8242936,4.9620786,5.0998635,5.237649,5.375434,4.3384194,3.299592,2.2625773,1.2255627,0.18673515,1.3506571,2.5127661,3.6748753,4.836984,6.000906,4.8750563,3.7492065,2.6251698,1.49932,0.37528324,7.3751316,14.37498,21.374828,28.374678,35.374527,29.500526,23.624716,17.750717,11.874905,6.000906,9.576068,13.149418,16.72458,20.299742,23.874905,21.637709,19.400513,17.163317,14.924308,12.687112,10.1870365,7.686961,5.186886,2.6868105,0.18673515,0.19942589,0.21211663,0.22480737,0.2374981,0.25018883,0.2374981,0.22480737,0.21211663,0.19942589,0.18673515,0.3245203,0.46230546,0.6000906,0.73787576,0.87566096,0.7995165,0.72518504,0.6508536,0.5747091,0.50037766,0.43692398,0.37528324,0.31182957,0.25018883,0.18673515,0.18673515,0.18673515,0.18673515,0.18673515,0.18673515,0.17585737,0.16316663,0.15047589,0.13778515,0.12509441,0.13778515,0.15047589,0.16316663,0.17585737,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.19942589,0.40066472,0.6000906,0.7995165,1.0007553,0.7995165,0.6000906,0.40066472,0.19942589,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.15047589,0.2374981,0.3245203,0.41335547,0.50037766,0.40066472,0.2991388,0.19942589,0.099712946,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.099712946,0.13778515,0.17585737,0.21211663,0.25018883,0.25018883,0.25018883,0.25018883,0.25018883,0.25018883,0.25018883,0.25018883,0.25018883,0.25018883,0.25018883,0.21211663,0.17585737,0.13778515,0.099712946,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.0870222,0.11240368,0.13778515,0.16316663,0.18673515,0.28826106,0.387974,0.48768693,0.5873999,0.6871128,0.5493277,0.41335547,0.2755703,0.13778515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.0870222,0.11240368,0.13778515,0.16316663,0.18673515,0.41335547,0.63816285,0.8629702,1.0877775,1.3125849,1.1131591,0.9119202,0.7124943,0.51306844,0.31182957,0.2991388,0.28826106,0.2755703,0.26287958,0.25018883,0.25018883,0.25018883,0.25018883,0.25018883,0.25018883,0.66173136,1.0750868,1.4866294,1.8999848,2.3133402,1.8619126,1.4122978,0.96268314,0.51306844,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.2374981,0.28826106,0.33721104,0.387974,0.43692398,0.36259252,0.28826106,0.21211663,0.13778515,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.17585737,0.28826106,0.40066472,0.51306844,0.62547207,0.87566096,1.1258497,1.3742256,1.6244144,1.8746033,1.5881553,1.2998942,1.0116332,0.72518504,0.43692398,0.34990177,0.26287958,0.17585737,0.0870222,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,2.8626678,2.4003625,1.938057,1.4757515,1.0116332,0.5493277,0.56927025,0.58921283,0.6091554,0.629098,0.6508536,0.968122,1.2853905,1.6026589,1.9199274,2.2371957,2.3677292,2.4982624,2.6269827,2.7575161,2.8880494,3.5932918,4.2967215,5.0019636,5.7072062,6.412449,7.268167,8.122072,8.977791,9.8316965,10.687414,10.190662,9.692098,9.195346,8.696781,8.200029,7.703278,7.2047133,6.7079616,6.209397,5.712645,5.964647,6.2166486,6.4704633,6.722465,6.9744673,8.997733,11.019187,13.042453,15.065719,17.087172,17.408066,17.727148,18.048042,18.367125,18.688019,15.198066,11.708113,8.21816,4.7282066,1.2382535,2.0722163,2.907992,3.7419548,4.5777307,5.411693,5.5077806,5.6020546,5.6981416,5.7924156,5.8866897,5.8341136,5.7833505,5.730775,5.678199,5.6256227,6.002719,6.379815,6.7569118,7.135821,7.512917,6.5647373,5.618371,4.670192,3.7220123,2.7756457,2.465629,2.1556125,1.845596,1.5355793,1.2255627,2.6324217,4.0392804,5.4479527,6.8548117,8.26167,7.665206,7.066928,6.4704633,5.8721857,5.275721,4.461701,3.6494937,2.8372865,2.0250793,1.2128719,2.335096,3.4573197,4.5795436,5.7017674,6.825804,6.057108,5.290225,4.5233417,3.7546456,2.9877625,2.5453994,2.1030366,1.6606737,1.2183108,0.774135,1.1167849,1.4594349,1.8020848,2.1447346,2.4873846,3.2705846,4.0519714,4.835171,5.618371,6.399758,6.588306,6.775041,6.9617763,7.1503243,7.3370595,7.7848616,8.232663,8.680465,9.128266,9.574255,9.072064,8.569874,8.067683,7.5654926,7.063302,10.419096,13.776703,17.13431,20.491917,23.849524,28.195194,32.540867,36.884724,41.230396,45.574253,41.145187,36.716118,32.285236,27.854357,23.42529,21.1609,18.894695,16.630306,14.364102,12.099712,11.184166,10.270433,9.354887,8.439341,7.5256076,9.023115,10.520622,12.018129,13.515636,15.013144,17.607492,20.201841,22.798004,25.392353,27.986704,22.400965,16.813416,11.224051,5.638314,0.05076295,1.6371052,3.2252605,4.8134155,6.399758,7.987913,6.92733,5.866747,4.8079767,3.7473936,2.6868105,2.6704938,2.6523643,2.6342347,2.617918,2.5997884,2.7919624,2.9841363,3.1781235,3.3702974,3.5624714,6.720652,9.87702,13.035201,16.193382,19.34975,17.60024,15.850732,14.09941,12.349901,10.600392,10.745429,10.890467,11.035503,11.18054,11.325577,10.857833,10.390089,9.922344,9.4546,8.9868555,7.6724577,6.35806,5.041849,3.727451,2.4130533,12.895603,23.378153,33.860703,44.34325,54.8258,59.709923,64.595856,69.47998,74.36591,79.25003,66.062546,52.875053,39.687565,26.500074,13.312584,15.522586,17.732588,19.942589,22.15259,24.36259,25.820213,27.277836,28.735456,30.193079,31.650702,30.347181,29.045473,27.741953,26.440247,25.136726,21.831696,18.528477,15.221634,11.916603,8.613385,11.880343,15.147303,18.41426,21.683033,24.949991,22.944855,20.939718,18.934582,16.929445,14.924308,12.790451,10.654781,8.519112,6.3852544,4.249584,5.177821,6.104245,7.0324817,7.9607186,8.887142,7.3497505,5.812358,4.274966,2.7375734,1.2001812,1.0007553,0.7995165,0.6000906,0.40066472,0.19942589,1.1530442,2.1048496,3.056655,4.0102735,4.9620786,6.7079616,8.452031,10.197914,11.941984,13.687867,11.862214,10.038374,8.212721,6.3870673,4.5632267,4.740897,4.9167547,5.0944247,5.272095,5.4497657,5.3573046,5.2648435,5.1723824,5.0799212,4.98746,6.836682,8.6877165,10.536939,12.387974,14.237195,11.715364,9.19172,6.6698895,4.1480584,1.6244144,7.2047133,12.785012,18.36531,23.94561,29.52591,25.272697,21.019487,16.768091,12.514881,8.26167,11.381779,14.501887,17.621996,20.742105,23.862213,21.96404,20.067682,18.169512,16.273151,14.37498,11.735307,9.0956335,6.454147,3.8144734,1.1747998,0.98443866,0.79589057,0.6055295,0.41516843,0.22480737,0.21936847,0.21574254,0.21030366,0.20486477,0.19942589,0.35534066,0.5094425,0.6653573,0.8194591,0.97537386,0.88291276,0.7904517,0.6979906,0.6055295,0.51306844,0.44961473,0.387974,0.3245203,0.26287958,0.19942589,0.19942589,0.19942589,0.19942589,0.19942589,0.19942589,0.18310922,0.16497959,0.14684997,0.13053331,0.11240368,0.11965553,0.12690738,0.13415924,0.14322405,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.14322405,0.17223145,0.2030518,0.23205921,0.26287958,0.36984438,0.47680917,0.5855869,0.69255173,0.7995165,0.6399758,0.48043507,0.3208944,0.15954071,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.52213323,0.9445535,1.3669738,1.789394,2.2118144,1.7694515,1.3270886,0.88472575,0.44236287,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.13959812,0.20486477,0.27013144,0.33539808,0.40066472,0.3770962,0.35534066,0.33177215,0.3100166,0.28826106,0.25925365,0.23205921,0.20486477,0.17767033,0.15047589,0.13959812,0.13053331,0.11965553,0.11059072,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.07977036,0.11059072,0.13959812,0.17041849,0.19942589,0.2030518,0.20486477,0.20667773,0.21030366,0.21211663,0.21755551,0.2229944,0.22662032,0.23205921,0.2374981,0.21755551,0.19761293,0.17767033,0.15772775,0.13778515,0.11059072,0.08339628,0.054388877,0.027194439,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.092461094,0.11059072,0.12690738,0.14503701,0.16316663,0.26469254,0.3680314,0.46955732,0.5728962,0.6744221,0.56020546,0.44417584,0.32995918,0.21574254,0.099712946,0.08520924,0.07070554,0.054388877,0.03988518,0.025381476,0.02175555,0.01994259,0.018129626,0.014503701,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.07433146,0.09427405,0.11421664,0.13415924,0.15410182,0.17585737,0.35171473,0.5293851,0.7070554,0.88472575,1.062396,0.9246109,0.7868258,0.6508536,0.51306844,0.37528324,0.35171473,0.32995918,0.30820364,0.28463513,0.26287958,0.25562772,0.24837588,0.23931105,0.23205921,0.22480737,0.55476654,0.88472575,1.214685,1.5446441,1.8746033,1.5101979,1.1457924,0.7795739,0.41516843,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.04169814,0.034446288,0.027194439,0.01994259,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.032633327,0.065266654,0.09789998,0.13053331,0.16316663,0.20486477,0.24837588,0.29007402,0.33177215,0.37528324,0.3100166,0.24474995,0.1794833,0.11421664,0.05076295,0.054388877,0.059827764,0.065266654,0.07070554,0.07433146,0.072518505,0.07070554,0.06707962,0.065266654,0.06164073,0.059827764,0.058014803,0.054388877,0.052575916,0.05076295,0.052575916,0.054388877,0.058014803,0.059827764,0.06164073,0.15047589,0.2374981,0.3245203,0.41335547,0.50037766,0.7106813,0.91917205,1.1294757,1.3397794,1.550083,1.3307146,1.1095331,0.8901646,0.67079616,0.44961473,0.36440548,0.27919623,0.19579996,0.11059072,0.025381476,0.03988518,0.054388877,0.07070554,0.08520924,0.099712946,2.5381477,2.1991236,1.8619126,1.5247015,1.1874905,0.85027945,0.90285534,0.9554313,1.0080072,1.0605831,1.1131591,1.3724127,1.6316663,1.892733,2.1519866,2.4130533,2.6469254,2.8826106,3.1182957,3.3521678,3.587853,4.273153,4.95664,5.6419396,6.3272395,7.0125394,7.75948,8.508233,9.255174,10.002114,10.750868,10.4045925,10.060129,9.715667,9.3693905,9.024928,8.729415,8.435715,8.140202,7.844689,7.549176,7.817495,8.0858135,8.352319,8.620637,8.887142,10.707357,12.527572,14.347786,16.168001,17.988214,17.803293,17.61837,17.431635,17.246714,17.06179,13.907236,10.752681,7.5981264,4.441758,1.2872034,1.9579996,2.6269827,3.2977788,3.966762,4.6375585,4.8641787,5.092612,5.319232,5.5476656,5.774286,5.482399,5.1905117,4.896812,4.604925,4.313038,4.8297324,5.3482394,5.864934,6.3816285,6.9001355,6.104245,5.3101673,4.514277,3.720199,2.9243085,2.617918,2.3097143,2.0033236,1.69512,1.3869164,2.6016014,3.8180993,5.032784,6.247469,7.462154,7.117691,6.773228,6.4269524,6.0824895,5.7380266,4.788034,3.8380418,2.8880494,1.938057,0.9880646,1.9326181,2.8771715,3.8217251,4.7680917,5.712645,5.2158933,4.7173285,4.220577,3.7220123,3.2252605,2.7031271,2.179181,1.6570477,1.1349145,0.61278135,1.1729867,1.7331922,2.2933977,2.8517902,3.4119956,4.4907084,5.567608,6.644508,7.723221,8.80012,9.287807,9.775495,10.263181,10.750868,11.236742,10.932164,10.627586,10.323009,10.016619,9.712041,9.119202,8.528176,7.935337,7.3424983,6.7496595,8.977791,11.204109,13.43224,15.660371,17.886688,21.402023,24.917358,28.432692,31.948027,35.461548,32.015106,28.56685,25.120409,21.672155,18.225714,18.133251,18.04079,17.94833,17.85587,17.763407,17.020092,16.276777,15.535276,14.791962,14.05046,13.531953,13.015259,12.496751,11.980057,11.463363,14.514579,17.567608,20.620636,23.671852,26.724882,21.40021,16.075539,10.749055,5.424384,0.099712946,1.2998942,2.5000753,3.7002566,4.900438,6.1006193,5.391751,4.6846952,3.97764,3.2705846,2.561716,2.465629,2.3677292,2.269829,2.1719291,2.0758421,2.5472124,3.0203958,3.491766,3.9649491,4.4381323,6.6644506,8.892582,11.120712,13.347031,15.575162,15.687565,15.799969,15.912373,16.024776,16.13718,14.726695,13.318023,11.907538,10.497053,9.088382,10.352016,11.617464,12.882912,14.14836,15.411995,12.84484,10.277685,7.71053,5.143375,2.5744069,10.46442,18.354433,26.244446,34.13446,42.02447,47.38178,52.739082,58.098198,63.4555,68.812805,58.038372,47.262123,36.487686,25.711435,14.936998,17.794228,20.653269,23.510498,26.367727,29.224957,28.815228,28.405499,27.995768,27.584227,27.174496,26.545399,25.914488,25.285389,24.654478,24.025381,20.676838,17.330109,13.981567,10.634838,7.28811,10.384649,13.483003,16.579542,19.677896,22.774435,21.965855,21.15546,20.345066,19.534672,18.724277,16.229641,13.735004,11.240368,8.745731,6.249282,6.4178877,6.58468,6.7532854,6.9200783,7.0868707,5.924762,4.762653,3.6005437,2.4366217,1.2745126,1.1004683,0.9246109,0.7505665,0.5747091,0.40066472,1.6425442,2.8844235,4.1281157,5.369995,6.6118746,7.851941,9.092008,10.332074,11.57214,12.812206,11.137029,9.461852,7.7866745,6.11331,4.4381323,4.655688,4.8732433,5.090799,5.3083544,5.524097,6.378002,7.230095,8.082188,8.934279,9.788185,12.32452,14.862667,17.400814,19.93715,22.475298,18.555672,14.636047,10.714609,6.794984,2.8753586,7.036108,11.195044,15.355793,19.514729,23.675478,21.04487,18.41426,15.785465,13.154857,10.524248,13.189302,15.854358,18.519413,21.184467,23.849524,22.292189,20.734854,19.177519,17.620184,16.062849,13.281764,10.502492,7.723221,4.942136,2.1628644,1.7694515,1.3778516,0.98443866,0.59283876,0.19942589,0.2030518,0.20486477,0.20667773,0.21030366,0.21211663,0.38434806,0.55839247,0.7306239,0.90285534,1.0750868,0.9644961,0.8557183,0.7451276,0.6345369,0.52575916,0.46230546,0.40066472,0.33721104,0.2755703,0.21211663,0.21211663,0.21211663,0.21211663,0.21211663,0.21211663,0.19036107,0.16679256,0.14503701,0.12328146,0.099712946,0.10333887,0.10515183,0.10696479,0.11059072,0.11240368,0.09064813,0.06707962,0.045324065,0.02175555,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.032633327,0.065266654,0.09789998,0.13053331,0.16316663,0.23568514,0.30820364,0.38072214,0.45324063,0.52575916,0.5402629,0.55476654,0.56927025,0.5855869,0.6000906,0.48043507,0.36077955,0.23931105,0.11965553,0.0,0.03988518,0.07977036,0.11965553,0.15954071,0.19942589,1.0442665,1.889107,2.7357605,3.5806012,4.4254417,3.540716,2.6541772,1.7694515,0.88472575,0.0,0.0,0.0,0.0,0.0,0.0,0.018129626,0.034446288,0.052575916,0.07070554,0.0870222,0.13053331,0.17223145,0.21574254,0.2574407,0.2991388,0.35534066,0.40972954,0.46411842,0.52032024,0.5747091,0.48224804,0.38978696,0.29732585,0.20486477,0.11240368,0.13053331,0.14684997,0.16497959,0.18310922,0.19942589,0.15954071,0.11965553,0.07977036,0.03988518,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.059827764,0.08339628,0.10515183,0.12690738,0.15047589,0.15410182,0.15954071,0.16497959,0.17041849,0.17585737,0.18492219,0.19579996,0.20486477,0.21574254,0.22480737,0.2229944,0.21936847,0.21755551,0.21574254,0.21211663,0.17041849,0.12690738,0.08520924,0.04169814,0.0,0.018129626,0.034446288,0.052575916,0.07070554,0.0870222,0.09789998,0.10696479,0.11784257,0.12690738,0.13778515,0.24293698,0.3480888,0.45324063,0.55839247,0.66173136,0.56927025,0.47680917,0.38434806,0.291887,0.19942589,0.17041849,0.13959812,0.11059072,0.07977036,0.05076295,0.045324065,0.03988518,0.034446288,0.030820364,0.025381476,0.038072214,0.05076295,0.06164073,0.07433146,0.0870222,0.10333887,0.11784257,0.13234627,0.14684997,0.16316663,0.291887,0.4224203,0.5529536,0.68167394,0.8122072,0.73787576,0.66173136,0.5873999,0.51306844,0.43692398,0.40429065,0.37165734,0.34083697,0.30820364,0.2755703,0.25925365,0.24474995,0.23024625,0.21574254,0.19942589,0.44780177,0.69436467,0.94274056,1.1893034,1.4376793,1.1566701,0.8774739,0.5982776,0.31726846,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.034446288,0.032633327,0.030820364,0.027194439,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.027194439,0.054388877,0.08339628,0.11059072,0.13778515,0.17223145,0.20667773,0.24293698,0.27738327,0.31182957,0.2574407,0.2030518,0.14684997,0.092461094,0.038072214,0.047137026,0.058014803,0.06707962,0.07795739,0.0870222,0.08339628,0.07795739,0.072518505,0.06707962,0.06164073,0.058014803,0.052575916,0.047137026,0.04169814,0.038072214,0.04169814,0.047137026,0.052575916,0.058014803,0.06164073,0.12509441,0.18673515,0.25018883,0.31182957,0.37528324,0.54570174,0.71430725,0.88472575,1.0551442,1.2255627,1.0732739,0.91917205,0.7668832,0.61459434,0.46230546,0.38072214,0.29732585,0.21574254,0.13234627,0.05076295,0.054388877,0.059827764,0.065266654,0.07070554,0.07433146,2.2118144,1.9996977,1.7875811,1.5754645,1.3633479,1.1494182,1.2346275,1.3198367,1.405046,1.4902552,1.5754645,1.7767034,1.9797552,2.182807,2.3858588,2.5870976,2.9279346,3.2669585,3.6077955,3.9468195,4.2876563,4.953014,5.618371,6.281915,6.947273,7.61263,8.252605,8.892582,9.5325575,10.172533,10.812509,10.620335,10.428161,10.234174,10.042,9.849826,9.757364,9.664904,9.572442,9.479981,9.38752,9.670342,9.953164,10.234174,10.516996,10.799818,12.416981,14.034143,15.653119,17.27028,18.887444,18.196705,17.50778,16.817041,16.128115,15.437376,12.618219,9.79725,6.978093,4.157123,1.3379664,1.84197,2.3477864,2.8517902,3.3576066,3.8616104,4.2223897,4.5831695,4.942136,5.3029156,5.661882,5.130684,4.597673,4.064662,3.531651,3.000453,3.6567454,4.314851,4.972956,5.6292486,6.2873545,5.6455655,5.0019636,4.360175,3.7183862,3.0747845,2.770207,2.465629,2.1592383,1.8546607,1.550083,2.572594,3.5951047,4.6176157,5.6401267,6.6626377,6.5701766,6.4777155,6.3852544,6.2927933,6.200332,5.1125546,4.024777,2.9369993,1.8492218,0.76325727,1.5301404,2.2970235,3.0657198,3.832603,4.599486,4.3728657,4.1444325,3.917812,3.6893787,3.4627585,2.8608549,2.2571385,1.6552348,1.0533313,0.44961473,1.2273756,2.0051367,2.7828975,3.5606585,4.3384194,5.710832,7.083245,8.455658,9.82807,11.200482,11.9873085,12.775948,13.562773,14.349599,15.138238,14.079468,13.022511,11.965553,10.906783,9.849826,9.168152,8.484665,7.802991,7.119504,6.43783,7.5346723,8.631515,9.73017,10.827013,11.925668,14.608852,17.29385,19.980661,22.665659,25.348843,22.885027,20.419397,17.955582,15.489952,13.024323,15.105604,17.185072,19.26454,21.345821,23.42529,22.85602,22.284937,21.715666,21.144583,20.575312,18.042604,15.509895,12.977186,10.444477,7.911769,11.421664,14.93156,18.443268,21.953163,25.46306,20.399454,15.337664,10.274059,5.2122674,0.15047589,0.96268314,1.7748904,2.5870976,3.3993049,4.213325,3.8579843,3.5026438,3.147303,2.7919624,2.4366217,2.2607644,2.0830941,1.9054236,1.7277533,1.550083,2.3024626,3.054842,3.8072214,4.559601,5.3119802,6.6100616,7.9081426,9.2044115,10.502492,11.800573,13.77489,15.749206,17.725336,19.699652,21.675781,18.709774,15.74558,12.779573,9.815379,6.849373,9.848013,12.84484,15.84348,18.840307,21.837133,18.017221,14.19731,10.377398,6.5574856,2.7375734,8.03505,13.332527,18.630003,23.92748,29.224957,35.05363,40.88412,46.714607,52.545094,58.375584,50.012386,41.64919,33.287807,24.92461,16.563227,20.067682,23.57214,27.07841,30.582867,34.087322,31.810242,29.533161,27.254267,24.977186,22.700104,22.741802,22.785315,22.827011,22.870523,22.912222,19.52198,16.13174,12.741501,9.353074,5.962834,8.890768,11.81689,14.744824,17.67276,20.600695,20.985043,21.36939,21.75555,22.139898,22.524246,19.670645,16.815228,13.959812,11.104396,8.2507925,7.6579537,7.065115,6.472276,5.8794374,5.2865987,4.499773,3.7129474,2.9243085,2.137483,1.3506571,1.2001812,1.0497054,0.89922947,0.7505665,0.6000906,2.132044,3.6658103,5.197764,6.7297173,8.26167,8.997733,9.731983,10.468046,11.202296,11.938358,10.411844,8.887142,7.362441,5.8377395,4.313038,4.5704784,4.8279195,5.08536,5.3428006,5.600241,7.3968873,9.195346,10.991992,12.790451,14.587097,17.812357,21.037619,24.262878,27.488138,30.7134,25.394167,20.07856,14.759329,9.441909,4.12449,6.8656893,9.605076,12.344462,15.085662,17.825048,16.817041,15.810846,14.802839,13.794832,12.786825,14.996826,17.206827,19.41683,21.626831,23.836832,22.620335,21.402023,20.185526,18.967215,17.750717,14.830034,11.909351,8.990481,6.069799,3.150929,2.5544643,1.9598125,1.3651608,0.7705091,0.17585737,0.18492219,0.19579996,0.20486477,0.21574254,0.22480737,0.41516843,0.6055295,0.79589057,0.98443866,1.1747998,1.0478923,0.91917205,0.79226464,0.6653573,0.53663695,0.4749962,0.41335547,0.34990177,0.28826106,0.22480737,0.22480737,0.22480737,0.22480737,0.22480737,0.22480737,0.19761293,0.17041849,0.14322405,0.11421664,0.0870222,0.08520924,0.08339628,0.07977036,0.07795739,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.04169814,0.08520924,0.12690738,0.17041849,0.21211663,0.32814622,0.44236287,0.55839247,0.6726091,0.7868258,0.7106813,0.6327239,0.55476654,0.47680917,0.40066472,0.3208944,0.23931105,0.15954071,0.07977036,0.0,0.059827764,0.11965553,0.1794833,0.23931105,0.2991388,1.5682126,2.8354735,4.102734,5.369995,6.637256,5.3101673,3.9830787,2.6541772,1.3270886,0.0,0.0,0.0,0.0,0.0,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.11965553,0.13959812,0.15954071,0.1794833,0.19942589,0.33177215,0.46411842,0.5982776,0.7306239,0.8629702,0.70524246,0.5475147,0.38978696,0.23205921,0.07433146,0.11965553,0.16497959,0.21030366,0.25562772,0.2991388,0.23931105,0.1794833,0.11965553,0.059827764,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.03988518,0.054388877,0.07070554,0.08520924,0.099712946,0.10696479,0.11421664,0.12328146,0.13053331,0.13778515,0.15228885,0.16679256,0.18310922,0.19761293,0.21211663,0.22662032,0.24293698,0.2574407,0.27194437,0.28826106,0.23024625,0.17223145,0.11421664,0.058014803,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.10333887,0.10515183,0.10696479,0.11059072,0.11240368,0.21936847,0.32814622,0.43511102,0.5420758,0.6508536,0.58014804,0.5094425,0.4405499,0.36984438,0.2991388,0.25562772,0.21030366,0.16497959,0.11965553,0.07433146,0.06707962,0.059827764,0.052575916,0.045324065,0.038072214,0.05076295,0.06164073,0.07433146,0.0870222,0.099712946,0.11059072,0.11965553,0.13053331,0.13959812,0.15047589,0.23205921,0.3154555,0.39703882,0.48043507,0.5620184,0.5493277,0.53663695,0.52575916,0.51306844,0.50037766,0.45686656,0.41516843,0.37165734,0.32995918,0.28826106,0.26469254,0.24293698,0.21936847,0.19761293,0.17585737,0.34083697,0.5058166,0.67079616,0.83577573,1.0007553,0.80495536,0.6091554,0.41516843,0.21936847,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.027194439,0.030820364,0.032633327,0.034446288,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.13959812,0.16679256,0.19579996,0.2229944,0.25018883,0.20486477,0.15954071,0.11421664,0.07070554,0.025381476,0.03988518,0.054388877,0.07070554,0.08520924,0.099712946,0.092461094,0.08520924,0.07795739,0.07070554,0.06164073,0.054388877,0.047137026,0.03988518,0.032633327,0.025381476,0.032633327,0.03988518,0.047137026,0.054388877,0.06164073,0.099712946,0.13778515,0.17585737,0.21211663,0.25018883,0.38072214,0.5094425,0.6399758,0.7705091,0.89922947,0.81583315,0.7306239,0.64541465,0.56020546,0.4749962,0.39522585,0.3154555,0.23568514,0.15410182,0.07433146,0.07070554,0.065266654,0.059827764,0.054388877,0.05076295,1.887294,1.8002719,1.7132497,1.6244144,1.5373923,1.4503701,1.5682126,1.6842422,1.8020848,1.9199274,2.03777,2.182807,2.327844,2.472881,2.617918,2.762955,3.207131,3.6531196,4.0972953,4.5432844,4.98746,5.632875,6.2782893,6.921891,7.567306,8.212721,8.745731,9.27693,9.80994,10.342952,10.874149,10.834265,10.794379,10.754494,10.714609,10.674724,10.785315,10.8959055,11.004683,11.115273,11.225864,11.5231905,11.820516,12.117842,12.415168,12.712494,14.126604,15.542528,16.958452,18.372562,19.786674,18.59193,17.397188,16.202446,15.007704,13.812962,11.327391,8.841819,6.35806,3.872488,1.3869164,1.7277533,2.0667772,2.4076142,2.7466383,3.0874753,3.5806012,4.071914,4.5650396,5.0581656,5.5494785,4.7771564,4.004834,3.2325122,2.4601903,1.6878681,2.4855716,3.2832751,4.079166,4.876869,5.674573,5.185073,4.695573,4.2042603,3.7147603,3.2252605,2.9224956,2.619731,2.3169663,2.0142014,1.7132497,2.5417736,3.3721104,4.2024474,5.032784,5.863121,6.0226617,6.1822023,6.341743,6.5030966,6.6626377,5.4370747,4.213325,2.9877625,1.7621996,0.53663695,1.1276628,1.7168756,2.3079014,2.8971143,3.48814,3.529838,3.5733492,3.6150475,3.6567454,3.7002566,3.0167696,2.335096,1.651609,0.969935,0.28826106,1.2817645,2.277081,3.2723975,4.267714,5.2630305,6.929143,8.597069,10.264994,11.9329195,13.600845,14.68681,15.774588,16.862366,17.950142,19.03792,17.22677,15.417434,13.608097,11.7969475,9.987611,9.215289,8.442966,7.6706448,6.8983226,6.1241875,6.093367,6.060734,6.0281005,5.995467,5.962834,7.817495,9.672155,11.526816,13.383289,15.23795,13.754947,12.271944,10.78894,9.30775,7.8247466,12.077957,16.329353,20.582563,24.835773,29.087172,28.690132,28.293095,27.894243,27.497204,27.100164,22.553255,18.004532,13.457622,8.910711,4.361988,8.330563,12.297325,16.2659,20.232662,24.199425,19.400513,14.599788,9.799063,5.0001507,0.19942589,0.62547207,1.0497054,1.4757515,1.8999848,2.324218,2.322405,2.3205922,2.3169663,2.3151531,2.3133402,2.0558996,1.7966459,1.5392052,1.2817645,1.0243238,2.0577126,3.0892882,4.122677,5.1542525,6.187641,6.5556726,6.921891,7.2899227,7.6579537,8.024173,11.862214,15.700256,19.538298,23.374527,27.212568,22.692852,18.173138,13.651608,9.131892,4.612177,9.342196,14.072216,18.802235,23.532255,28.262274,23.189604,18.116936,13.044266,7.9715962,2.9007401,5.6056805,8.31062,11.015561,13.720501,16.425442,22.727299,29.029158,35.33283,41.634686,47.936543,41.988213,36.03807,30.087927,24.137783,18.187641,22.339325,26.492823,30.644506,34.798004,38.949688,34.805256,30.660824,26.514578,22.370146,18.225714,18.94002,19.654327,20.370447,21.084755,21.800875,18.367125,14.935185,11.503247,8.069496,4.6375585,7.3950744,10.152591,12.910107,15.667623,18.425138,20.004229,21.585133,23.164223,24.745127,26.324217,23.109835,19.89545,16.679256,13.464873,10.25049,8.898021,7.5455503,6.19308,4.84061,3.48814,3.0747845,2.663242,2.2498865,1.8383441,1.4249886,1.2998942,1.1747998,1.0497054,0.9246109,0.7995165,2.6233568,4.445384,6.2674117,8.089439,9.91328,10.141713,10.371959,10.602205,10.832452,11.062697,9.686659,8.312433,6.9382076,5.562169,4.1879435,4.4852695,4.782595,5.0799212,5.377247,5.674573,8.417585,11.160598,13.901797,16.64481,19.387821,23.300196,27.212568,31.12494,35.037315,38.949688,32.234474,25.521074,18.804049,12.090648,5.375434,6.695271,8.015107,9.334945,10.654781,11.974618,12.589212,13.20562,13.820213,14.434808,15.049402,16.80435,18.559298,20.314245,22.069193,23.82414,22.946667,22.069193,21.19172,20.314245,19.436771,16.376492,13.318023,10.257742,7.1974616,4.137181,3.339477,2.5417736,1.745883,0.9481794,0.15047589,0.16679256,0.18492219,0.2030518,0.21936847,0.2374981,0.44417584,0.6526665,0.85934424,1.067835,1.2745126,1.1294757,0.98443866,0.83940166,0.69436467,0.5493277,0.48768693,0.42423326,0.36259252,0.2991388,0.2374981,0.2374981,0.2374981,0.2374981,0.2374981,0.2374981,0.20486477,0.17223145,0.13959812,0.10696479,0.07433146,0.06707962,0.059827764,0.052575916,0.045324065,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.052575916,0.10515183,0.15772775,0.21030366,0.26287958,0.42060733,0.57833505,0.73424983,0.8919776,1.0497054,0.8792868,0.7106813,0.5402629,0.36984438,0.19942589,0.15954071,0.11965553,0.07977036,0.03988518,0.0,0.07977036,0.15954071,0.23931105,0.3208944,0.40066472,2.0903459,3.780027,5.469708,7.159389,8.8508835,7.079619,5.3101673,3.540716,1.7694515,0.0,0.0,0.0,0.0,0.0,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.11059072,0.10696479,0.10515183,0.10333887,0.099712946,0.3100166,0.52032024,0.7306239,0.93911463,1.1494182,0.92823684,0.70524246,0.48224804,0.25925365,0.038072214,0.11059072,0.18310922,0.25562772,0.32814622,0.40066472,0.3208944,0.23931105,0.15954071,0.07977036,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.01994259,0.027194439,0.034446288,0.04169814,0.05076295,0.059827764,0.07070554,0.07977036,0.09064813,0.099712946,0.11965553,0.13959812,0.15954071,0.1794833,0.19942589,0.23205921,0.26469254,0.29732585,0.32995918,0.36259252,0.29007402,0.21755551,0.14503701,0.072518505,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.10696479,0.10333887,0.09789998,0.092461094,0.0870222,0.19761293,0.30820364,0.4169814,0.5275721,0.63816285,0.58921283,0.5420758,0.4949388,0.44780177,0.40066472,0.34083697,0.27919623,0.21936847,0.15954071,0.099712946,0.09064813,0.07977036,0.07070554,0.059827764,0.05076295,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.11784257,0.12328146,0.12690738,0.13234627,0.13778515,0.17223145,0.20667773,0.24293698,0.27738327,0.31182957,0.36259252,0.41335547,0.46230546,0.51306844,0.5620184,0.5094425,0.45686656,0.40429065,0.35171473,0.2991388,0.27013144,0.23931105,0.21030366,0.1794833,0.15047589,0.23205921,0.3154555,0.39703882,0.48043507,0.5620184,0.45324063,0.34264994,0.23205921,0.12328146,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.01994259,0.027194439,0.034446288,0.04169814,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.018129626,0.034446288,0.052575916,0.07070554,0.0870222,0.10696479,0.12690738,0.14684997,0.16679256,0.18673515,0.15228885,0.11784257,0.08339628,0.047137026,0.012690738,0.032633327,0.052575916,0.072518505,0.092461094,0.11240368,0.10333887,0.092461094,0.08339628,0.072518505,0.06164073,0.052575916,0.04169814,0.032633327,0.02175555,0.012690738,0.02175555,0.032633327,0.04169814,0.052575916,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.21574254,0.3045777,0.39522585,0.48587397,0.5747091,0.55839247,0.5402629,0.52213323,0.5058166,0.48768693,0.40972954,0.33177215,0.25562772,0.17767033,0.099712946,0.08520924,0.07070554,0.054388877,0.03988518,0.025381476,1.5627737,1.6008459,1.6371052,1.6751775,1.7132497,1.7495089,1.8999848,2.0504606,2.1991236,2.3495996,2.5000753,2.5870976,2.6741197,2.762955,2.8499773,2.9369993,3.48814,4.0374675,4.5867953,5.137936,5.6872635,6.3127356,6.9382076,7.5618668,8.187339,8.812811,9.237044,9.663091,10.087324,10.51337,10.937603,11.050007,11.162411,11.274815,11.3872175,11.499621,11.813264,12.125093,12.436923,12.750566,13.062395,13.374225,13.687867,13.999697,14.313339,14.625169,15.838041,17.0491,18.261972,19.474844,20.687716,18.987158,17.288412,15.5878525,13.887294,12.186734,10.038374,7.8882003,5.7380266,3.587853,1.4376793,1.6117238,1.7875811,1.9616255,2.137483,2.3133402,2.9369993,3.5624714,4.1879435,4.8134155,5.4370747,4.4254417,3.4119956,2.4003625,1.3869164,0.37528324,1.3125849,2.2498865,3.1871881,4.12449,5.0617914,4.7245803,4.3873696,4.0501585,3.7129474,3.3757362,3.0747845,2.7756457,2.474694,2.175555,1.8746033,2.5127661,3.149116,3.787279,4.4254417,5.0617914,5.475147,5.8866897,6.300045,6.7134004,7.124943,5.763408,4.40006,3.0367124,1.6751775,0.31182957,0.72518504,1.1367276,1.550083,1.9616255,2.374981,2.6868105,3.000453,3.3122826,3.6241121,3.9377546,3.1744974,2.4130533,1.649796,0.8883517,0.12509441,1.3379664,2.5508385,3.7618973,4.974769,6.187641,8.149267,10.112705,12.07433,14.037769,15.999394,17.388124,18.77504,20.161957,21.550686,22.937603,20.375887,17.812357,15.250641,12.687112,10.125396,9.262425,8.399456,7.5382986,6.6753283,5.812358,4.650249,3.48814,2.324218,1.162109,0.0,1.0243238,2.0504606,3.0747845,4.100921,5.125245,4.6248674,4.12449,3.6241121,3.1255474,2.6251698,9.050309,15.475449,21.900587,28.325727,34.750866,34.524246,34.29944,34.07463,33.849823,33.625015,27.062092,20.50098,13.938056,7.3751316,0.8122072,5.237649,9.663091,14.088532,18.512161,22.937603,18.399757,13.861912,9.324066,4.788034,0.25018883,0.28826106,0.3245203,0.36259252,0.40066472,0.43692398,0.7868258,1.1367276,1.4866294,1.8383441,2.1882458,1.8492218,1.5120108,1.1747998,0.8375887,0.50037766,1.8129625,3.1255474,4.4381323,5.750717,7.063302,6.4994707,5.9374523,5.375434,4.8116026,4.249584,9.949538,15.649493,21.349447,27.049402,32.749355,26.675932,20.600695,14.525456,8.450218,2.374981,8.838193,15.299591,21.762802,28.224201,34.687412,28.361986,22.038374,15.712947,9.38752,3.0620937,3.1744974,3.2869012,3.3993049,3.5117085,3.6241121,10.399154,17.174194,23.951048,30.724277,37.499317,33.962227,30.425138,26.888048,23.349146,19.812056,24.61278,29.411692,34.212418,39.01314,43.812054,37.80027,31.788486,25.774889,19.763105,13.749508,15.138238,16.525154,17.912071,19.3008,20.687716,17.212267,13.736817,10.263181,6.787732,3.3122826,5.89938,8.488291,11.075388,13.662486,16.249584,19.025229,21.799063,24.574707,27.350353,30.124186,26.550837,22.975676,19.400513,15.825351,12.250188,10.138086,8.024173,5.9120708,3.7999697,1.6878681,1.649796,1.6117238,1.5754645,1.5373923,1.49932,1.3996071,1.2998942,1.2001812,1.1004683,1.0007553,3.1128569,5.224958,7.3370595,9.449161,11.563075,11.287505,11.011934,10.738177,10.462607,10.1870365,8.963287,7.7377243,6.5121617,5.2865987,4.062849,4.40006,4.7372713,5.0744824,5.411693,5.750717,9.438283,13.124036,16.813416,20.499168,24.186733,28.788033,33.38752,37.987003,42.588303,47.18779,39.074783,30.963589,22.85058,14.737573,6.624565,6.5248523,6.4251394,6.3254266,6.2257137,6.1241875,8.363196,10.600392,12.837588,15.074784,17.31198,18.611874,19.911768,21.211662,22.513369,23.813263,23.274813,22.738176,22.199726,21.66309,21.12464,17.92476,14.724882,11.525003,8.325124,5.125245,4.12449,3.1255474,2.124792,1.1258497,0.12509441,0.15047589,0.17585737,0.19942589,0.22480737,0.25018883,0.4749962,0.69980353,0.9246109,1.1494182,1.3742256,1.2128719,1.0497054,0.8883517,0.72518504,0.5620184,0.50037766,0.43692398,0.37528324,0.31182957,0.25018883,0.25018883,0.25018883,0.25018883,0.25018883,0.25018883,0.21211663,0.17585737,0.13778515,0.099712946,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06164073,0.12509441,0.18673515,0.25018883,0.31182957,0.51306844,0.7124943,0.9119202,1.1131591,1.3125849,1.0497054,0.7868258,0.52575916,0.26287958,0.0,0.0,0.0,0.0,0.0,0.0,0.099712946,0.19942589,0.2991388,0.40066472,0.50037766,2.612479,4.7245803,6.836682,8.950596,11.062697,8.849071,6.637256,4.4254417,2.2118144,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.28826106,0.5747091,0.8629702,1.1494182,1.4376793,1.1494182,0.8629702,0.5747091,0.28826106,0.0,0.099712946,0.19942589,0.2991388,0.40066472,0.50037766,0.40066472,0.2991388,0.19942589,0.099712946,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.0870222,0.11240368,0.13778515,0.16316663,0.18673515,0.2374981,0.28826106,0.33721104,0.387974,0.43692398,0.34990177,0.26287958,0.17585737,0.0870222,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.17585737,0.28826106,0.40066472,0.51306844,0.62547207,0.6000906,0.5747091,0.5493277,0.52575916,0.50037766,0.42423326,0.34990177,0.2755703,0.19942589,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.17585737,0.28826106,0.40066472,0.51306844,0.62547207,0.5620184,0.50037766,0.43692398,0.37528324,0.31182957,0.2755703,0.2374981,0.19942589,0.16316663,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,0.2991388,0.34990177,0.40066472,0.44961473,0.50037766,0.42423326,0.34990177,0.2755703,0.19942589,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,1.9126755,1.983381,2.0522738,2.1229792,2.1918716,2.2625773,2.3205922,2.3767939,2.4348087,2.4928236,2.5508385,2.6704938,2.7901495,2.909805,3.0294604,3.149116,3.682127,4.215138,4.748149,5.279347,5.812358,6.397945,6.981719,7.567306,8.152893,8.736667,8.943344,9.14821,9.353074,9.557939,9.762803,9.904215,10.047439,10.190662,10.332074,10.475298,11.3056345,12.134158,12.964496,13.794832,14.625169,14.462003,14.300649,14.137483,13.974316,13.812962,14.875358,15.937754,17.00015,18.062546,19.124943,17.330109,15.535276,13.740443,11.94561,10.150778,8.437528,6.7242785,5.0128417,3.299592,1.5881553,1.9797552,2.373168,2.764768,3.1581807,3.5497808,3.7093215,3.870675,4.0302157,4.1897564,4.349297,3.8108473,3.2705846,2.7303216,2.1900587,1.649796,2.6396735,3.6295512,4.6194286,5.6093063,6.599184,6.341743,6.0843024,5.826862,5.569421,5.3119802,4.6792564,4.0483456,3.4156215,2.7828975,2.1501737,3.0693457,3.9903307,4.9095025,5.8304877,6.7496595,7.3733187,7.995165,8.617011,9.24067,9.862516,8.044115,6.2275267,4.409125,2.5925364,0.774135,1.114972,1.455809,1.794833,2.13567,2.474694,2.7883365,3.100166,3.4119956,3.7256382,4.0374675,4.229642,4.421816,4.615803,4.8079767,5.0001507,5.3446136,5.6890764,6.035352,6.379815,6.7242785,8.05318,9.380268,10.707357,12.034446,13.363347,14.3604765,15.357606,16.354736,17.351866,18.350807,19.268166,20.185526,21.102884,22.020243,22.937603,20.332375,17.727148,15.121921,12.516694,9.91328,8.000604,6.0879283,4.175253,2.2625773,0.34990177,1.2545701,2.1592383,3.0657198,3.9703882,4.8750563,4.3329806,3.7909048,3.247016,2.70494,2.1628644,7.2953615,12.427858,17.560356,22.692852,27.82535,27.64768,27.470009,27.29234,27.114668,26.936998,21.690285,16.443571,11.195044,5.9483304,0.69980353,4.2405195,7.7794223,11.320138,14.860854,18.399757,14.770206,11.1406555,7.509291,3.87974,0.25018883,0.28826106,0.3245203,0.36259252,0.40066472,0.43692398,0.72518504,1.0116332,1.2998942,1.5881553,1.8746033,1.5881553,1.2998942,1.0116332,0.72518504,0.43692398,1.5446441,2.6523643,3.7600844,4.8678045,5.975525,5.5929894,5.2104545,4.8279195,4.445384,4.062849,8.519112,12.977186,17.43526,21.893335,26.349598,21.474543,16.599485,11.724429,6.849373,1.9743162,7.130382,12.284635,17.4407,22.594954,27.749205,22.725487,17.699953,12.674421,7.650702,2.6251698,2.7248828,2.8245957,2.9243085,3.0258346,3.1255474,8.562622,13.999697,19.438585,24.87566,30.312735,28.148058,25.98338,23.816889,21.652212,19.487535,23.129776,26.772018,30.416073,34.058315,37.700558,35.47968,33.260612,31.039732,28.820665,26.599787,25.192928,23.784256,22.377398,20.97054,19.561867,18.069798,16.57773,15.085662,13.591781,12.099712,12.311829,12.525759,12.737875,12.949992,13.162108,15.428311,17.692701,19.957092,22.223295,24.487686,21.626831,18.767788,15.906934,13.047892,10.1870365,8.600695,7.0125394,5.424384,3.8380418,2.2498865,2.2118144,2.175555,2.137483,2.0994108,2.0631514,1.9308052,1.7966459,1.6642996,1.5319533,1.3996071,3.5008307,5.600241,7.699652,9.800876,11.900287,11.537694,11.175101,10.812509,10.449916,10.087324,9.518054,8.94697,8.3777,7.806617,7.2373466,7.9226465,8.607946,9.293246,9.976733,10.662033,12.462305,14.262577,16.062849,17.863121,19.663393,23.485117,27.306843,31.13038,34.952106,38.775642,32.74029,26.704939,20.669586,14.634234,8.600695,8.009668,7.420456,6.82943,6.240217,5.6491914,9.101072,12.549327,15.999394,19.449463,22.89953,22.34295,21.78456,21.22798,20.669586,20.113007,19.868258,19.621695,19.376944,19.132195,18.887444,16.05741,13.227375,10.397341,7.567306,4.7372713,3.8108473,2.8826106,1.9543737,1.0279498,0.099712946,0.11965553,0.13959812,0.15954071,0.1794833,0.19942589,0.40066472,0.6000906,0.7995165,1.0007553,1.2001812,1.0696479,0.93911463,0.8103943,0.67986095,0.5493277,0.49675176,0.44417584,0.39159992,0.34083697,0.28826106,0.27194437,0.2574407,0.24293698,0.22662032,0.21211663,0.19036107,0.16679256,0.14503701,0.12328146,0.099712946,0.0870222,0.07433146,0.06164073,0.05076295,0.038072214,0.032633327,0.027194439,0.02175555,0.018129626,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,0.42060733,0.58921283,0.75963134,0.9300498,1.1004683,1.1421664,1.1856775,1.2273756,1.2708868,1.3125849,1.1004683,0.8883517,0.6744221,0.46230546,0.25018883,0.28463513,0.3208944,0.35534066,0.38978696,0.42423326,2.1102884,3.7945306,5.480586,7.1648283,8.8508835,7.0868707,5.3246713,3.5624714,1.8002719,0.038072214,0.099712946,0.16316663,0.22480737,0.28826106,0.34990177,0.2991388,0.25018883,0.19942589,0.15047589,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.5855869,1.1693609,1.7549478,2.3405347,2.9243085,2.7031271,2.4801328,2.2571385,2.034144,1.8129625,1.5301404,1.2473183,0.9644961,0.68167394,0.40066472,0.3208944,0.23931105,0.15954071,0.07977036,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.072518505,0.09427405,0.11784257,0.13959812,0.16316663,0.23205921,0.30276474,0.37165734,0.44236287,0.51306844,0.4169814,0.32270733,0.22662032,0.13234627,0.038072214,0.052575916,0.06707962,0.08339628,0.09789998,0.11240368,0.10333887,0.092461094,0.08339628,0.072518505,0.06164073,0.15228885,0.24293698,0.33177215,0.4224203,0.51306844,0.52213323,0.533011,0.5420758,0.5529536,0.5620184,0.48224804,0.40247768,0.32270733,0.24293698,0.16316663,0.15228885,0.14322405,0.13234627,0.12328146,0.11240368,0.11240368,0.11240368,0.11240368,0.11240368,0.11240368,0.11059072,0.10696479,0.10515183,0.10333887,0.099712946,0.092461094,0.08520924,0.07795739,0.07070554,0.06164073,0.15228885,0.24293698,0.33177215,0.4224203,0.51306844,0.46230546,0.41335547,0.36259252,0.31182957,0.26287958,0.23205921,0.2030518,0.17223145,0.14322405,0.11240368,0.11784257,0.12328146,0.12690738,0.13234627,0.13778515,0.11059072,0.08339628,0.054388877,0.027194439,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.09064813,0.06707962,0.045324065,0.02175555,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.10333887,0.092461094,0.08339628,0.072518505,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.04169814,0.08520924,0.12690738,0.17041849,0.21211663,0.2520018,0.291887,0.33177215,0.37165734,0.41335547,0.35534066,0.29732585,0.23931105,0.18310922,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,2.2625773,2.3641033,2.467442,2.570781,2.6723068,2.7756457,2.7393866,2.70494,2.6704938,2.6342347,2.5997884,2.752077,2.904366,3.056655,3.2107568,3.3630457,3.877927,4.3928084,4.9076896,5.422571,5.9374523,6.4831543,7.027043,7.572745,8.116633,8.662335,8.647832,8.6333275,8.617011,8.602508,8.588004,8.760235,8.9324665,9.104698,9.27693,9.449161,10.798005,12.145037,13.492067,14.840912,16.187943,15.54978,14.91343,14.275268,13.637105,13.000754,13.912675,14.824595,15.738328,16.650248,17.562168,15.673061,13.782142,11.893035,10.002114,8.113008,6.836682,5.562169,4.2876563,3.0131438,1.7368182,2.3477864,2.956942,3.5679104,4.177066,4.788034,4.4816437,4.177066,3.872488,3.5679104,3.2633326,3.1944401,3.1273603,3.0602808,2.9932013,2.9243085,3.966762,5.009216,6.051669,7.0941224,8.138389,7.9607186,7.783048,7.605378,7.4277077,7.250037,6.285541,5.319232,4.3547363,3.39024,2.4257438,3.6277382,4.8297324,6.0317264,7.2355337,8.437528,9.269678,10.101828,10.93579,11.7679405,12.60009,10.328448,8.054993,5.7815375,3.5098956,1.2382535,1.504759,1.7730774,2.039583,2.3079014,2.5744069,2.8880494,3.199879,3.5117085,3.825351,4.137181,5.2847857,6.432391,7.5799966,8.727602,9.875207,9.353074,8.830941,8.306994,7.7848616,7.262728,7.95528,8.647832,9.340384,10.032935,10.725487,11.332829,11.940171,12.547514,13.154857,13.762199,18.160446,22.55688,26.955128,31.353374,35.74981,31.402325,27.05484,22.707355,18.359873,14.012388,11.350959,8.6877165,6.0244746,3.3630457,0.69980353,1.4848163,2.269829,3.054842,3.8398547,4.6248674,4.0392804,3.4555066,2.8699198,2.2843328,1.7005589,5.540414,9.380268,13.220123,17.059978,20.899832,20.769299,20.64058,20.510046,20.379513,20.250792,16.316664,12.384347,8.452031,4.519716,0.5873999,3.2415771,5.8975673,8.551744,11.207735,13.861912,11.1406555,8.417585,5.6945157,2.9732587,0.25018883,0.28826106,0.3245203,0.36259252,0.40066472,0.43692398,0.66173136,0.8883517,1.1131591,1.3379664,1.5627737,1.3252757,1.0877775,0.85027945,0.61278135,0.37528324,1.2781386,2.179181,3.0820365,3.9848917,4.8877473,4.6846952,4.4816437,4.2804046,4.077353,3.874301,7.0904965,10.304879,13.519262,16.735458,19.94984,16.274965,12.60009,8.925215,5.2503395,1.5754645,5.422571,9.269678,13.116784,16.965704,20.81281,17.087172,13.363347,9.637709,5.9120708,2.1882458,2.275268,2.3622901,2.4493124,2.5381477,2.6251698,6.7242785,10.825199,14.924308,19.025229,23.124338,22.332073,21.539808,20.747543,19.955278,19.163015,21.646772,24.132345,26.617916,29.101675,31.587248,33.159084,34.73274,36.304577,37.878227,39.450066,35.24762,31.045172,26.842724,22.640276,18.43783,18.92733,19.41683,19.908142,20.397642,20.887142,18.724277,16.563227,14.400362,12.237497,10.074633,11.829581,13.584529,15.339477,17.094423,18.849373,16.704638,14.559902,12.415168,10.270433,8.125698,7.063302,6.000906,4.936697,3.874301,2.811905,2.7756457,2.7375734,2.6995013,2.663242,2.6251698,2.4601903,2.2952106,2.1302311,1.9652514,1.8002719,3.8869917,5.975525,8.062244,10.150778,12.237497,11.787883,11.338268,10.88684,10.437225,9.987611,10.07282,10.15803,10.243238,10.326634,10.411844,11.445232,12.476809,13.510198,14.541773,15.575162,15.488139,15.399304,15.312282,15.22526,15.138238,18.182201,21.22798,24.271942,27.31772,30.361685,26.403988,22.448103,18.490406,14.532708,10.57501,9.494485,8.415772,7.3352466,6.2547207,5.1741953,9.837135,14.500074,19.163015,23.825954,28.487082,26.072214,23.657349,21.242483,18.827616,16.41275,16.459887,16.507025,16.554161,16.603111,16.650248,14.190058,11.729868,9.269678,6.8094873,4.349297,3.4953918,2.6396735,1.7857682,0.9300498,0.07433146,0.09064813,0.10515183,0.11965553,0.13415924,0.15047589,0.3245203,0.50037766,0.6744221,0.85027945,1.0243238,0.92823684,0.83033687,0.7324369,0.6345369,0.53663695,0.4949388,0.45324063,0.40972954,0.3680314,0.3245203,0.2955129,0.26469254,0.23568514,0.20486477,0.17585737,0.16679256,0.15954071,0.15228885,0.14503701,0.13778515,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.065266654,0.054388877,0.045324065,0.034446288,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.32814622,0.46774435,0.6073425,0.7469406,0.8883517,1.2346275,1.5827163,1.9308052,2.277081,2.6251698,2.1991236,1.7748904,1.3506571,0.9246109,0.50037766,0.46955732,0.4405499,0.40972954,0.38072214,0.34990177,1.6080978,2.864481,4.122677,5.3808727,6.637256,5.3246713,4.0120864,2.6995013,1.3869164,0.07433146,0.19942589,0.3245203,0.44961473,0.5747091,0.69980353,0.5747091,0.44961473,0.3245203,0.19942589,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.88291276,1.7658255,2.6469254,3.529838,4.4127507,4.255023,4.0972953,3.9395678,3.7818398,3.6241121,2.960568,2.2952106,1.6298534,0.9644961,0.2991388,0.23931105,0.1794833,0.11965553,0.059827764,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.058014803,0.07795739,0.09789998,0.11784257,0.13778515,0.22662032,0.31726846,0.40791658,0.49675176,0.5873999,0.48587397,0.3825351,0.27919623,0.17767033,0.07433146,0.07977036,0.08520924,0.09064813,0.09427405,0.099712946,0.092461094,0.08520924,0.07795739,0.07070554,0.06164073,0.13053331,0.19761293,0.26469254,0.33177215,0.40066472,0.44417584,0.4894999,0.53482395,0.58014804,0.62547207,0.5402629,0.4550536,0.36984438,0.28463513,0.19942589,0.19217403,0.18492219,0.17767033,0.17041849,0.16316663,0.15047589,0.13778515,0.12509441,0.11240368,0.099712946,0.09427405,0.09064813,0.08520924,0.07977036,0.07433146,0.072518505,0.07070554,0.06707962,0.065266654,0.06164073,0.13053331,0.19761293,0.26469254,0.33177215,0.40066472,0.36259252,0.3245203,0.28826106,0.25018883,0.21211663,0.19036107,0.16679256,0.14503701,0.12328146,0.099712946,0.11059072,0.11965553,0.13053331,0.13959812,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.05076295,0.06164073,0.07433146,0.0870222,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.092461094,0.08520924,0.07795739,0.07070554,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.034446288,0.07070554,0.10515183,0.13959812,0.17585737,0.20486477,0.23568514,0.26469254,0.2955129,0.3245203,0.28463513,0.24474995,0.20486477,0.16497959,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,2.612479,2.7466383,2.8826106,3.0167696,3.152742,3.2869012,3.159994,3.0330863,2.904366,2.7774587,2.6505513,2.8354735,3.0203958,3.2053177,3.39024,3.5751622,4.071914,4.5704784,5.06723,5.565795,6.0625467,6.5683637,7.072367,7.5781837,8.082188,8.588004,8.352319,8.116633,7.8827615,7.647076,7.413204,7.614443,7.817495,8.020547,8.221786,8.424837,10.290376,12.154101,14.01964,15.885179,17.750717,16.637558,15.524399,14.413053,13.299893,12.186734,12.949992,13.713249,14.474693,15.23795,15.999394,14.014201,12.03082,10.045626,8.0604315,6.0752378,5.237649,4.40006,3.5624714,2.7248828,1.887294,2.715818,3.5425289,4.36924,5.197764,6.0244746,5.2557783,4.4852695,3.7147603,2.9442513,2.175555,2.5798457,2.9841363,3.39024,3.7945306,4.2006345,5.295664,6.390693,7.4857225,8.580752,9.675781,9.577881,9.479981,9.382081,9.284182,9.188094,7.890013,6.591932,5.295664,3.9975824,2.6995013,4.1843176,5.669134,7.155763,8.640579,10.125396,11.16785,12.210303,13.252756,14.29521,15.337664,12.610968,9.882459,7.155763,4.4272547,1.7005589,1.8945459,2.0903459,2.2843328,2.4801328,2.6741197,2.9877625,3.299592,3.6132345,3.925064,4.2368937,6.33993,8.442966,10.546003,12.647227,14.750263,13.359721,11.970992,10.58045,9.189907,7.799365,7.85738,7.915395,7.9715962,8.029612,8.087626,8.3051815,8.5227375,8.740293,8.957849,9.175404,17.052727,24.930048,32.80737,40.684692,48.562016,42.472275,36.382534,30.292791,24.20305,18.11331,14.699501,11.287505,7.8755093,4.461701,1.0497054,1.7150626,2.38042,3.045777,3.7093215,4.3746786,3.7473936,3.1201086,2.4928236,1.8655385,1.2382535,3.785466,6.3326783,8.87989,11.427103,13.974316,13.892733,13.809336,13.727753,13.644357,13.562773,10.944855,8.326937,5.709019,3.092914,0.4749962,2.2444477,4.0157123,5.7851634,7.554615,9.324066,7.509291,5.6945157,3.87974,2.0649643,0.25018883,0.28826106,0.3245203,0.36259252,0.40066472,0.43692398,0.6000906,0.76325727,0.9246109,1.0877775,1.2491312,1.062396,0.87566096,0.6871128,0.50037766,0.31182957,1.0098201,1.7078108,2.4058013,3.101979,3.7999697,3.778214,3.7546456,3.73289,3.7093215,3.6875658,5.660069,7.6325727,9.605076,11.5775795,13.550082,11.075388,8.600695,6.1241875,3.6494937,1.1747998,3.7147603,6.2547207,8.794682,11.334642,13.874602,11.450671,9.024928,6.599184,4.175253,1.7495089,1.8256533,1.8999848,1.9743162,2.0504606,2.124792,4.8877473,7.650702,10.411844,13.174799,15.937754,16.517902,17.09805,17.678198,18.258347,18.836681,20.165583,21.492672,22.81976,24.146849,25.473938,30.840307,36.204865,41.57123,46.935787,52.300346,45.302307,38.306087,31.30805,24.310015,17.31198,19.78486,22.257742,24.730623,27.203503,29.674572,25.138538,20.600695,16.062849,11.525003,6.987158,8.232663,9.4781685,10.721861,11.967366,13.212872,11.782444,10.352016,8.921589,7.4929743,6.0625467,5.524097,4.98746,4.4508233,3.9123733,3.3757362,3.3376641,3.299592,3.2633326,3.2252605,3.1871881,2.9895754,2.7919624,2.5943494,2.3967366,2.1991236,4.274966,6.350808,8.424837,10.500679,12.574709,12.038072,11.499621,10.962985,10.424535,9.8878975,10.627586,11.367275,12.106964,12.848466,13.588155,14.967819,16.347483,17.727148,19.106813,20.48829,18.512161,16.537846,14.561715,12.5873995,10.613083,12.879286,15.147303,17.41532,19.681522,21.949537,20.069496,18.189453,16.309412,14.429369,12.549327,10.979301,9.409276,7.83925,6.2692246,4.699199,10.57501,16.449009,22.324821,28.200632,34.07463,29.80148,25.53014,21.256987,16.985647,12.712494,13.0515175,13.392355,13.7331915,14.072216,14.413053,12.322706,10.232361,8.1420145,6.051669,3.9631362,3.1799364,2.3967366,1.6153497,0.8321498,0.05076295,0.059827764,0.07070554,0.07977036,0.09064813,0.099712946,0.25018883,0.40066472,0.5493277,0.69980353,0.85027945,0.7850128,0.7197462,0.6544795,0.58921283,0.52575916,0.49312583,0.4604925,0.42785916,0.39522585,0.36259252,0.31726846,0.27194437,0.22662032,0.18310922,0.13778515,0.14503701,0.15228885,0.15954071,0.16679256,0.17585737,0.16316663,0.15047589,0.13778515,0.12509441,0.11240368,0.09789998,0.08339628,0.06707962,0.052575916,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.23568514,0.3444629,0.4550536,0.5656443,0.6744221,1.3270886,1.9797552,2.6324217,3.2850883,3.9377546,3.299592,2.663242,2.0250793,1.3869164,0.7505665,0.6544795,0.56020546,0.46411842,0.36984438,0.2755703,1.1059072,1.9344311,2.764768,3.5951047,4.4254417,3.5624714,2.6995013,1.8383441,0.97537386,0.11240368,0.2991388,0.48768693,0.6744221,0.8629702,1.0497054,0.85027945,0.6508536,0.44961473,0.25018883,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,1.1802386,2.3604772,3.540716,4.7209544,5.89938,5.806919,5.714458,5.621997,5.529536,5.4370747,4.3891826,3.343103,2.2952106,1.2473183,0.19942589,0.15954071,0.11965553,0.07977036,0.03988518,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.04169814,0.059827764,0.07795739,0.09427405,0.11240368,0.2229944,0.33177215,0.44236287,0.5529536,0.66173136,0.5529536,0.44236287,0.33177215,0.2229944,0.11240368,0.10696479,0.10333887,0.09789998,0.092461094,0.0870222,0.08339628,0.07795739,0.072518505,0.06707962,0.06164073,0.10696479,0.15228885,0.19761293,0.24293698,0.28826106,0.3680314,0.44780177,0.5275721,0.6073425,0.6871128,0.5982776,0.5076295,0.4169814,0.32814622,0.2374981,0.23205921,0.22662032,0.2229944,0.21755551,0.21211663,0.18673515,0.16316663,0.13778515,0.11240368,0.0870222,0.07977036,0.072518505,0.065266654,0.058014803,0.05076295,0.052575916,0.054388877,0.058014803,0.059827764,0.06164073,0.10696479,0.15228885,0.19761293,0.24293698,0.28826106,0.26287958,0.2374981,0.21211663,0.18673515,0.16316663,0.14684997,0.13234627,0.11784257,0.10333887,0.0870222,0.10333887,0.11784257,0.13234627,0.14684997,0.16316663,0.13053331,0.09789998,0.065266654,0.032633327,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.038072214,0.05076295,0.06164073,0.07433146,0.0870222,0.07070554,0.052575916,0.034446288,0.018129626,0.0,0.018129626,0.034446288,0.052575916,0.07070554,0.0870222,0.08339628,0.07795739,0.072518505,0.06707962,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.027194439,0.054388877,0.08339628,0.11059072,0.13778515,0.15772775,0.17767033,0.19761293,0.21755551,0.2374981,0.21574254,0.19217403,0.17041849,0.14684997,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,2.962381,3.1291735,3.2977788,3.4645715,3.633177,3.7999697,3.5806012,3.3594196,3.1400511,2.9206827,2.6995013,2.9170568,3.1346123,3.3521678,3.5697234,3.787279,4.267714,4.748149,5.2267714,5.7072062,6.187641,6.6517596,7.117691,7.5818095,8.047741,8.511859,8.056806,7.6017523,7.1466985,6.6916447,6.2365913,6.4704633,6.7025228,6.9345818,7.166641,7.400513,9.782746,12.164979,14.547212,16.929445,19.311678,17.725336,16.13718,14.5508375,12.962683,11.374527,11.9873085,12.60009,13.212872,13.825653,14.436621,12.357153,10.277685,8.198216,6.1169357,4.0374675,3.636803,3.2379513,2.8372865,2.4366217,2.03777,3.0820365,4.1281157,5.1723824,6.2166486,7.262728,6.0281005,4.7916603,3.5570326,2.322405,1.0877775,1.9652514,2.8427253,3.720199,4.597673,5.475147,6.622752,7.7703576,8.917963,10.065568,11.213174,11.195044,11.176914,11.160598,11.142468,11.124338,9.494485,7.8646317,6.2347784,4.604925,2.9750717,4.74271,6.510349,8.2779875,10.045626,11.813264,13.064208,14.316965,15.569723,16.82248,18.075237,14.893488,11.709926,8.528176,5.3446136,2.1628644,2.2843328,2.4076142,2.5308957,2.6523643,2.7756457,3.0874753,3.3993049,3.7129474,4.024777,4.3366065,7.3950744,10.451729,13.510198,16.566853,19.62532,17.368181,15.10923,12.852092,10.594954,8.337815,7.75948,7.1829576,6.604623,6.0281005,5.4497657,5.277534,5.105303,4.933071,4.76084,4.5867953,15.945006,27.301403,38.659615,50.017826,61.376034,53.542225,45.710224,37.878227,30.044416,22.212418,18.049856,13.887294,9.724731,5.562169,1.3996071,1.9453088,2.4891977,3.0348995,3.5806012,4.12449,3.4555066,2.7847104,2.1157274,1.4449311,0.774135,2.030518,3.2850883,4.539658,5.7942286,7.0506115,7.0143523,6.979906,6.94546,6.9092,6.874754,5.573047,4.269527,2.9678197,1.6642996,0.36259252,1.2473183,2.132044,3.0167696,3.9033084,4.788034,3.87974,2.9732587,2.0649643,1.1566701,0.25018883,0.28826106,0.3245203,0.36259252,0.40066472,0.43692398,0.53663695,0.63816285,0.73787576,0.8375887,0.93730164,0.7995165,0.66173136,0.52575916,0.387974,0.25018883,0.7433147,1.2346275,1.7277533,2.220879,2.712192,2.8699198,3.0276475,3.1853752,3.343103,3.5008307,4.229642,4.9602656,5.6890764,6.4197006,7.1503243,5.8758116,4.599486,3.3249733,2.0504606,0.774135,2.0069497,3.2397642,4.4725785,5.7053933,6.9382076,5.812358,4.688321,3.5624714,2.4366217,1.3125849,1.3742256,1.4376793,1.49932,1.5627737,1.6244144,3.049403,4.4743915,5.89938,7.324369,8.749357,10.701918,12.654479,14.607039,16.5596,18.512161,18.682579,18.852999,19.021603,19.192022,19.36244,28.519714,37.676987,46.836075,55.99335,65.15063,55.357,45.56519,35.771564,25.979753,16.187943,20.642391,25.096842,29.553102,34.007553,38.462,31.550987,24.63816,17.725336,10.812509,3.8996825,4.6357455,5.369995,6.104245,6.8403077,7.574558,6.8602505,6.14413,5.429823,4.7155156,3.9993954,3.9867048,3.975827,3.9631362,3.9504454,3.9377546,3.8996825,3.8616104,3.825351,3.787279,3.7492065,3.5207734,3.290527,3.0602808,2.8300345,2.5997884,4.6629395,6.7242785,8.78743,10.850581,12.91192,12.28826,11.662788,11.037316,10.411844,9.788185,11.182353,12.578335,13.972503,15.366671,16.762651,18.490406,20.218159,21.945911,23.671852,25.399607,21.537996,17.674572,13.812962,9.949538,6.0879283,7.5781837,9.066626,10.556881,12.047136,13.537392,13.735004,13.932617,14.13023,14.327844,14.525456,12.464118,10.4045925,8.345067,6.285541,4.2242026,11.312886,18.399757,25.488441,32.575314,39.66218,33.532555,27.40293,21.27149,15.141864,9.012237,9.644961,10.277685,10.910409,11.543133,12.175857,10.455356,8.734854,7.0143523,5.295664,3.5751622,2.864481,2.1556125,1.4449311,0.73424983,0.025381476,0.030820364,0.034446288,0.03988518,0.045324065,0.05076295,0.17585737,0.2991388,0.42423326,0.5493277,0.6744221,0.6417888,0.6091554,0.57833505,0.54570174,0.51306844,0.4894999,0.46774435,0.44417584,0.4224203,0.40066472,0.34083697,0.27919623,0.21936847,0.15954071,0.099712946,0.12328146,0.14503701,0.16679256,0.19036107,0.21211663,0.19942589,0.18673515,0.17585737,0.16316663,0.15047589,0.13053331,0.11059072,0.09064813,0.07070554,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.14322405,0.2229944,0.30276474,0.3825351,0.46230546,1.4195497,2.3767939,3.3358512,4.2930956,5.2503395,4.40006,3.5497808,2.6995013,1.8492218,1.0007553,0.83940166,0.67986095,0.52032024,0.36077955,0.19942589,0.60190356,1.0043813,1.4068589,1.8093367,2.2118144,1.8002719,1.3869164,0.97537386,0.5620184,0.15047589,0.40066472,0.6508536,0.89922947,1.1494182,1.3996071,1.1258497,0.85027945,0.5747091,0.2991388,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,1.4775645,2.955129,4.4326935,5.910258,7.3878226,7.360628,7.3316207,7.304426,7.2772317,7.250037,5.81961,4.3891826,2.960568,1.5301404,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.027194439,0.04169814,0.058014803,0.072518505,0.0870222,0.21755551,0.3480888,0.47680917,0.6073425,0.73787576,0.6200332,0.50219065,0.38434806,0.26831847,0.15047589,0.13415924,0.11965553,0.10515183,0.09064813,0.07433146,0.072518505,0.07070554,0.06707962,0.065266654,0.06164073,0.08520924,0.10696479,0.13053331,0.15228885,0.17585737,0.29007402,0.40429065,0.52032024,0.6345369,0.7505665,0.6544795,0.56020546,0.46411842,0.36984438,0.2755703,0.27194437,0.27013144,0.26831847,0.26469254,0.26287958,0.22480737,0.18673515,0.15047589,0.11240368,0.07433146,0.065266654,0.054388877,0.045324065,0.034446288,0.025381476,0.032633327,0.03988518,0.047137026,0.054388877,0.06164073,0.08520924,0.10696479,0.13053331,0.15228885,0.17585737,0.16316663,0.15047589,0.13778515,0.12509441,0.11240368,0.10515183,0.09789998,0.09064813,0.08339628,0.07433146,0.09427405,0.11421664,0.13415924,0.15410182,0.17585737,0.13959812,0.10515183,0.07070554,0.034446288,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.072518505,0.07070554,0.06707962,0.065266654,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.11059072,0.11965553,0.13053331,0.13959812,0.15047589,0.14503701,0.13959812,0.13415924,0.13053331,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,3.3122826,3.5117085,3.7129474,3.9123733,4.1117992,4.313038,3.9993954,3.6875658,3.3757362,3.0620937,2.7502642,3.000453,3.2506418,3.5008307,3.7492065,3.9993954,4.461701,4.9258194,5.388125,5.8504305,6.3127356,6.736969,7.1630154,7.5872483,8.013294,8.437528,7.763106,7.0868707,6.412449,5.7380266,5.0617914,5.3246713,5.5875506,5.8504305,6.11331,6.3743763,9.275117,12.174044,15.074784,17.975525,20.87445,18.813112,16.749962,14.68681,12.625471,10.56232,11.024626,11.486931,11.949236,12.413355,12.87566,10.700105,8.52455,6.350808,4.175253,1.9996977,2.03777,2.0758421,2.1121013,2.1501737,2.1882458,3.4500678,4.7118897,5.975525,7.2373466,8.499168,6.8004227,5.0998635,3.3993049,1.7005589,0.0,1.3506571,2.6995013,4.0501585,5.4008155,6.7496595,7.949841,9.1500225,10.3502035,11.5503845,12.750566,12.812206,12.87566,12.937301,13.000754,13.062395,11.10077,9.137331,7.175706,5.2122674,3.2506418,5.2992897,7.3497505,9.400211,11.450671,13.499319,14.96238,16.425442,17.886688,19.34975,20.81281,17.174194,13.537392,9.900589,6.261973,2.6251698,2.6741197,2.7248828,2.7756457,2.8245957,2.8753586,3.1871881,3.5008307,3.8126602,4.12449,4.4381323,8.450218,12.462305,16.474392,20.48829,24.500376,21.374828,18.24928,15.125546,11.999999,8.874452,7.663393,6.450521,5.237649,4.024777,2.811905,2.2498865,1.6878681,1.1258497,0.5620184,0.0,14.837286,29.674572,44.51367,59.350956,74.18824,64.612175,55.037918,45.46185,35.887596,26.31334,21.40021,16.487082,11.573953,6.6626377,1.7495089,2.175555,2.5997884,3.0258346,3.4500678,3.874301,3.1618068,2.4493124,1.7368182,1.0243238,0.31182957,0.2755703,0.2374981,0.19942589,0.16316663,0.12509441,0.13778515,0.15047589,0.16316663,0.17585737,0.18673515,0.19942589,0.21211663,0.22480737,0.2374981,0.25018883,0.25018883,0.25018883,0.25018883,0.25018883,0.25018883,0.25018883,0.25018883,0.25018883,0.25018883,0.25018883,0.28826106,0.3245203,0.36259252,0.40066472,0.43692398,0.4749962,0.51306844,0.5493277,0.5873999,0.62547207,0.53663695,0.44961473,0.36259252,0.2755703,0.18673515,0.4749962,0.76325727,1.0497054,1.3379664,1.6244144,1.9616255,2.3006494,2.6378605,2.9750717,3.3122826,2.7992141,2.2879589,1.7748904,1.261822,0.7505665,0.6744221,0.6000906,0.52575916,0.44961473,0.37528324,0.2991388,0.22480737,0.15047589,0.07433146,0.0,0.17585737,0.34990177,0.52575916,0.69980353,0.87566096,0.9246109,0.97537386,1.0243238,1.0750868,1.1258497,1.2128719,1.2998942,1.3869164,1.4757515,1.5627737,4.8877473,8.212721,11.537694,14.862667,18.187641,17.199575,16.213324,15.22526,14.237195,13.24913,26.199121,39.149113,52.100918,65.05091,78.0009,65.413506,52.826103,40.236893,27.649492,15.062093,21.499924,27.937754,34.375584,40.813416,47.24943,37.963436,28.675629,19.387821,10.100015,0.8122072,1.0370146,1.261822,1.4866294,1.7132497,1.938057,1.938057,1.938057,1.938057,1.938057,1.938057,2.4493124,2.962381,3.4754493,3.9867048,4.499773,4.461701,4.4254417,4.3873696,4.349297,4.313038,4.0501585,3.787279,3.5243993,3.2633326,3.000453,5.049101,7.0995617,9.1500225,11.200482,13.24913,12.536636,11.8241415,11.111648,10.399154,9.686659,11.73712,13.7875805,15.838041,17.886688,19.93715,22.01299,24.08702,26.162863,28.236893,30.312735,24.562017,18.813112,13.062395,7.311678,1.5627737,2.275268,2.9877625,3.7002566,4.4127507,5.125245,7.400513,9.675781,11.949236,14.224504,16.499773,13.9507475,11.399909,8.849071,6.300045,3.7492065,12.050762,20.350506,28.650248,36.94999,45.249733,37.26182,29.27572,21.287807,13.299893,5.3119802,6.2384043,7.1630154,8.087626,9.012237,9.936848,8.588004,7.2373466,5.8866897,4.537845,3.1871881,2.5508385,1.9126755,1.2745126,0.63816285,0.0,0.0,0.0,0.0,0.0,0.0,0.099712946,0.19942589,0.2991388,0.40066472,0.50037766,0.50037766,0.50037766,0.50037766,0.50037766,0.50037766,0.48768693,0.4749962,0.46230546,0.44961473,0.43692398,0.36259252,0.28826106,0.21211663,0.13778515,0.06164073,0.099712946,0.13778515,0.17585737,0.21211663,0.25018883,0.2374981,0.22480737,0.21211663,0.19942589,0.18673515,0.16316663,0.13778515,0.11240368,0.0870222,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,1.5120108,2.7756457,4.0374675,5.2992897,6.5629244,5.5005283,4.4381323,3.3757362,2.3133402,1.2491312,1.0243238,0.7995165,0.5747091,0.34990177,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.50037766,0.8122072,1.1258497,1.4376793,1.7495089,1.3996071,1.0497054,0.69980353,0.34990177,0.0,0.0,0.0,0.0,0.0,0.0,1.7748904,3.5497808,5.3246713,7.0995617,8.874452,8.912524,8.950596,8.9868555,9.024928,9.063,7.250037,5.4370747,3.6241121,1.8129625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.21211663,0.36259252,0.51306844,0.66173136,0.8122072,0.6871128,0.5620184,0.43692398,0.31182957,0.18673515,0.16316663,0.13778515,0.11240368,0.0870222,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.21211663,0.36259252,0.51306844,0.66173136,0.8122072,0.7124943,0.61278135,0.51306844,0.41335547,0.31182957,0.31182957,0.31182957,0.31182957,0.31182957,0.31182957,0.26287958,0.21211663,0.16316663,0.11240368,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.0870222,0.11240368,0.13778515,0.16316663,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,2.6505513,2.8608549,3.0693457,3.2796493,3.489953,3.7002566,3.4083695,3.1146698,2.8227828,2.5308957,2.2371957,2.42937,2.6233568,2.8155308,3.007705,3.199879,3.5697234,3.9395678,4.309412,4.6792564,5.050914,5.4407005,5.8304877,6.2202744,6.6100616,6.9998484,6.4233265,5.844991,5.2666564,4.690134,4.1117992,4.9675174,5.823236,6.677141,7.5328593,8.386765,10.616709,12.846653,15.07841,17.308353,19.538298,17.718082,15.897869,14.077655,12.25744,10.437225,10.622148,10.80707,10.991992,11.176914,11.361836,9.487233,7.61263,5.7380266,3.8616104,1.987007,2.0232663,2.0577126,2.0921588,2.126605,2.1628644,3.290527,4.41819,5.5458527,6.6717024,7.799365,6.599184,5.4008155,4.2006345,3.000453,1.8002719,2.7901495,3.780027,4.7699046,5.7597823,6.7496595,7.890013,9.030367,10.17072,11.30926,12.449615,12.937301,13.424988,13.912675,14.400362,14.888049,13.535579,12.183108,10.830639,9.4781685,8.125698,8.950596,9.775495,10.600392,11.42529,12.250188,13.167547,14.084907,15.002265,15.919624,16.836983,14.500074,12.163166,9.824444,7.4875355,5.1506267,5.7597823,6.3707504,6.979906,7.5890613,8.200029,7.476658,6.755099,6.0317264,5.3101673,4.5867953,10.990179,17.39175,23.795134,30.196705,36.60009,30.755096,24.910107,19.065115,13.220123,7.3751316,6.378002,5.3808727,4.3819304,3.3848011,2.3876717,2.0033236,1.6171626,1.2328146,0.8466535,0.46230546,12.23931,24.018127,35.79513,47.57214,59.350956,51.7347,44.12026,36.504,28.889559,21.275116,17.757969,14.240821,10.721861,7.2047133,3.6875658,3.6222992,3.5570326,3.491766,3.4283123,3.3630457,2.9206827,2.47832,2.034144,1.5917811,1.1494182,1.0805258,1.0098201,0.93911463,0.87022203,0.7995165,0.81764615,0.83577573,0.8520924,0.87022203,0.8883517,0.82671094,0.7668832,0.7070554,0.64722764,0.5873999,0.61278135,0.63816285,0.66173136,0.6871128,0.7124943,0.63816285,0.5620184,0.48768693,0.41335547,0.33721104,0.3444629,0.35171473,0.36077955,0.3680314,0.37528324,0.40066472,0.42423326,0.44961473,0.4749962,0.50037766,0.57833505,0.6544795,0.7324369,0.8103943,0.8883517,1.1403534,1.3923552,1.6443571,1.8981718,2.1501737,2.3767939,2.6052272,2.8318477,3.0602808,3.2869012,2.810092,2.333283,1.8546607,1.3778516,0.89922947,0.87566096,0.85027945,0.824898,0.7995165,0.774135,0.6345369,0.4949388,0.35534066,0.21574254,0.07433146,0.2030518,0.32995918,0.45686656,0.5855869,0.7124943,0.80676836,0.90285534,0.99712944,1.0932164,1.1874905,1.6117238,2.03777,2.4620032,2.8880494,3.3122826,5.9392653,8.568061,11.195044,13.822026,16.450823,15.283275,14.115726,12.948178,11.780631,10.613083,22.259554,33.90784,45.556126,57.202595,68.85088,57.55975,46.27043,34.9793,23.689981,12.400664,17.721708,23.044567,28.367426,33.690285,39.01314,32.147453,25.283577,18.417887,11.552197,4.688321,4.1480584,3.6077955,3.0675328,2.5272698,1.987007,1.8999848,1.8129625,1.7241274,1.6371052,1.550083,2.0722163,2.5943494,3.1182957,3.6404288,4.162562,4.0574102,3.9522583,3.8471067,3.7419548,3.636803,3.4047437,3.1726844,2.9406252,2.7067533,2.474694,4.4145637,6.354434,8.294304,10.234174,12.175857,11.978244,11.780631,11.583018,11.385405,11.187792,12.770509,14.353225,15.935941,17.516844,19.099562,20.827314,22.555067,24.282822,26.010574,27.738327,23.137028,18.537542,13.938056,9.336758,4.7372713,5.569421,6.401571,7.2355337,8.067683,8.899834,11.65735,14.4148655,17.172382,19.929897,22.687414,19.87007,17.052727,14.235382,11.418038,8.600695,14.19731,19.795738,25.392353,30.990782,36.5874,30.147755,23.70811,17.266655,10.827013,4.3873696,6.0480433,7.706904,9.367578,11.028252,12.687112,10.97205,9.256987,7.5419245,5.826862,4.1117992,3.290527,2.467442,1.6443571,0.823085,0.0,0.0,0.0,0.0,0.0,0.0,0.07977036,0.15954071,0.23931105,0.3208944,0.40066472,0.40247768,0.40429065,0.40791658,0.40972954,0.41335547,0.42060733,0.42785916,0.43511102,0.44236287,0.44961473,0.38434806,0.3208944,0.25562772,0.19036107,0.12509441,0.15228885,0.1794833,0.20667773,0.23568514,0.26287958,0.25562772,0.24837588,0.23931105,0.23205921,0.22480737,0.19579996,0.16497959,0.13415924,0.10515183,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03988518,0.07977036,0.11965553,0.15954071,0.19942589,1.209246,2.220879,3.2306993,4.2405195,5.2503395,4.655688,4.059223,3.4645715,2.8699198,2.275268,1.9706904,1.6642996,1.3597219,1.0551442,0.7505665,0.6544795,0.56020546,0.46411842,0.36984438,0.2755703,0.39522585,0.5148814,0.6345369,0.7541924,0.87566096,0.9808127,1.0841516,1.1893034,1.2944553,1.3996071,1.1204109,0.83940166,0.56020546,0.27919623,0.0,0.0,0.0,0.0,0.0,0.0,1.7730774,3.5443418,5.317419,7.0904965,8.861761,8.549932,8.238102,7.9244595,7.61263,7.3008003,6.109684,4.9203806,3.729264,2.5399606,1.3506571,1.0823387,0.81583315,0.5475147,0.27919623,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.17041849,0.29007402,0.40972954,0.5293851,0.6508536,0.57833505,0.5058166,0.43329805,0.36077955,0.28826106,0.2574407,0.22662032,0.19761293,0.16679256,0.13778515,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.07795739,0.07977036,0.08339628,0.08520924,0.0870222,0.21030366,0.33177215,0.4550536,0.57833505,0.69980353,0.6327239,0.5656443,0.49675176,0.42967212,0.36259252,0.35534066,0.3480888,0.34083697,0.33177215,0.3245203,0.28463513,0.24474995,0.20486477,0.16497959,0.12509441,0.10515183,0.08520924,0.065266654,0.045324065,0.025381476,0.034446288,0.045324065,0.054388877,0.065266654,0.07433146,0.072518505,0.07070554,0.06707962,0.065266654,0.06164073,0.065266654,0.06707962,0.07070554,0.072518505,0.07433146,0.08520924,0.09427405,0.10515183,0.11421664,0.12509441,0.13778515,0.15047589,0.16316663,0.17585737,0.18673515,0.15772775,0.12690738,0.09789998,0.06707962,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.04169814,0.034446288,0.027194439,0.01994259,0.012690738,0.01994259,0.027194439,0.034446288,0.04169814,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.059827764,0.058014803,0.054388877,0.052575916,0.05076295,0.059827764,0.07070554,0.07977036,0.09064813,0.099712946,0.0870222,0.07433146,0.06164073,0.05076295,0.038072214,1.987007,2.2081885,2.427557,2.6469254,2.8681068,3.0874753,2.8155308,2.5417736,2.269829,1.9978848,1.7241274,1.8600996,1.9942589,2.1302311,2.2643902,2.4003625,2.6777458,2.955129,3.2325122,3.5098956,3.787279,4.1426196,4.49796,4.853301,5.2068286,5.562169,5.081734,4.603112,4.122677,3.6422417,3.1618068,4.610364,6.057108,7.5056653,8.952409,10.399154,11.9601145,13.519262,15.080223,16.63937,18.20033,16.623055,15.045776,13.466686,11.889409,10.312131,10.21967,10.127209,10.034748,9.9422865,9.849826,8.274362,6.70071,5.125245,3.5497808,1.9743162,2.0069497,2.039583,2.0722163,2.1048496,2.137483,3.1291735,4.122677,5.1143675,6.107871,7.0995617,6.399758,5.6999545,5.0001507,4.3003473,3.6005437,4.229642,4.860553,5.4896507,6.1205616,6.7496595,7.8301854,8.910711,9.989424,11.069949,12.1504755,13.062395,13.974316,14.888049,15.799969,16.71189,15.970387,15.227073,14.485571,13.742256,13.000754,12.60009,12.199425,11.800573,11.399909,10.999244,11.372714,11.744371,12.117842,12.489499,12.862969,11.8241415,10.7871275,9.750113,8.713099,7.6742706,8.845445,10.014805,11.184166,12.35534,13.524701,11.7679405,10.009366,8.252605,6.495845,4.7372713,13.53014,22.323008,31.115877,39.906933,48.699802,40.135365,31.57093,23.004683,14.440247,5.8758116,5.092612,4.309412,3.5280252,2.7448254,1.9616255,1.7549478,1.54827,1.3397794,1.1331016,0.9246109,9.643148,18.359873,27.07841,35.79513,44.511856,38.857227,33.2026,27.547966,21.891523,16.236893,14.115726,11.992747,9.869768,7.746789,5.6256227,5.0708566,4.514277,3.9595103,3.4047437,2.8499773,2.6777458,2.5055144,2.333283,2.1592383,1.987007,1.8854811,1.7821422,1.6806163,1.5772774,1.4757515,1.4975071,1.5192627,1.5428312,1.5645868,1.5881553,1.455809,1.3216497,1.1893034,1.0569572,0.9246109,0.97537386,1.0243238,1.0750868,1.1258497,1.1747998,1.0243238,0.87566096,0.72518504,0.5747091,0.42423326,0.40247768,0.38072214,0.35715362,0.33539808,0.31182957,0.3245203,0.33721104,0.34990177,0.36259252,0.37528324,0.61822027,0.85934424,1.1022812,1.3452182,1.5881553,1.8057107,2.0232663,2.2408218,2.4583774,2.6741197,2.7919624,2.909805,3.0276475,3.1454902,3.2633326,2.819157,2.3767939,1.9344311,1.4920682,1.0497054,1.0750868,1.1004683,1.1258497,1.1494182,1.1747998,0.969935,0.7650702,0.56020546,0.35534066,0.15047589,0.23024625,0.3100166,0.38978696,0.46955732,0.5493277,0.69073874,0.83033687,0.969935,1.1095331,1.2491312,2.0123885,2.7756457,3.53709,4.3003473,5.0617914,6.9925966,8.921589,10.852394,12.783199,14.712192,13.36516,12.018129,10.669285,9.322253,7.9752226,18.319986,28.664751,39.009518,49.35428,59.699043,49.70781,39.71476,29.721708,19.730473,9.737422,13.945308,18.153194,22.359268,26.567154,30.77504,26.33328,21.88971,17.447952,13.00438,8.562622,7.2572894,5.9519563,4.646623,3.343103,2.03777,1.8619126,1.6878681,1.5120108,1.3379664,1.162109,1.69512,2.228131,2.759329,3.29234,3.825351,3.6531196,3.4808881,3.3068438,3.1346123,2.962381,2.759329,2.5580902,2.3550384,2.1519866,1.9507477,3.780027,5.6093063,7.440398,9.269678,11.10077,11.418038,11.735307,12.052575,12.3698435,12.687112,13.802084,14.917056,16.032028,17.147,18.261972,19.641636,21.023113,22.402779,23.782444,25.162107,21.71204,18.261972,14.811904,11.361836,7.911769,8.865387,9.817192,10.770811,11.722616,12.674421,15.915998,19.155762,22.395527,25.63529,28.875055,25.789392,22.705544,19.61988,16.534218,13.45037,16.34567,19.239159,22.13446,25.029762,27.925062,23.031878,18.140503,13.247317,8.354132,3.4627585,5.857682,8.252605,10.64753,13.042453,15.437376,13.357908,11.27844,9.197159,7.117691,5.038223,4.0302157,3.0222087,2.0142014,1.0080072,0.0,0.0,0.0,0.0,0.0,0.0,0.059827764,0.11965553,0.1794833,0.23931105,0.2991388,0.3045777,0.3100166,0.3154555,0.3208944,0.3245203,0.35171473,0.38072214,0.40791658,0.43511102,0.46230546,0.40791658,0.35171473,0.29732585,0.24293698,0.18673515,0.20486477,0.2229944,0.23931105,0.2574407,0.2755703,0.27194437,0.27013144,0.26831847,0.26469254,0.26287958,0.22662032,0.19217403,0.15772775,0.12328146,0.0870222,0.07070554,0.052575916,0.034446288,0.018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.90829426,1.6642996,2.422118,3.1799364,3.9377546,3.8108473,3.682127,3.5552197,3.4283123,3.299592,2.9152439,2.5308957,2.1447346,1.7603867,1.3742256,1.209246,1.0442665,0.8792868,0.71430725,0.5493277,0.7523795,0.9554313,1.1566701,1.3597219,1.5627737,1.4594349,1.357909,1.2545701,1.1530442,1.0497054,0.83940166,0.630911,0.42060733,0.21030366,0.0,0.0,0.0,0.0,0.0,0.0,1.7694515,3.540716,5.3101673,7.079619,8.8508835,8.187339,7.5256076,6.8620634,6.200332,5.5367875,4.9693303,4.401873,3.834416,3.2669585,2.6995013,2.1646774,1.6298534,1.0950294,0.56020546,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.12690738,0.21755551,0.30820364,0.39703882,0.48768693,0.46774435,0.44780177,0.42785916,0.40791658,0.387974,0.35171473,0.31726846,0.28282216,0.24837588,0.21211663,0.18673515,0.16316663,0.13778515,0.11240368,0.0870222,0.092461094,0.09789998,0.10333887,0.10696479,0.11240368,0.20667773,0.30276474,0.39703882,0.49312583,0.5873999,0.5529536,0.5166943,0.48224804,0.44780177,0.41335547,0.39703882,0.3825351,0.3680314,0.35171473,0.33721104,0.30820364,0.27738327,0.24837588,0.21755551,0.18673515,0.15954071,0.13234627,0.10515183,0.07795739,0.05076295,0.058014803,0.065266654,0.072518505,0.07977036,0.0870222,0.08339628,0.07795739,0.072518505,0.06707962,0.06164073,0.06707962,0.072518505,0.07795739,0.08339628,0.0870222,0.10696479,0.12690738,0.14684997,0.16679256,0.18673515,0.18673515,0.18673515,0.18673515,0.18673515,0.18673515,0.16497959,0.14322405,0.11965553,0.09789998,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.034446288,0.032633327,0.030820364,0.027194439,0.025381476,0.027194439,0.030820364,0.032633327,0.034446288,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.058014803,0.052575916,0.047137026,0.04169814,0.038072214,0.045324065,0.052575916,0.059827764,0.06707962,0.07433146,0.07433146,0.07433146,0.07433146,0.07433146,0.07433146,1.3252757,1.5555218,1.7857682,2.0142014,2.2444477,2.474694,2.222692,1.9706904,1.7168756,1.4648738,1.2128719,1.2908293,1.3669738,1.4449311,1.5228885,1.6008459,1.7857682,1.9706904,2.1556125,2.3405347,2.525457,2.8445382,3.1654327,3.484514,3.8054085,4.12449,3.7419548,3.3594196,2.9768846,2.5943494,2.2118144,4.25321,6.2927933,8.3323765,10.371959,12.413355,13.301706,14.191871,15.082036,15.9722,16.862366,15.528025,14.191871,12.857531,11.5231905,10.1870365,9.817192,9.447348,9.077503,8.70766,8.337815,7.063302,5.7869763,4.512464,3.2379513,1.9616255,1.9924458,2.0232663,2.0522738,2.0830941,2.1121013,2.9696326,3.827164,4.6846952,5.542227,6.399758,6.200332,6.000906,5.7996674,5.600241,5.4008155,5.669134,5.9392653,6.209397,6.4795284,6.7496595,7.7703576,8.789243,9.80994,10.830639,11.849524,13.1874895,14.525456,15.863422,17.199575,18.537542,18.405195,18.27285,18.140503,18.008158,17.87581,16.249584,14.625169,13.000754,11.374527,9.750113,9.577881,9.40565,9.231606,9.059374,8.887142,9.1500225,9.412902,9.675781,9.936848,10.199727,11.929294,13.660673,15.39024,17.119806,18.849373,16.05741,13.265448,10.471672,7.6797094,4.8877473,16.0701,27.252453,38.434807,49.61716,60.799515,49.515633,38.229942,26.94425,15.660371,4.3746786,3.8072214,3.2397642,2.6723068,2.1048496,1.5373923,1.5083848,1.4775645,1.4467441,1.4177368,1.3869164,7.0451727,12.701616,18.359873,24.018127,29.674572,25.979753,22.284937,18.590118,14.895301,11.200482,10.471672,9.744674,9.017676,8.290678,7.5618668,6.5176005,5.473334,4.4272547,3.3829882,2.3369088,2.4348087,2.5327086,2.6306088,2.7266958,2.8245957,2.6904364,2.5544643,2.420305,2.2843328,2.1501737,2.1773682,2.2045624,2.231757,2.2607644,2.2879589,2.0830941,1.8782293,1.6733645,1.4666867,1.261822,1.3379664,1.4122978,1.4866294,1.5627737,1.6371052,1.4122978,1.1874905,0.96268314,0.73787576,0.51306844,0.4604925,0.40791658,0.35534066,0.30276474,0.25018883,0.25018883,0.25018883,0.25018883,0.25018883,0.25018883,0.65810543,1.064209,1.4721256,1.8800422,2.2879589,2.469255,2.6523643,2.8354735,3.0167696,3.199879,3.207131,3.2143826,3.2216346,3.2306993,3.2379513,2.8300345,2.422118,2.0142014,1.6080978,1.2001812,1.2745126,1.3506571,1.4249886,1.49932,1.5754645,1.305333,1.0352017,0.7650702,0.4949388,0.22480737,0.2574407,0.29007402,0.32270733,0.35534066,0.387974,0.5728962,0.75781834,0.94274056,1.1276628,1.3125849,2.4130533,3.5117085,4.612177,5.712645,6.813113,8.044115,9.27693,10.509744,11.7425585,12.975373,11.447045,9.920531,8.392203,6.8656893,5.337362,14.380419,23.421663,32.46472,41.50778,50.549023,41.854053,33.1609,24.464117,15.769149,7.07418,10.167094,13.260008,16.352922,19.444023,22.536938,20.517298,18.497658,16.478018,14.458377,12.436923,10.368333,8.29793,6.2275267,4.157123,2.08672,1.8256533,1.5627737,1.2998942,1.0370146,0.774135,1.3180238,1.8600996,2.4021754,2.9442513,3.48814,3.247016,3.007705,2.7665808,2.5272698,2.2879589,2.1157274,1.9416829,1.7694515,1.5972201,1.4249886,3.1454902,4.8641787,6.58468,8.3051815,10.025683,10.857833,11.689982,12.522133,13.354282,14.188245,14.835473,15.4827,16.129929,16.777155,17.424383,18.457771,19.489347,20.522736,21.554312,22.5877,20.287052,17.988214,15.687565,13.386916,11.088079,12.15954,13.232814,14.304275,15.377548,16.450823,20.172834,23.894846,27.618671,31.340685,35.062695,31.71053,28.35836,25.00438,21.652212,18.300045,18.492218,18.684393,18.876566,19.070553,19.262728,15.917811,12.572895,9.22798,5.883064,2.5381477,5.667321,8.798307,11.927481,15.058467,18.187641,15.741954,13.29808,10.852394,8.406708,5.962834,4.7699046,3.576975,2.3858588,1.1929294,0.0,0.0,0.0,0.0,0.0,0.0,0.03988518,0.07977036,0.11965553,0.15954071,0.19942589,0.20667773,0.21574254,0.2229944,0.23024625,0.2374981,0.28463513,0.33177215,0.38072214,0.42785916,0.4749962,0.42967212,0.38434806,0.34083697,0.2955129,0.25018883,0.2574407,0.26469254,0.27194437,0.27919623,0.28826106,0.29007402,0.291887,0.2955129,0.29732585,0.2991388,0.25925365,0.21936847,0.1794833,0.13959812,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.6055295,1.1095331,1.6153497,2.1193533,2.6251698,2.9641938,3.3050308,3.6458678,3.9848917,4.325729,3.8597972,3.395679,2.9297476,2.465629,1.9996977,1.7658255,1.5301404,1.2944553,1.0605831,0.824898,1.1095331,1.3941683,1.6806163,1.9652514,2.2498865,1.93987,1.6298534,1.3198367,1.0098201,0.69980353,0.56020546,0.42060733,0.27919623,0.13959812,0.0,0.0,0.0,0.0,0.0,0.0,1.7676386,3.5352771,5.3029156,7.0705543,8.838193,7.8247466,6.813113,5.7996674,4.788034,3.774588,3.83079,3.8851788,3.9395678,3.9957695,4.0501585,3.247016,2.4456866,1.6425442,0.83940166,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.08520924,0.14503701,0.20486477,0.26469254,0.3245203,0.35715362,0.38978696,0.4224203,0.4550536,0.48768693,0.44780177,0.40791658,0.3680314,0.32814622,0.28826106,0.25018883,0.21211663,0.17585737,0.13778515,0.099712946,0.10696479,0.11421664,0.12328146,0.13053331,0.13778515,0.20486477,0.27194437,0.34083697,0.40791658,0.4749962,0.47318324,0.46955732,0.46774435,0.46411842,0.46230546,0.4405499,0.4169814,0.39522585,0.37165734,0.34990177,0.32995918,0.3100166,0.29007402,0.27013144,0.25018883,0.21574254,0.1794833,0.14503701,0.11059072,0.07433146,0.07977036,0.08520924,0.09064813,0.09427405,0.099712946,0.092461094,0.08520924,0.07795739,0.07070554,0.06164073,0.07070554,0.07795739,0.08520924,0.092461094,0.099712946,0.13053331,0.15954071,0.19036107,0.21936847,0.25018883,0.2374981,0.22480737,0.21211663,0.19942589,0.18673515,0.17223145,0.15772775,0.14322405,0.12690738,0.11240368,0.09064813,0.06707962,0.045324065,0.02175555,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.027194439,0.030820364,0.032633327,0.034446288,0.038072214,0.034446288,0.032633327,0.030820364,0.027194439,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.054388877,0.047137026,0.03988518,0.032633327,0.025381476,0.030820364,0.034446288,0.03988518,0.045324065,0.05076295,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.66173136,0.90285534,1.1421664,1.3832904,1.6226015,1.8619126,1.6298534,1.3977941,1.1657349,0.9318628,0.69980353,0.7197462,0.73968875,0.75963134,0.7795739,0.7995165,0.8919776,0.98443866,1.0768998,1.1693609,1.261822,1.54827,1.8329052,2.1175404,2.4021754,2.6868105,2.4021754,2.1175404,1.8329052,1.54827,1.261822,3.8942437,6.526665,9.1609,11.793322,14.425743,14.645112,14.86448,15.085662,15.30503,15.524399,14.432995,13.339779,12.246562,11.155159,10.061942,9.414715,8.767487,8.120259,7.473032,6.825804,5.8504305,4.8750563,3.8996825,2.9243085,1.9507477,1.9779422,2.0051367,2.032331,2.0595255,2.08672,2.810092,3.531651,4.255023,4.9783955,5.6999545,5.999093,6.300045,6.599184,6.9001355,7.1992745,7.1104393,7.019791,6.929143,6.8403077,6.7496595,7.71053,8.669587,9.630457,10.589515,11.5503845,13.312584,15.074784,16.836983,18.599184,20.363195,20.840004,21.316814,21.795437,22.272245,22.750868,19.90089,17.050913,14.199123,11.349146,8.499168,7.783048,7.065115,6.347182,5.6292486,4.9131284,6.474089,8.036863,9.599637,11.162411,12.725184,15.014956,17.304728,19.5945,21.884272,24.175856,20.34688,16.519714,12.692551,8.865387,5.038223,18.610062,32.1819,45.75555,59.32739,72.90104,58.8959,44.890766,30.883818,16.880495,2.8753586,2.521831,2.1701162,1.8165885,1.4648738,1.1131591,1.260009,1.4068589,1.5555218,1.7023718,1.8492218,4.4471974,7.0451727,9.643148,12.23931,14.837286,13.102281,11.367275,9.63227,7.897265,6.16226,6.82943,7.4966,8.165584,8.832754,9.499924,7.9643445,6.430578,4.894999,3.3594196,1.8256533,2.1918716,2.5599031,2.9279346,3.294153,3.6621845,3.4953918,3.3267863,3.159994,2.9932013,2.8245957,2.857229,2.8898623,2.9224956,2.955129,2.9877625,2.7103791,2.4329958,2.1556125,1.8782293,1.6008459,1.7005589,1.8002719,1.8999848,1.9996977,2.0994108,1.8002719,1.49932,1.2001812,0.89922947,0.6000906,0.5166943,0.43511102,0.35171473,0.27013144,0.18673515,0.17585737,0.16316663,0.15047589,0.13778515,0.12509441,0.6979906,1.2708868,1.84197,2.4148662,2.9877625,3.1346123,3.2832751,3.4301252,3.576975,3.7256382,3.6222992,3.5207734,3.4174345,3.3140955,3.2125697,2.8409123,2.467442,2.0957847,1.7223145,1.3506571,1.4757515,1.6008459,1.7241274,1.8492218,1.9743162,1.6407311,1.305333,0.969935,0.6345369,0.2991388,0.28463513,0.27013144,0.25562772,0.23931105,0.22480737,0.4550536,0.6852999,0.9155461,1.1457924,1.3742256,2.811905,4.249584,5.6872635,7.124943,8.562622,9.097446,9.63227,10.167094,10.701918,11.236742,9.530745,7.8229337,6.115123,4.407312,2.6995013,10.439038,18.18039,25.919926,33.659462,41.399002,34.002113,26.605227,19.206526,11.809638,4.4127507,6.390693,8.366822,10.344765,12.322706,14.300649,14.703127,15.105604,15.508082,15.91056,16.313038,13.477564,10.642091,7.806617,4.972956,2.137483,1.7875811,1.4376793,1.0877775,0.73787576,0.387974,0.93911463,1.4920682,2.0450218,2.5979755,3.149116,2.8427253,2.5345216,2.228131,1.9199274,1.6117238,1.4703126,1.3270886,1.1856775,1.0424535,0.89922947,2.5091403,4.119051,5.730775,7.3406854,8.950596,10.297627,11.644659,12.99169,14.340534,15.687565,15.867048,16.048346,16.227829,16.40731,16.586794,17.272095,17.957394,18.642694,19.327993,20.013294,18.862062,17.712645,16.563227,15.411995,14.262577,15.455506,16.646622,17.839552,19.03248,20.22541,24.42967,28.635744,32.840004,37.044266,41.25034,37.629852,34.009365,30.390692,26.770205,23.14972,20.64058,18.129625,15.620485,13.109532,10.600392,8.801933,7.0052876,5.2068286,3.4101827,1.6117238,5.47696,9.342196,13.207433,17.072668,20.937904,18.127813,15.31772,12.507628,9.697536,6.887445,5.5095935,4.1317415,2.7557032,1.3778516,0.0,0.0,0.0,0.0,0.0,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.11059072,0.11965553,0.13053331,0.13959812,0.15047589,0.21755551,0.28463513,0.35171473,0.42060733,0.48768693,0.45324063,0.4169814,0.3825351,0.3480888,0.31182957,0.3100166,0.30820364,0.3045777,0.30276474,0.2991388,0.30820364,0.3154555,0.32270733,0.32995918,0.33721104,0.291887,0.24837588,0.2030518,0.15772775,0.11240368,0.09064813,0.06707962,0.045324065,0.02175555,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.30276474,0.55476654,0.80676836,1.0605831,1.3125849,2.1193533,2.9279346,3.7347028,4.5432844,5.3500524,4.804351,4.2604623,3.7147603,3.1708715,2.6251698,2.3205922,2.0142014,1.7096237,1.405046,1.1004683,1.4666867,1.8347181,2.2027495,2.570781,2.9369993,2.420305,1.9017978,1.3851035,0.8665961,0.34990177,0.27919623,0.21030366,0.13959812,0.07070554,0.0,0.0,0.0,0.0,0.0,0.0,1.7658255,3.529838,5.295664,7.059676,8.825501,7.462154,6.1006193,4.7372713,3.3757362,2.0123885,2.6904364,3.3666716,4.0447197,4.7227674,5.4008155,4.329355,3.2597067,2.1900587,1.1204109,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.04169814,0.072518505,0.10333887,0.13234627,0.16316663,0.24837588,0.33177215,0.4169814,0.50219065,0.5873999,0.5420758,0.49675176,0.45324063,0.40791658,0.36259252,0.31182957,0.26287958,0.21211663,0.16316663,0.11240368,0.12328146,0.13234627,0.14322405,0.15228885,0.16316663,0.2030518,0.24293698,0.28282216,0.32270733,0.36259252,0.39159992,0.4224203,0.45324063,0.48224804,0.51306844,0.48224804,0.45324063,0.4224203,0.39159992,0.36259252,0.35171473,0.34264994,0.33177215,0.32270733,0.31182957,0.27013144,0.22662032,0.18492219,0.14322405,0.099712946,0.10333887,0.10515183,0.10696479,0.11059072,0.11240368,0.10333887,0.092461094,0.08339628,0.072518505,0.06164073,0.072518505,0.08339628,0.092461094,0.10333887,0.11240368,0.15228885,0.19217403,0.23205921,0.27194437,0.31182957,0.28826106,0.26287958,0.2374981,0.21211663,0.18673515,0.1794833,0.17223145,0.16497959,0.15772775,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.01994259,0.027194439,0.034446288,0.04169814,0.05076295,0.04169814,0.034446288,0.027194439,0.01994259,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.052575916,0.04169814,0.032633327,0.02175555,0.012690738,0.014503701,0.018129626,0.01994259,0.02175555,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.15047589,0.0,0.25018883,0.50037766,0.7505665,1.0007553,1.2491312,1.0370146,0.824898,0.61278135,0.40066472,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.0,0.0,0.0,0.0,0.0,0.25018883,0.50037766,0.7505665,1.0007553,1.2491312,1.062396,0.87566096,0.6871128,0.50037766,0.31182957,3.53709,6.7623506,9.987611,13.212872,16.438131,15.986704,15.537089,15.087475,14.63786,14.188245,13.337966,12.487686,11.637406,10.7871275,9.936848,9.012237,8.087626,7.1630154,6.2365913,5.3119802,4.6375585,3.9631362,3.2869012,2.612479,1.938057,1.9616255,1.987007,2.0123885,2.03777,2.0631514,2.6505513,3.2379513,3.825351,4.4127507,5.0001507,5.7996674,6.599184,7.400513,8.200029,8.999546,8.549932,8.100317,7.650702,7.1992745,6.7496595,7.650702,8.549932,9.449161,10.3502035,11.249433,13.437678,15.624111,17.812357,20.000603,22.187037,23.274813,24.36259,25.450369,26.538147,27.624111,23.550385,19.474844,15.399304,11.325577,7.250037,5.9882154,4.7245803,3.4627585,2.1991236,0.93730164,3.7999697,6.6626377,9.525306,12.387974,15.250641,18.100618,20.950596,23.800573,26.65055,29.500526,24.63816,19.775795,14.911617,10.049252,5.186886,21.15002,37.111343,53.076294,69.03761,85.00075,68.27436,51.549778,34.8252,18.100618,1.3742256,1.2382535,1.1004683,0.96268314,0.824898,0.6871128,1.0116332,1.3379664,1.6624867,1.987007,2.3133402,1.8492218,1.3869164,0.9246109,0.46230546,0.0,0.22480737,0.44961473,0.6744221,0.89922947,1.1258497,3.1871881,5.2503395,7.311678,9.374829,11.437981,9.412902,7.3878226,5.3627434,3.3376641,1.3125849,1.9507477,2.5870976,3.2252605,3.8616104,4.499773,4.3003473,4.099108,3.8996825,3.7002566,3.5008307,3.53709,3.5751622,3.6132345,3.6494937,3.6875658,3.3376641,2.9877625,2.6378605,2.2879589,1.938057,2.0631514,2.1882458,2.3133402,2.4366217,2.561716,2.1882458,1.8129625,1.4376793,1.062396,0.6871128,0.5747091,0.46230546,0.34990177,0.2374981,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.73787576,1.4757515,2.2118144,2.94969,3.6875658,3.7999697,3.9123733,4.024777,4.137181,4.249584,4.0374675,3.825351,3.6132345,3.3993049,3.1871881,2.8499773,2.5127661,2.175555,1.8383441,1.49932,1.6751775,1.8492218,2.0250793,2.1991236,2.374981,1.9743162,1.5754645,1.1747998,0.774135,0.37528324,0.31182957,0.25018883,0.18673515,0.12509441,0.06164073,0.33721104,0.61278135,0.8883517,1.162109,1.4376793,3.2125697,4.98746,6.7623506,8.537241,10.312131,10.150778,9.987611,9.824444,9.663091,9.499924,7.61263,5.7253356,3.8380418,1.9507477,0.06164073,6.4994707,12.937301,19.375132,25.812962,32.25079,26.150173,20.049553,13.948935,7.850128,1.7495089,2.612479,3.4754493,4.3384194,5.199577,6.0625467,8.887142,11.711739,14.538147,17.362743,20.187338,16.586794,12.988064,9.38752,5.7869763,2.1882458,1.7495089,1.3125849,0.87566096,0.43692398,0.0,0.5620184,1.1258497,1.6878681,2.2498865,2.811905,2.4366217,2.0631514,1.6878681,1.3125849,0.93730164,0.824898,0.7124943,0.6000906,0.48768693,0.37528324,1.8746033,3.3757362,4.8750563,6.3743763,7.8755093,9.737422,11.599335,13.46306,15.324973,17.186886,16.900436,16.612177,16.325727,16.037468,15.749206,16.08823,16.425442,16.762651,17.099863,17.437075,17.437075,17.437075,17.437075,17.437075,17.437075,18.749659,20.062244,21.374828,22.687414,23.999998,28.68832,33.37483,38.06315,42.749657,47.43798,43.549175,39.66218,35.775192,31.888199,27.999393,22.787127,17.57486,12.362592,7.1503243,1.938057,1.6878681,1.4376793,1.1874905,0.93730164,0.6871128,5.2884116,9.8878975,14.487384,19.08687,23.68817,20.511858,17.33736,14.162864,10.986553,7.8120556,6.249282,4.688321,3.1255474,1.5627737,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.15047589,0.2374981,0.3245203,0.41335547,0.50037766,0.4749962,0.44961473,0.42423326,0.40066472,0.37528324,0.36259252,0.34990177,0.33721104,0.3245203,0.31182957,0.3245203,0.33721104,0.34990177,0.36259252,0.37528324,0.3245203,0.2755703,0.22480737,0.17585737,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.2745126,2.5508385,3.825351,5.0998635,6.3743763,5.750717,5.125245,4.499773,3.874301,3.2506418,2.8753586,2.5000753,2.124792,1.7495089,1.3742256,1.8256533,2.275268,2.7248828,3.1744974,3.6241121,2.9007401,2.175555,1.4503701,0.72518504,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.7621996,3.5243993,5.2884116,7.0506115,8.812811,7.0995617,5.388125,3.6748753,1.9616255,0.25018883,1.550083,2.8499773,4.1498713,5.4497657,6.7496595,5.411693,4.07554,2.7375734,1.3996071,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13778515,0.2755703,0.41335547,0.5493277,0.6871128,0.63816285,0.5873999,0.53663695,0.48768693,0.43692398,0.37528324,0.31182957,0.25018883,0.18673515,0.12509441,0.13778515,0.15047589,0.16316663,0.17585737,0.18673515,0.19942589,0.21211663,0.22480737,0.2374981,0.25018883,0.31182957,0.37528324,0.43692398,0.50037766,0.5620184,0.52575916,0.48768693,0.44961473,0.41335547,0.37528324,0.37528324,0.37528324,0.37528324,0.37528324,0.37528324,0.3245203,0.2755703,0.22480737,0.17585737,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.17585737,0.22480737,0.2755703,0.3245203,0.37528324,0.33721104,0.2991388,0.26287958,0.22480737,0.18673515,0.18673515,0.18673515,0.18673515,0.18673515,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.0,0.20667773,0.41516843,0.62184614,0.83033687,1.0370146,0.8629702,0.6871128,0.51306844,0.33721104,0.16316663,0.13778515,0.11240368,0.0870222,0.06164073,0.038072214,0.10515183,0.17223145,0.23931105,0.30820364,0.37528324,0.5747091,0.774135,0.97537386,1.1747998,1.3742256,1.1874905,1.0007553,0.8122072,0.62547207,0.43692398,3.442816,6.446895,9.452786,12.456866,15.462758,15.087475,14.712192,14.336908,13.961625,13.588155,13.08959,12.592838,12.094274,11.597522,11.10077,9.954978,8.809185,7.665206,6.5194135,5.375434,4.612177,3.8507326,3.0874753,2.324218,1.5627737,1.6624867,1.7621996,1.8619126,1.9616255,2.0631514,2.6396735,3.2180085,3.7945306,4.3728657,4.949388,5.567608,6.185828,6.8022356,7.420456,8.036863,7.6797094,7.322556,6.965402,6.6082487,6.249282,7.0542374,7.859193,8.664148,9.470917,10.275872,11.847711,13.419549,14.9932,16.565039,18.136877,18.985344,19.831997,20.680464,21.527117,22.375584,20.950596,19.525606,18.100618,16.67563,15.250641,12.939114,10.629399,8.319685,6.009971,3.7002566,6.3707504,9.039432,11.709926,14.380419,17.0491,18.381628,19.714155,21.046682,22.37921,23.711737,19.948027,16.182505,12.416981,8.653271,4.8877473,17.779724,30.671701,43.56549,56.457466,69.34944,56.12751,42.90557,29.681824,16.459887,3.2379513,2.70494,2.1719291,1.6407311,1.1077201,0.5747091,0.89922947,1.2255627,1.550083,1.8746033,2.1991236,1.7730774,1.3452182,0.91735905,0.4894999,0.06164073,0.2755703,0.48768693,0.69980353,0.9119202,1.1258497,3.0620937,5.0001507,6.9382076,8.874452,10.812509,9.432844,8.05318,6.6717024,5.292038,3.9123733,3.9377546,3.9631362,3.9867048,4.0120864,4.0374675,3.827164,3.6168604,3.4083695,3.198066,2.9877625,3.0820365,3.1781235,3.2723975,3.3666716,3.4627585,3.4772623,3.491766,3.5080826,3.5225863,3.53709,4.2894692,5.041849,5.7942286,6.546608,7.3008003,6.604623,5.910258,5.2140803,4.519716,3.825351,3.2506418,2.6741197,2.0994108,1.5247015,0.9499924,0.78319985,0.61459434,0.44780177,0.27919623,0.11240368,0.6852999,1.258196,1.8292793,2.4021754,2.9750717,3.780027,4.5849824,5.389938,6.1948934,6.9998484,6.1278133,5.2557783,4.3819304,3.5098956,2.6378605,3.2125697,3.787279,4.361988,4.936697,5.5132194,5.727149,5.942891,6.156821,6.3725634,6.588306,5.774286,4.9620786,4.1498713,3.3376641,2.525457,2.126605,1.7295663,1.3325275,0.9354887,0.53663695,0.774135,1.0116332,1.2491312,1.4866294,1.7241274,3.435564,5.145188,6.8548117,8.564435,10.275872,9.775495,9.275117,8.774739,8.274362,7.7757964,7.454902,7.135821,6.814926,6.494032,6.1749506,10.101828,14.030518,17.957394,21.884272,25.812962,21.675781,17.536787,13.399607,9.262425,5.125245,5.237649,5.3500524,5.462456,5.57486,5.6872635,8.238102,10.7871275,13.337966,15.8869915,18.43783,15.107417,11.777005,8.446592,5.1179934,1.7875811,1.6352923,1.4830034,1.3307146,1.1766127,1.0243238,1.2998942,1.5754645,1.8492218,2.124792,2.4003625,2.175555,1.9507477,1.7241274,1.49932,1.2745126,1.4231756,1.5700256,1.7168756,1.8655385,2.0123885,3.2524548,4.4925213,5.732588,6.972654,8.212721,9.817192,11.421664,13.027949,14.632421,16.236893,15.877926,15.517147,15.15818,14.7974,14.436621,15.5878525,16.73727,17.886688,19.03792,20.187338,21.202597,22.217857,23.233116,24.246561,25.26182,24.75419,24.246561,23.740746,23.233116,22.725487,28.157122,33.590572,39.022205,44.455654,49.88729,44.519108,39.15274,33.784557,28.418188,23.050007,19.284483,15.520773,11.755249,7.989726,4.2242026,5.567608,6.9092,8.252605,9.594198,10.937603,13.464873,15.992143,18.519413,21.046682,23.575766,20.350506,17.125244,13.899984,10.674724,7.4494634,5.9882154,4.5251546,3.0620937,1.6008459,0.13778515,0.11059072,0.08339628,0.054388877,0.027194439,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.12328146,0.19579996,0.26831847,0.34083697,0.41335547,0.38978696,0.3680314,0.3444629,0.32270733,0.2991388,0.34990177,0.40066472,0.44961473,0.50037766,0.5493277,0.50219065,0.4550536,0.40791658,0.36077955,0.31182957,0.27013144,0.22662032,0.18492219,0.14322405,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,1.3434052,2.6849976,4.028403,5.369995,6.7134004,6.510349,6.3072968,6.104245,5.903006,5.6999545,5.219519,4.7390842,4.2604623,3.780027,3.299592,3.636803,3.975827,4.313038,4.650249,4.98746,4.0030212,3.0167696,2.032331,1.0478923,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,1.8220274,3.644055,5.467895,7.2899227,9.11195,7.3751316,5.638314,3.8996825,2.1628644,0.42423326,1.6352923,2.8445382,4.0555973,5.2648435,6.4759026,5.529536,4.5849824,3.6404288,2.6940625,1.7495089,1.4920682,1.2346275,0.97718686,0.7197462,0.46230546,0.36984438,0.27738327,0.18492219,0.092461094,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.11059072,0.21936847,0.32995918,0.4405499,0.5493277,0.52032024,0.4894999,0.4604925,0.42967212,0.40066472,0.3480888,0.2955129,0.24293698,0.19036107,0.13778515,0.15047589,0.16316663,0.17585737,0.18673515,0.19942589,0.2030518,0.20486477,0.20667773,0.21030366,0.21211663,0.27194437,0.33177215,0.39159992,0.45324063,0.51306844,0.49675176,0.48224804,0.46774435,0.45324063,0.43692398,0.42423326,0.41335547,0.40066472,0.387974,0.37528324,0.38434806,0.39522585,0.40429065,0.41516843,0.42423326,0.36984438,0.3154555,0.25925365,0.20486477,0.15047589,0.13778515,0.12509441,0.11240368,0.099712946,0.0870222,0.09427405,0.10333887,0.11059072,0.11784257,0.12509441,0.16497959,0.20486477,0.24474995,0.28463513,0.3245203,0.32814622,0.32995918,0.33177215,0.33539808,0.33721104,0.30276474,0.26831847,0.23205921,0.19761293,0.16316663,0.13778515,0.11240368,0.0870222,0.06164073,0.038072214,0.032633327,0.027194439,0.02175555,0.018129626,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.04169814,0.034446288,0.027194439,0.01994259,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.04169814,0.034446288,0.027194439,0.01994259,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.0,0.16497959,0.32995918,0.4949388,0.65991837,0.824898,0.6871128,0.5493277,0.41335547,0.2755703,0.13778515,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.21030366,0.3444629,0.48043507,0.61459434,0.7505665,0.89922947,1.0497054,1.2001812,1.3506571,1.49932,1.3125849,1.1258497,0.93730164,0.7505665,0.5620184,3.346729,6.1332526,8.917963,11.702674,14.487384,14.188245,13.887294,13.588155,13.287203,12.988064,12.843027,12.697989,12.552953,12.407916,12.262879,10.897718,9.5325575,8.167397,6.8022356,5.4370747,4.5867953,3.738329,2.8880494,2.03777,1.1874905,1.3633479,1.5373923,1.7132497,1.887294,2.0631514,2.6306088,3.198066,3.7655232,4.3329806,4.900438,5.335549,5.77066,6.205771,6.640882,7.07418,6.8094873,6.544795,6.2801023,6.01541,5.750717,6.4595857,7.170267,7.8791356,8.589817,9.300498,10.257742,11.214987,12.172231,13.129475,14.0867195,14.694061,15.303217,15.91056,16.517902,17.125244,18.350807,19.574556,20.80012,22.025682,23.249432,19.891825,16.536032,13.176612,9.820818,6.4632115,8.939718,11.418038,13.894546,16.372866,18.849373,18.66445,18.479528,18.294605,18.109684,17.92476,15.257894,12.589212,9.922344,7.2554765,4.5867953,14.409427,24.232058,34.054688,43.87732,53.69995,43.98066,34.259556,24.540262,14.819156,5.0998635,4.171627,3.245203,2.3169663,1.3905423,0.46230546,0.7868258,1.1131591,1.4376793,1.7621996,2.08672,1.69512,1.3017071,0.9101072,0.5166943,0.12509441,0.3245203,0.52575916,0.72518504,0.9246109,1.1258497,2.9369993,4.749962,6.5629244,8.375887,10.1870365,9.452786,8.716724,7.9824743,7.2482243,6.5121617,5.924762,5.337362,4.749962,4.162562,3.5751622,3.3557937,3.1346123,2.9152439,2.6958754,2.474694,2.6269827,2.7792716,2.9333735,3.0856624,3.2379513,3.6168604,3.9975824,4.3783045,4.7572136,5.137936,6.5176005,7.897265,9.27693,10.658407,12.038072,11.022813,10.007553,8.992294,7.9770355,6.9617763,5.924762,4.8877473,3.8507326,2.811905,1.7748904,1.4648738,1.1548572,0.8448406,0.53482395,0.22480737,0.6327239,1.0406405,1.4467441,1.8546607,2.2625773,3.7600844,5.2575917,6.755099,8.252605,9.750113,8.21816,6.684393,5.1524396,3.6204863,2.08672,3.5751622,5.0617914,6.550234,8.036863,9.525306,9.780933,10.034748,10.290376,10.54419,10.799818,9.574255,8.350506,7.124943,5.89938,4.6756306,3.9431937,3.2107568,2.47832,1.745883,1.0116332,1.2128719,1.4122978,1.6117238,1.8129625,2.0123885,3.6567454,5.3029156,6.947273,8.59163,10.2378,9.400211,8.562622,7.7250338,6.887445,6.049856,7.2971745,8.544493,9.791811,11.040942,12.28826,13.704185,15.121921,16.539658,17.957394,19.375132,17.199575,15.025834,12.850279,10.674724,8.499168,7.8628187,7.224656,6.588306,5.9501433,5.3119802,7.5872483,9.862516,12.137785,14.413053,16.68832,13.628039,10.567759,7.507478,4.4471974,1.3869164,1.5192627,1.651609,1.7857682,1.9181144,2.0504606,2.03777,2.0250793,2.0123885,1.9996977,1.987007,1.9126755,1.8383441,1.7621996,1.6878681,1.6117238,2.0196402,2.427557,2.8354735,3.24339,3.6494937,4.6303062,5.6093063,6.590119,7.569119,8.549932,9.896963,11.245807,12.592838,13.939869,15.2869005,14.855415,14.422117,13.990632,13.557334,13.125849,15.087475,17.0491,19.012539,20.974165,22.937603,24.96812,26.996826,29.027344,31.057861,33.08838,30.760536,28.432692,26.104849,23.777004,21.44916,27.627737,33.8045,39.983078,46.15984,52.338417,45.489044,38.6433,31.793924,24.948177,18.100618,15.781839,13.464873,11.147907,8.829127,6.5121617,9.447348,12.382534,15.31772,18.252907,21.188093,21.643147,22.098202,22.553255,23.008308,23.463362,20.187338,16.913128,13.637105,10.362894,7.0868707,5.7253356,4.361988,3.000453,1.6371052,0.2755703,0.21936847,0.16497959,0.11059072,0.054388877,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.09427405,0.15228885,0.21030366,0.26831847,0.3245203,0.3045777,0.28463513,0.26469254,0.24474995,0.22480737,0.33721104,0.44961473,0.5620184,0.6744221,0.7868258,0.67986095,0.5728962,0.46411842,0.35715362,0.25018883,0.21574254,0.1794833,0.14503701,0.11059072,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,1.4104849,2.819157,4.229642,5.6401267,7.0506115,7.26998,7.4893484,7.71053,7.9298983,8.149267,7.5654926,6.979906,6.394319,5.810545,5.224958,5.4497657,5.674573,5.89938,6.1241875,6.350808,5.105303,3.8597972,2.6142921,1.3705997,0.12509441,0.15047589,0.17585737,0.19942589,0.22480737,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,1.8818551,3.7655232,5.6473784,7.5292335,9.412902,7.650702,5.8866897,4.12449,2.3622901,0.6000906,1.7205015,2.8390994,3.9595103,5.0799212,6.200332,5.6473784,5.0944247,4.5432844,3.9903307,3.437377,2.9351864,2.4329958,1.9308052,1.4268016,0.9246109,0.73968875,0.55476654,0.36984438,0.18492219,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08339628,0.16497959,0.24837588,0.32995918,0.41335547,0.40247768,0.39159992,0.3825351,0.37165734,0.36259252,0.3208944,0.27738327,0.23568514,0.19217403,0.15047589,0.16316663,0.17585737,0.18673515,0.19942589,0.21211663,0.20486477,0.19761293,0.19036107,0.18310922,0.17585737,0.23205921,0.29007402,0.3480888,0.40429065,0.46230546,0.46955732,0.47680917,0.48587397,0.49312583,0.50037766,0.4749962,0.44961473,0.42423326,0.40066472,0.37528324,0.44417584,0.5148814,0.5855869,0.6544795,0.72518504,0.61459434,0.5058166,0.39522585,0.28463513,0.17585737,0.16316663,0.15047589,0.13778515,0.12509441,0.11240368,0.11421664,0.11784257,0.11965553,0.12328146,0.12509441,0.15410182,0.18492219,0.21574254,0.24474995,0.2755703,0.31726846,0.36077955,0.40247768,0.44417584,0.48768693,0.4169814,0.3480888,0.27738327,0.20667773,0.13778515,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.065266654,0.054388877,0.045324065,0.034446288,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.034446288,0.032633327,0.030820364,0.027194439,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.034446288,0.032633327,0.030820364,0.027194439,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.0,0.12328146,0.24474995,0.3680314,0.4894999,0.61278135,0.51306844,0.41335547,0.31182957,0.21211663,0.11240368,0.11240368,0.11240368,0.11240368,0.11240368,0.11240368,0.3154555,0.5166943,0.7197462,0.922798,1.1258497,1.2255627,1.3252757,1.4249886,1.5247015,1.6244144,1.4376793,1.2491312,1.062396,0.87566096,0.6871128,3.2524548,5.8177967,8.383139,10.946668,13.512011,13.287203,13.062395,12.837588,12.612781,12.387974,12.594651,12.803142,13.009819,13.21831,13.424988,11.840459,10.255929,8.669587,7.0850577,5.5005283,4.5632267,3.625925,2.6868105,1.7495089,0.8122072,1.062396,1.3125849,1.5627737,1.8129625,2.0631514,2.619731,3.1781235,3.7347028,4.2930956,4.8496747,5.101677,5.3554916,5.6074934,5.859495,6.11331,5.9392653,5.767034,5.5948024,5.422571,5.2503395,5.864934,6.4795284,7.0941224,7.71053,8.325124,8.667774,9.010424,9.353074,9.695724,10.036561,10.4045925,10.772624,11.1406555,11.506873,11.874905,15.749206,19.62532,23.49962,27.375734,31.250036,26.844538,22.440851,18.035353,13.629852,9.224354,11.510499,13.794832,16.080978,18.36531,20.649643,18.947271,17.2449,15.542528,13.840157,12.137785,10.567759,8.997733,7.4277077,5.857682,4.2876563,11.039129,17.792416,24.5457,31.297173,38.048645,31.831997,25.615349,19.396887,13.180238,6.9617763,5.6401267,4.3184767,2.9950142,1.6733645,0.34990177,0.6744221,1.0007553,1.3252757,1.649796,1.9743162,1.6171626,1.260009,0.90285534,0.54570174,0.18673515,0.37528324,0.5620184,0.7505665,0.93730164,1.1258497,2.811905,4.499773,6.187641,7.8755093,9.563377,9.47273,9.382081,9.293246,9.202598,9.11195,7.911769,6.7134004,5.5132194,4.313038,3.1128569,2.8826106,2.6523643,2.422118,2.1918716,1.9616255,2.1719291,2.382233,2.5925364,2.8028402,3.0131438,3.7582715,4.503399,5.2467136,5.9918413,6.736969,8.745731,10.752681,12.75963,14.7683935,16.775343,15.441002,14.104849,12.770509,11.434355,10.100015,8.600695,7.0995617,5.600241,4.100921,2.5997884,2.1483607,1.69512,1.2418793,0.7904517,0.33721104,0.58014804,0.823085,1.064209,1.3071461,1.550083,3.7401419,5.9302006,8.120259,10.310318,12.500377,10.306692,8.1148205,5.922949,3.729264,1.5373923,3.9377546,6.338117,8.73848,11.137029,13.537392,13.832905,14.128417,14.422117,14.71763,15.013144,13.376038,11.73712,10.100015,8.46291,6.825804,5.7579694,4.690134,3.6222992,2.5544643,1.4866294,1.649796,1.8129625,1.9743162,2.137483,2.3006494,3.87974,5.4606433,7.039734,8.620637,10.199727,9.024928,7.850128,6.6753283,5.5005283,4.325729,7.1394467,9.954978,12.770509,15.58604,18.399757,17.308353,16.215137,15.121921,14.030518,12.937301,12.725184,12.513068,12.299138,12.087022,11.874905,10.487988,9.099259,7.7123427,6.3254266,4.936697,6.9382076,8.937905,10.937603,12.937301,14.936998,12.14685,9.3567,6.5665503,3.778214,0.9880646,1.405046,1.8220274,2.2408218,2.657803,3.0747845,2.7756457,2.474694,2.175555,1.8746033,1.5754645,1.649796,1.7241274,1.8002719,1.8746033,1.9507477,2.617918,3.2850883,3.9522583,4.6194286,5.2884116,6.008158,6.7279043,7.4476504,8.167397,8.887142,9.976733,11.068136,12.157727,13.247317,14.336908,13.832905,13.327088,12.823084,12.317267,11.813264,14.587097,17.362743,20.138388,22.912222,25.687866,28.73183,31.777609,34.823387,37.867348,40.913128,36.765068,32.61701,28.470764,24.322706,20.174648,27.098352,34.020245,40.942135,47.865837,54.787727,46.45898,38.132042,29.805105,21.478168,13.149418,12.279196,11.410787,10.540565,9.670342,8.80012,13.327088,17.85587,22.382835,26.909803,31.438583,29.819609,28.202446,26.585283,24.96812,23.349146,20.024172,16.699198,13.374225,10.049252,6.7242785,5.462456,4.2006345,2.9369993,1.6751775,0.41335547,0.32995918,0.24837588,0.16497959,0.08339628,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.06707962,0.11059072,0.15228885,0.19579996,0.2374981,0.21936847,0.2030518,0.18492219,0.16679256,0.15047589,0.3245203,0.50037766,0.6744221,0.85027945,1.0243238,0.8575313,0.69073874,0.52213323,0.35534066,0.18673515,0.15954071,0.13234627,0.10515183,0.07795739,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.09064813,0.06707962,0.045324065,0.02175555,0.0,1.4775645,2.955129,4.4326935,5.910258,7.3878226,8.029612,8.673213,9.3150015,9.956791,10.600392,9.909654,9.220728,8.529989,7.83925,7.1503243,7.262728,7.3751316,7.4875355,7.5999393,7.7123427,6.207584,4.702825,3.198066,1.693307,0.18673515,0.22480737,0.26287958,0.2991388,0.33721104,0.37528324,0.2991388,0.22480737,0.15047589,0.07433146,0.0,1.9434959,3.8851788,5.826862,7.7703576,9.712041,7.9244595,6.1368785,4.349297,2.561716,0.774135,1.8057107,2.8354735,3.8652363,4.894999,5.924762,5.765221,5.6056805,5.4443264,5.2847857,5.125245,4.3783045,3.6295512,2.8826106,2.13567,1.3869164,1.1095331,0.8321498,0.55476654,0.27738327,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.054388877,0.11059072,0.16497959,0.21936847,0.2755703,0.28463513,0.2955129,0.3045777,0.3154555,0.3245203,0.291887,0.25925365,0.22662032,0.19579996,0.16316663,0.17585737,0.18673515,0.19942589,0.21211663,0.22480737,0.20667773,0.19036107,0.17223145,0.15410182,0.13778515,0.19217403,0.24837588,0.30276474,0.35715362,0.41335547,0.44236287,0.47318324,0.50219065,0.533011,0.5620184,0.52575916,0.48768693,0.44961473,0.41335547,0.37528324,0.5058166,0.6345369,0.7650702,0.89560354,1.0243238,0.85934424,0.69436467,0.5293851,0.36440548,0.19942589,0.18673515,0.17585737,0.16316663,0.15047589,0.13778515,0.13415924,0.13234627,0.13053331,0.12690738,0.12509441,0.14503701,0.16497959,0.18492219,0.20486477,0.22480737,0.30820364,0.38978696,0.47318324,0.55476654,0.63816285,0.533011,0.42785916,0.32270733,0.21755551,0.11240368,0.11240368,0.11240368,0.11240368,0.11240368,0.11240368,0.09789998,0.08339628,0.06707962,0.052575916,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.027194439,0.030820364,0.032633327,0.034446288,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.027194439,0.030820364,0.032633327,0.034446288,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.0,0.07977036,0.15954071,0.23931105,0.3208944,0.40066472,0.33721104,0.2755703,0.21211663,0.15047589,0.0870222,0.099712946,0.11240368,0.12509441,0.13778515,0.15047589,0.42060733,0.69073874,0.96087015,1.2291887,1.49932,1.550083,1.6008459,1.649796,1.7005589,1.7495089,1.5627737,1.3742256,1.1874905,1.0007553,0.8122072,3.1581807,5.5023413,7.8483152,10.192475,12.536636,12.387974,12.237497,12.087022,11.938358,11.787883,12.348088,12.908294,13.466686,14.026892,14.587097,12.783199,10.9774885,9.171778,7.36788,5.562169,4.537845,3.5117085,2.4873846,1.4630609,0.43692398,0.76325727,1.0877775,1.4122978,1.7368182,2.0631514,2.610666,3.1581807,3.7056956,4.25321,4.800725,4.8696175,4.940323,5.009216,5.0799212,5.1506267,5.0708566,4.989273,4.9095025,4.8297324,4.749962,5.2702823,5.7906027,6.3091097,6.82943,7.3497505,7.077806,6.8058615,6.532104,6.26016,5.9882154,6.115123,6.24203,6.3707504,6.497658,6.624565,13.149418,19.67427,26.200935,32.72579,39.25064,33.79725,28.34567,22.892279,17.4407,11.9873085,14.079468,16.171627,18.265598,20.357758,22.449915,19.230095,16.010273,12.790451,9.570629,6.350808,5.8776245,5.4044414,4.933071,4.459888,3.9867048,7.6706448,11.352772,15.034899,18.717026,22.399153,19.685148,16.96933,14.255324,11.539507,8.825501,7.1068134,5.389938,3.673062,1.9543737,0.2374981,0.5620184,0.8883517,1.2128719,1.5373923,1.8619126,1.5392052,1.2183108,0.89560354,0.5728962,0.25018883,0.42423326,0.6000906,0.774135,0.9499924,1.1258497,2.6868105,4.249584,5.812358,7.3751316,8.937905,9.492672,10.047439,10.602205,11.156972,11.711739,9.900589,8.087626,6.2746634,4.461701,2.6505513,2.4094272,2.1701162,1.9308052,1.6896812,1.4503701,1.7168756,1.9851941,2.2516994,2.520018,2.7883365,3.8978696,5.0074024,6.1169357,7.228282,8.337815,10.97205,13.608097,16.242332,18.87838,21.512613,19.85738,18.202145,16.54691,14.891675,13.238253,11.274815,9.313189,7.3497505,5.388125,3.4246864,2.8300345,2.2353828,1.6407311,1.0442665,0.44961473,0.5275721,0.6055295,0.68167394,0.75963134,0.8375887,3.720199,6.60281,9.48542,12.368031,15.250641,12.397038,9.545248,6.6916447,3.8398547,0.9880646,4.3003473,7.61263,10.924912,14.237195,17.549479,17.884876,18.220274,18.555672,18.889257,19.224655,17.174194,15.125546,13.075087,11.024626,8.974165,7.572745,6.169512,4.7680917,3.3648586,1.9616255,2.08672,2.2118144,2.3369088,2.4620032,2.5870976,4.102734,5.616558,7.132195,8.647832,10.161655,8.649645,7.137634,5.6256227,4.1117992,2.5997884,6.981719,11.365462,15.747393,20.129324,24.513067,20.910711,17.308353,13.704185,10.101828,6.4994707,8.2507925,10.000301,11.74981,13.499319,15.250641,13.113158,10.975676,8.838193,6.70071,4.5632267,6.2873545,8.013294,9.737422,11.463363,13.1874895,10.667472,8.147454,5.6274357,3.1074178,0.5873999,1.2908293,1.9924458,2.6958754,3.397492,4.100921,3.5117085,2.9243085,2.3369088,1.7495089,1.162109,1.3869164,1.6117238,1.8383441,2.0631514,2.2879589,3.2143826,4.1426196,5.0708566,5.99728,6.925517,7.3841968,7.844689,8.3051815,8.765674,9.224354,10.058316,10.890467,11.722616,12.554766,13.386916,12.810393,12.232059,11.655537,11.077202,10.500679,14.0867195,17.674572,21.262424,24.850279,28.438131,32.497353,36.556576,40.617615,44.676838,48.737873,42.7696,36.80314,30.834867,24.866594,18.900135,26.567154,34.234173,41.903004,49.570023,57.23704,47.428913,37.6226,27.814472,18.008158,8.200029,8.778365,9.354887,9.933222,10.509744,11.088079,17.208641,23.327389,29.44795,35.568512,41.687263,37.997883,34.308502,30.617311,26.927933,23.236742,19.862818,16.487082,13.113158,9.737422,6.3616858,5.199577,4.0374675,2.8753586,1.7132497,0.5493277,0.4405499,0.32995918,0.21936847,0.11059072,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.03988518,0.06707962,0.09427405,0.12328146,0.15047589,0.13415924,0.11965553,0.10515183,0.09064813,0.07433146,0.31182957,0.5493277,0.7868258,1.0243238,1.261822,1.0352017,0.80676836,0.58014804,0.35171473,0.12509441,0.10515183,0.08520924,0.065266654,0.045324065,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,1.5446441,3.0892882,4.6357455,6.1803894,7.7250338,8.789243,9.855265,10.919474,11.985496,13.049705,12.255627,11.459737,10.665659,9.869768,9.07569,9.07569,9.07569,9.07569,9.07569,9.07569,7.309865,5.5458527,3.780027,2.0142014,0.25018883,0.2991388,0.34990177,0.40066472,0.44961473,0.50037766,0.40066472,0.2991388,0.19942589,0.099712946,0.0,2.0033236,4.004834,6.008158,8.009668,10.012992,8.200029,6.3870673,4.574105,2.762955,0.9499924,1.8909199,2.8300345,3.7691493,4.710077,5.6491914,5.883064,6.115123,6.347182,6.5792413,6.813113,5.81961,4.8279195,3.834416,2.8427253,1.8492218,1.4793775,1.1095331,0.73968875,0.36984438,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.027194439,0.054388877,0.08339628,0.11059072,0.13778515,0.16679256,0.19761293,0.22662032,0.2574407,0.28826106,0.26469254,0.24293698,0.21936847,0.19761293,0.17585737,0.18673515,0.19942589,0.21211663,0.22480737,0.2374981,0.21030366,0.18310922,0.15410182,0.12690738,0.099712946,0.15228885,0.20486477,0.2574407,0.3100166,0.36259252,0.41516843,0.46774435,0.52032024,0.5728962,0.62547207,0.5747091,0.52575916,0.4749962,0.42423326,0.37528324,0.5656443,0.7541924,0.9445535,1.1349145,1.3252757,1.1040943,0.88472575,0.6653573,0.44417584,0.22480737,0.21211663,0.19942589,0.18673515,0.17585737,0.16316663,0.15410182,0.14684997,0.13959812,0.13234627,0.12509441,0.13415924,0.14503701,0.15410182,0.16497959,0.17585737,0.29732585,0.42060733,0.5420758,0.6653573,0.7868258,0.64722764,0.5076295,0.3680314,0.22662032,0.0870222,0.099712946,0.11240368,0.12509441,0.13778515,0.15047589,0.13053331,0.11059072,0.09064813,0.07070554,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.01994259,0.027194439,0.034446288,0.04169814,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.01994259,0.027194439,0.034446288,0.04169814,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.16316663,0.13778515,0.11240368,0.0870222,0.06164073,0.0870222,0.11240368,0.13778515,0.16316663,0.18673515,0.52575916,0.8629702,1.2001812,1.5373923,1.8746033,1.8746033,1.8746033,1.8746033,1.8746033,1.8746033,1.6878681,1.49932,1.3125849,1.1258497,0.93730164,3.0620937,5.186886,7.311678,9.438283,11.563075,11.486931,11.4126,11.338268,11.262123,11.187792,12.099712,13.011633,13.925365,14.837286,15.749206,13.724127,11.700861,9.675781,7.650702,5.6256227,4.512464,3.3993049,2.2879589,1.1747998,0.06164073,0.46230546,0.8629702,1.261822,1.6624867,2.0631514,2.5997884,3.1382382,3.6748753,4.213325,4.749962,4.6375585,4.5251546,4.4127507,4.3003473,4.1879435,4.2006345,4.213325,4.2242026,4.2368937,4.249584,4.6756306,5.0998635,5.52591,5.9501433,6.3743763,5.487838,4.599486,3.7129474,2.8245957,1.938057,1.8256533,1.7132497,1.6008459,1.4866294,1.3742256,10.549629,19.725033,28.900436,38.07584,47.24943,40.74996,34.25049,27.749205,21.249735,14.750263,16.650248,18.550234,20.450218,22.350203,24.250187,19.512917,14.775645,10.036561,5.2992897,0.5620184,1.1874905,1.8129625,2.4366217,3.0620937,3.6875658,4.3003473,4.9131284,5.52591,6.1368785,6.7496595,7.5382986,8.325124,9.11195,9.900589,10.687414,8.575313,6.4632115,4.349297,2.2371957,0.12509441,0.44961473,0.774135,1.1004683,1.4249886,1.7495089,1.4630609,1.1747998,0.8883517,0.6000906,0.31182957,0.4749962,0.63816285,0.7995165,0.96268314,1.1258497,2.561716,3.9993954,5.4370747,6.874754,8.312433,9.512614,10.712796,11.912977,13.113158,14.313339,11.887595,9.461852,7.037921,4.612177,2.1882458,1.938057,1.6878681,1.4376793,1.1874905,0.93730164,1.261822,1.5881553,1.9126755,2.2371957,2.561716,4.0374675,5.5132194,6.987158,8.46291,9.936848,13.200181,16.4617,19.725033,22.988365,26.249886,24.27557,22.29944,20.325123,18.350807,16.374678,13.9507475,11.525003,9.099259,6.6753283,4.249584,3.5117085,2.7756457,2.03777,1.2998942,0.5620184,0.4749962,0.387974,0.2991388,0.21211663,0.12509441,3.7002566,7.2754188,10.850581,14.425743,18.000906,14.487384,10.975676,7.462154,3.9504454,0.43692398,4.6629395,8.887142,13.113158,17.33736,21.563377,21.936848,22.31213,22.687414,23.062696,23.43798,20.974165,18.512161,16.050158,13.588155,11.124338,9.38752,7.650702,5.9120708,4.175253,2.4366217,2.525457,2.612479,2.6995013,2.7883365,2.8753586,4.325729,5.774286,7.224656,8.675026,10.125396,8.274362,6.4251394,4.574105,2.7248828,0.87566096,6.825804,12.774135,18.724277,24.674421,30.624563,24.513067,18.399757,12.286448,6.1749506,0.06164073,3.774588,7.4875355,11.200482,14.91343,18.624565,15.738328,12.850279,9.96223,7.07418,4.1879435,5.638314,7.0868707,8.537241,9.987611,11.437981,9.188094,6.9382076,4.688321,2.4366217,0.18673515,1.1747998,2.1628644,3.150929,4.137181,5.125245,4.249584,3.3757362,2.5000753,1.6244144,0.7505665,1.1258497,1.49932,1.8746033,2.2498865,2.6251698,3.8126602,5.0001507,6.187641,7.3751316,8.562622,8.762048,8.963287,9.162713,9.362139,9.563377,10.138086,10.712796,11.287505,11.862214,12.436923,11.787883,11.137029,10.487988,9.837135,9.188094,13.588155,17.988214,22.388275,26.788336,31.188395,36.26288,41.33736,46.411842,51.488136,56.56262,48.77413,40.987457,33.19897,25.412296,17.625622,26.03777,34.449917,42.86206,51.27602,59.688168,48.39885,37.113155,25.82384,14.538147,3.2506418,5.275721,7.3008003,9.325879,11.349146,13.374225,21.08838,28.79891,36.513065,44.22541,51.93775,46.174343,40.41275,34.64934,28.887745,23.124338,19.699652,16.274965,12.850279,9.425592,6.000906,4.936697,3.874301,2.811905,1.7495089,0.6871128,0.5493277,0.41335547,0.2755703,0.13778515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.2991388,0.6000906,0.89922947,1.2001812,1.49932,1.2128719,0.9246109,0.63816285,0.34990177,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,1.6117238,3.2252605,4.836984,6.450521,8.062244,9.550687,11.037316,12.525759,14.012388,15.50083,14.599788,13.700559,12.799516,11.900287,10.999244,10.88684,10.774437,10.662033,10.549629,10.437225,8.412147,6.3870673,4.361988,2.3369088,0.31182957,0.37528324,0.43692398,0.50037766,0.5620184,0.62547207,0.50037766,0.37528324,0.25018883,0.12509441,0.0,2.0631514,4.12449,6.187641,8.2507925,10.312131,8.4756,6.637256,4.800725,2.962381,1.1258497,1.9743162,2.8245957,3.6748753,4.5251546,5.375434,6.000906,6.624565,7.250037,7.8755093,8.499168,7.262728,6.0244746,4.788034,3.5497808,2.3133402,1.8492218,1.3869164,0.9246109,0.46230546,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,0.2374981,0.22480737,0.21211663,0.19942589,0.18673515,0.19942589,0.21211663,0.22480737,0.2374981,0.25018883,0.21211663,0.17585737,0.13778515,0.099712946,0.06164073,0.11240368,0.16316663,0.21211663,0.26287958,0.31182957,0.387974,0.46230546,0.53663695,0.61278135,0.6871128,0.62547207,0.5620184,0.50037766,0.43692398,0.37528324,0.62547207,0.87566096,1.1258497,1.3742256,1.6244144,1.3506571,1.0750868,0.7995165,0.52575916,0.25018883,0.2374981,0.22480737,0.21211663,0.19942589,0.18673515,0.17585737,0.16316663,0.15047589,0.13778515,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.28826106,0.44961473,0.61278135,0.774135,0.93730164,0.76325727,0.5873999,0.41335547,0.2374981,0.06164073,0.0870222,0.11240368,0.13778515,0.16316663,0.18673515,0.16316663,0.13778515,0.11240368,0.0870222,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.13053331,0.11059072,0.09064813,0.07070554,0.05076295,0.07070554,0.09064813,0.11059072,0.13053331,0.15047589,0.5402629,0.9300498,1.3198367,1.7096237,2.0994108,2.1175404,2.13567,2.1519866,2.1701162,2.1882458,1.9217403,1.6570477,1.3923552,1.1276628,0.8629702,2.7919624,4.7227674,6.6517596,8.582565,10.51337,10.825199,11.137029,11.450671,11.762501,12.07433,12.797703,13.519262,14.242634,14.964193,15.687565,13.600845,11.512312,9.425592,7.3370595,5.2503395,4.267714,3.2850883,2.3024626,1.3198367,0.33721104,0.6399758,0.94274056,1.2455053,1.54827,1.8492218,2.4474995,3.045777,3.6422417,4.2405195,4.836984,4.6393714,4.441758,4.2441454,4.0483456,3.8507326,3.925064,3.9993954,4.07554,4.1498713,4.2242026,4.507025,4.7898474,5.0726695,5.3554916,5.638314,5.2702823,4.902251,4.5342193,4.168001,3.7999697,4.650249,5.5005283,6.350808,7.1992745,8.049554,14.059525,20.069496,26.079466,32.08944,38.099407,32.840004,27.580599,22.319382,17.059978,11.800573,13.332527,14.86448,16.398247,17.9302,19.462152,16.731833,14.003323,11.273002,8.54268,5.812358,5.6256227,5.4370747,5.2503395,5.0617914,4.8750563,4.9802084,5.08536,5.1905117,5.295664,5.4008155,6.037165,6.6753283,7.311678,7.949841,8.588004,6.892884,5.197764,3.5026438,1.8075237,0.11240368,0.38072214,0.64722764,0.9155461,1.1820517,1.4503701,1.2491312,1.0497054,0.85027945,0.6508536,0.44961473,1.3705997,2.2897718,3.2107568,4.1299286,5.049101,6.9925966,8.934279,10.877775,12.819458,14.762955,14.989574,15.218008,15.444629,15.673061,15.899682,13.258195,10.614896,7.9715962,5.33011,2.6868105,2.3568513,2.0268922,1.696933,1.3669738,1.0370146,1.2998942,1.5627737,1.8256533,2.08672,2.3495996,3.5171473,4.6846952,5.8522434,7.019791,8.187339,11.644659,15.101978,18.559298,22.01843,25.47575,23.782444,22.09095,20.397642,18.704334,17.01284,14.558089,12.103338,9.646774,7.192023,4.7372713,4.1498713,3.5624714,2.9750717,2.3876717,1.8002719,2.0250793,2.2498865,2.474694,2.6995013,2.9243085,5.388125,7.850128,10.312131,12.775948,15.23795,12.699803,10.163468,7.6253204,5.087173,2.5508385,5.859495,9.169965,12.480434,15.790904,19.099562,19.15939,19.219215,19.280857,19.340685,19.400513,17.609306,15.819912,14.030518,12.23931,10.449916,8.80012,7.1503243,5.5005283,3.8507326,2.1991236,2.2643902,2.3296568,2.3949237,2.4601903,2.525457,3.787279,5.049101,6.3127356,7.574558,8.838193,7.592687,6.347182,5.101677,3.8579843,2.612479,7.1031876,11.592083,16.08279,20.5735,25.062395,20.258043,15.45188,10.64753,5.8431783,1.0370146,4.006647,6.978093,9.947725,12.917358,15.8869915,13.488441,11.088079,8.6877165,6.2873545,3.8869917,5.027345,6.167699,7.308052,8.448405,9.5869465,7.8102427,6.0317264,4.255023,2.47832,0.69980353,1.3905423,2.079468,2.770207,3.4591327,4.1498713,3.8851788,3.6204863,3.3557937,3.0892882,2.8245957,2.8898623,2.955129,3.0203958,3.0856624,3.149116,4.6846952,6.2202744,7.755854,9.28962,10.825199,10.970237,11.115273,11.26031,11.405348,11.5503845,12.175857,12.799516,13.424988,14.05046,14.674119,13.260008,11.845898,10.429974,9.015862,7.5999393,11.399909,15.199879,18.999847,22.799818,26.599787,30.644506,34.689224,38.73576,42.78048,46.8252,40.313038,33.800873,27.2869,20.774738,14.262577,21.385706,28.507023,35.630154,42.753284,49.8746,41.33192,32.791054,24.246561,15.705695,7.1630154,8.98323,10.801631,12.621845,14.4420595,16.262274,22.098202,27.932314,33.76824,39.602356,45.438282,41.15425,36.872032,32.589817,28.307598,24.025381,20.22541,16.425442,12.625471,8.825501,5.0255322,4.1299286,3.2343252,2.3405347,1.4449311,0.5493277,0.4405499,0.32995918,0.21936847,0.11059072,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.28463513,0.52032024,0.7541924,0.9898776,1.2255627,0.99531645,0.7650702,0.53482395,0.3045777,0.07433146,0.12328146,0.17041849,0.21755551,0.26469254,0.31182957,0.30820364,0.30276474,0.29732585,0.291887,0.28826106,0.23024625,0.17223145,0.11421664,0.058014803,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.034446288,0.07070554,0.10515183,0.13959812,0.17585737,0.19036107,0.20486477,0.21936847,0.23568514,0.25018883,1.9598125,3.6694362,5.3808727,7.0904965,8.80012,10.107266,11.4144125,12.7233715,14.030518,15.337664,15.0693445,14.802839,14.534521,14.268016,13.999697,13.207433,12.415168,11.622903,10.830639,10.038374,9.882459,9.728357,9.572442,9.416528,9.262425,7.560054,5.857682,4.15531,2.4529383,0.7505665,1.1222239,1.4956942,1.8673514,2.2408218,2.612479,4.9203806,7.228282,9.53437,11.842272,14.150173,12.612781,11.075388,9.537996,8.000604,6.4632115,6.794984,7.1267557,7.460341,7.7921133,8.125698,9.169965,10.2142315,11.26031,12.304577,13.3506565,11.447045,9.545248,7.6416373,5.7398396,3.8380418,3.105605,2.373168,1.6407311,0.90829426,0.17585737,0.13959812,0.10515183,0.07070554,0.034446288,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.03988518,0.06707962,0.09427405,0.12328146,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.059827764,0.09427405,0.13053331,0.16497959,0.19942589,0.2574407,0.3154555,0.37165734,0.42967212,0.48768693,0.47680917,0.46774435,0.45686656,0.44780177,0.43692398,0.36984438,0.30276474,0.23568514,0.16679256,0.099712946,0.13234627,0.16497959,0.19761293,0.23024625,0.26287958,0.3444629,0.42785916,0.5094425,0.59283876,0.6744221,0.6327239,0.58921283,0.5475147,0.5058166,0.46230546,0.6544795,0.8466535,1.0406405,1.2328146,1.4249886,1.3923552,1.3597219,1.3270886,1.2944553,1.261822,1.2527572,1.2418793,1.2328146,1.2219368,1.2128719,1.0315757,0.8520924,0.6726091,0.49312583,0.31182957,0.27738327,0.24293698,0.20667773,0.17223145,0.13778515,0.26287958,0.387974,0.51306844,0.63816285,0.76325727,0.6399758,0.5166943,0.39522585,0.27194437,0.15047589,0.16497959,0.1794833,0.19579996,0.21030366,0.22480737,0.19036107,0.15410182,0.11965553,0.08520924,0.05076295,0.04169814,0.034446288,0.027194439,0.01994259,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.02175555,0.032633327,0.04169814,0.052575916,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.052575916,0.04169814,0.032633327,0.02175555,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.09789998,0.08339628,0.06707962,0.052575916,0.038072214,0.052575916,0.06707962,0.08339628,0.09789998,0.11240368,0.55476654,0.99712944,1.4394923,1.8818551,2.324218,2.3604772,2.3949237,2.42937,2.465629,2.5000753,2.1574254,1.8147756,1.4721256,1.1294757,0.7868258,2.521831,4.256836,5.9918413,7.7268467,9.461852,10.161655,10.863272,11.563075,12.262879,12.962683,13.495693,14.026892,14.559902,15.092914,15.624111,13.475751,11.325577,9.175404,7.02523,4.8750563,4.022964,3.1708715,2.3169663,1.4648738,0.61278135,0.81764615,1.0225109,1.2273756,1.4322405,1.6371052,2.2952106,2.953316,3.6096084,4.267714,4.9258194,4.6429973,4.360175,4.077353,3.7945306,3.5117085,3.6494937,3.787279,3.925064,4.062849,4.2006345,4.3402324,4.4798307,4.6194286,4.76084,4.900438,5.0527267,5.2050157,5.3573046,5.5095935,5.661882,7.474845,9.287807,11.10077,12.91192,14.724882,17.56942,20.415771,23.26031,26.104849,28.949387,24.930048,20.910711,16.889559,12.870221,8.8508835,10.014805,11.18054,12.344462,13.510198,14.674119,13.95256,13.229188,12.507628,11.784257,11.062697,10.061942,9.063,8.062244,7.063302,6.0625467,5.660069,5.2575917,4.855114,4.4526362,4.0501585,4.537845,5.0255322,5.5132194,5.999093,6.48678,5.2104545,3.9323158,2.6541772,1.3778516,0.099712946,0.3100166,0.52032024,0.7306239,0.93911463,1.1494182,1.0370146,0.9246109,0.8122072,0.69980353,0.5873999,2.2643902,3.9431937,5.620184,7.2971745,8.974165,11.421664,13.8691635,16.318476,18.765976,21.211662,20.468348,19.72322,18.978092,18.232965,17.487837,14.626982,11.7679405,8.907085,6.0480433,3.1871881,2.7774587,2.3677292,1.9579996,1.54827,1.1367276,1.3379664,1.5373923,1.7368182,1.938057,2.137483,2.9968271,3.8579843,4.7173285,5.576673,6.43783,10.089137,13.742256,17.395376,21.046682,24.699802,23.289318,21.880646,20.470161,19.059675,17.64919,15.165432,12.67986,10.194288,7.71053,5.224958,4.788034,4.349297,3.9123733,3.4754493,3.0367124,3.5751622,4.1117992,4.650249,5.186886,5.7253356,7.07418,8.424837,9.775495,11.124338,12.474996,10.912222,9.349448,7.7866745,6.2257137,4.6629395,7.057863,9.452786,11.847711,14.242634,16.637558,16.38193,16.128115,15.872487,15.616859,15.363045,14.244447,13.127662,12.009064,10.89228,9.775495,8.212721,6.6499467,5.087173,3.5243993,1.9616255,2.0051367,2.0468347,2.0903459,2.132044,2.175555,3.2506418,4.325729,5.4008155,6.4759026,7.549176,6.9092,6.2692246,5.6292486,4.989273,4.349297,7.380571,10.410031,13.439491,16.470764,19.500225,16.003021,12.5058155,9.006798,5.5095935,2.0123885,4.2405195,6.4668374,8.694968,10.9230995,13.149418,11.236742,9.325879,7.413204,5.5005283,3.587853,4.41819,5.2467136,6.0770507,6.9073873,7.7377243,6.432391,5.127058,3.8217251,2.518205,1.2128719,1.6044719,1.9978848,2.3894846,2.7828975,3.1744974,3.5207734,3.8652363,4.209699,4.554162,4.900438,4.655688,4.409125,4.164375,3.919625,3.6748753,5.5567303,7.440398,9.322253,11.205922,13.087777,13.176612,13.267261,13.357908,13.446743,13.537392,14.211814,14.888049,15.56247,16.236893,16.913128,14.732134,12.552953,10.371959,8.192778,6.011784,9.211663,12.411542,15.613234,18.813112,22.01299,25.027948,28.042906,31.057861,34.07282,37.087776,31.850126,26.612478,21.374828,16.13718,10.899531,16.733644,22.564133,28.398247,34.230545,40.062847,34.26499,28.467138,22.669285,16.873243,11.075388,12.690738,14.304275,15.919624,17.534973,19.150324,23.10802,27.065718,31.023417,34.9793,38.936996,36.13416,33.33313,30.53029,27.72745,24.92461,20.749357,16.575916,12.400664,8.225411,4.0501585,3.3231604,2.5943494,1.8673514,1.1403534,0.41335547,0.32995918,0.24837588,0.16497959,0.08339628,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.05076295,0.06164073,0.07433146,0.0870222,0.099712946,0.27013144,0.4405499,0.6091554,0.7795739,0.9499924,0.7777609,0.6055295,0.43329805,0.25925365,0.0870222,0.19579996,0.30276474,0.40972954,0.5166943,0.62547207,0.61459434,0.6055295,0.5946517,0.5855869,0.5747091,0.4604925,0.3444629,0.23024625,0.11421664,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.032633327,0.065266654,0.09789998,0.13053331,0.16316663,0.23024625,0.29732585,0.36440548,0.43329805,0.50037766,2.3079014,4.115425,5.922949,7.7304726,9.537996,10.665659,11.793322,12.919171,14.046834,15.174497,15.540715,15.905121,16.269526,16.635744,17.00015,15.528025,14.055899,12.581961,11.109835,9.637709,11.352772,13.067834,14.782897,16.49796,18.213022,14.744824,11.27844,7.8102427,4.3420453,0.87566096,1.745883,2.6142921,3.484514,4.3547363,5.224958,7.7776093,10.330261,12.882912,15.435563,17.988214,16.749962,15.511708,14.275268,13.037014,11.800573,11.615651,11.430729,11.245807,11.060884,10.874149,12.340837,13.80571,15.270584,16.735458,18.20033,15.633177,13.064208,10.497053,7.9298983,5.3627434,4.360175,3.3576066,2.3550384,1.35247,0.34990177,0.27919623,0.21030366,0.13959812,0.07070554,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.07977036,0.13415924,0.19036107,0.24474995,0.2991388,0.23931105,0.1794833,0.11965553,0.059827764,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.07070554,0.09064813,0.11059072,0.13053331,0.15047589,0.27738327,0.40429065,0.533011,0.65991837,0.7868258,0.7541924,0.72337204,0.69073874,0.65810543,0.62547207,0.5275721,0.42967212,0.33177215,0.23568514,0.13778515,0.15228885,0.16679256,0.18310922,0.19761293,0.21211663,0.30276474,0.39159992,0.48224804,0.5728962,0.66173136,0.6399758,0.61822027,0.5946517,0.5728962,0.5493277,0.6852999,0.8194591,0.9554313,1.0895905,1.2255627,1.4358664,1.6443571,1.8546607,2.0649643,2.275268,2.268016,2.2607644,2.2516994,2.2444477,2.2371957,1.889107,1.5428312,1.1947423,0.8466535,0.50037766,0.42967212,0.36077955,0.29007402,0.21936847,0.15047589,0.2374981,0.3245203,0.41335547,0.50037766,0.5873999,0.5166943,0.44780177,0.3770962,0.30820364,0.2374981,0.24293698,0.24837588,0.2520018,0.2574407,0.26287958,0.21755551,0.17223145,0.12690738,0.08339628,0.038072214,0.034446288,0.032633327,0.030820364,0.027194439,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.032633327,0.03988518,0.047137026,0.054388877,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.054388877,0.047137026,0.03988518,0.032633327,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.065266654,0.054388877,0.045324065,0.034446288,0.025381476,0.034446288,0.045324065,0.054388877,0.065266654,0.07433146,0.56927025,1.064209,1.5591478,2.0558996,2.5508385,2.6016014,2.6541772,2.7067533,2.759329,2.811905,2.3931105,1.9725033,1.551896,1.1331016,0.7124943,2.2516994,3.7927177,5.331923,6.872941,8.412147,9.499924,10.587702,11.675479,12.763257,13.849221,14.191871,14.534521,14.877171,15.219821,15.56247,13.3506565,11.137029,8.925215,6.7115874,4.499773,3.778214,3.054842,2.333283,1.6099107,0.8883517,0.99531645,1.1022812,1.209246,1.3180238,1.4249886,2.1429217,2.8608549,3.576975,4.2949085,5.0128417,4.64481,4.2767787,3.9105604,3.5425289,3.1744974,3.3757362,3.5751622,3.774588,3.975827,4.175253,4.171627,4.169814,4.168001,4.164375,4.162562,4.835171,5.5077806,6.1803894,6.8529987,7.5256076,10.29944,13.075087,15.850732,18.624565,21.40021,21.079315,20.760235,20.43934,20.120258,19.799364,17.020092,14.239008,11.459737,8.680465,5.89938,6.697084,7.494787,8.292491,9.090195,9.8878975,11.173288,12.456866,13.742256,15.027647,16.313038,14.500074,12.687112,10.874149,9.063,7.250037,6.33993,5.429823,4.519716,3.6096084,2.6995013,3.0367124,3.3757362,3.7129474,4.0501585,4.3873696,3.5280252,2.666868,1.8075237,0.9481794,0.0870222,0.23931105,0.39159992,0.54570174,0.6979906,0.85027945,0.824898,0.7995165,0.774135,0.7505665,0.72518504,3.159994,5.5948024,8.029612,10.46442,12.899229,15.852545,18.80586,21.757364,24.71068,27.662184,25.945307,24.228432,22.509743,20.792868,19.074179,15.9975815,12.920984,9.842574,6.7641635,3.6875658,3.198066,2.7067533,2.2172532,1.7277533,1.2382535,1.3742256,1.5120108,1.649796,1.7875811,1.9253663,2.47832,3.0294604,3.5824142,4.135368,4.688321,8.535428,12.382534,16.229641,20.076748,23.925667,22.798004,21.670341,20.542679,19.415016,18.287354,15.772775,13.258195,10.741803,8.227224,5.712645,5.424384,5.137936,4.8496747,4.5632267,4.274966,5.125245,5.975525,6.825804,7.6742706,8.52455,8.762048,8.999546,9.237044,9.474543,9.712041,9.12464,8.537241,7.949841,7.362441,6.775041,8.254418,9.735609,11.214987,12.694364,14.175554,13.604471,13.035201,12.464118,11.894848,11.325577,10.879588,10.435412,9.989424,9.545248,9.099259,7.6253204,6.149569,4.6756306,3.199879,1.7241274,1.745883,1.7658255,1.7857682,1.8057107,1.8256533,2.712192,3.6005437,4.4870825,5.375434,6.261973,6.2275267,6.19308,6.156821,6.1223745,6.0879283,7.6579537,9.22798,10.798005,12.368031,13.938056,11.747997,9.557939,7.36788,5.177821,2.9877625,4.4725785,5.957395,7.4422116,8.927028,10.411844,8.9868555,7.5618668,6.1368785,4.7118897,3.2869012,3.8072214,4.327542,4.847862,5.368182,5.8866897,5.0545397,4.2223897,3.39024,2.5580902,1.7241274,1.8202144,1.9144884,2.0105755,2.1048496,2.1991236,3.1545548,4.1099863,5.0654173,6.0208488,6.9744673,6.4197006,5.864934,5.3101673,4.7554007,4.2006345,6.430578,8.660522,10.890467,13.12041,15.350354,15.384801,15.419247,15.455506,15.489952,15.524399,16.249584,16.97477,17.699953,18.425138,19.150324,16.20426,13.260008,10.315757,7.369693,4.4254417,7.02523,9.625018,12.224807,14.824595,17.424383,19.409578,21.394772,23.379965,25.36516,27.350353,23.387217,19.424082,15.462758,11.499621,7.5382986,12.07977,16.623055,21.164526,25.70781,30.24928,27.19625,24.145035,21.092007,18.04079,14.9877615,16.398247,17.80692,19.217403,20.627888,22.038374,24.117842,26.19731,28.276777,30.358059,32.437527,31.114063,29.792414,28.470764,27.147303,25.825651,21.275116,16.72458,12.174044,7.6253204,3.0747845,2.514579,1.9543737,1.3941683,0.83577573,0.2755703,0.21936847,0.16497959,0.11059072,0.054388877,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.15047589,0.25562772,0.36077955,0.46411842,0.56927025,0.6744221,0.56020546,0.44417584,0.32995918,0.21574254,0.099712946,0.26831847,0.43511102,0.60190356,0.7705091,0.93730164,0.922798,0.90829426,0.8919776,0.8774739,0.8629702,0.69073874,0.5166943,0.3444629,0.17223145,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.27013144,0.38978696,0.5094425,0.630911,0.7505665,2.6559901,4.559601,6.4650245,8.370448,10.275872,11.222239,12.170418,13.116784,14.064963,15.013144,16.010273,17.007402,18.004532,19.003473,20.000603,17.846804,15.694818,13.54283,11.390844,9.237044,12.823084,16.40731,19.993351,23.577578,27.163618,21.929596,16.697386,11.465176,6.2329655,1.0007553,2.3677292,3.7347028,5.10349,6.4704633,7.837437,10.634838,13.43224,16.229641,19.027042,21.824444,20.887142,19.94984,19.012539,18.075237,17.137936,16.434505,15.732889,15.02946,14.327844,13.6244135,15.509895,17.395376,19.280857,21.164526,23.050007,19.817493,16.584982,13.352469,10.119957,6.887445,5.614745,4.3420453,3.0693457,1.7966459,0.52575916,0.42060733,0.3154555,0.21030366,0.10515183,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.11965553,0.2030518,0.28463513,0.3680314,0.44961473,0.36077955,0.27013144,0.1794833,0.09064813,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.07977036,0.08520924,0.09064813,0.09427405,0.099712946,0.29732585,0.4949388,0.69255173,0.8901646,1.0877775,1.0333886,0.97718686,0.922798,0.8684091,0.8122072,0.6852999,0.55839247,0.42967212,0.30276474,0.17585737,0.17223145,0.17041849,0.16679256,0.16497959,0.16316663,0.25925365,0.35715362,0.4550536,0.5529536,0.6508536,0.64722764,0.64541465,0.6417888,0.6399758,0.63816285,0.71430725,0.79226464,0.87022203,0.9481794,1.0243238,1.4775645,1.9308052,2.382233,2.8354735,3.2869012,3.2832751,3.2778363,3.2723975,3.2669585,3.2633326,2.7466383,2.231757,1.7168756,1.2019942,0.6871128,0.581961,0.47680917,0.37165734,0.26831847,0.16316663,0.21211663,0.26287958,0.31182957,0.36259252,0.41335547,0.39522585,0.3770962,0.36077955,0.34264994,0.3245203,0.3208944,0.3154555,0.3100166,0.3045777,0.2991388,0.24474995,0.19036107,0.13415924,0.07977036,0.025381476,0.027194439,0.030820364,0.032633327,0.034446288,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.04169814,0.047137026,0.052575916,0.058014803,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.058014803,0.052575916,0.047137026,0.04169814,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.032633327,0.027194439,0.02175555,0.018129626,0.012690738,0.018129626,0.02175555,0.027194439,0.032633327,0.038072214,0.5855869,1.1331016,1.6806163,2.228131,2.7756457,2.8445382,2.9152439,2.9841363,3.054842,3.1255474,2.6269827,2.1302311,1.6316663,1.1349145,0.63816285,1.983381,3.3267863,4.6720047,6.017223,7.362441,8.838193,10.312131,11.787883,13.261822,14.737573,14.889862,15.0421505,15.194439,15.346728,15.50083,13.225562,10.950294,8.675026,6.399758,4.12449,3.531651,2.9406252,2.3477864,1.7549478,1.162109,1.1729867,1.1820517,1.1929294,1.2019942,1.2128719,1.9906329,2.7665808,3.5443418,4.322103,5.0998635,4.646623,4.195195,3.7419548,3.290527,2.8372865,3.100166,3.3630457,3.6241121,3.8869917,4.1498713,4.004834,3.8597972,3.7147603,3.5697234,3.4246864,4.6176157,5.810545,7.0016613,8.194591,9.38752,13.125849,16.862366,20.600695,24.33721,28.075539,24.589212,21.104698,17.620184,14.13567,10.649343,9.110137,7.569119,6.0299134,4.4907084,2.94969,3.3793623,3.8090343,4.2405195,4.670192,5.0998635,8.392203,11.684544,14.976884,18.269224,21.563377,18.938208,16.313038,13.687867,11.062697,8.437528,7.019791,5.6020546,4.1843176,2.7665808,1.3506571,1.5373923,1.7241274,1.9126755,2.0994108,2.2879589,1.845596,1.403233,0.96087015,0.5166943,0.07433146,0.17041849,0.26469254,0.36077955,0.4550536,0.5493277,0.61278135,0.6744221,0.73787576,0.7995165,0.8629702,4.0555973,7.2482243,10.440851,13.633478,16.824293,20.281612,23.740746,27.198065,30.655384,34.112705,31.422268,28.73183,26.043207,23.352772,20.662334,17.368181,14.072216,10.778063,7.4820967,4.1879435,3.6168604,3.04759,2.47832,1.9072367,1.3379664,1.4122978,1.4866294,1.5627737,1.6371052,1.7132497,1.9579996,2.2027495,2.4474995,2.6922495,2.9369993,6.979906,11.022813,15.065719,19.106813,23.14972,22.304878,21.460037,20.615198,19.770357,18.925516,16.380117,13.834718,11.289318,8.745731,6.200332,6.0625467,5.924762,5.7869763,5.6491914,5.5132194,6.6753283,7.837437,8.999546,10.161655,11.325577,10.449916,9.574255,8.700407,7.8247466,6.9490857,7.3370595,7.7250338,8.113008,8.499168,8.887142,9.452786,10.016619,10.582263,11.147907,11.711739,10.827013,9.9422865,9.057561,8.172835,7.28811,7.51473,7.743163,7.9697833,8.198216,8.424837,7.037921,5.6491914,4.262275,2.8753586,1.4866294,1.4848163,1.4830034,1.4793775,1.4775645,1.4757515,2.175555,2.8753586,3.5751622,4.274966,4.974769,5.5458527,6.115123,6.684393,7.2554765,7.8247466,7.935337,8.044115,8.154706,8.265296,8.374074,7.4929743,6.6100616,5.727149,4.844236,3.9631362,4.704638,5.4479527,6.189454,6.932769,7.6742706,6.736969,5.7996674,4.8623657,3.925064,2.9877625,3.198066,3.4083695,3.6168604,3.827164,4.0374675,3.6766882,3.3177216,2.956942,2.5979755,2.2371957,2.034144,1.8329052,1.6298534,1.4268016,1.2255627,2.7901495,4.3547363,5.919323,7.4857225,9.050309,8.185526,7.320743,6.454147,5.5893636,4.7245803,7.3026133,9.880646,12.456866,15.034899,17.612932,17.592989,17.573046,17.553104,17.533161,17.513218,18.287354,19.063301,19.837437,20.613384,21.38752,17.678198,13.967064,10.257742,6.546608,2.8372865,4.836984,6.836682,8.838193,10.837891,12.837588,13.793019,14.746637,15.702069,16.6575,17.612932,14.924308,12.237497,9.550687,6.8620634,4.175253,7.4277077,10.680162,13.932617,17.185072,20.437527,20.129324,19.822933,19.514729,19.208338,18.900135,20.105755,21.309563,22.515182,23.720802,24.92461,25.12766,25.330713,25.531952,25.735004,25.938055,26.095783,26.251698,26.409426,26.567154,26.724882,21.799063,16.875055,11.949236,7.02523,2.0994108,1.7078108,1.3143979,0.922798,0.5293851,0.13778515,0.11059072,0.08339628,0.054388877,0.027194439,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.05076295,0.0870222,0.12509441,0.16316663,0.19942589,0.23931105,0.27919623,0.3208944,0.36077955,0.40066472,0.34264994,0.28463513,0.22662032,0.17041849,0.11240368,0.34083697,0.56745726,0.79589057,1.0225109,1.2491312,1.2291887,1.209246,1.1893034,1.1693609,1.1494182,0.91917205,0.69073874,0.4604925,0.23024625,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.027194439,0.054388877,0.08339628,0.11059072,0.13778515,0.3100166,0.48224804,0.6544795,0.82671094,1.0007553,3.002266,5.0055895,7.0071006,9.010424,11.011934,11.780631,12.547514,13.314397,14.083094,14.849977,16.47983,18.109684,19.739536,21.36939,22.999243,20.167397,17.335548,14.501887,11.67004,8.838193,14.293397,19.746788,25.201992,30.657198,36.1124,29.114367,22.118143,15.120108,8.122072,1.1258497,2.9895754,4.855114,6.720652,8.584378,10.449916,13.492067,16.534218,19.578182,22.620335,25.662485,25.024323,24.387972,23.74981,23.11346,22.475298,21.255173,20.03505,18.814926,17.5948,16.374678,18.680767,20.985043,23.289318,25.595406,27.899681,24.001812,20.105755,16.207886,12.310016,8.412147,6.869315,5.328297,3.785466,2.2426348,0.69980353,0.56020546,0.42060733,0.27919623,0.13959812,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.15954071,0.27013144,0.38072214,0.4894999,0.6000906,0.48043507,0.36077955,0.23931105,0.11965553,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.09064813,0.07977036,0.07070554,0.059827764,0.05076295,0.31726846,0.5855869,0.8520924,1.1204109,1.3869164,1.310772,1.2328146,1.1548572,1.0768998,1.0007553,0.8430276,0.6852999,0.5275721,0.36984438,0.21211663,0.19217403,0.17223145,0.15228885,0.13234627,0.11240368,0.21755551,0.32270733,0.42785916,0.533011,0.63816285,0.6544795,0.6726091,0.69073874,0.7070554,0.72518504,0.7451276,0.7650702,0.7850128,0.80495536,0.824898,1.5192627,2.2154403,2.909805,3.6041696,4.3003473,4.2967215,4.2949085,4.2930956,4.2894692,4.2876563,3.6041696,2.9224956,2.2408218,1.5573349,0.87566096,0.73424983,0.5946517,0.4550536,0.3154555,0.17585737,0.18673515,0.19942589,0.21211663,0.22480737,0.2374981,0.27194437,0.30820364,0.34264994,0.3770962,0.41335547,0.39703882,0.3825351,0.3680314,0.35171473,0.33721104,0.27194437,0.20667773,0.14322405,0.07795739,0.012690738,0.01994259,0.027194439,0.034446288,0.04169814,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.052575916,0.054388877,0.058014803,0.059827764,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.059827764,0.058014803,0.054388877,0.052575916,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06164073,0.12509441,0.18673515,0.25018883,0.31182957,0.25018883,0.18673515,0.12509441,0.06164073,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.6000906,1.2001812,1.8002719,2.4003625,3.000453,3.0874753,3.1744974,3.2633326,3.350355,3.437377,2.8626678,2.2879589,1.7132497,1.1367276,0.5620184,1.7132497,2.8626678,4.0120864,5.163317,6.3127356,8.174648,10.036561,11.900287,13.762199,15.624111,15.5878525,15.54978,15.511708,15.475449,15.437376,13.100468,10.761745,8.424837,6.0879283,3.7492065,3.2869012,2.8245957,2.3622901,1.8999848,1.4376793,1.3506571,1.261822,1.1747998,1.0877775,1.0007553,1.8383441,2.6741197,3.5117085,4.349297,5.186886,4.650249,4.1117992,3.5751622,3.0367124,2.5000753,2.8245957,3.149116,3.4754493,3.7999697,4.12449,3.8380418,3.5497808,3.2633326,2.9750717,2.6868105,4.40006,6.11331,7.8247466,9.537996,11.249433,15.950445,20.649643,25.350657,30.049854,34.750866,28.10092,21.450974,14.799213,8.149267,1.49932,1.2001812,0.89922947,0.6000906,0.2991388,0.0,0.06164073,0.12509441,0.18673515,0.25018883,0.31182957,5.612932,10.912222,16.213324,21.512613,26.811903,23.374527,19.93715,16.499773,13.062395,9.625018,7.699652,5.774286,3.8507326,1.9253663,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.16316663,0.13778515,0.11240368,0.0870222,0.06164073,0.099712946,0.13778515,0.17585737,0.21211663,0.25018883,0.40066472,0.5493277,0.69980353,0.85027945,1.0007553,4.949388,8.899834,12.850279,16.800724,20.749357,24.712494,28.675629,32.63695,36.60009,40.563225,36.899227,33.23704,29.574858,25.912674,22.25049,18.736969,15.22526,11.711739,8.200029,4.688321,4.0374675,3.386614,2.7375734,2.08672,1.4376793,1.4503701,1.4630609,1.4757515,1.4866294,1.49932,1.4376793,1.3742256,1.3125849,1.2491312,1.1874905,5.424384,9.663091,13.899984,18.136877,22.375584,21.811752,21.249735,20.687716,20.125698,19.561867,16.98746,14.413053,11.836833,9.262425,6.688019,6.70071,6.7134004,6.7242785,6.736969,6.7496595,8.225411,9.699349,11.175101,12.650853,14.124791,12.137785,10.150778,8.161958,6.1749506,4.1879435,5.5494785,6.9128265,8.274362,9.637709,10.999244,10.649343,10.29944,9.949538,9.599637,9.249735,8.049554,6.849373,5.6491914,4.4508233,3.2506418,4.1498713,5.049101,5.9501433,6.849373,7.750415,6.450521,5.1506267,3.8507326,2.5508385,1.2491312,1.2255627,1.2001812,1.1747998,1.1494182,1.1258497,1.6371052,2.1501737,2.663242,3.1744974,3.6875658,4.8623657,6.037165,7.211965,8.386765,9.563377,8.212721,6.8620634,5.5132194,4.162562,2.811905,3.2379513,3.6621845,4.0882306,4.512464,4.936697,4.936697,4.936697,4.936697,4.936697,4.936697,4.4870825,4.0374675,3.587853,3.1382382,2.6868105,2.5870976,2.4873846,2.3876717,2.2879589,2.1882458,2.3006494,2.4130533,2.525457,2.6378605,2.7502642,2.2498865,1.7495089,1.2491312,0.7505665,0.25018883,2.4257438,4.599486,6.775041,8.950596,11.124338,9.949538,8.774739,7.5999393,6.4251394,5.2503395,8.174648,11.10077,14.025079,16.949387,19.87551,19.799364,19.725033,19.650702,19.574556,19.500225,20.325123,21.15002,21.97492,22.799818,23.624716,19.150324,14.675932,10.199727,5.7253356,1.2491312,2.6505513,4.0501585,5.4497657,6.849373,8.2507925,8.174648,8.100317,8.024173,7.949841,7.8755093,6.4632115,5.050914,3.636803,2.2245052,0.8122072,2.7756457,4.7372713,6.70071,8.662335,10.625773,13.062395,15.50083,17.937452,20.375887,22.812508,23.813263,24.812206,25.812962,26.811903,27.812658,26.137482,24.462305,22.787127,21.11195,19.436771,21.07569,22.712795,24.349901,25.987005,27.624111,22.324821,17.025532,11.724429,6.4251394,1.1258497,0.89922947,0.6744221,0.44961473,0.22480737,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,0.22480737,0.19942589,0.17585737,0.15047589,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.41335547,0.69980353,0.9880646,1.2745126,1.5627737,1.5373923,1.5120108,1.4866294,1.4630609,1.4376793,1.1494182,0.8629702,0.5747091,0.28826106,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.34990177,0.5747091,0.7995165,1.0243238,1.2491312,3.350355,5.4497657,7.549176,9.6504,11.74981,12.337211,12.92461,13.512011,14.09941,14.68681,16.949387,19.211964,21.474543,23.73712,25.999697,22.487988,18.974466,15.462758,11.949236,8.437528,15.76371,23.088078,30.412447,37.736816,45.063,36.299137,27.537088,18.77504,10.012992,1.2491312,3.6132345,5.975525,8.337815,10.700105,13.062395,16.349297,19.63801,22.924911,26.211813,29.500526,29.163317,28.824291,28.487082,28.14987,27.812658,26.074028,24.33721,22.600391,20.861761,19.124943,21.849825,24.574707,27.299591,30.024473,32.749355,28.187943,23.624716,19.06149,14.500074,9.936848,8.125698,6.3127356,4.499773,2.6868105,0.87566096,0.69980353,0.52575916,0.34990177,0.17585737,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.19942589,0.33721104,0.4749962,0.61278135,0.7505665,0.6000906,0.44961473,0.2991388,0.15047589,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.33721104,0.6744221,1.0116332,1.3506571,1.6878681,1.5881553,1.4866294,1.3869164,1.2872034,1.1874905,1.0007553,0.8122072,0.62547207,0.43692398,0.25018883,0.21211663,0.17585737,0.13778515,0.099712946,0.06164073,0.17585737,0.28826106,0.40066472,0.51306844,0.62547207,0.66173136,0.69980353,0.73787576,0.774135,0.8122072,0.774135,0.73787576,0.69980353,0.66173136,0.62547207,1.5627737,2.5000753,3.437377,4.3746786,5.3119802,5.3119802,5.3119802,5.3119802,5.3119802,5.3119802,4.461701,3.6132345,2.762955,1.9126755,1.062396,0.8883517,0.7124943,0.53663695,0.36259252,0.18673515,0.16316663,0.13778515,0.11240368,0.0870222,0.06164073,0.15047589,0.2374981,0.3245203,0.41335547,0.50037766,0.4749962,0.44961473,0.42423326,0.40066472,0.37528324,0.2991388,0.22480737,0.15047589,0.07433146,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07433146,0.15047589,0.22480737,0.2991388,0.37528324,0.2991388,0.22480737,0.15047589,0.07433146,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.48587397,0.969935,1.455809,1.93987,2.4257438,2.4891977,2.5544643,2.619731,2.6849976,2.7502642,2.333283,1.9144884,1.4975071,1.0805258,0.66173136,1.7241274,2.7883365,3.8507326,4.9131284,5.975525,7.46578,8.954222,10.444477,11.934732,13.424988,13.406858,13.390542,13.372412,13.354282,13.337966,11.483305,9.626831,7.7721705,5.91751,4.062849,3.5932918,3.1219215,2.6523643,2.182807,1.7132497,1.6026589,1.4920682,1.3832904,1.2726997,1.162109,1.9670644,2.7720199,3.576975,4.3819304,5.186886,4.708264,4.227829,3.7473936,3.2669585,2.7883365,2.9007401,3.0131438,3.1255474,3.2379513,3.350355,3.8199122,4.2894692,4.76084,5.230397,5.6999545,6.755099,7.8102427,8.865387,9.920531,10.975676,14.340534,17.705393,21.070251,24.43511,27.799969,22.489801,17.179634,11.869466,6.5592985,1.2491312,1.5972201,1.9453088,2.2915847,2.6396735,2.9877625,2.467442,1.9471219,1.4268016,0.90829426,0.387974,4.604925,8.821876,13.04064,17.257591,21.474543,18.889257,16.305786,13.720501,11.135216,8.549932,6.869315,5.1905117,3.5098956,1.8292793,0.15047589,0.15047589,0.15047589,0.15047589,0.15047589,0.15047589,0.19942589,0.25018883,0.2991388,0.34990177,0.40066472,0.3770962,0.35534066,0.33177215,0.3100166,0.28826106,0.533011,0.7777609,1.0225109,1.2672608,1.5120108,4.762653,8.013294,11.262123,14.512766,17.763407,21.104698,24.4478,27.790903,31.132193,34.475296,31.309864,28.144432,24.980812,21.815378,18.649946,16.207886,13.765825,11.321951,8.87989,6.43783,5.9483304,5.4570174,4.9675174,4.478018,3.9867048,3.4482548,2.907992,2.3677292,1.8274662,1.2872034,1.3017071,1.3180238,1.3325275,1.3470312,1.3633479,5.282973,9.202598,13.122223,17.04185,20.963285,20.664148,20.366821,20.069496,19.77217,19.474844,17.545853,15.6150465,13.684241,11.755249,9.824444,10.297627,10.770811,11.242181,11.715364,12.186734,12.681673,13.176612,13.673364,14.168303,14.663241,13.466686,12.271944,11.077202,9.882459,8.6877165,9.255174,9.822631,10.390089,10.957546,11.525003,11.452485,11.379966,11.307447,11.234929,11.162411,10.15803,9.151835,8.147454,7.1430726,6.1368785,6.4704633,6.8022356,7.135821,7.4675927,7.799365,7.1050005,6.4106355,5.714458,5.0200934,4.325729,4.360175,4.3946214,4.4290676,4.465327,4.499773,4.2405195,3.9794528,3.720199,3.4591327,3.199879,4.856927,6.5157876,8.172835,9.829884,11.486931,10.203354,8.917963,7.6325727,6.347182,5.0617914,5.1941376,5.328297,5.4606433,5.5929894,5.7253356,5.529536,5.335549,5.139749,4.945762,4.749962,4.233268,3.7147603,3.198066,2.6795588,2.1628644,2.6016014,3.0421512,3.482701,3.923251,4.361988,4.077353,3.7927177,3.5080826,3.2216346,2.9369993,2.5852847,2.231757,1.8800422,1.5283275,1.1747998,3.6531196,6.1296263,8.607946,11.084454,13.562773,12.460492,11.358211,10.254116,9.151835,8.049554,10.40278,12.754191,15.107417,17.460642,19.812056,19.942589,20.073122,20.201841,20.332375,20.462908,20.865387,21.267864,21.670341,22.072819,22.475298,18.57924,14.684997,10.790753,6.8946967,3.000453,3.9051213,4.8097897,5.714458,6.6191263,7.5256076,7.2844834,7.0451727,6.8058615,6.5647373,6.3254266,5.4443264,4.5650396,3.6857529,2.8046532,1.9253663,3.5951047,5.2648435,6.9345818,8.604321,10.275872,12.565643,14.855415,17.145187,19.43496,21.724731,22.810696,23.894846,24.980812,26.064962,27.149115,25.390541,23.630154,21.869768,20.10938,18.350807,19.920834,21.490858,23.060884,24.630909,26.199121,21.634083,17.070856,12.504003,7.9407763,3.3757362,2.7303216,2.084907,1.4394923,0.79407763,0.15047589,0.12690738,0.10515183,0.08339628,0.059827764,0.038072214,0.56745726,1.0968424,1.6280404,2.1574254,2.6868105,2.3133402,1.938057,1.5627737,1.1874905,0.8122072,0.6508536,0.48768693,0.3245203,0.16316663,0.0,0.11965553,0.23931105,0.36077955,0.48043507,0.6000906,0.97174793,1.3452182,1.7168756,2.0903459,2.4620032,2.0268922,1.5917811,1.1566701,0.72337204,0.28826106,0.48043507,0.6726091,0.86478317,1.0569572,1.2491312,1.2382535,1.2255627,1.2128719,1.2001812,1.1874905,1.4576219,1.7277533,1.9978848,2.268016,2.5381477,2.3024626,2.0667772,1.8329052,1.5972201,1.3633479,1.2908293,1.2183108,1.1457924,1.0732739,1.0007553,0.85934424,0.7197462,0.58014804,0.4405499,0.2991388,0.29007402,0.27919623,0.27013144,0.25925365,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.06707962,0.13415924,0.2030518,0.27013144,0.33721104,0.33721104,0.33721104,0.33721104,0.33721104,0.33721104,0.27919623,0.2229944,0.16497959,0.10696479,0.05076295,0.14684997,0.24474995,0.34264994,0.4405499,0.53663695,0.7668832,0.99712944,1.2273756,1.4576219,1.6878681,1.7875811,1.887294,1.987007,2.08672,2.1882458,4.3728657,6.5574856,8.7421055,10.926725,13.113158,13.4050455,13.696932,13.990632,14.282519,14.574407,16.880495,19.18477,21.490858,23.795134,26.09941,23.470613,20.840004,18.209396,15.580601,12.949992,17.980963,23.01012,28.041092,33.07025,38.099407,32.437527,26.775644,21.11195,15.4500675,9.788185,10.1054535,10.422722,10.73999,11.057259,11.374527,14.432995,17.48965,20.548119,23.604773,26.66324,26.955128,27.247015,27.540714,27.832602,28.124489,26.617916,25.109531,23.60296,22.094576,20.588003,22.649342,24.712494,26.775644,28.836983,30.900135,27.693003,24.485872,21.276928,18.069798,14.862667,12.375282,9.8878975,7.400513,4.9131284,2.4257438,2.124792,1.8256533,1.5247015,1.2255627,0.9246109,1.2128719,1.49932,1.7875811,2.0758421,2.3622901,2.277081,2.1918716,2.1066625,2.0232663,1.938057,1.5718386,1.2074331,0.8430276,0.47680917,0.11240368,0.15954071,0.20667773,0.25562772,0.30276474,0.34990177,0.3100166,0.27013144,0.23024625,0.19036107,0.15047589,0.38978696,0.629098,0.87022203,1.1095331,1.3506571,1.2980812,1.2455053,1.1929294,1.1403534,1.0877775,0.95180535,0.81764615,0.68167394,0.5475147,0.41335547,0.34990177,0.28826106,0.22480737,0.16316663,0.099712946,0.18673515,0.2755703,0.36259252,0.44961473,0.53663695,0.5982776,0.65810543,0.7179332,0.7777609,0.8375887,0.8103943,0.78319985,0.7541924,0.726998,0.69980353,1.5573349,2.4148662,3.2723975,4.1299286,4.98746,4.8678045,4.748149,4.6266804,4.507025,4.3873696,3.6948178,3.002266,2.3097143,1.6171626,0.9246109,0.79770356,0.67079616,0.5420758,0.41516843,0.28826106,0.24837588,0.20667773,0.16679256,0.12690738,0.0870222,0.15228885,0.21755551,0.28282216,0.3480888,0.41335547,0.38978696,0.3680314,0.3444629,0.32270733,0.2991388,0.24293698,0.18492219,0.12690738,0.07070554,0.012690738,0.02175555,0.032633327,0.04169814,0.052575916,0.06164073,0.059827764,0.058014803,0.054388877,0.052575916,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.059827764,0.07070554,0.07977036,0.09064813,0.099712946,0.09789998,0.09427405,0.092461094,0.09064813,0.0870222,0.08339628,0.07795739,0.072518505,0.06707962,0.06164073,0.065266654,0.06707962,0.07070554,0.072518505,0.07433146,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.059827764,0.11965553,0.1794833,0.23931105,0.2991388,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.36984438,0.73968875,1.1095331,1.4793775,1.8492218,1.892733,1.9344311,1.9779422,2.0196402,2.0631514,1.8020848,1.5428312,1.2817645,1.0225109,0.76325727,1.7368182,2.712192,3.6875658,4.6629395,5.638314,6.755099,7.8718834,8.990481,10.107266,11.225864,11.227677,11.22949,11.233116,11.234929,11.236742,9.864329,8.491917,7.119504,5.7470913,4.3746786,3.8978696,3.4192474,2.9424384,2.465629,1.987007,1.8546607,1.7223145,1.5899682,1.4576219,1.3252757,2.0975976,2.8699198,3.6422417,4.4145637,5.186886,4.764466,4.3420453,3.919625,3.4972048,3.0747845,2.9750717,2.8753586,2.7756457,2.6741197,2.5744069,3.8017826,5.029158,6.258347,7.4857225,8.713099,9.110137,9.507175,9.904215,10.303066,10.700105,12.730623,14.759329,16.789846,18.820364,20.84907,16.880495,12.910107,8.939718,4.9693303,1.0007553,1.9942589,2.9895754,3.9848917,4.9802084,5.975525,4.8732433,3.7691493,2.666868,1.5645868,0.46230546,3.5969179,6.73153,9.867955,13.002567,16.13718,14.405801,12.672608,10.939416,9.208037,7.474845,6.0407915,4.604925,3.1690586,1.7350051,0.2991388,0.26287958,0.22480737,0.18673515,0.15047589,0.11240368,0.2374981,0.36259252,0.48768693,0.61278135,0.73787576,0.6544795,0.5728962,0.4894999,0.40791658,0.3245203,0.6653573,1.0043813,1.3452182,1.6842422,2.0250793,4.574105,7.124943,9.675781,12.224807,14.775645,17.496902,20.219973,22.94304,25.664299,28.387367,25.7205,23.051819,20.38495,17.718082,15.049402,13.67699,12.304577,10.932164,9.5597515,8.187339,7.85738,7.5274205,7.1974616,6.867502,6.5375433,5.4443264,4.3529234,3.2597067,2.1683033,1.0750868,1.167548,1.260009,1.35247,1.4449311,1.5373923,5.139749,8.7421055,12.344462,15.946819,19.549175,19.518354,19.485722,19.453089,19.420456,19.387821,18.102432,16.817041,15.531651,14.248073,12.962683,13.894546,14.828221,15.760084,16.691946,17.625622,17.139748,16.655687,16.169813,15.685752,15.199879,14.7974,14.394923,13.992445,13.589968,13.1874895,12.96087,12.732436,12.5058155,12.277383,12.050762,12.255627,12.460492,12.665357,12.870221,13.075087,12.264692,11.454298,10.645717,9.835322,9.024928,8.789243,8.55537,8.319685,8.0858135,7.850128,7.75948,7.6706448,7.5799966,7.4893484,7.400513,7.494787,7.590874,7.6851482,7.7794223,7.8755093,6.8421206,5.810545,4.7771564,3.7455807,2.712192,4.853301,6.9925966,9.131892,11.273002,13.412297,12.192173,10.97205,9.751925,8.531802,7.311678,7.1521373,6.9925966,6.833056,6.6717024,6.5121617,6.1223745,5.732588,5.3428006,4.953014,4.5632267,3.97764,3.392053,2.808279,2.222692,1.6371052,2.617918,3.5969179,4.5777307,5.5567303,6.5375433,5.8558693,5.1723824,4.4907084,3.8072214,3.1255474,2.9206827,2.715818,2.5091403,2.3042755,2.0994108,4.880495,7.6597667,10.440851,13.220123,15.999394,14.969632,13.939869,12.910107,11.880343,10.850581,12.629097,14.409427,16.189756,17.970085,19.750414,20.085812,20.419397,20.754795,21.090193,21.425592,21.40565,21.385706,21.365765,21.345821,21.325878,18.00997,14.695875,11.379966,8.064057,4.749962,5.1596913,5.569421,5.979151,6.390693,6.8004227,6.394319,5.9900284,5.5857377,5.179634,4.7753434,4.4272547,4.079166,3.73289,3.3848011,3.0367124,4.4145637,5.7924156,7.170267,8.548119,9.924157,12.067079,14.210001,16.352922,18.495844,20.636953,21.808126,22.977488,24.146849,25.318022,26.487383,24.641787,22.798004,20.952408,19.106813,17.26303,18.765976,20.267109,21.770054,23.273,24.774134,20.945156,17.114367,13.28539,9.4546,5.6256227,4.559601,3.4953918,2.42937,1.3651608,0.2991388,0.25562772,0.21030366,0.16497959,0.11965553,0.07433146,1.1349145,2.1954978,3.254268,4.314851,5.375434,4.6248674,3.874301,3.1255474,2.374981,1.6244144,1.2998942,0.97537386,0.6508536,0.3245203,0.0,0.19036107,0.38072214,0.56927025,0.75963134,0.9499924,1.7205015,2.4891977,3.2597067,4.0302157,4.800725,3.930503,3.0602808,2.1900587,1.3198367,0.44961473,0.5475147,0.64541465,0.7433147,0.83940166,0.93730164,0.93730164,0.93730164,0.93730164,0.93730164,0.93730164,1.7658255,2.5925364,3.4192474,4.2477713,5.0744824,4.592234,4.1099863,3.6277382,3.1454902,2.663242,2.5308957,2.3967366,2.2643902,2.132044,1.9996977,1.7205015,1.4394923,1.1602961,0.8792868,0.6000906,0.58014804,0.56020546,0.5402629,0.52032024,0.50037766,0.40066472,0.2991388,0.19942589,0.099712946,0.0,0.13415924,0.27013144,0.40429065,0.5402629,0.6744221,0.6744221,0.6744221,0.6744221,0.6744221,0.6744221,0.56020546,0.44417584,0.32995918,0.21574254,0.099712946,0.2955129,0.4894999,0.6852999,0.8792868,1.0750868,1.5101979,1.9453088,2.38042,2.8155308,3.2506418,3.2252605,3.199879,3.1744974,3.149116,3.1255474,5.3953767,7.665206,9.935035,12.2048645,14.474693,14.47288,14.4692545,14.467442,14.465629,14.462003,16.80979,19.157576,21.505362,23.85315,26.199121,24.45324,22.705544,20.957848,19.210152,17.462456,20.198215,22.932163,25.667925,28.401873,31.137632,28.574102,26.012386,23.45067,20.887142,18.325426,16.597672,14.869919,13.142166,11.4144125,9.686659,12.514881,15.343102,18.169512,20.997732,23.82414,24.746939,25.669737,26.592535,27.515333,28.438131,27.159992,25.881853,24.605528,23.327389,22.049252,23.45067,24.850279,26.249886,27.649492,29.049099,27.198065,25.345217,23.492369,21.63952,19.786674,16.624866,13.46306,10.29944,7.137634,3.975827,3.5497808,3.1255474,2.6995013,2.275268,1.8492218,2.4130533,2.9750717,3.53709,4.100921,4.6629395,4.3547363,4.0483456,3.7401419,3.4319382,3.1255474,2.5453994,1.9652514,1.3851035,0.80495536,0.22480737,0.2955129,0.36440548,0.43511102,0.5058166,0.5747091,0.52032024,0.46411842,0.40972954,0.35534066,0.2991388,0.44236287,0.5855869,0.726998,0.87022203,1.0116332,1.0080072,1.0025684,0.99712944,0.9916905,0.9880646,0.90466833,0.823085,0.73968875,0.65810543,0.5747091,0.48768693,0.40066472,0.31182957,0.22480737,0.13778515,0.19942589,0.26287958,0.3245203,0.387974,0.44961473,0.533011,0.61459434,0.6979906,0.7795739,0.8629702,0.8448406,0.82671094,0.8103943,0.79226464,0.774135,1.551896,2.3296568,3.1074178,3.8851788,4.6629395,4.421816,4.1825047,3.9431937,3.7020695,3.4627585,2.9279346,2.3931105,1.8582866,1.3216497,0.7868258,0.7070554,0.62728506,0.5475147,0.46774435,0.387974,0.33177215,0.27738327,0.2229944,0.16679256,0.11240368,0.15410182,0.19761293,0.23931105,0.28282216,0.3245203,0.3045777,0.28463513,0.26469254,0.24474995,0.22480737,0.18492219,0.14503701,0.10515183,0.065266654,0.025381476,0.032633327,0.03988518,0.047137026,0.054388877,0.06164073,0.058014803,0.052575916,0.047137026,0.04169814,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.058014803,0.07795739,0.09789998,0.11784257,0.13778515,0.13234627,0.12690738,0.12328146,0.11784257,0.11240368,0.10333887,0.092461094,0.08339628,0.072518505,0.06164073,0.06707962,0.072518505,0.07795739,0.08339628,0.0870222,0.07433146,0.06164073,0.05076295,0.038072214,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.045324065,0.09064813,0.13415924,0.1794833,0.22480737,0.19942589,0.17585737,0.15047589,0.12509441,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.25562772,0.5094425,0.7650702,1.020698,1.2745126,1.2944553,1.3143979,1.3343405,1.3542831,1.3742256,1.2726997,1.1693609,1.067835,0.9644961,0.8629702,1.7495089,2.6378605,3.5243993,4.4127507,5.2992897,6.0444174,6.789545,7.5346723,8.2798,9.024928,9.046683,9.070251,9.092008,9.115576,9.137331,8.247167,7.3570023,6.4668374,5.576673,4.688321,4.2024474,3.7183862,3.2325122,2.7466383,2.2625773,2.1066625,1.9525607,1.7966459,1.6425442,1.4866294,2.228131,2.9678197,3.7075086,4.4471974,5.186886,4.8224807,4.458075,4.0918565,3.727451,3.3630457,3.049403,2.7375734,2.4257438,2.1121013,1.8002719,3.785466,5.77066,7.755854,9.739235,11.724429,11.465176,11.205922,10.944855,10.685601,10.424535,11.120712,11.815077,12.509441,13.20562,13.899984,11.269376,8.640579,6.009971,3.3793623,0.7505665,2.3931105,4.0356545,5.678199,7.320743,8.963287,7.2772317,5.5929894,3.9069343,2.222692,0.53663695,2.5907235,4.6429973,6.695271,8.747544,10.799818,9.920531,9.039432,8.160145,7.2790446,6.399758,5.2104545,4.019338,2.8300345,1.6407311,0.44961473,0.37528324,0.2991388,0.22480737,0.15047589,0.07433146,0.2755703,0.4749962,0.6744221,0.87566096,1.0750868,0.9318628,0.7904517,0.64722764,0.5058166,0.36259252,0.79770356,1.2328146,1.6679256,2.1030366,2.5381477,4.3873696,6.2365913,8.087626,9.936848,11.787883,13.889107,15.992143,18.095179,20.198215,22.29944,20.129324,17.959208,15.789091,13.618975,11.450671,11.147907,10.845142,10.542377,10.239613,9.936848,9.768243,9.597824,9.427405,9.256987,9.088382,7.4422116,5.7978544,4.1516843,2.5073273,0.8629702,1.0333886,1.2019942,1.3724127,1.5428312,1.7132497,4.9983377,8.281613,11.566701,14.851789,18.136877,18.37075,18.60281,18.834867,19.066927,19.3008,18.660824,18.020847,17.380873,16.740896,16.100922,17.493277,18.885632,20.277987,21.670341,23.062696,21.597824,20.13295,18.668076,17.203201,15.738328,16.128115,16.517902,16.907688,17.297476,17.687263,16.664753,15.6422415,14.61973,13.597219,12.574709,13.056956,13.539205,14.023266,14.505513,14.9877615,14.373167,13.75676,13.142166,12.527572,11.912977,11.109835,10.306692,9.5053625,8.70222,7.900891,8.415772,8.930654,9.445535,9.960417,10.475298,10.629399,10.785315,10.939416,11.095331,11.249433,9.445535,7.6398244,5.8341136,4.0302157,2.2245052,4.847862,7.4694057,10.092763,12.714307,15.337664,14.182806,13.027949,11.873092,10.718235,9.563377,9.110137,8.656897,8.205468,7.752228,7.3008003,6.7152133,6.1296263,5.5458527,4.9602656,4.3746786,3.7220123,3.0693457,2.4166791,1.7658255,1.1131591,2.6324217,4.1516843,5.67276,7.192023,8.713099,7.6325727,6.552047,5.473334,4.3928084,3.3122826,3.254268,3.198066,3.1400511,3.0820365,3.0258346,6.107871,9.189907,12.271944,15.355793,18.43783,17.480585,16.52334,15.564283,14.607039,13.649796,14.857228,16.064661,17.272095,18.479528,19.68696,20.227224,20.767487,21.307749,21.848013,22.388275,21.945911,21.501736,21.059374,20.61701,20.174648,17.4407,14.70494,11.969179,9.235231,6.4994707,6.414262,6.3308654,6.245656,6.1604466,6.0752378,5.504154,4.934884,4.365614,3.7945306,3.2252605,3.4101827,3.5951047,3.780027,3.9649491,4.1498713,5.235836,6.319988,7.404139,8.490104,9.574255,11.570327,13.564586,15.5606575,17.554916,19.549175,20.80556,22.06013,23.3147,24.56927,25.825651,23.894846,21.965855,20.03505,18.104244,16.175253,17.609306,19.045172,20.479225,21.915092,23.349146,20.254417,17.15969,14.064963,10.970237,7.8755093,6.390693,4.9058766,3.4192474,1.9344311,0.44961473,0.3825351,0.3154555,0.24837588,0.1794833,0.11240368,1.7023718,3.29234,4.882308,6.472276,8.062244,6.9382076,5.812358,4.688321,3.5624714,2.4366217,1.9507477,1.4630609,0.97537386,0.48768693,0.0,0.25925365,0.52032024,0.7795739,1.0406405,1.2998942,2.467442,3.63499,4.802538,5.9700856,7.137634,5.8323007,4.5269675,3.2216346,1.9181144,0.61278135,0.61459434,0.61822027,0.6200332,0.62184614,0.62547207,0.63816285,0.6508536,0.66173136,0.6744221,0.6871128,2.0722163,3.4573197,4.842423,6.2275267,7.61263,6.882006,6.153195,5.422571,4.691947,3.9631362,3.7691493,3.576975,3.3848011,3.1926272,3.000453,2.5798457,2.1592383,1.7404441,1.3198367,0.89922947,0.87022203,0.83940166,0.8103943,0.7795739,0.7505665,0.6000906,0.44961473,0.2991388,0.15047589,0.0,0.2030518,0.40429065,0.6073425,0.8103943,1.0116332,1.0116332,1.0116332,1.0116332,1.0116332,1.0116332,0.83940166,0.6671702,0.4949388,0.32270733,0.15047589,0.44236287,0.73424983,1.0279498,1.3198367,1.6117238,2.2516994,2.8916752,3.531651,4.17344,4.8134155,4.6629395,4.512464,4.361988,4.213325,4.062849,6.4178877,8.772926,11.127964,13.483003,15.838041,15.540715,15.243389,14.94425,14.646925,14.349599,16.740896,19.13038,21.519865,23.909351,26.300648,25.435865,24.56927,23.704485,22.839703,21.97492,22.41547,22.854206,23.294756,23.735306,24.174044,24.712494,25.24913,25.78758,26.326029,26.862667,23.089891,19.317116,15.544341,11.771566,8.000604,10.596766,13.194741,15.792717,18.390692,20.986855,22.540564,24.09246,25.644356,27.198065,28.74996,27.702068,26.654177,25.608097,24.560204,23.512312,24.250187,24.988064,25.724127,26.462002,27.199877,26.703125,26.204561,25.70781,25.209244,24.712494,20.87445,17.038223,13.200181,9.362139,5.52591,4.974769,4.4254417,3.874301,3.3249733,2.7756457,3.6132345,4.4508233,5.2884116,6.1241875,6.9617763,6.432391,5.903006,5.371808,4.842423,4.313038,3.5171473,2.72307,1.9271792,1.1331016,0.33721104,0.42967212,0.52213323,0.61459434,0.7070554,0.7995165,0.7306239,0.65991837,0.58921283,0.52032024,0.44961473,0.4949388,0.5402629,0.5855869,0.629098,0.6744221,0.7179332,0.75963134,0.8031424,0.8448406,0.8883517,0.8575313,0.82671094,0.79770356,0.7668832,0.73787576,0.62547207,0.51306844,0.40066472,0.28826106,0.17585737,0.21211663,0.25018883,0.28826106,0.3245203,0.36259252,0.46774435,0.5728962,0.678048,0.78319985,0.8883517,0.8792868,0.872035,0.86478317,0.8575313,0.85027945,1.54827,2.2444477,2.9424384,3.6404288,4.3366065,3.97764,3.6168604,3.2578938,2.8971143,2.5381477,2.1592383,1.7821422,1.405046,1.0279498,0.6508536,0.61822027,0.5855869,0.5529536,0.52032024,0.48768693,0.4169814,0.3480888,0.27738327,0.20667773,0.13778515,0.15772775,0.17767033,0.19761293,0.21755551,0.2374981,0.21936847,0.2030518,0.18492219,0.16679256,0.15047589,0.12690738,0.10515183,0.08339628,0.059827764,0.038072214,0.04169814,0.047137026,0.052575916,0.058014803,0.06164073,0.054388877,0.047137026,0.03988518,0.032633327,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.054388877,0.08520924,0.11421664,0.14503701,0.17585737,0.16679256,0.15954071,0.15228885,0.14503701,0.13778515,0.12328146,0.10696479,0.092461094,0.07795739,0.06164073,0.07070554,0.07795739,0.08520924,0.092461094,0.099712946,0.0870222,0.07433146,0.06164073,0.05076295,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.15047589,0.15047589,0.15047589,0.15047589,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13959812,0.27919623,0.42060733,0.56020546,0.69980353,0.6979906,0.69436467,0.69255173,0.69073874,0.6871128,0.7433147,0.79770356,0.8520924,0.90829426,0.96268314,1.7621996,2.561716,3.3630457,4.162562,4.9620786,5.335549,5.7072062,6.0806766,6.452334,6.825804,6.867502,6.9092,6.9527116,6.9944096,7.037921,6.630004,6.2220874,5.814171,5.408067,5.0001507,4.507025,4.0157123,3.5225863,3.0294604,2.5381477,2.3604772,2.182807,2.0051367,1.8274662,1.649796,2.3568513,3.0657198,3.7727752,4.4798307,5.186886,4.880495,4.572292,4.264088,3.9576974,3.6494937,3.1255474,2.5997884,2.0758421,1.550083,1.0243238,3.7673361,6.510349,9.253361,11.99456,14.737573,13.820213,12.902855,11.985496,11.068136,10.150778,9.510801,8.870826,8.229037,7.5890613,6.9490857,5.660069,4.36924,3.0802233,1.789394,0.50037766,2.7901495,5.0799212,7.369693,9.659465,11.949236,9.683033,7.415017,5.147001,2.8807976,0.61278135,1.5827163,2.5526514,3.5225863,4.4925213,5.462456,5.4352617,5.408067,5.37906,5.351866,5.3246713,4.3801174,3.435564,2.4891977,1.5446441,0.6000906,0.48768693,0.37528324,0.26287958,0.15047589,0.038072214,0.31182957,0.5873999,0.8629702,1.1367276,1.4122978,1.209246,1.0080072,0.80495536,0.60190356,0.40066472,0.9300498,1.4594349,1.9906329,2.520018,3.049403,4.2006345,5.3500524,6.4994707,7.650702,8.80012,10.283124,11.764315,13.247317,14.730321,16.211512,14.53996,12.866595,11.195044,9.52168,7.850128,8.617011,9.385707,10.152591,10.919474,11.6881695,11.677292,11.668227,11.65735,11.648285,11.637406,9.440096,7.2427855,5.045475,2.8481643,0.6508536,0.8974165,1.1457924,1.3923552,1.6407311,1.887294,4.855114,7.8229337,10.790753,13.75676,16.72458,17.223145,17.719896,18.216648,18.715212,19.211964,19.217403,19.222843,19.228281,19.231907,19.237347,21.090193,22.94304,24.795889,26.646925,28.499771,26.055899,23.610212,21.164526,18.720652,16.274965,17.457016,18.64088,19.822933,21.004984,22.187037,20.370447,18.552046,16.735458,14.917056,13.100468,13.860099,14.61973,15.379361,16.140806,16.900436,16.47983,16.059223,15.640429,15.219821,14.799213,13.430427,12.059827,10.689227,9.32044,7.949841,9.070251,10.190662,11.30926,12.429671,13.550082,13.765825,13.979754,14.195497,14.409427,14.625169,12.047136,9.470917,6.892884,4.314851,1.7368182,4.842423,7.948028,11.05182,14.157425,17.26303,16.173439,15.082036,13.992445,12.902855,11.813264,11.068136,10.323009,9.577881,8.832754,8.087626,7.308052,6.526665,5.7470913,4.9675174,4.1879435,3.4681973,2.7466383,2.0268922,1.3071461,0.5873999,2.6469254,4.708264,6.7677894,8.827314,10.88684,9.409276,7.931711,6.454147,4.976582,3.5008307,3.589666,3.680314,3.7691493,3.8597972,3.9504454,7.3352466,10.720048,14.104849,17.48965,20.87445,19.989725,19.105,18.220274,17.335548,16.450823,17.08536,17.719896,18.354433,18.990784,19.62532,20.370447,21.115576,21.860703,22.605831,23.349146,22.484362,21.61958,20.754795,19.890013,19.025229,16.869617,14.715817,12.5602045,10.4045925,8.2507925,7.6706448,7.0904965,6.510349,5.9302006,5.3500524,4.615803,3.87974,3.1454902,2.4094272,1.6751775,2.3931105,3.1092308,3.827164,4.5450974,5.2630305,6.055295,6.8475595,7.6398244,8.432089,9.224354,11.071762,12.919171,14.7683935,16.615803,18.463211,19.80299,21.142769,22.48255,23.822329,25.162107,23.147905,21.131891,19.117691,17.101677,15.087475,16.454449,17.823235,19.190208,20.557182,21.924156,19.565493,17.205015,14.844538,12.485873,10.125396,8.219973,6.3145485,4.409125,2.5055144,0.6000906,0.5094425,0.42060733,0.32995918,0.23931105,0.15047589,2.269829,4.3891826,6.510349,8.629702,10.750868,9.249735,7.750415,6.249282,4.749962,3.2506418,2.5997884,1.9507477,1.2998942,0.6508536,0.0,0.32995918,0.65991837,0.9898776,1.3198367,1.649796,3.2143826,4.780782,6.345369,7.909956,9.474543,7.7340984,5.995467,4.255023,2.514579,0.774135,0.68167394,0.58921283,0.49675176,0.40429065,0.31182957,0.33721104,0.36259252,0.387974,0.41335547,0.43692398,2.38042,4.322103,6.265599,8.207282,10.150778,9.171778,8.194591,7.217404,6.240217,5.2630305,5.009216,4.7572136,4.505212,4.25321,3.9993954,3.43919,2.8807976,2.3205922,1.7603867,1.2001812,1.1602961,1.1204109,1.0805258,1.0406405,1.0007553,0.7995165,0.6000906,0.40066472,0.19942589,0.0,0.27013144,0.5402629,0.8103943,1.0805258,1.3506571,1.3506571,1.3506571,1.3506571,1.3506571,1.3506571,1.1204109,0.8901646,0.65991837,0.42967212,0.19942589,0.58921283,0.9808127,1.3705997,1.7603867,2.1501737,2.9950142,3.8398547,4.6846952,5.529536,6.3743763,6.1006193,5.825049,5.5494785,5.275721,5.0001507,7.440398,9.880646,12.320893,14.759329,17.199575,16.606737,16.01571,15.422873,14.830034,14.237195,16.67019,19.103188,21.53437,23.967365,26.400362,26.416677,26.434807,26.452936,26.469254,26.487383,24.632723,22.778063,20.921589,19.066927,17.212267,20.850883,24.487686,28.124489,31.763105,35.399906,29.582111,23.766127,17.946516,12.130532,6.3127356,8.680465,11.048194,13.415923,15.781839,18.149569,20.332375,22.515182,24.697989,26.880796,29.06179,28.244144,27.42831,26.610664,25.793018,24.975372,25.049704,25.125849,25.20018,25.274511,25.350657,26.208187,27.065718,27.92325,28.78078,29.638311,25.124035,20.613384,16.099108,11.586644,7.07418,6.399758,5.7253356,5.049101,4.3746786,3.7002566,4.8134155,5.924762,7.037921,8.149267,9.262425,8.510046,7.757667,7.0052876,6.2529078,5.5005283,4.4907084,3.4808881,2.469255,1.4594349,0.44961473,0.5656443,0.67986095,0.79589057,0.9101072,1.0243238,0.93911463,0.8557183,0.7705091,0.6852999,0.6000906,0.5475147,0.4949388,0.44236287,0.38978696,0.33721104,0.42785916,0.5166943,0.6073425,0.6979906,0.7868258,0.8103943,0.8321498,0.8557183,0.8774739,0.89922947,0.76325727,0.62547207,0.48768693,0.34990177,0.21211663,0.22480737,0.2374981,0.25018883,0.26287958,0.2755703,0.40247768,0.5293851,0.65810543,0.7850128,0.9119202,0.9155461,0.91735905,0.91917205,0.922798,0.9246109,1.5428312,2.1592383,2.7774587,3.395679,4.0120864,3.531651,3.053029,2.572594,2.0921588,1.6117238,1.3923552,1.1729867,0.95180535,0.7324369,0.51306844,0.5275721,0.5420758,0.55839247,0.5728962,0.5873999,0.50219065,0.4169814,0.33177215,0.24837588,0.16316663,0.15954071,0.15772775,0.15410182,0.15228885,0.15047589,0.13415924,0.11965553,0.10515183,0.09064813,0.07433146,0.07070554,0.065266654,0.059827764,0.054388877,0.05076295,0.052575916,0.054388877,0.058014803,0.059827764,0.06164073,0.052575916,0.04169814,0.032633327,0.02175555,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.052575916,0.092461094,0.13234627,0.17223145,0.21211663,0.2030518,0.19217403,0.18310922,0.17223145,0.16316663,0.14322405,0.12328146,0.10333887,0.08339628,0.06164073,0.072518505,0.08339628,0.092461094,0.10333887,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.099712946,0.12509441,0.15047589,0.17585737,0.19942589,0.15954071,0.11965553,0.07977036,0.03988518,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.21211663,0.42423326,0.63816285,0.85027945,1.062396,1.7748904,2.4873846,3.199879,3.9123733,4.6248674,4.6248674,4.6248674,4.6248674,4.6248674,4.6248674,4.688321,4.749962,4.8116026,4.8750563,4.936697,5.0128417,5.087173,5.163317,5.237649,5.3119802,4.8116026,4.313038,3.8126602,3.3122826,2.811905,2.612479,2.4130533,2.2118144,2.0123885,1.8129625,2.4873846,3.1618068,3.8380418,4.512464,5.186886,4.936697,4.688321,4.4381323,4.1879435,3.9377546,3.199879,2.4620032,1.7241274,0.9880646,0.25018883,3.7492065,7.250037,10.750868,14.249886,17.750717,16.175253,14.599788,13.024323,11.450671,9.875207,7.900891,5.924762,3.9504454,1.9743162,0.0,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,3.1871881,6.1241875,9.063,11.999999,14.936998,12.087022,9.237044,6.3870673,3.53709,0.6871128,0.5747091,0.46230546,0.34990177,0.2374981,0.12509441,0.9499924,1.7748904,2.5997884,3.4246864,4.249584,3.5497808,2.8499773,2.1501737,1.4503701,0.7505665,0.6000906,0.44961473,0.2991388,0.15047589,0.0,0.34990177,0.69980353,1.0497054,1.3996071,1.7495089,1.4866294,1.2255627,0.96268314,0.69980353,0.43692398,1.062396,1.6878681,2.3133402,2.9369993,3.5624714,4.0120864,4.461701,4.9131284,5.3627434,5.812358,6.6753283,7.5382986,8.399456,9.262425,10.125396,8.950596,7.7757964,6.599184,5.424384,4.249584,6.0879283,7.9244595,9.762803,11.599335,13.437678,13.588155,13.736817,13.887294,14.037769,14.188245,11.437981,8.6877165,5.9374523,3.1871881,0.43692398,0.76325727,1.0877775,1.4122978,1.7368182,2.0631514,4.7118897,7.362441,10.012992,12.661731,15.312282,16.075539,16.836983,17.60024,18.361685,19.124943,19.775795,20.424837,21.07569,21.724731,22.375584,24.68711,27.000452,29.31198,31.625319,33.936848,30.51216,27.087475,23.662788,20.238102,16.811602,18.787731,20.762047,22.738176,24.712494,26.68681,24.07433,21.461851,18.849373,16.236893,13.6244135,14.663241,15.700256,16.73727,17.774284,18.813112,18.588305,18.361685,18.136877,17.912071,17.687263,15.749206,13.812962,11.874905,9.936848,8.000604,9.724731,11.450671,13.174799,14.90074,16.624866,16.900436,17.174194,17.449764,17.725336,18.000906,14.650551,11.300196,7.949841,4.599486,1.2491312,4.836984,8.424837,12.012691,15.600543,19.188396,18.16226,17.137936,16.1118,15.087475,14.06315,13.024323,11.9873085,10.950294,9.91328,8.874452,7.900891,6.925517,5.9501433,4.974769,3.9993954,3.2125697,2.4257438,1.6371052,0.85027945,0.06164073,2.663242,5.2630305,7.8628187,10.462607,13.062395,11.187792,9.313189,7.4367723,5.562169,3.6875658,3.925064,4.162562,4.40006,4.6375585,4.8750563,8.562622,12.250188,15.937754,19.62532,23.312885,22.500679,21.686659,20.87445,20.062244,19.250036,19.311678,19.375132,19.436771,19.500225,19.561867,20.511858,21.461851,22.411844,23.361835,24.311829,23.024624,21.737421,20.450218,19.163015,17.87581,16.300346,14.724882,13.149418,11.575767,10.000301,8.925215,7.850128,6.775041,5.6999545,4.6248674,3.7256382,2.8245957,1.9253663,1.0243238,0.12509441,1.3742256,2.6251698,3.874301,5.125245,6.3743763,6.874754,7.3751316,7.8755093,8.375887,8.874452,10.57501,12.27557,13.974316,15.674874,17.375433,18.800423,20.22541,21.650398,23.075388,24.500376,22.399153,20.299742,18.20033,16.099108,13.999697,15.299591,16.599485,17.89938,19.199274,20.499168,18.874754,17.25034,15.624111,13.999697,12.375282,10.049252,7.7250338,5.4008155,3.0747845,0.7505665,0.63816285,0.52575916,0.41335547,0.2991388,0.18673515,2.8372865,5.487838,8.138389,10.7871275,13.437678,11.563075,9.686659,7.8120556,5.9374523,4.062849,3.2506418,2.4366217,1.6244144,0.8122072,0.0,0.40066472,0.7995165,1.2001812,1.6008459,1.9996977,3.9631362,5.924762,7.8882003,9.849826,11.813264,9.637709,7.462154,5.2865987,3.1128569,0.93730164,0.7505665,0.5620184,0.37528324,0.18673515,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,2.6868105,5.186886,7.686961,10.1870365,12.687112,11.46155,10.2378,9.012237,7.7866745,6.5629244,6.249282,5.9374523,5.6256227,5.3119802,5.0001507,4.3003473,3.6005437,2.9007401,2.1991236,1.49932,1.4503701,1.3996071,1.3506571,1.2998942,1.2491312,1.0007553,0.7505665,0.50037766,0.25018883,0.0,0.33721104,0.6744221,1.0116332,1.3506571,1.6878681,1.6878681,1.6878681,1.6878681,1.6878681,1.6878681,1.3996071,1.1131591,0.824898,0.53663695,0.25018883,0.73787576,1.2255627,1.7132497,2.1991236,2.6868105,3.738329,4.788034,5.8377395,6.887445,7.93715,7.5382986,7.137634,6.736969,6.338117,5.9374523,8.46291,10.986553,13.512011,16.037468,18.562923,17.674572,16.788034,15.899682,15.013144,14.124791,16.599485,19.074179,21.550686,24.025381,26.500074,27.399303,28.300346,29.199575,30.100618,30.999847,26.849976,22.700104,18.550234,14.400362,10.25049,16.98746,23.724428,30.463211,37.20018,43.93715,36.07433,28.213324,20.350506,12.487686,4.6248674,6.7623506,8.899834,11.037316,13.174799,15.312282,18.126,20.937904,23.74981,26.561714,29.375433,28.788033,28.200632,27.613234,27.025833,26.43662,25.84922,25.26182,24.674421,24.08702,23.49962,25.71325,27.925062,30.136877,32.350506,34.562317,29.375433,24.188547,18.999847,13.812962,8.624263,7.8247466,7.02523,6.2257137,5.424384,4.6248674,6.011784,7.400513,8.78743,10.174346,11.563075,10.587702,9.612328,8.636953,7.66158,6.688019,5.462456,4.2368937,3.0131438,1.7875811,0.5620184,0.69980353,0.8375887,0.97537386,1.1131591,1.2491312,1.1494182,1.0497054,0.9499924,0.85027945,0.7505665,0.6000906,0.44961473,0.2991388,0.15047589,0.0,0.13778515,0.2755703,0.41335547,0.5493277,0.6871128,0.76325727,0.8375887,0.9119202,0.9880646,1.062396,0.89922947,0.73787576,0.5747091,0.41335547,0.25018883,0.2374981,0.22480737,0.21211663,0.19942589,0.18673515,0.33721104,0.48768693,0.63816285,0.7868258,0.93730164,0.9499924,0.96268314,0.97537386,0.9880646,1.0007553,1.5373923,2.0758421,2.612479,3.149116,3.6875658,3.0874753,2.4873846,1.887294,1.2872034,0.6871128,0.62547207,0.5620184,0.50037766,0.43692398,0.37528324,0.43692398,0.50037766,0.5620184,0.62547207,0.6871128,0.5873999,0.48768693,0.387974,0.28826106,0.18673515,0.16316663,0.13778515,0.11240368,0.0870222,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,0.2374981,0.22480737,0.21211663,0.19942589,0.18673515,0.16316663,0.13778515,0.11240368,0.0870222,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.27738327,0.55476654,0.8321498,1.1095331,1.3869164,1.8818551,2.3767939,2.8717327,3.3666716,3.8616104,3.917812,3.972201,4.028403,4.082792,4.137181,4.207886,4.2767787,4.347484,4.41819,4.4870825,4.5668526,4.646623,4.7282066,4.8079767,4.8877473,4.5632267,4.2368937,3.9123733,3.587853,3.2633326,3.5044568,3.7473936,3.9903307,4.233268,4.4743915,4.5795436,4.6846952,4.7898474,4.894999,5.0001507,5.7833505,6.5647373,7.3479376,8.129324,8.912524,7.8120556,6.7115874,5.612932,4.512464,3.4119956,5.569421,7.7268467,9.884272,12.0416975,14.200936,13.327088,12.455053,11.583018,10.70917,9.837135,8.009668,6.1822023,4.3547363,2.5272698,0.69980353,1.4122978,2.124792,2.8372865,3.5497808,4.262275,5.8304877,7.3968873,8.9651,10.533313,12.099712,9.789998,7.4802837,5.1705694,2.8608549,0.5493277,0.4604925,0.36984438,0.27919623,0.19036107,0.099712946,0.7668832,1.4358664,2.1030366,2.770207,3.437377,2.8717327,2.3079014,1.742257,1.1766127,0.61278135,0.7505665,0.8883517,1.0243238,1.162109,1.2998942,1.3977941,1.4956942,1.5917811,1.6896812,1.7875811,1.6371052,1.4866294,1.3379664,1.1874905,1.0370146,1.4177368,1.7966459,2.1773682,2.5580902,2.9369993,3.303218,3.6676233,4.0320287,4.3982472,4.762653,5.482399,6.202145,6.921891,7.6416373,8.363196,7.5945,6.827617,6.060734,5.292038,4.5251546,6.6100616,8.694968,10.779876,12.864782,14.94969,14.347786,13.745882,13.142166,12.540262,11.938358,9.626831,7.317117,5.0074024,2.6976883,0.387974,0.6726091,0.9572442,1.2418793,1.5283275,1.8129625,4.3946214,6.978093,9.5597515,12.143224,14.724882,14.98051,15.234324,15.489952,15.74558,15.999394,16.659313,17.319231,17.980963,18.64088,19.3008,20.9651,22.629398,24.295511,25.959812,27.625923,25.087776,22.54963,20.013294,17.475147,14.936998,16.519714,18.102432,19.685148,21.267864,22.85058,20.656897,18.465023,16.273151,14.079468,11.887595,13.41411,14.942437,16.470764,17.99728,19.525606,19.235533,18.94546,18.655384,18.36531,18.075237,16.38737,14.699501,13.011633,11.325577,9.637709,10.959359,12.282822,13.604471,14.927934,16.249584,16.316664,16.385555,16.452635,16.519714,16.586794,13.9507475,11.312886,8.675026,6.037165,3.3993049,6.430578,9.460039,12.489499,15.520773,18.550234,17.369995,16.189756,15.009518,13.829279,12.650853,11.764315,10.879588,9.994863,9.110137,8.225411,7.420456,6.6155005,5.810545,5.0055895,4.2006345,3.6748753,3.149116,2.6251698,2.0994108,1.5754645,3.5824142,5.5893636,7.5981264,9.605076,11.612025,10.174346,8.736667,7.3008003,5.863121,4.4254417,5.087173,5.750717,6.412449,7.07418,7.7377243,11.024626,14.311526,17.60024,20.887142,24.175856,24.146849,24.119654,24.09246,24.065266,24.03807,23.414412,22.792566,22.17072,21.54706,20.925215,21.788185,22.649342,23.512312,24.375282,25.238253,24.509441,23.782444,23.055445,22.326633,21.599636,19.68696,17.774284,15.861609,13.9507475,12.038072,10.843329,9.646774,8.452031,7.2572894,6.0625467,4.95664,3.8525455,2.7466383,1.6425442,0.53663695,1.452183,2.3677292,3.2832751,4.1970086,5.1125546,5.924762,6.736969,7.549176,8.363196,9.175404,10.197914,11.220426,12.242936,13.265448,14.287958,15.455506,16.623055,17.790602,18.958149,20.125698,20.042301,19.960718,19.877321,19.795738,19.712341,19.099562,18.48678,17.87581,17.26303,16.650248,15.40293,14.155612,12.908294,11.6591625,10.411844,8.55537,6.697084,4.84061,2.9823234,1.1258497,0.969935,0.81583315,0.65991837,0.5058166,0.34990177,2.4384346,4.5251546,6.6118746,8.700407,10.7871275,9.353074,7.9172077,6.4831543,5.047288,3.6132345,3.3322253,3.053029,2.7720199,2.4928236,2.2118144,2.5816586,2.953316,3.3231604,3.6930048,4.062849,5.235836,6.4070096,7.5799966,8.752983,9.924157,8.089439,6.2547207,4.420003,2.5852847,0.7505665,0.6000906,0.44961473,0.2991388,0.15047589,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,2.9678197,5.7851634,8.602508,11.419851,14.237195,13.446743,12.658105,11.867653,11.077202,10.28675,9.271491,8.258044,7.2427855,6.2275267,5.2122674,4.6248674,4.0374675,3.4500678,2.8626678,2.275268,2.182807,2.0903459,1.9978848,1.9054236,1.8129625,1.455809,1.0968424,0.73968875,0.3825351,0.025381476,0.3245203,0.62547207,0.9246109,1.2255627,1.5247015,2.030518,2.5345216,3.0403383,3.5443418,4.0501585,4.3982472,4.744523,5.092612,5.4407005,5.7869763,6.3852544,6.981719,7.5799966,8.178274,8.774739,9.251548,9.73017,10.20698,10.685601,11.162411,11.418038,11.671853,11.927481,12.183108,12.436923,13.301706,14.168303,15.033086,15.897869,16.762651,17.047287,17.331923,17.61837,17.903006,18.187641,19.92446,21.66309,23.399908,25.136726,26.875357,28.2659,29.654629,31.045172,32.435715,33.824444,30.740593,27.654932,24.56927,21.48542,18.399757,23.233116,28.064661,32.898018,37.729565,42.562923,35.626526,28.691946,21.757364,14.8227825,7.8882003,10.1054535,12.322706,14.53996,16.757214,18.974466,21.438282,23.900286,26.36229,28.824291,31.288109,30.880192,30.472275,30.064358,29.658255,29.250338,28.929443,28.610363,28.289469,27.970387,27.649492,29.460642,31.26998,33.079315,34.890465,36.699802,31.80299,26.904366,22.007553,17.11074,12.212116,11.784257,11.358211,10.930351,10.502492,10.074633,11.557636,13.04064,14.521831,16.004833,17.487837,15.926876,14.367728,12.806767,11.24762,9.686659,8.345067,7.0016613,5.660069,4.3166637,2.9750717,3.2180085,3.4591327,3.7020695,3.9450066,4.1879435,3.874301,3.5624714,3.2506418,2.9369993,2.6251698,2.1719291,1.7205015,1.2672608,0.81583315,0.36259252,0.40429065,0.44780177,0.4894999,0.533011,0.5747091,0.65810543,0.73968875,0.823085,0.90466833,0.9880646,0.86478317,0.7433147,0.6200332,0.49675176,0.37528324,0.4749962,0.5747091,0.6744221,0.774135,0.87566096,0.872035,0.87022203,0.8665961,0.86478317,0.8629702,0.8665961,0.872035,0.8774739,0.88291276,0.8883517,1.4757515,2.0631514,2.6505513,3.2379513,3.825351,3.5642843,3.3050308,3.045777,2.7847104,2.525457,2.6269827,2.7303216,2.8318477,2.9351864,3.0367124,2.764768,2.4928236,2.2190661,1.9471219,1.6751775,1.3796645,1.0841516,0.7904517,0.4949388,0.19942589,0.22662032,0.25562772,0.28282216,0.3100166,0.33721104,0.2755703,0.21211663,0.15047589,0.0870222,0.025381476,0.030820364,0.034446288,0.03988518,0.045324065,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.04169814,0.034446288,0.027194439,0.01994259,0.012690738,0.014503701,0.018129626,0.01994259,0.02175555,0.025381476,0.065266654,0.10515183,0.14503701,0.18492219,0.22480737,0.24474995,0.26469254,0.28463513,0.3045777,0.3245203,0.3208944,0.3154555,0.3100166,0.3045777,0.2991388,0.26831847,0.23568514,0.2030518,0.17041849,0.13778515,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03988518,0.07977036,0.11965553,0.15954071,0.19942589,0.15954071,0.11965553,0.07977036,0.03988518,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.34264994,0.6852999,1.0279498,1.3705997,1.7132497,1.9906329,2.268016,2.5453994,2.8227828,3.100166,3.2107568,3.3195345,3.4301252,3.540716,3.6494937,3.727451,3.8054085,3.8833659,3.9595103,4.0374675,4.122677,4.207886,4.2930956,4.3783045,4.461701,4.313038,4.162562,4.0120864,3.8616104,3.7129474,4.3982472,5.081734,5.767034,6.452334,7.137634,6.6717024,6.207584,5.7416525,5.277534,4.8116026,6.628191,8.442966,10.257742,12.072517,13.887294,12.4242325,10.962985,9.499924,8.036863,6.5756154,7.3896356,8.205468,9.019489,9.835322,10.649343,10.480737,10.310318,10.139899,9.969481,9.800876,8.120259,6.439643,4.76084,3.0802233,1.3996071,2.7756457,4.1498713,5.52591,6.9001355,8.274362,8.471974,8.669587,8.8672,9.064813,9.262425,7.4929743,5.7217097,3.9522583,2.182807,0.41335547,0.3444629,0.27738327,0.21030366,0.14322405,0.07433146,0.5855869,1.0950294,1.6044719,2.1157274,2.6251698,2.1954978,1.7658255,1.3343405,0.90466833,0.4749962,0.89922947,1.3252757,1.7495089,2.175555,2.5997884,2.4456866,2.2897718,2.13567,1.9797552,1.8256533,1.7875811,1.7495089,1.7132497,1.6751775,1.6371052,1.7730774,1.9072367,2.0432088,2.1773682,2.3133402,2.5925364,2.8717327,3.152742,3.4319382,3.7129474,4.2894692,4.8678045,5.4443264,6.0226617,6.599184,6.240217,5.8794374,5.520471,5.1596913,4.800725,7.132195,9.465478,11.7969475,14.13023,16.4617,15.107417,13.753134,12.397038,11.042755,9.686659,7.817495,5.9483304,4.077353,2.2081885,0.33721104,0.581961,0.82671094,1.0732739,1.3180238,1.5627737,4.077353,6.591932,9.108324,11.622903,14.137483,13.885481,13.631665,13.379663,13.127662,12.87566,13.544643,14.21544,14.884423,15.555219,16.224201,17.243088,18.260159,19.277231,20.294304,21.313189,19.66158,18.011784,16.361988,14.712192,13.062395,14.2516985,15.442815,16.632118,17.823235,19.012539,17.239462,15.468197,13.695119,11.922042,10.150778,12.166792,14.184619,16.202446,18.220274,20.238102,19.882761,19.52742,19.17208,18.816738,18.463211,17.025532,15.5878525,14.150173,12.712494,11.274815,12.195799,13.114971,14.034143,14.955129,15.8743,15.734702,15.595104,15.455506,15.314095,15.174497,13.24913,11.325577,9.400211,7.474845,5.5494785,8.02236,10.49524,12.968122,15.439189,17.912071,16.57773,15.243389,13.907236,12.572895,11.236742,10.504305,9.771869,9.039432,8.306994,7.574558,6.9400206,6.305484,5.669134,5.034597,4.40006,4.137181,3.874301,3.6132345,3.350355,3.0874753,4.501586,5.91751,7.3334336,8.747544,10.161655,9.162713,8.161958,7.1630154,6.16226,5.163317,6.249282,7.3370595,8.424837,9.512614,10.600392,13.486629,16.374678,19.262728,22.150776,25.037014,25.794832,26.55265,27.310469,28.068287,28.824291,27.517145,26.210001,24.902855,23.595709,22.286749,23.062696,23.836832,24.61278,25.386915,26.162863,25.994257,25.827465,25.660673,25.492067,25.325274,23.075388,20.8255,18.575615,16.325727,14.075842,12.75963,11.445232,10.130835,8.814624,7.500226,6.189454,4.880495,3.5697234,2.2607644,0.9499924,1.5301404,2.1102884,2.6904364,3.2705846,3.8507326,4.974769,6.1006193,7.224656,8.350506,9.474543,9.820818,10.165281,10.509744,10.854207,11.200482,12.11059,13.020698,13.930804,14.839099,15.749206,17.68545,19.61988,21.554312,23.490557,25.424988,22.89953,20.375887,17.85043,15.324973,12.799516,11.929294,11.060884,10.190662,9.32044,8.450218,7.059676,5.669134,4.2804046,2.8898623,1.49932,1.3017071,1.1059072,0.90829426,0.7106813,0.51306844,2.03777,3.5624714,5.087173,6.6118746,8.136576,7.1430726,6.147756,5.1524396,4.157123,3.1618068,3.4156215,3.6676233,3.919625,4.171627,4.4254417,4.764466,5.105303,5.4443264,5.7851634,6.1241875,6.506723,6.889258,7.271793,7.654328,8.036863,6.542982,5.047288,3.5515938,2.0577126,0.5620184,0.44961473,0.33721104,0.22480737,0.11240368,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,3.247016,6.3816285,9.518054,12.652666,15.787278,15.431937,15.07841,14.723069,14.367728,14.012388,12.295512,10.576823,8.859948,7.1430726,5.424384,4.949388,4.4743915,3.9993954,3.5243993,3.049403,2.9152439,2.7792716,2.6451125,2.5091403,2.374981,1.9108626,1.4449311,0.9808127,0.5148814,0.05076295,0.31182957,0.5747091,0.8375887,1.1004683,1.3633479,2.373168,3.3829882,4.3928084,5.4026284,6.412449,7.3950744,8.3777,9.360326,10.342952,11.325577,12.032633,12.739688,13.446743,14.155612,14.862667,14.7683935,14.672306,14.5780325,14.481945,14.387671,15.297778,16.207886,17.117992,18.0281,18.938208,18.142317,17.34824,16.55235,15.758271,14.96238,16.420002,17.877625,19.335245,20.792868,22.25049,23.249432,24.250187,25.250942,26.249886,27.25064,29.130682,31.010725,32.890766,34.77081,36.650852,34.6294,32.609756,30.590118,28.570477,26.550837,29.47696,32.404892,35.33283,38.26076,41.186886,35.178726,29.17238,23.164223,17.157877,11.14972,13.448557,15.74558,18.042604,20.339626,22.63665,24.750565,26.862667,28.974768,31.08687,33.200783,32.97235,32.74573,32.517296,32.290676,32.062244,32.009666,31.957092,31.904516,31.85194,31.799364,33.208035,34.614895,36.021755,37.430424,38.837284,34.230545,29.621996,25.015257,20.406708,15.799969,15.74558,15.689378,15.63499,15.580601,15.524399,17.103489,18.680767,20.258043,21.835321,23.4126,21.267864,19.123129,16.976582,14.831847,12.687112,11.227677,9.768243,8.306994,6.8475595,5.388125,5.7344007,6.0824895,6.430578,6.776854,7.124943,6.599184,6.0752378,5.5494785,5.0255322,4.499773,3.7455807,2.9895754,2.2353828,1.4793775,0.72518504,0.6726091,0.6200332,0.56745726,0.5148814,0.46230546,0.5529536,0.6417888,0.7324369,0.823085,0.9119202,0.83033687,0.7469406,0.6653573,0.581961,0.50037766,0.7124943,0.9246109,1.1367276,1.3506571,1.5627737,1.4068589,1.2527572,1.0968424,0.94274056,0.7868258,0.7850128,0.78319985,0.7795739,0.7777609,0.774135,1.4122978,2.0504606,2.6868105,3.3249733,3.9631362,4.0429068,4.122677,4.2024474,4.2822175,4.361988,4.6303062,4.896812,5.1651306,5.431636,5.6999545,5.092612,4.4852695,3.877927,3.2705846,2.663242,2.1719291,1.6824293,1.1929294,0.70342946,0.21211663,0.291887,0.37165734,0.45324063,0.533011,0.61278135,0.50037766,0.387974,0.2755703,0.16316663,0.05076295,0.047137026,0.045324065,0.04169814,0.03988518,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.034446288,0.032633327,0.030820364,0.027194439,0.025381476,0.030820364,0.034446288,0.03988518,0.045324065,0.05076295,0.07977036,0.11059072,0.13959812,0.17041849,0.19942589,0.2520018,0.3045777,0.35715362,0.40972954,0.46230546,0.47680917,0.49312583,0.5076295,0.52213323,0.53663695,0.4604925,0.3825351,0.3045777,0.22662032,0.15047589,0.13778515,0.12509441,0.11240368,0.099712946,0.0870222,0.07070554,0.052575916,0.034446288,0.018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.40791658,0.81583315,1.2219368,1.6298534,2.03777,2.0975976,2.1574254,2.2172532,2.277081,2.3369088,2.5018883,2.666868,2.8318477,2.9968271,3.1618068,3.247016,3.3322253,3.4174345,3.5026438,3.587853,3.6766882,3.7673361,3.8579843,3.9468195,4.0374675,4.062849,4.0882306,4.1117992,4.137181,4.162562,5.290225,6.4178877,7.5455503,8.673213,9.800876,8.765674,7.7304726,6.695271,5.660069,4.6248674,7.473032,10.319383,13.167547,16.01571,18.862062,17.038223,15.212569,13.386916,11.563075,9.737422,9.20985,8.682278,8.154706,7.6271334,7.0995617,7.6325727,8.165584,8.696781,9.229793,9.762803,8.23085,6.697084,5.1651306,3.633177,2.0994108,4.137181,6.1749506,8.212721,10.25049,12.28826,11.115273,9.9422865,8.7693,7.5981264,6.4251394,5.1941376,3.9649491,2.7357605,1.504759,0.2755703,0.23024625,0.18492219,0.13959812,0.09427405,0.05076295,0.40247768,0.7541924,1.1077201,1.4594349,1.8129625,1.5174497,1.2219368,0.92823684,0.6327239,0.33721104,1.0497054,1.7621996,2.474694,3.1871881,3.8996825,3.491766,3.0856624,2.6777458,2.269829,1.8619126,1.938057,2.0123885,2.08672,2.1628644,2.2371957,2.128418,2.0178273,1.9072367,1.7966459,1.6878681,1.8818551,2.077655,2.2716422,2.467442,2.663242,3.0983531,3.531651,3.966762,4.401873,4.836984,4.8841214,4.933071,4.9802084,5.027345,5.0744824,7.654328,10.234174,12.815832,15.3956785,17.975525,15.867048,13.760386,11.651911,9.545248,7.4367723,6.008158,4.5777307,3.147303,1.7168756,0.28826106,0.49312583,0.6979906,0.90285534,1.1077201,1.3125849,3.7600844,6.207584,8.655084,11.102583,13.550082,12.790451,12.03082,11.269376,10.509744,9.750113,10.429974,11.109835,11.789696,12.469557,13.149418,13.519262,13.889107,14.260764,14.630608,15.000452,14.237195,13.475751,12.712494,11.949236,11.187792,11.985496,12.783199,13.57909,14.376793,15.174497,13.822026,12.469557,11.117086,9.764616,8.412147,10.919474,13.426801,15.935941,18.443268,20.950596,20.529987,20.10938,19.690586,19.26998,18.849373,17.661882,16.474392,15.2869005,14.09941,12.91192,13.430427,13.947122,14.465629,14.982323,15.50083,15.152741,14.804652,14.456564,14.110288,13.762199,12.549327,11.338268,10.125396,8.912524,7.699652,9.6141405,11.530442,13.44493,15.359419,17.27572,15.785465,14.29521,12.804955,11.314699,9.824444,9.244296,8.664148,8.0858135,7.5056653,6.925517,6.4595857,5.995467,5.529536,5.0654173,4.599486,4.599486,4.599486,4.599486,4.599486,4.599486,5.422571,6.245656,7.066928,7.890013,8.713099,8.149267,7.5872483,7.02523,6.4632115,5.89938,7.413204,8.925215,10.437225,11.949236,13.46306,15.950445,18.43783,20.925215,23.4126,25.899984,27.442814,28.985645,30.528477,32.069496,33.612328,31.61988,29.627434,27.634989,25.642542,23.650097,24.33721,25.024323,25.71325,26.400362,27.087475,27.480886,27.872486,28.2659,28.6575,29.050913,26.462002,23.874905,21.287807,18.700708,16.1118,14.677745,13.2418785,11.807825,10.371959,8.937905,7.422269,5.908445,4.3928084,2.8771715,1.3633479,1.6080978,1.8528478,2.0975976,2.3423476,2.5870976,4.024777,5.462456,6.9001355,8.337815,9.775495,9.441909,9.110137,8.776552,8.444779,8.113008,8.765674,9.416528,10.069194,10.721861,11.374527,15.326786,19.279043,23.233116,27.185373,31.137632,26.6995,22.26318,17.825048,13.386916,8.950596,8.457471,7.9643445,7.473032,6.979906,6.48678,5.565795,4.6429973,3.720199,2.7974012,1.8746033,1.6352923,1.3941683,1.1548572,0.9155461,0.6744221,1.6371052,2.5997884,3.5624714,4.5251546,5.487838,4.933071,4.3783045,3.8217251,3.2669585,2.712192,3.4972048,4.2822175,5.06723,5.8522434,6.637256,6.947273,7.2572894,7.567306,7.877322,8.187339,7.7794223,7.3733187,6.965402,6.5574856,6.149569,4.994712,3.8398547,2.6849976,1.5301404,0.37528324,0.2991388,0.22480737,0.15047589,0.07433146,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,3.5280252,6.979906,10.431787,13.885481,17.33736,17.417131,17.496902,17.578485,17.658255,17.738026,15.31772,12.897416,10.477111,8.056806,5.638314,5.275721,4.9131284,4.550536,4.1879435,3.825351,3.6476808,3.4700103,3.29234,3.1146698,2.9369993,2.3641033,1.79302,1.2201238,0.64722764,0.07433146,0.2991388,0.52575916,0.7505665,0.97537386,1.2001812,2.715818,4.229642,5.7452784,7.2609153,8.774739,10.391902,12.010877,13.628039,15.245202,16.862366,17.680012,18.497658,19.315304,20.13295,20.950596,20.283426,19.614443,18.947271,18.280102,17.612932,19.177519,20.742105,22.308504,23.87309,25.437677,22.982927,20.528175,18.071611,15.616859,13.162108,15.792717,18.423326,21.052122,23.68273,26.31334,26.574406,26.837286,27.100164,27.363045,27.624111,29.995466,32.36501,34.73455,37.105904,39.47545,38.520016,37.564583,36.610966,35.655537,34.700104,35.722614,36.745125,37.767635,38.790146,39.812656,34.73274,29.652817,24.572895,19.492973,14.413053,16.789846,19.166641,21.545248,23.92204,26.300648,28.062847,29.825047,31.587248,33.349445,35.11346,35.06451,35.017372,34.970234,34.9231,34.87596,35.08989,35.305634,35.51956,35.735306,35.949234,36.95543,37.959812,38.966003,39.970387,40.974766,36.658104,32.339626,28.022963,23.704485,19.387821,19.70509,20.022358,20.339626,20.656897,20.975977,22.647528,24.320892,25.992445,27.66581,29.33736,26.607038,23.87853,21.148209,18.417887,15.687565,14.110288,12.5330105,10.955733,9.378455,7.799365,8.252605,8.705847,9.157274,9.610515,10.061942,9.325879,8.588004,7.850128,7.112252,6.3743763,5.317419,4.2604623,3.2016919,2.1447346,1.0877775,0.93911463,0.79226464,0.64541465,0.49675176,0.34990177,0.44780177,0.54570174,0.6417888,0.73968875,0.8375887,0.79589057,0.7523795,0.7106813,0.6671702,0.62547207,0.9499924,1.2745126,1.6008459,1.9253663,2.2498865,1.9416829,1.6352923,1.3270886,1.020698,0.7124943,0.7016165,0.69255173,0.68167394,0.6726091,0.66173136,1.3506571,2.03777,2.7248828,3.4119956,4.099108,4.519716,4.940323,5.3609304,5.7797246,6.200332,6.6318173,7.065115,7.498413,7.9298983,8.363196,7.420456,6.4777155,5.5349746,4.592234,3.6494937,2.9641938,2.280707,1.5954071,0.9101072,0.22480737,0.35715362,0.4894999,0.62184614,0.7541924,0.8883517,0.72518504,0.5620184,0.40066472,0.2374981,0.07433146,0.065266654,0.054388877,0.045324065,0.034446288,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.027194439,0.030820364,0.032633327,0.034446288,0.038072214,0.045324065,0.052575916,0.059827764,0.06707962,0.07433146,0.09427405,0.11421664,0.13415924,0.15410182,0.17585737,0.25925365,0.3444629,0.42967212,0.5148814,0.6000906,0.6345369,0.67079616,0.70524246,0.73968875,0.774135,0.6526665,0.5293851,0.40791658,0.28463513,0.16316663,0.15047589,0.13778515,0.12509441,0.11240368,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.47318324,0.9445535,1.4177368,1.889107,2.3622901,2.2045624,2.0468347,1.889107,1.7331922,1.5754645,1.794833,2.0142014,2.2353828,2.4547513,2.6741197,2.7683938,2.8608549,2.953316,3.045777,3.1382382,3.2325122,3.3267863,3.4228733,3.5171473,3.6132345,3.8126602,4.0120864,4.213325,4.4127507,4.612177,6.1822023,7.752228,9.322253,10.89228,12.462305,10.857833,9.253361,7.647076,6.0426044,4.4381323,8.317872,12.197612,16.077353,19.957092,23.836832,21.650398,19.462152,17.27572,15.087475,12.899229,11.030065,9.1609,7.2899227,5.4207582,3.5497808,4.784408,6.019036,7.2554765,8.490104,9.724731,8.339628,6.9545245,5.569421,4.1843176,2.7992141,5.5005283,8.200029,10.899531,13.600845,16.300346,13.75676,11.214987,8.673213,6.1296263,3.587853,2.8971143,2.2081885,1.5174497,0.82671094,0.13778515,0.11421664,0.092461094,0.07070554,0.047137026,0.025381476,0.21936847,0.41516843,0.6091554,0.80495536,1.0007553,0.83940166,0.67986095,0.52032024,0.36077955,0.19942589,1.2001812,2.1991236,3.199879,4.2006345,5.199577,4.539658,3.87974,3.2198215,2.5599031,1.8999848,2.08672,2.275268,2.4620032,2.6505513,2.8372865,2.4819458,2.128418,1.7730774,1.4177368,1.062396,1.1729867,1.2817645,1.3923552,1.502946,1.6117238,1.9054236,2.1973107,2.4891977,2.7828975,3.0747845,3.529838,3.9848917,4.439945,4.894999,5.3500524,8.178274,11.004683,13.832905,16.659313,19.487535,16.62668,13.767638,10.906783,8.047741,5.186886,4.1970086,3.207131,2.2172532,1.2273756,0.2374981,0.40247768,0.56745726,0.7324369,0.8974165,1.062396,3.442816,5.823236,8.201842,10.582263,12.962683,11.695421,10.428161,9.159087,7.891826,6.624565,7.315304,8.00423,8.694968,9.385707,10.074633,9.79725,9.519867,9.242483,8.9651,8.6877165,8.812811,8.937905,9.063,9.188094,9.313189,9.71748,10.12177,10.527874,10.932164,11.338268,10.4045925,9.47273,8.539054,7.607191,6.6753283,9.672155,12.670795,15.667623,18.66445,21.66309,21.177216,20.693155,20.207281,19.72322,19.237347,18.300045,17.362743,16.425442,15.488139,14.5508375,14.665054,14.779271,14.895301,15.009518,15.125546,14.57078,14.014201,13.4594345,12.904668,12.349901,11.849524,11.349146,10.850581,10.3502035,9.849826,11.207735,12.565643,13.92174,15.279649,16.637558,14.9932,13.347031,11.702674,10.058316,8.412147,7.9842873,7.558241,7.130382,6.7025228,6.2746634,5.979151,5.6854506,5.389938,5.0944247,4.800725,5.0617914,5.3246713,5.5875506,5.8504305,6.11331,6.341743,6.5719895,6.8022356,7.0324817,7.262728,7.137634,7.0125394,6.887445,6.7623506,6.637256,8.575313,10.51337,12.449615,14.387671,16.325727,18.412449,20.499168,22.5877,24.674421,26.762953,29.090797,31.416828,33.74467,36.072517,38.40036,35.722614,33.04487,30.367123,27.689377,25.011631,25.611723,26.211813,26.811903,27.411995,28.012085,28.965704,29.91751,30.869314,31.822931,32.77474,29.85043,26.924307,23.999998,21.07569,18.149569,16.59586,15.040338,13.484816,11.929294,10.375585,8.655084,6.9345818,5.2140803,3.4953918,1.7748904,1.6842422,1.5954071,1.504759,1.4141108,1.3252757,3.0747845,4.8242936,6.5756154,8.325124,10.074633,9.064813,8.054993,7.0451727,6.035352,5.0255322,5.4207582,5.814171,6.209397,6.604623,6.9998484,12.969934,18.94002,24.910107,30.880192,36.850277,30.49947,24.150475,17.799667,11.450671,5.0998635,4.985647,4.8696175,4.7554007,4.6393714,4.5251546,4.070101,3.6150475,3.159994,2.70494,2.2498865,1.9670644,1.6842422,1.403233,1.1204109,0.8375887,1.2382535,1.6371052,2.03777,2.4366217,2.8372865,2.72307,2.6070402,2.4928236,2.3767939,2.2625773,3.5806012,4.896812,6.2148356,7.5328593,8.8508835,9.130079,9.409276,9.690285,9.969481,10.25049,9.052122,7.855567,6.6571984,5.4606433,4.262275,3.4482548,2.6324217,1.8165885,1.0025684,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,3.8072214,7.5781837,11.347333,15.118295,18.887444,19.402325,19.917208,20.432089,20.94697,21.461851,18.33993,15.218008,12.094274,8.972352,5.8504305,5.600241,5.3500524,5.0998635,4.8496747,4.599486,4.3801174,4.160749,3.9395678,3.720199,3.5008307,2.819157,2.1392958,1.4594349,0.7795739,0.099712946,0.28826106,0.4749962,0.66173136,0.85027945,1.0370146,3.0584679,5.0781083,7.0977483,9.117389,11.137029,13.390542,15.6422415,17.895754,20.147453,22.400965,23.327389,24.255627,25.18205,26.110287,27.03671,25.796644,24.558392,23.318325,22.078259,20.838192,23.057259,25.278137,27.497204,29.718082,31.93715,27.821724,23.70811,19.592686,15.477262,11.361836,15.165432,18.967215,22.77081,26.572592,30.374374,29.89938,29.424383,28.949387,28.47439,27.999393,30.860249,33.71929,36.580147,39.43919,42.30004,42.410633,42.519413,42.63,42.740593,42.84937,41.96827,41.085358,40.202446,39.319534,38.43662,34.284935,30.133251,25.979753,21.82807,17.674572,20.13295,22.589514,25.047892,27.504456,29.962833,31.37513,32.78743,34.199726,35.612022,37.024323,37.15667,37.29083,37.423172,37.55552,37.687866,38.170113,38.652363,39.13461,39.61686,40.100918,40.702824,41.304726,41.908443,42.510345,43.11225,39.08566,35.05726,31.030668,27.002264,22.975676,23.6646,24.35534,25.044266,25.735004,26.425743,28.19338,29.959208,31.726845,33.494484,35.262123,31.948027,28.632118,25.318022,22.002113,18.688019,16.992899,15.297778,13.602658,11.907538,10.212419,10.770811,11.327391,11.885782,12.442362,13.000754,12.050762,11.10077,10.150778,9.200785,8.2507925,6.889258,5.529536,4.169814,2.810092,1.4503701,1.2074331,0.9644961,0.72337204,0.48043507,0.2374981,0.34264994,0.44780177,0.5529536,0.65810543,0.76325727,0.75963134,0.75781834,0.7541924,0.7523795,0.7505665,1.1874905,1.6244144,2.0631514,2.5000753,2.9369993,2.47832,2.0178273,1.5573349,1.0968424,0.63816285,0.6200332,0.60190356,0.5855869,0.56745726,0.5493277,1.2872034,2.0250793,2.762955,3.5008307,4.2368937,4.9983377,5.7579694,6.5176005,7.2772317,8.036863,8.63514,9.233418,9.829884,10.428161,11.024626,9.7483,8.470161,7.192023,5.915697,4.6375585,3.7582715,2.8771715,1.9978848,1.1167849,0.2374981,0.4224203,0.6073425,0.79226464,0.97718686,1.162109,0.9499924,0.73787576,0.52575916,0.31182957,0.099712946,0.08339628,0.065266654,0.047137026,0.030820364,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.01994259,0.027194439,0.034446288,0.04169814,0.05076295,0.059827764,0.07070554,0.07977036,0.09064813,0.099712946,0.11059072,0.11965553,0.13053331,0.13959812,0.15047589,0.26831847,0.38434806,0.50219065,0.6200332,0.73787576,0.79226464,0.8466535,0.90285534,0.9572442,1.0116332,0.8448406,0.678048,0.5094425,0.34264994,0.17585737,0.16316663,0.15047589,0.13778515,0.12509441,0.11240368,0.09064813,0.06707962,0.045324065,0.02175555,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.53663695,1.0750868,1.6117238,2.1501737,2.6868105,2.3133402,1.938057,1.5627737,1.1874905,0.8122072,1.0877775,1.3633479,1.6371052,1.9126755,2.1882458,2.2879589,2.3876717,2.4873846,2.5870976,2.6868105,2.7883365,2.8880494,2.9877625,3.0874753,3.1871881,3.5624714,3.9377546,4.313038,4.688321,5.0617914,7.07418,9.086569,11.10077,13.113158,15.125546,12.949992,10.774437,8.600695,6.4251394,4.249584,9.162713,14.074029,18.987158,23.900286,28.811602,26.262575,23.711737,21.162712,18.611874,16.062849,12.850279,9.637709,6.4251394,3.2125697,0.0,1.938057,3.874301,5.812358,7.750415,9.686659,8.450218,7.211965,5.975525,4.7372713,3.5008307,6.8620634,10.225109,13.588155,16.949387,20.312433,16.400059,12.487686,8.575313,4.6629395,0.7505665,0.6000906,0.44961473,0.2991388,0.15047589,0.0,0.0,0.0,0.0,0.0,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.16316663,0.13778515,0.11240368,0.0870222,0.06164073,1.3506571,2.6378605,3.925064,5.2122674,6.4994707,5.5875506,4.6756306,3.7618973,2.8499773,1.938057,2.2371957,2.5381477,2.8372865,3.1382382,3.437377,2.8372865,2.2371957,1.6371052,1.0370146,0.43692398,0.46230546,0.48768693,0.51306844,0.53663695,0.5620184,0.7124943,0.8629702,1.0116332,1.162109,1.3125849,2.175555,3.0367124,3.8996825,4.762653,5.6256227,8.700407,11.775192,14.849977,17.92476,20.999546,17.388124,13.77489,10.161655,6.550234,2.9369993,2.3876717,1.8383441,1.2872034,0.73787576,0.18673515,0.31182957,0.43692398,0.5620184,0.6871128,0.8122072,3.1255474,5.4370747,7.750415,10.061942,12.375282,10.600392,8.825501,7.0506115,5.275721,3.5008307,4.2006345,4.900438,5.600241,6.300045,6.9998484,6.0752378,5.1506267,4.2242026,3.299592,2.374981,3.386614,4.40006,5.411693,6.4251394,7.4367723,7.4494634,7.462154,7.474845,7.4875355,7.500226,6.987158,6.4759026,5.962834,5.4497657,4.936697,8.424837,11.912977,15.399304,18.887444,22.375584,21.824444,21.275116,20.725788,20.174648,19.62532,18.938208,18.24928,17.562168,16.875055,16.187943,15.899682,15.613234,15.324973,15.036712,14.750263,13.987006,13.225562,12.462305,11.700861,10.937603,11.14972,11.361836,11.575767,11.787883,11.999999,12.799516,13.600845,14.400362,15.199879,15.999394,14.199123,12.400664,10.600392,8.80012,6.9998484,6.7242785,6.450521,6.1749506,5.89938,5.6256227,5.5005283,5.375434,5.2503395,5.125245,5.0001507,5.524097,6.049856,6.5756154,7.0995617,7.6253204,7.262728,6.9001355,6.5375433,6.1749506,5.812358,6.1241875,6.43783,6.7496595,7.063302,7.3751316,9.737422,12.099712,14.462003,16.824293,19.188396,20.87445,22.562319,24.250187,25.938055,27.624111,30.736967,33.849823,36.96268,40.07554,43.188396,39.825348,36.462303,33.09926,29.738026,26.374979,26.888048,27.399303,27.912373,28.42544,28.936695,30.45052,31.96253,33.47454,34.988365,36.500374,33.23704,29.975523,26.71219,23.45067,20.187338,18.512161,16.836983,15.161806,13.486629,11.813264,9.8878975,7.9625316,6.037165,4.1117992,2.1882458,1.7621996,1.3379664,0.9119202,0.48768693,0.06164073,2.124792,4.1879435,6.249282,8.312433,10.375585,8.6877165,6.9998484,5.3119802,3.6241121,1.938057,2.0758421,2.2118144,2.3495996,2.4873846,2.6251698,10.613083,18.599184,26.587097,34.57501,42.562923,34.29944,26.03777,17.774284,9.512614,1.2491312,1.5120108,1.7748904,2.03777,2.3006494,2.561716,2.5744069,2.5870976,2.5997884,2.612479,2.6251698,2.3006494,1.9743162,1.649796,1.3252757,1.0007553,0.8375887,0.6744221,0.51306844,0.34990177,0.18673515,0.51306844,0.8375887,1.162109,1.4866294,1.8129625,3.6621845,5.5132194,7.362441,9.211663,11.062697,11.312886,11.563075,11.813264,12.06164,12.311829,10.324821,8.337815,6.350808,4.361988,2.374981,1.8999848,1.4249886,0.9499924,0.4749962,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,4.0882306,8.174648,12.262879,16.349297,20.437527,21.38752,22.337511,23.287504,24.237497,25.187489,21.362139,17.536787,13.713249,9.8878975,6.0625467,5.924762,5.7869763,5.6491914,5.5132194,5.375434,5.1125546,4.8496747,4.5867953,4.325729,4.062849,3.2742105,2.4873846,1.7005589,0.9119202,0.12509441,0.2755703,0.42423326,0.5747091,0.72518504,0.87566096,3.3993049,5.924762,8.450218,10.975676,13.499319,16.38737,19.275417,22.163467,25.049704,27.937754,28.974768,30.011782,31.05061,32.087624,33.124638,31.311676,29.500526,27.687565,25.874601,24.06164,26.936998,29.812357,32.687714,35.563072,38.43662,32.662334,26.888048,21.11195,15.337664,9.563377,14.538147,19.512917,24.487686,29.462456,34.437225,33.224354,32.013294,30.80042,29.58755,28.374678,31.725033,35.075386,38.425743,41.774284,45.124638,46.29944,47.47424,48.650852,49.82565,51.00045,48.212112,45.42559,42.637253,39.85073,37.062393,33.837135,30.611874,27.386612,24.163166,20.937904,23.476053,26.012386,28.550535,31.08687,33.625015,34.687412,35.74981,36.812206,37.8746,38.936996,39.25064,39.56247,39.8743,40.187943,40.49977,41.25034,41.999092,42.749657,43.500225,44.25079,44.45022,44.649643,44.85088,45.05031,45.249733,41.511406,37.774887,34.03656,30.300043,26.561714,27.625923,28.68832,29.750715,30.813112,31.875507,33.73742,35.599335,37.46306,39.32497,41.186886,37.2872,33.38752,29.487837,25.588154,21.686659,19.87551,18.062546,16.249584,14.436621,12.625471,13.287203,13.9507475,14.612478,15.27421,15.937754,14.775645,13.611723,12.449615,11.287505,10.125396,8.46291,6.8004227,5.137936,3.4754493,1.8129625,1.4757515,1.1367276,0.7995165,0.46230546,0.12509441,0.2374981,0.34990177,0.46230546,0.5747091,0.6871128,0.72518504,0.76325727,0.7995165,0.8375887,0.87566096,1.4249886,1.9743162,2.525457,3.0747845,3.6241121,3.0131438,2.4003625,1.7875811,1.1747998,0.5620184,0.53663695,0.51306844,0.48768693,0.46230546,0.43692398,1.2255627,2.0123885,2.7992141,3.587853,4.3746786,5.475147,6.5756154,7.6742706,8.774739,9.875207,10.636651,11.399909,12.163166,12.92461,13.687867,12.07433,10.462607,8.849071,7.2373466,5.6256227,4.550536,3.4754493,2.4003625,1.3252757,0.25018883,0.48768693,0.72518504,0.96268314,1.2001812,1.4376793,1.1747998,0.9119202,0.6508536,0.387974,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.2755703,0.42423326,0.5747091,0.72518504,0.87566096,0.9499924,1.0243238,1.1004683,1.1747998,1.2491312,1.0370146,0.824898,0.61278135,0.40066472,0.18673515,0.17585737,0.16316663,0.15047589,0.13778515,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.42967212,0.85934424,1.2908293,1.7205015,2.1501737,1.8981718,1.6443571,1.3923552,1.1403534,0.8883517,1.1874905,1.4866294,1.7875811,2.08672,2.3876717,2.3641033,2.3423476,2.3205922,2.2970235,2.275268,2.6142921,2.955129,3.294153,3.63499,3.975827,4.4145637,4.855114,5.295664,5.7344007,6.1749506,7.817495,9.460039,11.102583,12.745127,14.387671,12.87566,11.361836,9.849826,8.337815,6.825804,11.300196,15.774588,20.250792,24.725183,29.199575,25.997883,22.794378,19.592686,16.389181,13.1874895,10.573197,7.957093,5.3428006,2.7266958,0.11240368,1.6606737,3.207131,4.7554007,6.301858,7.850128,6.867502,5.8848767,4.902251,3.919625,2.9369993,5.614745,8.292491,10.970237,13.647983,16.325727,13.200181,10.074633,6.9490857,3.825351,0.69980353,0.56020546,0.42060733,0.27919623,0.13959812,0.0,0.0,0.0,0.0,0.0,0.0,0.032633327,0.065266654,0.09789998,0.13053331,0.16316663,0.25018883,0.33721104,0.42423326,0.51306844,0.6000906,1.5772774,2.5544643,3.531651,4.510651,5.487838,4.7699046,4.0519714,3.3358512,2.617918,1.8999848,2.3550384,2.810092,3.2651455,3.720199,4.175253,3.4174345,2.659616,1.9017978,1.1457924,0.387974,0.40429065,0.4224203,0.4405499,0.45686656,0.4749962,0.8194591,1.1657349,1.5101979,1.8546607,2.1991236,2.9877625,3.774588,4.5632267,5.3500524,6.1368785,8.562622,10.986553,13.412297,15.838041,18.261972,15.40293,12.542075,9.683033,6.8221784,3.9631362,3.4301252,2.8971143,2.3641033,1.8329052,1.2998942,1.3452182,1.3905423,1.4358664,1.4793775,1.5247015,3.4645715,5.4044414,7.344311,9.284182,11.225864,9.80994,8.39583,6.979906,5.565795,4.1498713,4.559601,4.9693303,5.3808727,5.7906027,6.200332,5.674573,5.1506267,4.6248674,4.099108,3.5751622,4.195195,4.8152285,5.4352617,6.055295,6.6753283,6.7152133,6.755099,6.794984,6.834869,6.874754,6.5194135,6.165886,5.810545,5.4552045,5.0998635,8.178274,11.254871,14.333282,17.40988,20.48829,20.138388,19.786674,19.436771,19.08687,18.736969,18.002718,17.266655,16.532406,15.798156,15.062093,14.458377,13.852847,13.247317,12.6417885,12.038072,11.845898,11.651911,11.459737,11.267563,11.075388,11.807825,12.540262,13.272699,14.005136,14.737573,15.332225,15.926876,16.52334,17.117992,17.712645,16.104548,14.498261,12.890164,11.282066,9.675781,8.966913,8.259857,7.552802,6.8457465,6.1368785,5.959208,5.7833505,5.6056805,5.42801,5.2503395,5.719897,6.189454,6.6608243,7.130382,7.5999393,7.2971745,6.9944096,6.6916447,6.390693,6.0879283,6.430578,6.773228,7.115878,7.456715,7.799365,9.6504,11.499621,13.3506565,15.199879,17.050913,18.367125,19.685148,21.003172,22.319382,23.637405,26.269827,28.90225,31.534672,34.16709,36.799515,34.45717,32.11482,29.772472,27.430124,25.087776,25.290829,25.492067,25.695118,25.89817,26.09941,27.310469,28.519714,29.730774,30.94002,32.149265,29.84499,27.540714,25.234627,22.930351,20.624262,18.894695,17.16513,15.435563,13.704185,11.974618,9.953164,7.9298983,5.906632,3.8851788,1.8619126,2.08672,2.3133402,2.5381477,2.762955,2.9877625,4.122677,5.2575917,6.392506,7.5274205,8.662335,7.3479376,6.0317264,4.7173285,3.4029307,2.08672,4.855114,7.6216946,10.390089,13.15667,15.925063,19.72322,23.519564,27.31772,31.115877,34.91222,28.467138,22.022057,15.576975,9.131892,2.6868105,2.619731,2.5526514,2.4855716,2.4166791,2.3495996,2.3006494,2.2498865,2.1991236,2.1501737,2.0994108,1.8782293,1.6552348,1.4322405,1.209246,0.9880646,0.8901646,0.79226464,0.69436467,0.5982776,0.50037766,0.88291276,1.2654479,1.647983,2.030518,2.4130533,4.505212,6.5973706,8.689529,10.781689,12.87566,12.757817,12.639976,12.522133,12.40429,12.28826,11.99456,11.702674,11.410787,11.117086,10.825199,9.171778,7.520169,5.866747,4.215138,2.561716,3.870675,5.177821,6.484967,7.7921133,9.099259,10.64753,12.193986,13.742256,15.290526,16.836983,17.922949,19.0071,20.093063,21.177216,22.26318,24.9373,27.613234,30.287354,32.963287,35.637405,30.057106,24.476809,18.89651,13.318023,7.7377243,7.569119,7.402326,7.2355337,7.066928,6.9001355,8.580752,10.259555,11.940171,13.620788,15.299591,12.752378,10.205167,7.6579537,5.1107416,2.561716,2.6795588,2.7974012,2.9152439,3.0330863,3.149116,6.882006,10.614896,14.347786,18.080675,21.811752,26.132042,30.452332,34.77262,39.09291,43.41139,42.222084,41.032784,39.841667,38.652363,37.46306,35.525,33.586945,31.650702,29.712645,27.774588,29.377245,30.979904,32.582565,34.185223,35.78788,31.2029,26.617916,22.032934,17.447952,12.862969,16.873243,20.881702,24.891975,28.90225,32.91252,32.682278,32.45203,32.221783,31.993351,31.763105,35.33464,38.90799,42.479527,46.052876,49.624413,50.329655,51.034897,51.74014,52.44538,53.150623,50.1121,47.075386,44.03686,41.00015,37.961624,36.206676,34.45173,32.69678,30.941832,29.186884,31.291735,33.396584,35.503246,37.608097,39.712944,40.452633,41.19232,41.93201,42.6717,43.4132,43.935337,44.45747,44.979603,45.501736,46.02568,46.464417,46.90497,47.345516,47.784256,48.224804,48.08702,47.949234,47.813263,47.675476,47.537693,44.06043,40.583168,37.10409,33.62683,30.149569,30.856623,31.56549,32.27255,32.979603,33.686657,35.619274,37.551895,39.484512,41.41713,43.349747,40.35292,37.354282,34.357452,31.360626,28.361986,26.63242,24.902855,23.171474,21.441908,19.712341,19.672457,19.632572,19.592686,19.552801,19.512917,18.459585,17.408066,16.354736,15.303217,14.249886,13.258195,12.264692,11.273002,10.279498,9.287807,8.977791,8.667774,8.357758,8.047741,7.7377243,6.8094873,5.883064,4.954827,4.02659,3.100166,2.7176309,2.335096,1.9525607,1.5700256,1.1874905,1.6171626,2.0468347,2.47832,2.907992,3.3376641,2.953316,2.5671551,2.182807,1.7966459,1.4122978,1.2074331,1.0025684,0.79770356,0.59283876,0.387974,1.2056202,2.0232663,2.8409123,3.6567454,4.4743915,5.4044414,6.3344913,7.264541,8.194591,9.12464,9.525306,9.924157,10.324821,10.725487,11.124338,9.989424,8.854509,7.7195945,6.58468,5.4497657,4.64481,3.8398547,3.0348995,2.229944,1.4249886,1.4358664,1.4449311,1.455809,1.4648738,1.4757515,1.2056202,0.9354887,0.6653573,0.39522585,0.12509441,0.10333887,0.07977036,0.058014803,0.034446288,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.018129626,0.034446288,0.052575916,0.07070554,0.0870222,0.15954071,0.23205921,0.3045777,0.3770962,0.44961473,0.38434806,0.3208944,0.25562772,0.19036107,0.12509441,0.24837588,0.36984438,0.49312583,0.61459434,0.73787576,0.8194591,0.90285534,0.98443866,1.067835,1.1494182,1.0025684,0.8557183,0.7070554,0.56020546,0.41335547,0.41516843,0.4169814,0.42060733,0.4224203,0.42423326,0.35534066,0.28463513,0.21574254,0.14503701,0.07433146,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.32270733,0.64541465,0.968122,1.2908293,1.6117238,1.4830034,1.35247,1.2219368,1.0932164,0.96268314,1.2872034,1.6117238,1.938057,2.2625773,2.5870976,2.4420607,2.2970235,2.1519866,2.0069497,1.8619126,2.4420607,3.0222087,3.6023567,4.1825047,4.762653,5.2666564,5.772473,6.2782893,6.782293,7.28811,8.560809,9.8316965,11.104396,12.377095,13.649796,12.799516,11.949236,11.10077,10.25049,9.400211,13.437678,17.475147,21.512613,25.550081,29.58755,25.73319,21.87702,18.022661,14.168303,10.312131,8.294304,6.2782893,4.2604623,2.2426348,0.22480737,1.3832904,2.5399606,3.6966307,4.855114,6.011784,5.2847857,4.557788,3.83079,3.101979,2.374981,4.367427,6.359873,8.352319,10.344765,12.337211,10.000301,7.663393,5.3246713,2.9877625,0.6508536,0.52032024,0.38978696,0.25925365,0.13053331,0.0,0.0,0.0,0.0,0.0,0.0,0.027194439,0.054388877,0.08339628,0.11059072,0.13778515,0.33721104,0.53663695,0.73787576,0.93730164,1.1367276,1.8057107,2.472881,3.1400511,3.8072214,4.4743915,3.9522583,3.4301252,2.907992,2.3858588,1.8619126,2.472881,3.0820365,3.6930048,4.3021603,4.9131284,3.9975824,3.0820365,2.1683033,1.2527572,0.33721104,0.3480888,0.35715362,0.3680314,0.3770962,0.387974,0.92823684,1.4666867,2.0069497,2.5472124,3.0874753,3.7999697,4.512464,5.224958,5.9374523,6.6499467,8.424837,10.199727,11.974618,13.749508,15.524399,13.417736,11.30926,9.202598,7.0941224,4.98746,4.4725785,3.9576974,3.442816,2.9279346,2.4130533,2.3767939,2.3423476,2.3079014,2.2716422,2.2371957,3.8054085,5.371808,6.9400206,8.508233,10.074633,9.019489,7.9643445,6.9092,5.8558693,4.800725,4.9203806,5.040036,5.1596913,5.279347,5.4008155,5.275721,5.1506267,5.0255322,4.900438,4.7753434,5.0019636,5.230397,5.4570174,5.6854506,5.9120708,5.979151,6.0480433,6.115123,6.1822023,6.249282,6.051669,5.8558693,5.658256,5.4606433,5.2630305,7.9298983,10.596766,13.265448,15.932315,18.599184,18.45052,18.300045,18.149569,17.999092,17.85043,17.06723,16.285843,15.502643,14.719443,13.938056,13.015259,12.092461,11.169662,10.246864,9.325879,9.702975,10.080072,10.457169,10.834265,11.213174,12.464118,13.716875,14.969632,16.22239,17.475147,17.864933,18.25472,18.644506,19.034294,19.425894,18.00997,16.59586,15.179935,13.765825,12.349901,11.209548,10.069194,8.930654,7.7903004,6.6499467,6.4197006,6.189454,5.959208,5.730775,5.5005283,5.915697,6.3308654,6.7442207,7.159389,7.574558,7.3316207,7.0904965,6.8475595,6.604623,6.3616858,6.735156,7.1068134,7.4802837,7.851941,8.225411,9.563377,10.899531,12.237497,13.575464,14.911617,15.859797,16.807976,17.754343,18.702522,19.650702,21.802689,23.954674,26.10666,28.26046,30.412447,29.090797,27.767334,26.445684,25.122223,23.800573,23.691795,23.58483,23.477865,23.369087,23.262123,24.170418,25.076899,25.985193,26.891674,27.799969,26.452936,25.105906,23.757061,22.41003,21.063,19.277231,17.493277,15.707508,13.92174,12.137785,10.018432,7.897265,5.7779117,3.6567454,1.5373923,2.4130533,3.2869012,4.162562,5.038223,5.9120708,6.1205616,6.3272395,6.53573,6.742408,6.9490857,6.008158,5.0654173,4.122677,3.1799364,2.2371957,7.6361985,13.031575,18.430578,23.827766,29.224957,28.833357,28.439943,28.048344,27.654932,27.26333,22.634838,18.008158,13.379663,8.752983,4.12449,3.727451,3.3304121,2.9333735,2.5345216,2.137483,2.0250793,1.9126755,1.8002719,1.6878681,1.5754645,1.455809,1.3343405,1.214685,1.0950294,0.97537386,0.94274056,0.9101072,0.8774739,0.8448406,0.8122072,1.2527572,1.693307,2.132044,2.572594,3.0131438,5.3482394,7.6833353,10.018432,12.351714,14.68681,14.202749,13.716875,13.232814,12.74694,12.262879,13.664299,15.067532,16.470764,17.872185,19.275417,16.445383,13.615349,10.785315,7.95528,5.125245,7.7395372,10.355642,12.969934,15.584227,18.20033,21.29506,24.389786,27.484512,30.581053,33.67578,31.757666,29.839552,27.92325,26.005135,24.08702,28.487082,32.887142,37.2872,41.687263,46.087322,38.752075,31.418642,24.081581,16.748148,9.412902,9.215289,9.017676,8.820063,8.62245,8.424837,12.047136,15.6694355,19.293549,22.915848,26.538147,22.230547,17.922949,13.615349,9.30775,5.0001507,5.08536,5.1705694,5.2557783,5.3391747,5.424384,10.364707,15.30503,20.245354,25.185677,30.124186,35.87853,41.629246,47.38359,53.134308,58.886837,55.469402,52.051968,48.634533,45.2171,41.799664,39.736515,37.675175,35.612022,33.550686,31.487534,31.817493,32.147453,32.477413,32.80737,33.13733,29.741652,26.347786,22.952106,19.55824,16.162561,19.208338,22.252302,25.29808,28.342045,31.387821,32.1402,32.892582,33.64496,34.39734,35.14972,38.946064,42.740593,46.535122,50.329655,54.124184,54.35987,54.595554,54.829426,55.065113,55.300797,52.012085,48.72518,45.438282,42.149567,38.862667,38.57803,38.293396,38.006947,37.722313,37.437675,39.111042,40.782593,42.45596,44.12751,45.800873,46.217854,46.63484,47.05182,47.47061,47.887592,48.62003,49.352467,50.084904,50.81734,51.549778,51.680313,51.810844,51.939564,52.0701,52.20063,51.725636,51.25064,50.775642,50.300648,49.82565,46.607643,43.389633,40.171623,36.95543,33.73742,34.09095,34.44266,34.794376,35.147907,35.49962,37.502945,39.504456,41.50778,43.50929,45.51261,43.41683,41.322857,39.22707,37.1331,35.037315,33.38933,31.743162,30.095179,28.447195,26.799213,26.05771,25.314396,24.572895,23.82958,23.088078,22.145338,21.202597,20.259857,19.317116,18.374376,18.051668,17.730774,17.408066,17.08536,16.762651,16.47983,16.197008,15.914186,15.633177,15.350354,13.383289,11.4144125,9.447348,7.4802837,5.5132194,4.710077,3.9069343,3.105605,2.3024626,1.49932,1.8093367,2.1193533,2.42937,2.7393866,3.049403,2.8916752,2.7357605,2.5780327,2.420305,2.2625773,1.8782293,1.4920682,1.1077201,0.72337204,0.33721104,1.1856775,2.032331,2.8807976,3.727451,4.574105,5.335549,6.09518,6.8548117,7.614443,8.375887,8.412147,8.450218,8.488291,8.52455,8.562622,7.9045167,7.2482243,6.590119,5.9320135,5.275721,4.7390842,4.2042603,3.6694362,3.1346123,2.5997884,2.382233,2.1646774,1.9471219,1.7295663,1.5120108,1.2346275,0.9572442,0.67986095,0.40247768,0.12509441,0.10515183,0.08520924,0.065266654,0.045324065,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.24474995,0.3770962,0.5094425,0.6417888,0.774135,0.64541465,0.5148814,0.38434806,0.25562772,0.12509441,0.21936847,0.3154555,0.40972954,0.5058166,0.6000906,0.69073874,0.7795739,0.87022203,0.96087015,1.0497054,0.968122,0.88472575,0.8031424,0.7197462,0.63816285,0.6544795,0.6726091,0.69073874,0.7070554,0.72518504,0.6091554,0.4949388,0.38072214,0.26469254,0.15047589,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.21574254,0.42967212,0.64541465,0.85934424,1.0750868,1.067835,1.0605831,1.0533313,1.0442665,1.0370146,1.3869164,1.7368182,2.08672,2.4366217,2.7883365,2.520018,2.2516994,1.9851941,1.7168756,1.4503701,2.269829,3.0892882,3.9105604,4.7300196,5.5494785,6.1205616,6.6898317,7.2609153,7.8301854,8.399456,9.302311,10.205167,11.108022,12.010877,12.91192,12.725184,12.536636,12.349901,12.163166,11.974618,15.575162,19.175705,22.774435,26.374979,29.975523,25.466686,20.95966,16.452635,11.94561,7.4367723,6.017223,4.597673,3.1781235,1.7567607,0.33721104,1.1040943,1.8727903,2.6396735,3.4083695,4.175253,3.7020695,3.2306993,2.7575161,2.2843328,1.8129625,3.1201086,4.4272547,5.7344007,7.041547,8.350506,6.8004227,5.2503395,3.7002566,2.1501737,0.6000906,0.48043507,0.36077955,0.23931105,0.11965553,0.0,0.0,0.0,0.0,0.0,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.42423326,0.73787576,1.0497054,1.3633479,1.6751775,2.032331,2.3894846,2.7466383,3.105605,3.4627585,3.1346123,2.808279,2.4801328,2.1519866,1.8256533,2.5907235,3.3557937,4.120864,4.8859344,5.6491914,4.5777307,3.5044568,2.4329958,1.3597219,0.28826106,0.29007402,0.291887,0.2955129,0.29732585,0.2991388,1.0352017,1.7694515,2.5055144,3.2397642,3.975827,4.612177,5.2503395,5.8866897,6.5248523,7.1630154,8.287052,9.412902,10.536939,11.662788,12.786825,11.432542,10.078259,8.722163,7.36788,6.011784,5.5150323,5.0182805,4.519716,4.022964,3.5243993,3.4101827,3.294153,3.1799364,3.0657198,2.94969,4.1444325,5.3391747,6.53573,7.7304726,8.925215,8.23085,7.5346723,6.8403077,6.14413,5.4497657,5.279347,5.1107416,4.940323,4.7699046,4.599486,4.8750563,5.1506267,5.424384,5.6999545,5.975525,5.810545,5.6455655,5.480586,5.315606,5.1506267,5.2449007,5.3391747,5.4352617,5.529536,5.6256227,5.5857377,5.5458527,5.504154,5.464269,5.424384,7.6833353,9.940474,12.197612,14.454751,16.71189,16.762651,16.811602,16.862366,16.913128,16.962078,16.13174,15.303217,14.47288,13.642544,12.812206,11.57214,10.332074,9.092008,7.851941,6.6118746,7.560054,8.508233,9.4546,10.40278,11.349146,13.122223,14.895301,16.668379,18.439642,20.212719,20.397642,20.582563,20.767487,20.952408,21.137331,19.915394,18.693457,17.469707,16.24777,15.025834,13.452183,11.880343,10.306692,8.734854,7.1630154,6.880193,6.5973706,6.3145485,6.0317264,5.750717,6.109684,6.4704633,6.82943,7.1902094,7.549176,7.36788,7.1847706,7.0016613,6.8203654,6.637256,7.039734,7.4422116,7.844689,8.247167,8.649645,9.474543,10.29944,11.124338,11.949236,12.774135,13.352469,13.928991,14.507326,15.085662,15.662184,17.335548,19.0071,20.680464,22.352016,24.025381,23.722616,23.419851,23.117086,22.814322,22.511557,22.094576,21.677593,21.260612,20.841818,20.424837,21.030367,21.634083,22.239613,22.845142,23.45067,23.05907,22.669285,22.279497,21.88971,21.499924,19.659767,17.819609,15.979452,14.139296,12.299138,10.081885,7.8646317,5.6473784,3.4301252,1.2128719,2.7375734,4.262275,5.7869763,7.313491,8.838193,8.116633,7.3968873,6.677141,5.957395,5.237649,4.666566,4.0972953,3.5280252,2.956942,2.3876717,10.41547,18.443268,26.471067,34.49705,42.52485,37.94168,33.360325,28.777155,24.193985,19.612629,16.802538,13.992445,11.182353,8.372261,5.562169,4.835171,4.1081734,3.3793623,2.6523643,1.9253663,1.7495089,1.5754645,1.3996071,1.2255627,1.0497054,1.0333886,1.015259,0.99712944,0.9808127,0.96268314,0.99531645,1.0279498,1.0605831,1.0932164,1.1258497,1.6226015,2.1193533,2.617918,3.1146698,3.6132345,6.189454,8.767487,11.34552,13.92174,16.499773,15.64768,14.795588,13.941682,13.08959,12.237497,15.335851,18.43239,21.530745,24.627283,27.725637,23.717176,19.71053,15.702069,11.695421,7.686961,11.610212,15.531651,19.4549,23.378153,27.299591,31.942587,36.585587,41.22858,45.869766,50.512764,45.592384,40.673817,35.753433,30.833055,25.912674,32.038673,38.16286,44.28705,50.41305,56.53724,47.447044,38.35866,29.266655,20.178274,11.088079,10.859646,10.633025,10.4045925,10.177972,9.949538,15.515334,21.079315,26.645111,32.210907,37.774887,31.706903,25.64073,19.572744,13.504758,7.4367723,7.4893484,7.5419245,7.5945,7.647076,7.699652,13.847408,19.995165,26.14292,32.290676,38.43843,45.623203,52.807976,59.992744,67.17751,74.36229,68.71672,63.072968,57.427402,51.781837,46.138084,43.94984,41.763405,39.57516,37.386913,35.20048,34.25774,33.315,32.37226,31.42952,30.486778,28.282217,26.077654,23.87309,21.666716,19.462152,21.543434,23.622902,25.70237,27.78184,29.86312,31.598125,33.33313,35.068134,36.80314,38.538147,42.55567,46.573196,50.59072,54.608246,58.62577,58.390087,58.1544,57.92053,57.684845,57.45097,53.912067,50.374977,46.837887,43.300797,39.761894,40.947575,42.13325,43.317116,44.502792,45.68847,46.928535,48.16679,49.406857,50.646923,51.88699,51.983078,52.07735,52.17344,52.26771,52.361984,53.304726,54.247467,55.19021,56.132946,57.075687,56.89439,56.71491,56.535423,56.35594,56.174644,55.36244,54.550232,53.738026,52.925816,52.111797,49.154854,46.197914,43.23916,40.282215,37.325275,37.32346,37.319836,37.318024,37.314396,37.312584,39.3848,41.457016,43.529232,45.60326,47.675476,46.482548,45.28962,44.098503,42.90557,41.712643,40.148056,38.58347,37.01707,35.452484,33.887897,32.442966,30.998034,29.553102,28.108171,26.66324,25.829277,24.997128,24.164978,23.332829,22.500679,22.846954,23.195044,23.543133,23.889408,24.237497,23.981869,23.728054,23.472427,23.218613,22.962984,19.955278,16.947575,13.939869,10.932164,7.9244595,6.7025228,5.480586,4.256836,3.0348995,1.8129625,2.0033236,2.1918716,2.382233,2.572594,2.762955,2.8318477,2.902553,2.9732587,3.0421512,3.1128569,2.5472124,1.983381,1.4177368,0.8520924,0.28826106,1.1657349,2.0432088,2.9206827,3.7981565,4.6756306,5.2648435,5.8558693,6.445082,7.0342946,7.6253204,7.3008003,6.9744673,6.6499467,6.3254266,5.999093,5.81961,5.6401267,5.4606433,5.279347,5.0998635,4.835171,4.5704784,4.305786,4.0392804,3.774588,3.3304121,2.8844235,2.4402475,1.9942589,1.550083,1.2654479,0.9808127,0.69436467,0.40972954,0.12509441,0.10696479,0.09064813,0.072518505,0.054388877,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.027194439,0.054388877,0.08339628,0.11059072,0.13778515,0.32995918,0.52213323,0.71430725,0.90829426,1.1004683,0.90466833,0.7106813,0.5148814,0.3208944,0.12509441,0.19217403,0.25925365,0.32814622,0.39522585,0.46230546,0.56020546,0.65810543,0.7541924,0.8520924,0.9499924,0.9318628,0.9155461,0.8974165,0.8792868,0.8629702,0.89560354,0.92823684,0.96087015,0.9916905,1.0243238,0.86478317,0.70524246,0.54570174,0.38434806,0.22480737,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.10696479,0.21574254,0.32270733,0.42967212,0.53663695,0.6526665,0.7668832,0.88291276,0.99712944,1.1131591,1.4866294,1.8619126,2.2371957,2.612479,2.9877625,2.5979755,2.2081885,1.8165885,1.4268016,1.0370146,2.0975976,3.1581807,4.216951,5.277534,6.338117,6.972654,7.607191,8.241728,8.8780775,9.512614,10.045626,10.576823,11.109835,11.642846,12.175857,12.650853,13.125849,13.600845,14.075842,14.5508375,17.712645,20.87445,24.03807,27.199877,30.361685,25.201992,20.042301,14.882609,9.7229185,4.5632267,3.7401419,2.9170568,2.0957847,1.2726997,0.44961473,0.82671094,1.2056202,1.5827163,1.9598125,2.3369088,2.1193533,1.9017978,1.6842422,1.4666867,1.2491312,1.8727903,2.4946365,3.1182957,3.7401419,4.361988,3.6005437,2.8372865,2.0758421,1.3125849,0.5493277,0.4405499,0.32995918,0.21936847,0.11059072,0.0,0.0,0.0,0.0,0.0,0.0,0.018129626,0.034446288,0.052575916,0.07070554,0.0870222,0.51306844,0.93730164,1.3633479,1.7875811,2.2118144,2.2607644,2.3079014,2.3550384,2.4021754,2.4493124,2.3169663,2.18462,2.0522738,1.9199274,1.7875811,2.7067533,3.6277382,4.5469103,5.467895,6.3870673,5.1578784,3.926877,2.6976883,1.4666867,0.2374981,0.23205921,0.22662032,0.2229944,0.21755551,0.21211663,1.1421664,2.0722163,3.002266,3.9323158,4.8623657,5.424384,5.9882154,6.550234,7.112252,7.6742706,8.149267,8.624263,9.099259,9.574255,10.049252,9.447348,8.845445,8.241728,7.6398244,7.037921,6.5574856,6.0770507,5.5966153,5.1179934,4.6375585,4.441758,4.2477713,4.0519714,3.8579843,3.6621845,4.4852695,5.3083544,6.1296263,6.9527116,7.7757964,7.440398,7.1050005,6.7696023,6.434204,6.1006193,5.6401267,5.179634,4.7191415,4.2604623,3.7999697,4.4743915,5.1506267,5.825049,6.4994707,7.175706,6.6173134,6.060734,5.5023413,4.945762,4.3873696,4.510651,4.632119,4.7554007,4.876869,5.0001507,5.1179934,5.235836,5.351866,5.469708,5.5875506,7.4349594,9.282369,11.129777,12.977186,14.824595,15.074784,15.324973,15.575162,15.825351,16.075539,15.198066,14.320591,13.443117,12.565643,11.6881695,10.130835,8.571687,7.0143523,5.4570174,3.8996825,5.4171324,6.9345818,8.452031,9.969481,11.486931,13.780329,16.071913,18.36531,20.656897,22.950293,22.930351,22.910408,22.890465,22.870523,22.85058,21.820818,20.789242,19.75948,18.729717,17.699953,15.694818,13.68968,11.684544,9.679407,7.6742706,7.3406854,7.0052876,6.6698895,6.3344913,6.000906,6.305484,6.6100616,6.9146395,7.219217,7.5256076,7.402326,7.2808576,7.157576,7.0342946,6.9128265,7.344311,7.7776093,8.210908,8.642392,9.07569,9.38752,9.699349,10.012992,10.324821,10.636651,10.845142,11.05182,11.26031,11.466989,11.675479,12.866595,14.059525,15.252454,16.445383,17.6365,18.354433,19.072367,19.7903,20.508232,21.224354,20.497355,19.770357,19.041546,18.314548,17.58755,17.890314,18.193079,18.495844,18.796797,19.099562,19.667019,20.234476,20.801933,21.36939,21.936848,20.042301,18.147755,16.25321,14.356851,12.462305,10.147152,7.8319983,5.516845,3.2016919,0.8883517,3.0620937,5.237649,7.413204,9.5869465,11.762501,10.114518,8.4683485,6.8203654,5.1723824,3.5243993,3.3267863,3.1291735,2.9333735,2.7357605,2.5381477,13.196554,23.85315,34.509743,45.168148,55.824745,47.05182,38.280704,29.507778,20.734854,11.961927,10.970237,9.976733,8.985043,7.993352,6.9998484,5.942891,4.8859344,3.827164,2.770207,1.7132497,1.4757515,1.2382535,1.0007553,0.76325727,0.52575916,0.6091554,0.69436467,0.7795739,0.86478317,0.9499924,1.0478923,1.1457924,1.2418793,1.3397794,1.4376793,1.9924458,2.5472124,3.101979,3.6567454,4.213325,7.0324817,9.851639,12.672608,15.491765,18.312735,17.092611,15.872487,14.652364,13.43224,12.212116,17.005589,21.797249,26.590723,31.382381,36.175854,30.98897,25.80571,20.620636,15.435563,10.25049,15.480887,20.70947,25.939869,31.170265,36.40066,42.59012,48.77957,54.970837,61.160294,67.34975,59.4271,51.506268,43.581806,35.65916,27.738327,35.588455,43.43677,51.28871,59.137028,66.98715,56.142014,45.298683,34.45173,23.606586,12.763257,12.5058155,12.248375,11.989121,11.731681,11.47424,18.983532,26.489197,33.998486,41.505966,49.013443,41.18507,33.358513,25.53014,17.701767,9.875207,9.89515,9.915092,9.935035,9.954978,9.97492,17.330109,24.685299,32.04049,39.395676,46.750866,55.367878,63.98489,72.603714,81.220726,89.83774,81.964035,74.092155,66.22027,58.34839,50.47469,48.163162,45.849823,43.538296,41.224957,38.91343,36.69799,34.482548,32.26711,30.051668,27.838041,26.82278,25.807522,24.792263,23.777004,22.761745,23.876717,24.99169,26.10666,27.221634,28.336605,31.05605,33.771866,36.4895,39.20713,41.92476,46.16528,50.4058,54.644505,58.885025,63.125546,62.420303,61.715057,61.009815,60.304573,59.59933,55.812054,52.024773,48.237495,44.45022,40.662937,43.317116,45.973106,48.62728,51.28327,53.93745,54.746033,55.5528,56.35957,57.168148,57.97492,57.7483,57.519863,57.293243,57.06481,56.83819,57.98942,59.142464,60.29551,61.44674,62.599785,62.110287,61.620785,61.12947,60.639973,60.15047,58.99924,57.849823,56.700405,55.549175,54.399754,51.70207,49.00438,46.30669,43.610813,40.913128,40.55416,40.197006,39.83985,39.4827,39.125546,41.268467,43.409576,45.552498,47.69542,49.83834,49.548267,49.258194,48.96812,48.678047,48.38797,46.90497,45.421963,43.940773,42.45777,40.974766,38.82822,36.67986,34.53331,32.38495,30.238403,29.51503,28.793472,28.070099,27.346727,26.625168,27.64224,28.659313,29.678198,30.695269,31.712341,31.485722,31.257288,31.030668,30.802235,30.575613,26.52727,22.480736,18.43239,14.385859,10.337513,8.694968,7.0524244,5.40988,3.7673361,2.124792,2.1954978,2.2643902,2.335096,2.4058013,2.474694,2.7720199,3.0693457,3.3666716,3.6658103,3.9631362,3.2180085,2.472881,1.7277533,0.9826257,0.2374981,1.1457924,2.0522738,2.960568,3.8670492,4.7753434,5.1941376,5.614745,6.035352,6.454147,6.874754,6.187641,5.5005283,4.8116026,4.12449,3.437377,3.7347028,4.0320287,4.329355,4.6266804,4.9258194,4.9294453,4.934884,4.940323,4.945762,4.949388,4.2767787,3.6041696,2.9333735,2.2607644,1.5881553,1.2944553,1.0025684,0.7106813,0.4169814,0.12509441,0.11059072,0.09427405,0.07977036,0.065266654,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.032633327,0.065266654,0.09789998,0.13053331,0.16316663,0.41516843,0.6671702,0.91917205,1.1729867,1.4249886,1.1657349,0.90466833,0.64541465,0.38434806,0.12509441,0.16497959,0.20486477,0.24474995,0.28463513,0.3245203,0.42967212,0.53482395,0.6399758,0.7451276,0.85027945,0.8974165,0.9445535,0.9916905,1.0406405,1.0877775,1.1349145,1.1820517,1.2291887,1.2781386,1.3252757,1.1204109,0.9155461,0.7106813,0.5058166,0.2991388,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.2374981,0.4749962,0.7124943,0.9499924,1.1874905,1.5881553,1.987007,2.3876717,2.7883365,3.1871881,2.6741197,2.1628644,1.649796,1.1367276,0.62547207,1.9253663,3.2252605,4.5251546,5.825049,7.124943,7.8247466,8.52455,9.224354,9.924157,10.625773,10.7871275,10.950294,11.111648,11.274815,11.437981,12.574709,13.713249,14.849977,15.986704,17.125244,19.850128,22.57501,25.299892,28.024776,30.749659,24.9373,19.124943,13.312584,7.500226,1.6878681,1.4630609,1.2382535,1.0116332,0.7868258,0.5620184,0.5493277,0.53663695,0.52575916,0.51306844,0.50037766,0.53663695,0.5747091,0.61278135,0.6508536,0.6871128,0.62547207,0.5620184,0.50037766,0.43692398,0.37528324,0.40066472,0.42423326,0.44961473,0.4749962,0.50037766,0.40066472,0.2991388,0.19942589,0.099712946,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.6000906,1.1367276,1.6751775,2.2118144,2.7502642,2.4873846,2.2245052,1.9616255,1.7005589,1.4376793,1.49932,1.5627737,1.6244144,1.6878681,1.7495089,2.8245957,3.8996825,4.974769,6.049856,7.124943,5.7380266,4.349297,2.962381,1.5754645,0.18673515,0.17585737,0.16316663,0.15047589,0.13778515,0.12509441,1.2491312,2.374981,3.5008307,4.6248674,5.750717,6.2365913,6.7242785,7.211965,7.699652,8.187339,8.013294,7.837437,7.663393,7.4875355,7.311678,7.462154,7.61263,7.763106,7.911769,8.062244,7.5999393,7.137634,6.6753283,6.2130227,5.750717,5.475147,5.199577,4.9258194,4.650249,4.3746786,4.8242936,5.275721,5.7253356,6.1749506,6.624565,6.6499467,6.6753283,6.70071,6.7242785,6.7496595,6.000906,5.2503395,4.499773,3.7492065,3.000453,4.07554,5.1506267,6.2257137,7.3008003,8.375887,7.4258947,6.4759026,5.524097,4.574105,3.6241121,3.774588,3.925064,4.07554,4.2242026,4.3746786,4.650249,4.9258194,5.199577,5.475147,5.750717,7.1865835,8.624263,10.061942,11.499621,12.937301,13.386916,13.838344,14.287958,14.737573,15.187187,14.262577,13.337966,12.413355,11.486931,10.56232,8.6877165,6.813113,4.936697,3.0620937,1.1874905,3.2742105,5.3627434,7.4494634,9.537996,11.624716,14.436621,17.25034,20.062244,22.87415,25.687866,25.46306,25.238253,25.011631,24.786825,24.562017,23.724428,22.886839,22.049252,21.211662,20.375887,17.937452,15.50083,13.062395,10.625773,8.187339,7.799365,7.413204,7.02523,6.637256,6.249282,6.4994707,6.7496595,6.9998484,7.250037,7.500226,7.4367723,7.3751316,7.311678,7.250037,7.1883965,7.650702,8.113008,8.575313,9.037619,9.499924,9.300498,9.099259,8.899834,8.700407,8.499168,8.337815,8.174648,8.013294,7.850128,7.686961,8.399456,9.11195,9.824444,10.536939,11.249433,12.988064,14.724882,16.4617,18.20033,19.93715,18.900135,17.863121,16.824293,15.787278,14.750263,14.750263,14.750263,14.750263,14.750263,14.750263,16.274965,17.799667,19.324368,20.850883,22.375584,20.424837,18.475903,16.525154,14.574407,12.625471,10.212419,7.799365,5.388125,2.9750717,0.5620184,3.388427,6.2130227,9.037619,11.862214,14.68681,12.112403,9.537996,6.9617763,4.3873696,1.8129625,1.987007,2.1628644,2.3369088,2.5127661,2.6868105,15.975826,29.261215,42.550232,55.837433,69.12463,56.161953,43.201084,30.23659,17.273907,4.313038,5.137936,5.962834,6.787732,7.61263,8.437528,7.0506115,5.661882,4.274966,2.8880494,1.49932,1.2001812,0.89922947,0.6000906,0.2991388,0.0,0.18673515,0.37528324,0.5620184,0.7505665,0.93730164,1.1004683,1.261822,1.4249886,1.5881553,1.7495089,2.3622901,2.9750717,3.587853,4.2006345,4.8116026,7.8755093,10.937603,13.999697,17.06179,20.125698,18.537542,16.949387,15.363045,13.77489,12.186734,18.675327,25.162107,31.650702,38.13748,44.62426,38.262577,31.90089,25.537392,19.175705,12.812206,19.34975,25.887293,32.424835,38.96238,45.499924,53.237648,60.975372,68.7131,76.45082,84.18673,73.26182,62.33872,51.41199,40.48708,29.562168,39.138237,48.71249,58.28856,67.862816,77.43707,64.83698,52.238705,39.636803,27.03671,14.436621,14.150173,13.861912,13.575464,13.287203,13.000754,22.449915,31.899076,41.35005,50.801025,60.250187,50.661427,41.074482,31.487534,21.900587,12.311829,12.299138,12.28826,12.27557,12.262879,12.250188,20.81281,29.375433,37.938053,46.50068,55.0633,65.11255,75.161804,85.21287,95.262115,105.31319,95.21136,85.11315,75.01133,64.913124,54.81311,52.374676,49.938053,47.49962,45.063,42.624565,39.136425,35.650097,32.161957,28.675629,25.187489,25.363346,25.537392,25.71325,25.887293,26.06315,26.211813,26.36229,26.512764,26.66324,26.811903,30.51216,34.212418,37.912674,41.61293,45.313187,49.774887,54.236588,58.700104,63.161804,67.62532,66.450516,65.27572,64.099106,62.924305,61.749504,57.712036,53.674572,49.637104,45.599636,41.56217,45.68847,49.81296,53.93745,58.06194,62.188244,62.561714,62.936996,63.31228,63.68756,64.06284,63.511703,62.962376,62.41305,61.861908,61.31258,62.67593,64.03747,65.40081,66.762344,68.125694,67.32436,66.52485,65.725334,64.92582,64.12449,62.637856,61.149414,59.662785,58.174343,56.687714,54.24928,51.812656,49.37422,46.937603,44.49917,43.78667,43.074177,42.361683,41.64919,40.936695,43.150322,45.362137,47.575764,49.78758,51.999393,52.612175,53.224957,53.837738,54.45052,55.0633,53.66188,52.26227,50.862667,49.46306,48.061638,45.211662,42.361683,39.511707,36.661728,33.811752,33.200783,32.588,31.975222,31.36244,30.749659,32.437527,34.125393,35.813263,37.499317,39.187187,38.98776,38.788334,38.587097,38.38767,38.188244,33.09926,28.012085,22.924911,17.837738,12.750566,10.687414,8.624263,6.5629244,4.499773,2.4366217,2.3876717,2.3369088,2.2879589,2.2371957,2.1882458,2.712192,3.2379513,3.7618973,4.2876563,4.8116026,3.8869917,2.962381,2.03777,1.1131591,0.18673515,1.1258497,2.0631514,3.000453,3.9377546,4.8750563,5.125245,5.375434,5.6256227,5.8758116,6.1241875,5.0744824,4.024777,2.9750717,1.9253663,0.87566096,1.649796,2.4257438,3.199879,3.975827,4.749962,5.0255322,5.2992897,5.57486,5.8504305,6.1241875,5.224958,4.325729,3.4246864,2.525457,1.6244144,1.3252757,1.0243238,0.72518504,0.42423326,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.50037766,0.8122072,1.1258497,1.4376793,1.7495089,1.4249886,1.1004683,0.774135,0.44961473,0.12509441,0.13778515,0.15047589,0.16316663,0.17585737,0.18673515,0.2991388,0.41335547,0.52575916,0.63816285,0.7505665,0.8629702,0.97537386,1.0877775,1.2001812,1.3125849,1.3742256,1.4376793,1.49932,1.5627737,1.6244144,1.3742256,1.1258497,0.87566096,0.62547207,0.37528324,0.31182957,0.25018883,0.18673515,0.12509441,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.19579996,0.38978696,0.5855869,0.7795739,0.97537386,1.2944553,1.6153497,1.9344311,2.2553256,2.5744069,2.1646774,1.7549478,1.3452182,0.9354887,0.52575916,1.9108626,3.294153,4.6792564,6.0643597,7.4494634,7.8247466,8.200029,8.575313,8.950596,9.325879,9.7773075,10.230548,10.681975,11.135216,11.586644,12.032633,12.476809,12.922797,13.366973,13.812962,16.091856,18.372562,20.653269,22.932163,25.212872,20.45203,15.693004,10.932164,6.1731377,1.4122978,1.2255627,1.0370146,0.85027945,0.66173136,0.4749962,0.4604925,0.44417584,0.42967212,0.41516843,0.40066472,0.45324063,0.5058166,0.55839247,0.6091554,0.66173136,0.58921283,0.5166943,0.44417584,0.37165734,0.2991388,0.3208944,0.34083697,0.36077955,0.38072214,0.40066472,0.32814622,0.25562772,0.18310922,0.11059072,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.4894999,0.91735905,1.3452182,1.7730774,2.1991236,2.1882458,2.175555,2.1628644,2.1501737,2.137483,2.124792,2.1121013,2.0994108,2.08672,2.0758421,2.808279,3.540716,4.273153,5.0055895,5.7380266,4.6194286,3.5026438,2.3858588,1.2672608,0.15047589,0.13959812,0.13053331,0.11965553,0.11059072,0.099712946,1.0007553,1.8999848,2.7992141,3.7002566,4.599486,5.0019636,5.4044414,5.806919,6.209397,6.6118746,6.4795284,6.347182,6.2148356,6.0824895,5.9501433,6.0643597,6.1803894,6.294606,6.4106355,6.5248523,6.2728505,6.0208488,5.767034,5.5150323,5.2630305,5.0200934,4.7771564,4.5342193,4.2930956,4.0501585,4.599486,5.1506267,5.6999545,6.249282,6.8004227,6.736969,6.6753283,6.6118746,6.550234,6.48678,5.7597823,5.032784,4.305786,3.576975,2.8499773,3.7256382,4.599486,5.475147,6.350808,7.224656,6.742408,6.26016,5.7779117,5.295664,4.8116026,5.4552045,6.096993,6.740595,7.382384,8.024173,7.7322855,7.440398,7.1466985,6.8548117,6.5629244,8.029612,9.498111,10.964798,12.433297,13.899984,15.484513,17.069042,18.655384,20.239914,21.824444,19.730473,17.634687,15.540715,13.44493,11.349146,9.655839,7.9607186,6.265599,4.5704784,2.8753586,5.275721,7.6742706,10.074633,12.474996,14.875358,17.400814,19.92446,22.449915,24.975372,27.50083,27.212568,26.924307,26.63786,26.349598,26.06315,24.60009,23.137028,21.675781,20.212719,18.749659,16.788034,14.824595,12.862969,10.899531,8.937905,8.178274,7.41683,6.6571984,5.8975673,5.137936,5.6056805,6.071612,6.539356,7.0071006,7.474845,7.2754188,7.07418,6.874754,6.6753283,6.4759026,7.224656,7.9752226,8.725789,9.474543,10.225109,10.223296,10.21967,10.217857,10.2142315,10.212419,9.815379,9.418341,9.019489,8.62245,8.225411,9.050309,9.875207,10.700105,11.525003,12.349901,13.318023,14.284332,15.252454,16.220575,17.186886,16.52334,15.857984,15.192626,14.527269,13.861912,13.832905,13.802084,13.773077,13.742256,13.713249,14.924308,16.13718,17.350052,18.562923,19.775795,18.410635,17.045475,15.680313,14.315152,12.949992,10.662033,8.375887,6.0879283,3.7999697,1.5120108,4.365614,7.217404,10.069194,12.922797,15.774588,13.143979,10.515183,7.8845744,5.2557783,2.6251698,2.9841363,3.3449159,3.7056956,4.064662,4.4254417,14.978697,25.53014,36.083393,46.63484,57.18809,47.65191,38.11754,28.581356,19.046986,9.512614,10.07282,10.633025,11.193231,11.751623,12.311829,10.471672,8.6333275,6.793171,4.953014,3.1128569,3.4228733,3.73289,4.0429068,4.3529234,4.6629395,3.972201,3.2832751,2.5925364,1.9017978,1.2128719,2.2879589,3.3630457,4.4381323,5.5132194,6.588306,6.4577727,6.3272395,6.1967063,6.0679855,5.9374523,8.337815,10.738177,13.136727,15.537089,17.937452,16.574104,15.212569,13.849221,12.487686,11.124338,16.757214,22.390087,28.022963,33.655838,39.2869,36.29551,33.30231,30.309109,27.31772,24.324518,26.868105,29.40988,31.953466,34.49524,37.037014,43.253662,49.466682,55.683334,61.898167,68.11301,59.439793,50.76839,42.095177,33.421967,24.750565,34.27587,43.799362,53.32467,62.849976,72.37528,60.53845,48.70524,36.87022,25.0352,13.200181,13.472125,13.745882,14.017827,14.289771,14.561715,21.49811,28.432692,35.367275,42.301857,49.23825,41.745277,34.2523,26.759327,19.268166,11.775192,12.380721,12.984438,13.589968,14.195497,14.799213,21.315,27.828976,34.344765,40.86055,47.374527,56.290676,65.20501,74.12116,83.0355,91.94984,83.26937,74.59072,65.910255,57.22979,48.549324,46.326633,44.105755,41.88306,39.66037,37.437675,34.83064,32.221783,29.614744,27.007704,24.400663,24.344461,24.290073,24.235683,24.179482,24.125093,23.912977,23.70086,23.48693,23.274813,23.062696,26.45475,29.846804,33.24067,36.63272,40.024776,44.07312,48.11965,52.168,56.21453,60.262875,59.40172,58.542374,57.68303,56.821873,55.96253,52.982018,50.003323,47.02281,44.0423,41.06179,44.557182,48.052574,51.547966,55.043358,58.536938,58.689224,58.843327,58.995617,59.147903,59.300194,59.28569,59.26937,59.254868,59.240364,59.22586,60.43692,61.64979,62.862663,64.07554,65.28841,64.367424,63.44825,62.527267,61.608093,60.68711,59.265747,57.84257,56.419395,54.99803,53.574856,51.40474,49.234623,47.06451,44.894394,42.724277,41.638313,40.550533,39.462757,38.374977,37.2872,38.84091,40.392807,41.944702,43.498413,45.05031,45.74286,46.43541,47.127964,47.820515,48.513065,48.183105,47.853146,47.52319,47.19323,46.86327,44.952408,43.043358,41.132496,39.221634,37.312584,35.876717,34.44266,33.006798,31.572742,30.136877,31.208338,32.277985,33.347633,34.417282,35.48693,35.76069,36.03263,36.304577,36.578335,36.850277,32.780178,28.710075,24.639975,20.569874,16.499773,14.025079,11.5503845,9.07569,6.599184,4.12449,4.0356545,3.9450066,3.8543584,3.7655232,3.6748753,4.1444325,4.615803,5.08536,5.5549173,6.0244746,5.5893636,5.1542525,4.7191415,4.2858434,3.8507326,4.699199,5.5494785,6.399758,7.250037,8.100317,7.989726,7.8791356,7.7703576,7.6597667,7.549176,6.2873545,5.0255322,3.7618973,2.5000753,1.2382535,1.7603867,2.2825198,2.8046532,3.3267863,3.8507326,4.5867953,5.3246713,6.0625467,6.8004227,7.5382986,6.6082487,5.678199,4.748149,3.8180993,2.8880494,2.3495996,1.8129625,1.2745126,0.73787576,0.19942589,0.2955129,0.38978696,0.48587397,0.58014804,0.6744221,0.54570174,0.41516843,0.28463513,0.15410182,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.15047589,0.40066472,0.6508536,0.89922947,1.1494182,1.3996071,1.1693609,0.93911463,0.7106813,0.48043507,0.25018883,0.26831847,0.28463513,0.30276474,0.3208944,0.33721104,0.4550536,0.5728962,0.69073874,0.80676836,0.9246109,0.99531645,1.064209,1.1349145,1.2056202,1.2745126,1.2980812,1.3198367,1.3434052,1.3651608,1.3869164,1.1802386,0.97174793,0.7650702,0.55839247,0.34990177,0.2991388,0.25018883,0.19942589,0.15047589,0.099712946,0.08339628,0.065266654,0.047137026,0.030820364,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.15228885,0.3045777,0.45686656,0.6091554,0.76325727,1.0025684,1.2418793,1.4830034,1.7223145,1.9616255,1.6552348,1.3470312,1.0406405,0.7324369,0.42423326,1.8945459,3.3648586,4.835171,6.305484,7.7757964,7.8247466,7.8755093,7.9244595,7.9752226,8.024173,8.767487,9.510801,10.252303,10.995618,11.73712,11.490557,11.242181,10.995618,10.747242,10.500679,12.335398,14.170115,16.004833,17.839552,19.67427,15.966762,12.259253,8.551744,4.844236,1.1367276,0.9880646,0.8375887,0.6871128,0.53663695,0.387974,0.36984438,0.35171473,0.33539808,0.31726846,0.2991388,0.3680314,0.43511102,0.50219065,0.56927025,0.63816285,0.55476654,0.47318324,0.38978696,0.30820364,0.22480737,0.23931105,0.25562772,0.27013144,0.28463513,0.2991388,0.25562772,0.21030366,0.16497959,0.11965553,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.38072214,0.6979906,1.015259,1.3325275,1.649796,1.887294,2.124792,2.3622901,2.5997884,2.8372865,2.7502642,2.663242,2.5744069,2.4873846,2.4003625,2.7901495,3.1799364,3.5697234,3.9595103,4.349297,3.5026438,2.6541772,1.8075237,0.96087015,0.11240368,0.10515183,0.09789998,0.09064813,0.08339628,0.07433146,0.7505665,1.4249886,2.0994108,2.7756457,3.4500678,3.7673361,4.0846047,4.401873,4.7191415,5.038223,4.947575,4.856927,4.7680917,4.6774435,4.5867953,4.668379,4.748149,4.8279195,4.9076896,4.98746,4.945762,4.902251,4.860553,4.8170414,4.7753434,4.5650396,4.3547363,4.1444325,3.9341288,3.7256382,4.3746786,5.0255322,5.674573,6.3254266,6.9744673,6.825804,6.6753283,6.5248523,6.3743763,6.2257137,5.520471,4.8152285,4.1099863,3.4047437,2.6995013,3.3757362,4.0501585,4.7245803,5.4008155,6.0752378,6.060734,6.0444174,6.0299134,6.01541,6.000906,7.135821,8.270736,9.40565,10.540565,11.675479,10.8143215,9.954978,9.0956335,8.234476,7.3751316,8.872639,10.370146,11.867653,13.36516,14.862667,17.582111,20.301556,23.022812,25.742256,28.4617,25.198366,21.933222,18.668076,15.40293,12.137785,10.622148,9.108324,7.592687,6.0770507,4.5632267,7.2754188,9.987611,12.699803,15.411995,18.124187,20.363195,22.600391,24.837587,27.074783,29.31198,28.962078,28.612175,28.262274,27.912373,27.56247,25.47575,23.387217,21.300497,19.211964,17.125244,15.636803,14.150173,12.661731,11.175101,9.686659,8.55537,7.422269,6.2891674,5.1578784,4.024777,4.710077,5.3953767,6.0806766,6.7641635,7.4494634,7.112252,6.775041,6.43783,6.1006193,5.7615952,6.8004227,7.837437,8.874452,9.91328,10.950294,11.144281,11.340081,11.535881,11.729868,11.925668,11.292944,10.66022,10.027496,9.394773,8.762048,9.699349,10.636651,11.575767,12.513068,13.45037,13.647983,13.845595,14.043208,14.240821,14.436621,14.144734,13.852847,13.559147,13.267261,12.975373,12.915545,12.855718,12.79589,12.734249,12.674421,13.575464,14.474693,15.375735,16.274965,17.174194,16.39462,15.6150465,14.835473,14.054086,13.274512,11.111648,8.950596,6.787732,4.6248674,2.4620032,5.3428006,8.221786,11.102583,13.98338,16.862366,14.177367,11.49237,8.807372,6.1223745,3.437377,3.9830787,4.5269675,5.0726695,5.618371,6.16226,13.979754,21.797249,29.614744,37.43224,45.249733,39.14186,33.035805,26.927933,20.820063,14.712192,15.007704,15.303217,15.596917,15.89243,16.187943,13.894546,11.602961,9.309563,7.017978,4.7245803,5.6455655,6.5647373,7.4857225,8.404895,9.325879,7.757667,6.189454,4.6230545,3.054842,1.4866294,3.4754493,5.462456,7.4494634,9.438283,11.42529,10.553255,9.679407,8.807372,7.935337,7.063302,8.80012,10.536939,12.27557,14.012388,15.749206,14.612478,13.475751,12.337211,11.200482,10.061942,14.840912,19.618069,24.395224,29.17238,33.94954,34.326633,34.705544,35.082638,35.459736,35.83683,34.384647,32.932465,31.480282,30.0281,28.574102,33.267864,37.959812,42.651756,47.345516,52.037464,45.617764,39.198063,32.77655,26.35685,19.93715,29.413506,38.888046,48.36259,57.83713,67.311676,56.241726,45.173588,34.101826,23.031878,11.961927,12.79589,13.628039,14.46019,15.292339,16.124489,20.544493,24.964495,29.384497,33.8045,38.224503,32.827312,27.430124,22.032934,16.635744,11.236742,12.460492,13.682428,14.904366,16.128115,17.350052,21.817192,26.284332,30.753284,35.220425,39.687565,47.4688,55.24641,63.027645,70.80707,78.5883,71.327385,64.06828,56.80737,49.546455,42.287354,40.280403,38.27164,36.26469,34.25774,32.25079,30.523039,28.795284,27.067532,25.339779,23.612024,23.327389,23.042755,22.75812,22.471672,22.187037,21.612328,21.037619,20.462908,19.888199,19.311678,22.397339,25.483002,28.56685,31.652514,34.738174,38.36954,42.002716,45.635895,49.267258,52.900436,52.354733,51.810844,51.265144,50.71944,50.175552,48.252,46.330257,44.406704,42.484966,40.563225,43.427704,46.292187,49.156666,52.02296,54.887444,54.81674,54.747845,54.67714,54.608246,54.53754,55.05786,55.578182,56.096687,56.61701,57.13733,58.199726,59.26212,60.324516,61.386913,62.44931,61.41048,60.369843,59.3292,58.290375,57.249733,55.891823,54.53573,53.17782,51.81991,50.462,48.560204,46.658405,44.754795,42.852997,40.949387,39.488136,38.025078,36.562016,35.10077,33.637707,34.529686,35.42166,36.315453,37.20743,38.099407,38.87173,39.644054,40.418186,41.19051,41.962833,42.702522,43.44221,44.1819,44.9234,45.66309,44.693153,43.723217,42.753284,41.783348,40.813416,38.554462,36.297325,34.040184,31.783047,29.524096,29.977337,30.430576,30.882004,31.335245,31.786673,32.5318,33.276928,34.022057,34.767185,35.51231,32.459282,29.408066,26.355038,23.302008,20.250792,17.362743,14.474693,11.586644,8.700407,5.812358,5.6818247,5.5531044,5.422571,5.292038,5.163317,5.576673,5.9918413,6.4070096,6.8221784,7.2373466,7.2917356,7.3479376,7.402326,7.456715,7.512917,8.274362,9.037619,9.800876,10.56232,11.325577,10.854207,10.384649,9.915092,9.445535,8.974165,7.500226,6.0244746,4.550536,3.0747845,1.6008459,1.8691645,2.1392958,2.4094272,2.6795588,2.94969,4.1498713,5.3500524,6.550234,7.750415,8.950596,7.989726,7.0306687,6.069799,5.1107416,4.1498713,3.3757362,2.5997884,1.8256533,1.0497054,0.2755703,0.47680917,0.67986095,0.88291276,1.0841516,1.2872034,1.0406405,0.79226464,0.54570174,0.29732585,0.05076295,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.2991388,0.48768693,0.6744221,0.8629702,1.0497054,0.9155461,0.7795739,0.64541465,0.5094425,0.37528324,0.39703882,0.42060733,0.44236287,0.46411842,0.48768693,0.6091554,0.7324369,0.8557183,0.97718686,1.1004683,1.1276628,1.1548572,1.1820517,1.209246,1.2382535,1.2201238,1.2019942,1.1856775,1.167548,1.1494182,0.98443866,0.8194591,0.6544795,0.4894999,0.3245203,0.28826106,0.25018883,0.21211663,0.17585737,0.13778515,0.11421664,0.092461094,0.07070554,0.047137026,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.11059072,0.21936847,0.32995918,0.4405499,0.5493277,0.7106813,0.87022203,1.0297627,1.1893034,1.3506571,1.1457924,0.93911463,0.73424983,0.5293851,0.3245203,1.8800422,3.435564,4.989273,6.544795,8.100317,7.8247466,7.549176,7.2754188,6.9998484,6.7242785,7.757667,8.789243,9.822631,10.854207,11.887595,10.946668,10.007553,9.066626,8.127511,7.1865835,8.577126,9.967669,11.358211,12.74694,14.137483,11.483305,8.827314,6.1731377,3.5171473,0.8629702,0.7505665,0.63816285,0.52575916,0.41335547,0.2991388,0.27919623,0.25925365,0.23931105,0.21936847,0.19942589,0.28282216,0.36440548,0.44780177,0.5293851,0.61278135,0.52032024,0.42785916,0.33539808,0.24293698,0.15047589,0.15954071,0.17041849,0.1794833,0.19036107,0.19942589,0.18310922,0.16497959,0.14684997,0.13053331,0.11240368,0.09064813,0.06707962,0.045324065,0.02175555,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.27013144,0.47680917,0.6852999,0.8919776,1.1004683,1.5881553,2.0758421,2.561716,3.049403,3.53709,3.3757362,3.2125697,3.049403,2.8880494,2.7248828,2.7720199,2.819157,2.8681068,2.9152439,2.962381,2.3858588,1.8075237,1.2291887,0.6526665,0.07433146,0.07070554,0.065266654,0.059827764,0.054388877,0.05076295,0.50037766,0.9499924,1.3996071,1.8492218,2.3006494,2.5327086,2.764768,2.9968271,3.2306993,3.4627585,3.4156215,3.3666716,3.3195345,3.2723975,3.2252605,3.2705846,3.3140955,3.3594196,3.4047437,3.4500678,3.6168604,3.785466,3.9522583,4.120864,4.2876563,4.1099863,3.9323158,3.7546456,3.576975,3.3993049,4.1498713,4.900438,5.6491914,6.399758,7.1503243,6.9128265,6.6753283,6.43783,6.200332,5.962834,5.279347,4.597673,3.9141862,3.2325122,2.5508385,3.0258346,3.5008307,3.975827,4.4508233,4.9258194,5.377247,5.8304877,6.281915,6.735156,7.1883965,8.814624,10.442664,12.070704,13.696932,15.324973,13.898171,12.469557,11.042755,9.6141405,8.187339,9.715667,11.242181,12.770509,14.297023,15.825351,19.679708,23.535881,27.390238,31.244596,35.10077,30.66445,26.229942,21.795437,17.359118,12.92461,11.59027,10.255929,8.919776,7.5854354,6.249282,9.275117,12.299138,15.324973,18.350807,21.374828,23.325577,25.274511,27.22526,29.174194,31.12494,30.7134,30.300043,29.886688,29.475145,29.06179,26.349598,23.637405,20.925215,18.213022,15.50083,14.487384,13.475751,12.462305,11.450671,10.437225,8.9324665,7.4277077,5.922949,4.41819,2.911618,3.8144734,4.7173285,5.620184,6.5230393,7.4258947,6.9508986,6.4759026,5.999093,5.524097,5.049101,6.3743763,7.699652,9.024928,10.3502035,11.675479,12.067079,12.460492,12.852092,13.245504,13.637105,12.770509,11.9021,11.035503,10.167094,9.300498,10.3502035,11.399909,12.449615,13.499319,14.5508375,13.9779415,13.4050455,12.8321495,12.259253,11.6881695,11.7679405,11.847711,11.927481,12.007251,12.087022,11.998186,11.907538,11.81689,11.728055,11.637406,12.224807,12.812206,13.399607,13.987006,14.574407,14.380419,14.184619,13.990632,13.794832,13.600845,11.563075,9.525306,7.4875355,5.4497657,3.4119956,6.319988,9.22798,12.135971,15.0421505,17.950142,15.210756,12.469557,9.73017,6.9907837,4.249584,4.9802084,5.710832,6.439643,7.170267,7.900891,12.982625,18.06436,23.147905,28.229641,33.311375,30.631815,27.952257,25.272697,22.59314,19.911768,19.942589,19.97341,20.002417,20.033237,20.062244,17.31742,14.572594,11.827768,9.082943,6.338117,7.8682575,9.398398,10.928538,12.456866,13.987006,11.543133,9.097446,6.6517596,4.207886,1.7621996,4.6629395,7.5618668,10.462607,13.363347,16.262274,14.646925,13.033388,11.418038,9.802689,8.187339,9.262425,10.337513,11.4126,12.487686,13.562773,12.64904,11.73712,10.825199,9.91328,8.999546,12.922797,16.844234,20.767487,24.690737,28.612175,32.35957,36.106964,39.854355,43.60356,47.350956,41.903004,36.45505,31.0071,25.559147,20.113007,23.282066,26.452936,29.621996,32.792866,35.961926,31.793924,27.627737,23.459736,19.291735,15.125546,24.55114,33.97492,43.400513,52.82429,62.24988,51.945004,41.640125,31.335245,21.030367,10.725487,12.117842,13.510198,14.902553,16.294909,17.687263,19.592686,21.49811,23.401722,25.307144,27.212568,23.909351,20.607946,17.304728,14.00151,10.700105,12.540262,14.380419,16.220575,18.060734,19.90089,22.319382,24.739687,27.159992,29.580297,32.000603,38.64511,45.28962,51.934128,58.58045,65.22495,59.38359,53.544037,47.704483,41.864933,36.02538,34.23236,32.43934,30.648132,28.855112,27.062092,26.215439,25.366972,24.520319,23.671852,22.8252,22.310318,21.795437,21.280556,20.765673,20.250792,19.311678,18.374376,17.437075,16.499773,15.56247,18.33993,21.117388,23.894846,26.672306,29.449764,32.667774,35.88397,39.10198,42.319984,45.537994,45.307747,45.077503,44.847256,44.61701,44.386765,43.52198,42.657196,41.79241,40.92763,40.062847,42.29823,44.5318,46.76718,49.002567,51.23795,50.94425,50.652363,50.360474,50.066776,49.774887,50.830032,51.885178,52.94032,53.995464,55.05061,55.96253,56.87445,57.78818,58.700104,59.612022,58.451725,57.293243,56.132946,54.972652,53.812355,52.519714,51.22707,49.93443,48.641785,47.349144,45.715664,44.08037,42.44508,40.809788,39.174496,37.337963,35.49962,33.66309,31.824745,29.988214,30.220274,30.452332,30.684391,30.91645,31.150324,32.002415,32.854507,33.7066,34.560505,35.412598,37.221935,39.033085,40.842422,42.651756,44.462906,44.432087,44.40308,44.37226,44.34325,44.31243,41.23221,38.151985,35.071762,31.993351,28.913128,28.748148,28.583168,28.418188,28.253208,28.08823,29.304728,30.523039,31.739536,32.957848,34.174343,32.1402,30.104244,28.070099,26.035955,23.999998,20.700407,17.400814,14.09941,10.799818,7.500226,7.3298078,7.159389,6.9907837,6.8203654,6.6499467,7.0107265,7.369693,7.7304726,8.089439,8.450218,8.99592,9.539809,10.085511,10.629399,11.175101,11.849524,12.525759,13.200181,13.874602,14.5508375,13.720501,12.890164,12.059827,11.22949,10.399154,8.713099,7.02523,5.337362,3.6494937,1.9616255,1.9797552,1.9978848,2.0142014,2.032331,2.0504606,3.7129474,5.375434,7.037921,8.700407,10.362894,9.373016,8.383139,7.3932614,6.4033837,5.411693,4.40006,3.388427,2.374981,1.3633479,0.34990177,0.65991837,0.969935,1.2799516,1.5899682,1.8999848,1.5355793,1.1693609,0.80495536,0.4405499,0.07433146,0.07433146,0.07433146,0.07433146,0.07433146,0.07433146,0.19942589,0.3245203,0.44961473,0.5747091,0.69980353,0.65991837,0.6200332,0.58014804,0.5402629,0.50037766,0.5275721,0.55476654,0.581961,0.6091554,0.63816285,0.7650702,0.8919776,1.020698,1.1476053,1.2745126,1.260009,1.2455053,1.2291887,1.214685,1.2001812,1.1421664,1.0841516,1.0279498,0.969935,0.9119202,0.7904517,0.6671702,0.54570174,0.4224203,0.2991388,0.2755703,0.25018883,0.22480737,0.19942589,0.17585737,0.14684997,0.11965553,0.092461094,0.065266654,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06707962,0.13415924,0.2030518,0.27013144,0.33721104,0.4169814,0.49675176,0.57833505,0.65810543,0.73787576,0.6345369,0.533011,0.42967212,0.32814622,0.22480737,1.8655385,3.5044568,5.145188,6.7859187,8.424837,7.8247466,7.224656,6.624565,6.0244746,5.424384,6.7478466,8.069496,9.39296,10.714609,12.038072,10.4045925,8.772926,7.1394467,5.5077806,3.874301,4.8206677,5.765221,6.7097745,7.654328,8.600695,6.9980354,5.3953767,3.7927177,2.1900587,0.5873999,0.51306844,0.43692398,0.36259252,0.28826106,0.21211663,0.19036107,0.16679256,0.14503701,0.12328146,0.099712946,0.19761293,0.2955129,0.39159992,0.4894999,0.5873999,0.48587397,0.3825351,0.27919623,0.17767033,0.07433146,0.07977036,0.08520924,0.09064813,0.09427405,0.099712946,0.11059072,0.11965553,0.13053331,0.13959812,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.15954071,0.2574407,0.35534066,0.45324063,0.5493277,1.2872034,2.0250793,2.762955,3.5008307,4.2368937,3.9993954,3.7618973,3.5243993,3.2869012,3.049403,2.7557032,2.4601903,2.1646774,1.8691645,1.5754645,1.2672608,0.96087015,0.6526665,0.3444629,0.038072214,0.034446288,0.032633327,0.030820364,0.027194439,0.025381476,0.25018883,0.4749962,0.69980353,0.9246109,1.1494182,1.2980812,1.4449311,1.5917811,1.7404441,1.887294,1.8818551,1.8782293,1.8727903,1.8673514,1.8619126,1.8727903,1.8818551,1.892733,1.9017978,1.9126755,2.2897718,2.666868,3.045777,3.4228733,3.7999697,3.6549325,3.5098956,3.3648586,3.2198215,3.0747845,3.925064,4.7753434,5.6256227,6.4759026,7.324369,6.9998484,6.6753283,6.350808,6.0244746,5.6999545,5.040036,4.3801174,3.720199,3.0602808,2.4003625,2.6741197,2.94969,3.2252605,3.5008307,3.774588,4.695573,5.614745,6.53573,7.454902,8.375887,10.49524,12.6145935,14.73576,16.855114,18.974466,16.980207,14.985949,12.989877,10.995618,8.999546,10.556881,12.114216,13.673364,15.230699,16.788034,21.777306,26.766579,31.757666,36.746937,41.738026,36.132343,30.528477,24.922796,19.317116,13.713249,12.558392,11.401722,10.246864,9.092008,7.93715,11.274815,14.612478,17.950142,21.287807,24.625471,26.287958,27.950443,29.61293,31.275417,32.937904,32.46291,31.987911,31.512915,31.03792,30.562923,27.22526,23.887594,20.54993,17.212267,13.874602,13.337966,12.799516,12.262879,11.724429,11.187792,9.309563,7.4331465,5.5549173,3.6766882,1.8002719,2.9206827,4.0392804,5.1596913,6.2801023,7.400513,6.787732,6.1749506,5.562169,4.949388,4.3366065,5.9501433,7.5618668,9.175404,10.7871275,12.400664,12.989877,13.580903,14.170115,14.759329,15.350354,14.248073,13.145792,12.0416975,10.939416,9.837135,10.999244,12.163166,13.325275,14.487384,15.649493,14.3079,12.964496,11.622903,10.279498,8.937905,9.389333,9.842574,10.2958145,10.747242,11.200482,11.080828,10.959359,10.839704,10.720048,10.600392,10.874149,11.14972,11.42529,11.700861,11.974618,12.364405,12.754191,13.145792,13.535579,13.925365,12.012691,10.100015,8.187339,6.2746634,4.361988,7.2971745,10.232361,13.167547,16.102734,19.03792,16.242332,13.446743,10.652968,7.85738,5.0617914,5.977338,6.892884,7.8084297,8.722163,9.637709,11.985496,14.33147,16.679256,19.027042,21.374828,22.121769,22.870523,23.617464,24.364405,25.113157,24.877472,24.641787,24.407915,24.17223,23.938358,20.740292,17.542227,14.34416,11.147907,7.949841,10.09095,12.230246,14.369541,16.51065,18.649946,15.326786,12.005438,8.682278,5.3591175,2.03777,5.8504305,9.663091,13.475751,17.288412,21.099258,18.742407,16.385555,14.026892,11.67004,9.313189,9.724731,10.138086,10.549629,10.962985,11.374527,10.687414,10.000301,9.313189,8.624263,7.93715,11.004683,14.072216,17.139748,20.207281,23.274813,30.392506,37.510197,44.627888,51.74558,58.86327,49.419548,39.97764,30.533916,21.092007,11.650098,13.29808,14.94425,16.592234,18.240217,19.886387,17.971897,16.05741,14.142921,12.22662,10.312131,19.688774,29.06179,38.43843,47.813263,57.18809,47.64647,38.108475,28.56685,19.027042,9.487233,11.439794,13.392355,15.344915,17.297476,19.250036,18.639069,18.029913,17.420757,16.80979,16.200634,14.991387,13.785768,12.576522,11.369088,10.161655,12.620032,15.076597,17.534973,19.993351,22.449915,22.823385,23.195044,23.5667,23.94017,24.311829,29.823235,35.33283,40.842422,46.352013,51.861607,47.441605,43.021603,38.6016,34.181595,29.761593,28.184317,26.607038,25.029762,23.452484,21.875206,21.90784,21.940474,21.973106,22.00574,22.038374,21.293245,20.548119,19.80299,19.057863,18.312735,17.01284,15.712947,14.413053,13.113158,11.813264,14.282519,16.751774,19.222843,21.692097,24.163166,26.964193,29.767033,32.569874,35.37271,38.175552,38.26076,38.34416,38.429367,38.514576,38.599785,38.79196,38.984135,39.17812,39.370296,39.56247,41.166943,42.773228,44.377697,45.98217,47.586643,47.071762,46.55688,46.041996,45.527115,45.012234,46.602203,48.192173,49.78214,51.37211,52.962074,53.725334,54.48678,55.250034,56.01329,56.774734,55.494785,54.214832,52.934883,51.65493,50.374977,49.147602,47.920227,46.692852,45.465477,44.2381,42.869312,41.50234,40.135365,38.76658,37.399605,35.18779,32.974163,30.762348,28.550535,26.336908,25.909048,25.483002,25.055143,24.627283,24.199425,25.1331,26.064962,26.996826,27.930502,28.862364,31.743162,34.622147,37.502945,40.381927,43.262726,44.172832,45.08294,45.99305,46.903156,47.813263,43.909954,40.008457,36.10515,32.201843,28.300346,27.517145,26.73576,25.952559,25.16936,24.387972,26.077654,27.767334,29.457016,31.146698,32.838192,31.819305,30.802235,29.785162,28.768091,27.749205,24.03807,20.325123,16.612177,12.899229,9.188094,8.977791,8.767487,8.557183,8.34688,8.138389,8.442966,8.747544,9.052122,9.3567,9.663091,10.698292,11.731681,12.766883,13.802084,14.837286,15.4246855,16.012085,16.599485,17.186886,17.774284,16.584982,15.3956785,14.204562,13.015259,11.8241415,9.924157,8.024173,6.1241875,4.2260156,2.324218,2.0903459,1.8546607,1.6207886,1.3851035,1.1494182,3.2760234,5.4008155,7.5256076,9.6504,11.775192,10.754494,9.735609,8.714911,7.6942134,6.6753283,5.424384,4.175253,2.9243085,1.6751775,0.42423326,0.8430276,1.260009,1.6769904,2.0957847,2.5127661,2.030518,1.54827,1.064209,0.581961,0.099712946,0.0870222,0.07433146,0.06164073,0.05076295,0.038072214,0.099712946,0.16316663,0.22480737,0.28826106,0.34990177,0.40429065,0.4604925,0.5148814,0.56927025,0.62547207,0.65810543,0.69073874,0.72337204,0.7541924,0.7868258,0.91917205,1.0533313,1.1856775,1.3180238,1.4503701,1.3923552,1.3343405,1.2781386,1.2201238,1.162109,1.064209,0.968122,0.87022203,0.77232206,0.6744221,0.5946517,0.5148814,0.43511102,0.35534066,0.2755703,0.26287958,0.25018883,0.2374981,0.22480737,0.21211663,0.1794833,0.14684997,0.11421664,0.08339628,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,1.8492218,3.5751622,5.2992897,7.02523,8.749357,7.8247466,6.9001355,5.975525,5.049101,4.12449,5.7380266,7.3497505,8.963287,10.57501,12.186734,9.862516,7.5382986,5.2122674,2.8880494,0.5620184,1.062396,1.5627737,2.0631514,2.561716,3.0620937,2.5127661,1.9616255,1.4122978,0.8629702,0.31182957,0.2755703,0.2374981,0.19942589,0.16316663,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.11240368,0.22480737,0.33721104,0.44961473,0.5620184,0.44961473,0.33721104,0.22480737,0.11240368,0.0,0.0,0.0,0.0,0.0,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.9880646,1.9743162,2.962381,3.9504454,4.936697,4.6248674,4.313038,3.9993954,3.6875658,3.3757362,2.7375734,2.0994108,1.4630609,0.824898,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06164073,0.12509441,0.18673515,0.25018883,0.31182957,0.34990177,0.387974,0.42423326,0.46230546,0.50037766,0.4749962,0.44961473,0.42423326,0.40066472,0.37528324,0.96268314,1.550083,2.137483,2.7248828,3.3122826,3.199879,3.0874753,2.9750717,2.8626678,2.7502642,3.7002566,4.650249,5.600241,6.550234,7.500226,7.0868707,6.6753283,6.261973,5.8504305,5.4370747,4.800725,4.162562,3.5243993,2.8880494,2.2498865,2.324218,2.4003625,2.474694,2.5508385,2.6251698,4.0120864,5.4008155,6.787732,8.174648,9.563377,12.175857,14.786523,17.400814,20.013294,22.625772,20.062244,17.500528,14.936998,12.375282,9.811753,11.399909,12.988064,14.574407,16.162561,17.750717,23.874905,29.999092,36.12509,42.24928,48.375282,41.60024,34.8252,28.050158,21.275116,14.500074,13.524701,12.549327,11.575767,10.600392,9.625018,13.274512,16.924006,20.575312,24.224806,27.8743,29.250338,30.624563,32.000603,33.37483,34.750866,34.212418,33.67578,33.13733,32.600693,32.062244,28.10092,24.137783,20.174648,16.213324,12.250188,12.186734,12.125093,12.06164,11.999999,11.938358,9.686659,7.4367723,5.186886,2.9369993,0.6871128,2.0250793,3.3630457,4.699199,6.037165,7.3751316,6.624565,5.8758116,5.125245,4.3746786,3.6241121,5.524097,7.424082,9.325879,11.225864,13.125849,13.912675,14.699501,15.488139,16.274965,17.06179,15.725637,14.387671,13.049705,11.711739,10.375585,11.650098,12.92461,14.200936,15.475449,16.749962,14.63786,12.525759,10.411844,8.299743,6.187641,7.0125394,7.837437,8.662335,9.487233,10.312131,10.161655,10.012992,9.862516,9.712041,9.563377,9.525306,9.487233,9.449161,9.412902,9.374829,10.3502035,11.325577,12.299138,13.274512,14.249886,12.462305,10.674724,8.887142,7.0995617,5.3119802,8.274362,11.236742,14.200936,17.163317,20.125698,17.27572,14.425743,11.575767,8.725789,5.8758116,6.9744673,8.074935,9.175404,10.275872,11.374527,10.988366,10.600392,10.212419,9.824444,9.438283,13.613536,17.786976,21.962229,26.137482,30.312735,29.812357,29.31198,28.811602,28.313036,27.812658,24.163166,20.511858,16.862366,13.212872,9.563377,12.311829,15.062093,17.812357,20.562622,23.312885,19.112251,14.91343,10.712796,6.5121617,2.3133402,7.037921,11.762501,16.487082,21.213474,25.938055,22.837889,19.737724,16.637558,13.537392,10.437225,10.1870365,9.936848,9.686659,9.438283,9.188094,8.725789,8.26167,7.799365,7.3370595,6.874754,9.088382,11.300196,13.512011,15.725637,17.937452,28.42544,38.911617,49.399605,59.887592,70.37558,56.93609,43.500225,30.062546,16.624866,3.1871881,3.3122826,3.437377,3.5624714,3.6875658,3.8126602,4.1498713,4.4870825,4.8242936,5.163317,5.5005283,14.826408,24.150475,33.47454,42.80042,52.12449,43.349747,34.57501,25.80027,17.025532,8.2507925,10.763558,13.274512,15.787278,18.300045,20.81281,17.687263,14.561715,11.437981,8.312433,5.186886,6.0752378,6.9617763,7.850128,8.736667,9.625018,12.699803,15.774588,18.849373,21.924156,25.000753,23.325577,21.650398,19.975222,18.300045,16.624866,20.999546,25.374224,29.750715,34.125393,38.500072,35.49962,32.50098,29.500526,26.500074,23.49962,22.138086,20.774738,19.413204,18.049856,16.68832,17.60024,18.512161,19.425894,20.337814,21.249735,20.27436,19.3008,18.325426,17.350052,16.374678,14.712192,13.049705,11.3872175,9.724731,8.062244,10.225109,12.387974,14.5508375,16.71189,18.874754,21.262424,23.650097,26.03777,28.42544,30.813112,31.211964,31.612629,32.013294,32.412144,32.81281,34.06194,35.312885,36.562016,37.81296,39.06209,40.037464,41.01284,41.988213,42.961773,43.93715,43.199272,42.46321,41.725334,40.987457,40.24958,42.374374,44.49917,46.62577,48.750565,50.875355,51.488136,52.099106,52.711887,53.32467,53.93745,52.53784,51.138237,49.736816,48.337208,46.937603,45.775494,44.613384,43.449463,42.287354,41.125244,40.024776,38.924305,37.825653,36.72518,35.624714,33.037617,30.45052,27.861609,25.274511,22.687414,21.599636,20.511858,19.424082,18.338116,17.25034,18.261972,19.275417,20.287052,21.300497,22.31213,26.262575,30.213022,34.163467,38.1121,42.062546,43.911766,45.762802,47.612022,49.46306,51.31228,46.5877,41.863117,37.136726,32.412144,27.687565,26.287958,24.88835,23.48693,22.087322,20.687716,22.85058,25.011631,27.174496,29.33736,31.500225,31.500225,31.500225,31.500225,31.500225,31.500225,27.373922,23.249432,19.124943,15.000452,10.874149,10.625773,10.375585,10.125396,9.875207,9.625018,9.875207,10.125396,10.375585,10.625773,10.874149,12.400664,13.925365,15.4500675,16.97477,18.49947,18.999847,19.500225,20.000603,20.499168,20.999546,19.449463,17.89938,16.349297,14.799213,13.24913,11.137029,9.024928,6.9128265,4.800725,2.6868105,2.1991236,1.7132497,1.2255627,0.73787576,0.25018883,2.8372865,5.424384,8.013294,10.600392,13.1874895,12.137785,11.088079,10.038374,8.9868555,7.93715,6.450521,4.9620786,3.4754493,1.987007,0.50037766,1.0243238,1.550083,2.0758421,2.5997884,3.1255474,2.525457,1.9253663,1.3252757,0.72518504,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.15047589,0.2991388,0.44961473,0.6000906,0.7505665,0.7868258,0.824898,0.8629702,0.89922947,0.93730164,1.0750868,1.2128719,1.3506571,1.4866294,1.6244144,1.5247015,1.4249886,1.3252757,1.2255627,1.1258497,0.9880646,0.85027945,0.7124943,0.5747091,0.43692398,0.40066472,0.36259252,0.3245203,0.28826106,0.25018883,0.25018883,0.25018883,0.25018883,0.25018883,0.25018883,0.21211663,0.17585737,0.13778515,0.099712946,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.099712946,0.099712946,0.099712946,0.099712946,0.099712946,0.10515183,0.11059072,0.11421664,0.11965553,0.12509441,1.6697385,3.2143826,4.76084,6.305484,7.850128,6.9508986,6.049856,5.1506267,4.249584,3.350355,4.6303062,5.910258,7.1902094,8.470161,9.750113,8.160145,6.5701766,4.9802084,3.39024,1.8002719,2.465629,3.1291735,3.7945306,4.459888,5.125245,4.233268,3.339477,2.4474995,1.5555218,0.66173136,0.5620184,0.46230546,0.36259252,0.26287958,0.16316663,0.13959812,0.11784257,0.09427405,0.072518505,0.05076295,0.14322405,0.23568514,0.32814622,0.42060733,0.51306844,0.44780177,0.3825351,0.31726846,0.2520018,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.7904517,1.5790904,2.3695421,3.159994,3.9504454,3.7002566,3.4500678,3.199879,2.94969,2.6995013,2.1900587,1.6806163,1.1693609,0.65991837,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.034446288,0.07070554,0.10515183,0.13959812,0.17585737,0.18673515,0.19942589,0.21211663,0.22480737,0.2374981,0.32814622,0.4169814,0.5076295,0.5982776,0.6871128,0.64541465,0.60190356,0.56020546,0.5166943,0.4749962,0.5728962,0.67079616,0.7668832,0.86478317,0.96268314,1.5899682,2.2172532,2.8445382,3.4718235,4.100921,3.9830787,3.8652363,3.7473936,3.6295512,3.5117085,4.327542,5.143375,5.957395,6.773228,7.5872483,7.1466985,6.7079616,6.2674117,5.826862,5.388125,5.139749,4.893186,4.64481,4.3982472,4.1498713,4.1825047,4.215138,4.2477713,4.2804046,4.313038,5.7597823,7.208339,8.655084,10.101828,11.5503845,14.485571,17.420757,20.355944,23.289318,26.224504,23.273,20.319685,17.368181,14.4148655,11.463363,12.772322,14.083094,15.392053,16.702824,18.011784,22.970236,27.926876,32.885326,37.84197,42.80042,37.15667,31.514729,25.87279,20.229036,14.587097,13.918114,13.247317,12.578335,11.907538,11.236742,14.440247,17.64194,20.845444,24.047136,27.25064,28.151684,29.054539,29.957394,30.860249,31.763105,30.999847,30.23659,29.475145,28.71189,27.950443,25.000753,22.049252,19.099562,16.14987,13.200181,13.055143,12.910107,12.76507,12.620032,12.474996,10.364707,8.254418,6.14413,4.0356545,1.9253663,2.9841363,4.0447197,5.105303,6.165886,7.224656,7.0451727,6.8656893,6.684393,6.5049095,6.3254266,7.3841968,8.444779,9.5053625,10.564133,11.624716,12.114216,12.605529,13.095029,13.584529,14.074029,13.149418,12.224807,11.300196,10.375585,9.449161,10.56232,11.675479,12.786825,13.899984,15.013144,13.589968,12.166792,10.745429,9.322253,7.900891,8.350506,8.80012,9.249735,9.699349,10.150778,10.022058,9.89515,9.768243,9.639522,9.512614,9.449161,9.38752,9.325879,9.262425,9.200785,10.127209,11.055446,11.98187,12.910107,13.838344,12.299138,10.761745,9.224354,7.686961,6.149569,8.740293,11.329204,13.919927,16.51065,19.099562,16.80435,14.510953,12.215742,9.920531,7.6253204,8.007855,8.39039,8.772926,9.155461,9.537996,9.501737,9.467291,9.432844,9.396585,9.362139,13.082338,16.802538,20.522736,24.242935,27.963135,27.92325,27.883364,27.841667,27.80178,27.761896,24.752378,21.74286,18.733343,15.722012,12.712494,15.464571,18.216648,20.97054,23.722616,26.474693,23.011934,19.55099,16.08823,12.625471,9.162713,12.360779,15.557032,18.755098,21.953163,25.149418,22.687414,20.22541,17.761595,15.299591,12.837588,12.348088,11.856775,11.367275,10.877775,10.388275,9.414715,8.442966,7.4694057,6.497658,5.524097,7.402326,9.280556,11.156972,13.035201,14.911617,25.773077,36.63272,47.492367,58.352013,69.21166,60.310013,51.408367,42.50491,33.60326,24.699802,20.934278,17.170568,13.4050455,9.639522,5.8758116,5.7017674,5.529536,5.3573046,5.185073,5.0128417,12.7233715,20.432089,28.142618,35.85315,43.561867,36.49131,29.42257,22.352016,15.281462,8.212721,9.935035,11.65735,13.379663,15.101978,16.824293,14.394923,11.965553,9.53437,7.1050005,4.6756306,5.469708,6.265599,7.059676,7.855567,8.649645,11.18054,13.709623,16.240519,18.769602,21.300497,19.864632,18.430578,16.99471,15.5606575,14.124791,17.792416,21.460037,25.12766,28.795284,32.46291,30.051668,27.64224,25.232813,22.821573,20.412146,19.250036,18.087927,16.924006,15.761897,14.599788,15.314095,16.030214,16.744522,17.460642,18.17495,17.379059,16.584982,15.789091,14.995013,14.199123,12.859344,11.519565,10.179785,8.840006,7.500226,9.788185,12.07433,14.362289,16.650248,18.938208,21.367577,23.796947,26.22813,28.6575,31.08687,31.509289,31.93171,32.35413,32.778362,33.200783,35.287502,37.37422,39.462757,41.549477,43.63801,44.74573,45.85345,46.95936,48.067078,49.174797,48.25925,47.345516,46.429974,45.514427,44.600693,46.199726,47.80057,49.399605,51.00045,52.599483,52.90225,53.205013,53.50778,53.810543,54.113308,52.11542,50.11754,48.11965,46.12177,44.125698,42.840305,41.554916,40.269524,38.984135,37.700558,36.596462,35.494183,34.3919,33.28962,32.187336,30.091553,27.997581,25.901796,23.807825,21.71204,20.629702,19.547363,18.465023,17.382685,16.300346,17.224958,18.149569,19.074179,20.000603,20.925215,23.898472,26.869919,29.843178,32.81462,35.78788,38.06496,40.342045,42.619125,44.898018,47.1751,44.792866,42.410633,40.02659,37.644356,35.262123,34.022057,32.78199,31.541924,30.301857,29.06179,30.24203,31.422268,32.602505,33.782745,34.962982,34.516994,34.07282,33.62683,33.182655,32.736664,28.586794,24.436922,20.287052,16.13718,11.9873085,11.584831,11.182353,10.779876,10.377398,9.97492,10.061942,10.150778,10.2378,10.324821,10.411844,12.295512,14.177367,16.059223,17.94289,19.824745,20.83094,21.835321,22.839703,23.845898,24.850279,22.390087,19.929897,17.469707,15.009518,12.549327,10.765372,8.979604,7.1956487,5.40988,3.625925,2.9406252,2.2553256,1.5700256,0.88472575,0.19942589,2.2734551,4.345671,6.4178877,8.490104,10.56232,10.448103,10.332074,10.217857,10.101828,9.987611,8.910711,7.8319983,6.755099,5.678199,4.599486,4.459888,4.3202896,4.1806917,4.0392804,3.8996825,3.2053177,2.5091403,1.8147756,1.1204109,0.42423326,0.35534066,0.28463513,0.21574254,0.14503701,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.11965553,0.23931105,0.36077955,0.48043507,0.6000906,0.629098,0.65991837,0.69073874,0.7197462,0.7505665,0.85934424,0.969935,1.0805258,1.1893034,1.2998942,1.2418793,1.1856775,1.1276628,1.0696479,1.0116332,0.8883517,0.76325727,0.63816285,0.51306844,0.387974,0.4224203,0.45686656,0.49312583,0.5275721,0.5620184,0.5076295,0.45324063,0.39703882,0.34264994,0.28826106,0.24474995,0.2030518,0.15954071,0.11784257,0.07433146,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.07433146,0.07433146,0.07433146,0.07433146,0.07433146,0.08520924,0.09427405,0.10515183,0.11421664,0.12509441,1.4902552,2.855416,4.220577,5.5857377,6.9508986,6.0752378,5.199577,4.325729,3.4500678,2.5744069,3.5225863,4.4707656,5.4171324,6.3653116,7.311678,6.4577727,5.6020546,4.748149,3.8924308,3.0367124,3.8670492,4.6973863,5.527723,6.35806,7.1883965,5.9519563,4.7173285,3.482701,2.2480736,1.0116332,0.85027945,0.6871128,0.52575916,0.36259252,0.19942589,0.1794833,0.15954071,0.13959812,0.11965553,0.099712946,0.17223145,0.24474995,0.31726846,0.38978696,0.46230546,0.44417584,0.42785916,0.40972954,0.39159992,0.37528324,0.2991388,0.22480737,0.15047589,0.07433146,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.09064813,0.06707962,0.045324065,0.02175555,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.59283876,1.1856775,1.7767034,2.3695421,2.962381,2.7756457,2.5870976,2.4003625,2.2118144,2.0250793,1.6425442,1.260009,0.8774739,0.4949388,0.11240368,0.09064813,0.06707962,0.045324065,0.02175555,0.0,0.07070554,0.13959812,0.21030366,0.27919623,0.34990177,0.37528324,0.40066472,0.42423326,0.44961473,0.4749962,0.59283876,0.7106813,0.82671094,0.9445535,1.062396,0.93911463,0.81764615,0.69436467,0.5728962,0.44961473,0.67079616,0.8901646,1.1095331,1.3307146,1.550083,2.2172532,2.8844235,3.5534067,4.220577,4.8877473,4.764466,4.6429973,4.519716,4.3982472,4.274966,4.954827,5.634688,6.3145485,6.9944096,7.6742706,7.208339,6.740595,6.2728505,5.805106,5.337362,5.480586,5.621997,5.765221,5.906632,6.049856,6.0407915,6.0299134,6.0208488,6.009971,6.000906,7.507478,9.015862,10.522435,12.03082,13.537392,16.795286,20.053179,23.30926,26.567154,29.825047,26.481945,23.140654,19.797552,16.454449,13.113158,14.144734,15.1781225,16.209698,17.243088,18.274662,22.065567,25.85466,29.645565,33.434654,37.22556,32.71491,28.204258,23.695421,19.18477,14.674119,14.309713,13.945308,13.580903,13.2146845,12.850279,15.604169,18.359873,21.115576,23.869465,26.625168,27.05484,27.484512,27.914185,28.34567,28.775343,27.787277,26.799213,25.812962,24.824896,23.836832,21.900587,19.96253,18.024473,16.08823,14.150173,13.92174,13.695119,13.466686,13.240066,13.011633,11.042755,9.072064,7.1031876,5.132497,3.1618068,3.9450066,4.7282066,5.5095935,6.2927933,7.07418,7.46578,7.855567,8.245354,8.63514,9.024928,9.244296,9.465478,9.684846,9.904215,10.125396,10.31757,10.509744,10.701918,10.894093,11.088079,10.57501,10.061942,9.550687,9.037619,8.52455,9.474543,10.424535,11.374527,12.32452,13.274512,12.542075,11.809638,11.077202,10.344765,9.612328,9.686659,9.762803,9.837135,9.91328,9.987611,9.882459,9.7773075,9.672155,9.567003,9.461852,9.374829,9.287807,9.200785,9.11195,9.024928,9.904215,10.785315,11.664601,12.545701,13.424988,12.137785,10.850581,9.561564,8.274362,6.987158,9.2044115,11.421664,13.640731,15.857984,18.075237,16.334793,14.594349,12.855718,11.115273,9.374829,9.039432,8.705847,8.370448,8.03505,7.699652,8.01692,8.334189,8.653271,8.970539,9.287807,12.552953,15.818098,19.083244,22.34839,25.611723,26.03233,26.452936,26.87173,27.29234,27.712946,25.34159,22.97205,20.602507,18.232965,15.863422,18.617313,21.373016,24.126905,26.882608,29.638311,26.911617,24.186733,21.461851,18.736969,16.012085,17.681824,19.353376,21.023113,22.692852,24.36259,22.536938,20.713097,18.887444,17.06179,15.23795,14.507326,13.776703,13.047892,12.317267,11.586644,10.1054535,8.62245,7.1394467,5.658256,4.175253,5.718084,7.2591023,8.801933,10.344765,11.887595,23.120712,34.352016,45.585133,56.81825,68.04955,63.682125,59.314697,54.94727,50.57984,46.212418,38.556274,30.901947,23.24762,15.593291,7.93715,7.2554765,6.5719895,5.8903155,5.2068286,4.5251546,10.620335,16.715515,22.810696,28.905876,34.99924,29.634686,24.27013,18.905573,13.539205,8.174648,9.108324,10.040187,10.97205,11.9057255,12.837588,11.102583,9.367578,7.6325727,5.8975673,4.162562,4.8641787,5.567608,6.2692246,6.972654,7.6742706,9.659465,11.644659,13.629852,15.6150465,17.60024,16.405499,15.210756,14.014201,12.819458,11.624716,14.585284,17.544039,20.504606,23.465176,26.425743,24.605528,22.785315,20.9651,19.144884,17.32467,16.361988,15.399304,14.436621,13.475751,12.513068,13.029762,13.548269,14.064963,14.581658,15.100165,14.485571,13.8691635,13.254569,12.639976,12.025381,11.008308,9.989424,8.972352,7.95528,6.9382076,9.349448,11.762501,14.175554,16.586794,18.999847,21.472729,23.94561,26.416677,28.889559,31.36244,31.808428,32.252605,32.69678,33.14277,33.586945,36.513065,39.437374,42.363495,45.287804,48.212112,49.45218,50.692245,51.932312,53.17238,54.412445,53.31923,52.227825,51.13461,50.043205,48.94999,50.025078,51.100163,52.17525,53.250336,54.325424,54.318172,54.30911,54.301857,54.294605,54.28735,51.693,49.09684,46.50249,43.908142,41.311977,39.90512,38.49826,37.08959,35.682728,34.27587,33.169964,32.06587,30.959963,29.854055,28.74996,27.147303,25.544643,23.941984,22.339325,20.736666,19.659767,18.582867,17.504154,16.427254,15.350354,16.187943,17.025532,17.863121,18.700708,19.538298,21.532557,23.526815,25.522888,27.517145,29.513218,32.21816,34.9231,37.628036,40.332977,43.037918,42.998035,42.95815,42.918262,42.87838,42.83668,41.75797,40.67744,39.596916,38.518204,37.437675,37.635292,37.832905,38.030518,38.22813,38.425743,37.535576,36.645412,35.75525,34.86508,33.97492,29.799665,25.624413,21.44916,17.27572,13.100468,12.545701,11.989121,11.434355,10.879588,10.324821,10.25049,10.174346,10.100015,10.025683,9.949538,12.19036,14.429369,16.67019,18.9092,21.15002,22.66022,24.170418,25.680614,27.190813,28.699198,25.330713,21.960415,18.590118,15.219821,11.849524,10.391902,8.934279,7.476658,6.0208488,4.5632267,3.680314,2.7974012,1.9144884,1.0333886,0.15047589,1.7078108,3.2651455,4.8224807,6.379815,7.93715,8.758422,9.577881,10.397341,11.2168,12.038072,11.369088,10.701918,10.034748,9.367578,8.700407,7.895452,7.0904965,6.285541,5.480586,4.6756306,3.8851788,3.094727,2.3042755,1.5156367,0.72518504,0.6091554,0.4949388,0.38072214,0.26469254,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.09064813,0.1794833,0.27013144,0.36077955,0.44961473,0.47318324,0.4949388,0.5166943,0.5402629,0.5620184,0.64541465,0.726998,0.8103943,0.8919776,0.97537386,0.96087015,0.9445535,0.9300498,0.9155461,0.89922947,0.7868258,0.6744221,0.5620184,0.44961473,0.33721104,0.44417584,0.5529536,0.65991837,0.7668832,0.87566096,0.7650702,0.6544795,0.54570174,0.43511102,0.3245203,0.27738327,0.23024625,0.18310922,0.13415924,0.0870222,0.07433146,0.06164073,0.05076295,0.038072214,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.065266654,0.07977036,0.09427405,0.11059072,0.12509441,1.310772,2.4946365,3.680314,4.8641787,6.049856,5.199577,4.349297,3.5008307,2.6505513,1.8002719,2.4148662,3.0294604,3.6458678,4.2604623,4.8750563,4.7554007,4.6357455,4.514277,4.3946214,4.274966,5.2702823,6.265599,7.2609153,8.254418,9.249735,7.6724577,6.09518,4.517903,2.9406252,1.3633479,1.1367276,0.9119202,0.6871128,0.46230546,0.2374981,0.21936847,0.2030518,0.18492219,0.16679256,0.15047589,0.2030518,0.25562772,0.30820364,0.36077955,0.41335547,0.44236287,0.47318324,0.50219065,0.533011,0.5620184,0.44961473,0.33721104,0.22480737,0.11240368,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.39522585,0.7904517,1.1856775,1.5809034,1.9743162,1.8492218,1.7241274,1.6008459,1.4757515,1.3506571,1.0950294,0.83940166,0.5855869,0.32995918,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.10515183,0.21030366,0.3154555,0.42060733,0.52575916,0.5620184,0.6000906,0.63816285,0.6744221,0.7124943,0.8575313,1.0025684,1.1476053,1.2926424,1.4376793,1.2346275,1.0333886,0.83033687,0.62728506,0.42423326,0.7668832,1.1095331,1.452183,1.794833,2.137483,2.8445382,3.5515938,4.2604623,4.9675174,5.674573,5.5476656,5.4207582,5.292038,5.1651306,5.038223,5.582112,6.1278133,6.6717024,7.217404,7.763106,7.268167,6.773228,6.2782893,5.7833505,5.2865987,5.81961,6.352621,6.885632,7.41683,7.949841,7.897265,7.844689,7.7921133,7.7395372,7.686961,9.255174,10.821573,12.389787,13.957999,15.524399,19.105,22.6856,26.264389,29.84499,33.42559,29.692701,25.959812,22.226921,18.494032,14.762955,15.517147,16.273151,17.027344,17.78335,18.537542,21.159086,23.782444,26.4058,29.027344,31.650702,28.273151,24.895601,21.518053,18.140503,14.762955,14.703127,14.643299,14.581658,14.521831,14.462003,16.769903,19.077805,21.385706,23.691795,25.999697,25.957998,25.914488,25.87279,25.829277,25.78758,24.574707,23.361835,22.150776,20.937904,19.725033,18.800423,17.87581,16.949387,16.024776,15.100165,14.790149,14.480132,14.170115,13.860099,13.550082,11.720803,9.88971,8.0604315,6.2293396,4.40006,4.9058766,5.40988,5.915697,6.4197006,6.925517,7.8845744,8.845445,9.804502,10.765372,11.724429,11.104396,10.484363,9.864329,9.244296,8.624263,8.519112,8.415772,8.31062,8.205468,8.100317,8.000604,7.900891,7.799365,7.699652,7.5999393,8.386765,9.175404,9.96223,10.750868,11.537694,11.494183,11.452485,11.410787,11.367275,11.325577,11.024626,10.725487,10.424535,10.125396,9.824444,9.742861,9.659465,9.577881,9.494485,9.412902,9.300498,9.188094,9.07569,8.963287,8.8508835,9.683033,10.515183,11.347333,12.179482,13.011633,11.974618,10.937603,9.900589,8.861761,7.8247466,9.670342,11.514126,13.359721,15.2053175,17.050913,15.865235,14.679558,13.495693,12.310016,11.124338,10.07282,9.019489,7.9679704,6.9146395,5.863121,6.532104,7.2029004,7.8718834,8.54268,9.211663,12.023568,14.831847,17.64194,20.45203,23.262123,24.143223,25.022509,25.901796,26.782896,27.662184,25.932617,24.20305,22.471672,20.742105,19.012539,21.770054,24.52757,27.285088,30.042603,32.800117,30.813112,28.824291,26.837286,24.850279,22.863272,23.004683,23.147905,23.289318,23.43254,23.575766,22.388275,21.200785,20.013294,18.825804,17.638313,16.666565,15.6966305,14.726695,13.75676,12.786825,10.794379,8.801933,6.8094873,4.8170414,2.8245957,4.0320287,5.239462,6.446895,7.654328,8.861761,20.468348,32.07131,43.677895,55.28267,66.88744,67.05424,67.22284,67.38963,67.558235,67.72503,56.178272,44.63514,33.090195,21.545248,10.000301,8.807372,7.614443,6.4233265,5.230397,4.0374675,8.517298,12.9971285,17.47696,21.956789,26.438433,22.778063,19.117691,15.457319,11.7969475,8.138389,8.2798,8.423024,8.564435,8.70766,8.8508835,7.8102427,6.7696023,5.730775,4.690134,3.6494937,4.2604623,4.8696175,5.480586,6.089741,6.70071,8.140202,9.579695,11.019187,12.460492,13.899984,12.944552,11.990934,11.035503,10.080072,9.12464,11.378153,13.629852,15.883366,18.135065,20.386765,19.157576,17.928387,16.697386,15.468197,14.237195,13.475751,12.712494,11.949236,11.187792,10.424535,10.745429,11.06451,11.385405,11.704487,12.025381,11.59027,11.155159,10.720048,10.284937,9.849826,9.155461,8.459284,7.764919,7.0705543,6.3743763,8.912524,11.450671,13.987006,16.525154,19.063301,21.57788,24.09246,26.607038,29.12343,31.63801,32.105755,32.571686,33.03943,33.507175,33.97492,37.736816,41.500526,45.262424,49.024323,52.788033,54.160442,55.532856,56.90527,58.277683,59.650093,58.379208,57.110134,55.83925,54.570175,53.299286,53.850426,54.399754,54.950897,55.500225,56.049553,55.732285,55.415016,55.097744,54.780476,54.463207,51.27058,48.077953,44.885326,41.6927,38.500072,36.969933,35.439793,33.909653,32.379513,30.849371,29.741652,28.635744,27.528025,26.420303,25.312584,24.20305,23.091705,21.982172,20.872639,19.763105,18.68983,17.61837,16.545097,15.471823,14.400362,15.1509285,15.899682,16.650248,17.400814,18.149569,19.168453,20.185526,21.202597,22.21967,23.236742,26.369541,29.50234,32.63514,35.76794,38.900738,41.2032,43.505665,45.808125,48.110588,50.41305,49.492065,48.572895,47.65191,46.732735,45.811752,45.026737,44.241726,43.456715,42.6717,41.88669,40.552345,39.218006,37.881855,36.547512,35.213173,31.012537,26.811903,22.613083,18.412449,14.211814,13.504758,12.797703,12.090648,11.381779,10.674724,10.437225,10.199727,9.96223,9.724731,9.487233,12.085209,14.683184,17.279346,19.877321,22.475298,24.489498,26.505512,28.519714,30.535728,32.54993,28.269526,23.990934,19.71053,15.430124,11.14972,10.020245,8.890768,7.75948,6.630004,5.5005283,4.420003,3.339477,2.2607644,1.1802386,0.099712946,1.1421664,2.18462,3.2270734,4.269527,5.3119802,7.066928,8.821876,10.576823,12.331772,14.0867195,13.829279,13.571837,13.314397,13.056956,12.799516,11.329204,9.860703,8.39039,6.9200783,5.4497657,4.5650396,3.680314,2.7955883,1.9108626,1.0243238,0.86478317,0.70524246,0.54570174,0.38434806,0.22480737,0.1794833,0.13415924,0.09064813,0.045324065,0.0,0.059827764,0.11965553,0.1794833,0.23931105,0.2991388,0.3154555,0.32995918,0.3444629,0.36077955,0.37528324,0.42967212,0.48587397,0.5402629,0.5946517,0.6508536,0.678048,0.70524246,0.7324369,0.75963134,0.7868258,0.6871128,0.5873999,0.48768693,0.387974,0.28826106,0.46774435,0.64722764,0.82671094,1.0080072,1.1874905,1.0225109,0.8575313,0.69255173,0.5275721,0.36259252,0.3100166,0.2574407,0.20486477,0.15228885,0.099712946,0.0870222,0.07433146,0.06164073,0.05076295,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.045324065,0.065266654,0.08520924,0.10515183,0.12509441,1.1294757,2.13567,3.1400511,4.1444325,5.1506267,4.325729,3.5008307,2.6741197,1.8492218,1.0243238,1.3071461,1.5899682,1.8727903,2.1556125,2.4366217,3.053029,3.6676233,4.2822175,4.896812,5.5132194,6.6717024,7.8319983,8.992294,10.152591,11.312886,9.39296,7.473032,5.5531044,3.633177,1.7132497,1.4249886,1.1367276,0.85027945,0.5620184,0.2755703,0.25925365,0.24474995,0.23024625,0.21574254,0.19942589,0.23205921,0.26469254,0.29732585,0.32995918,0.36259252,0.4405499,0.5166943,0.5946517,0.6726091,0.7505665,0.6000906,0.44961473,0.2991388,0.15047589,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.19761293,0.39522585,0.59283876,0.7904517,0.9880646,0.9246109,0.8629702,0.7995165,0.73787576,0.6744221,0.5475147,0.42060733,0.291887,0.16497959,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.13959812,0.27919623,0.42060733,0.56020546,0.69980353,0.7505665,0.7995165,0.85027945,0.89922947,0.9499924,1.1222239,1.2944553,1.4666867,1.6407311,1.8129625,1.5301404,1.2473183,0.9644961,0.68167394,0.40066472,0.86478317,1.3307146,1.794833,2.2607644,2.7248828,3.4718235,4.220577,4.9675174,5.714458,6.4632115,6.3308654,6.1967063,6.0643597,5.9320135,5.7996674,6.209397,6.6191263,7.0306687,7.440398,7.850128,7.327995,6.8058615,6.281915,5.7597823,5.237649,6.1604466,7.083245,8.00423,8.927028,9.849826,9.755551,9.659465,9.56519,9.470917,9.374829,11.00287,12.629097,14.257137,15.885179,17.513218,21.414715,25.318022,29.219519,33.122826,37.024323,32.903458,28.78078,24.658104,20.535427,16.41275,16.889559,17.368181,17.84499,18.3218,18.800423,20.254417,21.710226,23.164223,24.620031,26.074028,23.82958,21.585133,19.340685,17.094423,14.849977,15.094727,15.339477,15.584227,15.83079,16.075539,17.935638,19.795738,21.655838,23.514124,25.374224,24.859343,24.344461,23.82958,23.3147,22.799818,21.362139,19.92446,18.48678,17.0491,15.613234,15.700256,15.787278,15.8743,15.963136,16.050158,15.656745,15.265145,14.871732,14.480132,14.0867195,12.397038,10.707357,9.017676,7.327995,5.638314,5.864934,6.093367,6.319988,6.546608,6.775041,8.3051815,9.835322,11.365462,12.895603,14.425743,12.964496,11.50506,10.045626,8.584378,7.124943,6.722465,6.319988,5.91751,5.5150323,5.1125546,5.424384,5.7380266,6.049856,6.3616858,6.6753283,7.3008003,7.9244595,8.549932,9.175404,9.800876,10.448103,11.095331,11.7425585,12.389787,13.037014,12.362592,11.6881695,11.011934,10.337513,9.663091,9.603263,9.541622,9.481794,9.421967,9.362139,9.224354,9.088382,8.950596,8.812811,8.675026,9.460039,10.245051,11.030065,11.815077,12.60009,11.813264,11.024626,10.2378,9.449161,8.662335,10.13446,11.606586,13.080525,14.55265,16.024776,15.3956785,14.764768,14.13567,13.504758,12.87566,11.104396,9.334945,7.5654926,5.7942286,4.024777,5.047288,6.069799,7.0923095,8.1148205,9.137331,11.49237,13.847408,16.202446,18.557486,20.912523,22.252302,23.592083,24.931862,26.27164,27.613234,26.52183,25.43224,24.34265,23.253057,22.161655,24.922796,27.682125,30.443268,33.2026,35.961926,34.712795,33.46185,32.21272,30.961775,29.712645,28.32754,26.942436,25.557333,24.17223,22.787127,22.237799,21.686659,21.137331,20.588003,20.036863,18.827616,17.61837,16.40731,15.198066,13.987006,11.485118,8.98323,6.4795284,3.97764,1.4757515,2.3477864,3.2198215,4.0918565,4.9657044,5.8377395,17.815983,29.792414,41.770657,53.74709,65.725334,70.428154,75.129166,79.83199,84.53482,89.23765,73.80208,58.368332,42.932766,27.497204,12.06164,10.359268,8.656897,6.9545245,5.2521524,3.5497808,6.414262,9.280556,12.145037,15.009518,17.873999,15.919624,13.965251,12.009064,10.05469,8.100317,7.453089,6.8058615,6.156821,5.5095935,4.8623657,4.517903,4.171627,3.827164,3.482701,3.1382382,3.6549325,4.171627,4.690134,5.2068286,5.7253356,6.6191263,7.51473,8.410334,9.304124,10.199727,9.48542,8.7693,8.054993,7.3406854,6.624565,8.1692095,9.715667,11.26031,12.804955,14.349599,13.709623,13.069647,12.429671,11.789696,11.14972,10.587702,10.025683,9.461852,8.899834,8.337815,8.459284,8.582565,8.705847,8.827314,8.950596,8.694968,8.439341,8.185526,7.9298983,7.6742706,7.3026133,6.929143,6.5574856,6.185828,5.812358,8.4756,11.137029,13.800271,16.4617,19.124943,21.683033,24.23931,26.7974,29.35549,31.911768,32.40308,32.892582,33.38208,33.873394,34.362892,38.96238,43.561867,48.163162,52.76265,57.362137,58.866894,60.371655,61.878227,63.382984,64.88774,63.439186,61.992443,60.5457,59.09714,57.6504,57.675777,57.69935,57.724728,57.75011,57.77549,57.148205,56.52092,55.891823,55.264538,54.637253,50.84816,47.05726,43.268166,39.47726,35.688168,34.034748,32.383137,30.729715,29.078106,27.424685,26.315151,25.205618,24.094273,22.98474,21.875206,21.256987,20.64058,20.022358,19.404139,18.787731,17.719896,16.652061,15.584227,14.518205,13.45037,14.112101,14.775645,15.437376,16.099108,16.762651,16.802538,16.842422,16.882307,16.922194,16.962078,20.522736,24.081581,27.64224,31.2029,34.761745,39.408367,44.053177,48.697987,53.342796,57.98761,57.227978,56.468346,55.7069,54.94727,54.187637,52.420002,50.652363,48.884724,47.117085,45.349445,43.56912,41.7906,40.010273,38.229942,36.44961,32.22541,27.999393,23.77519,19.549175,15.324973,14.465629,13.604471,12.745127,11.885782,11.024626,10.625773,10.225109,9.824444,9.425592,9.024928,11.980057,14.935185,17.890314,20.845444,23.800573,26.320591,28.840609,31.360626,33.880646,36.40066,31.210152,26.019638,20.829126,15.640429,10.449916,9.646774,8.845445,8.042302,7.2391596,6.43783,5.1596913,3.8833659,2.6052272,1.3270886,0.05076295,0.57833505,1.1040943,1.6316663,2.1592383,2.6868105,5.377247,8.067683,10.75812,13.446743,16.13718,16.289469,16.441757,16.59586,16.748148,16.900436,14.764768,12.63091,10.49524,8.3595705,6.2257137,5.2449007,4.265901,3.2850883,2.3042755,1.3252757,1.1204109,0.9155461,0.7106813,0.5058166,0.2991388,0.23931105,0.1794833,0.11965553,0.059827764,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.15772775,0.16497959,0.17223145,0.1794833,0.18673515,0.21574254,0.24293698,0.27013144,0.29732585,0.3245203,0.39522585,0.46411842,0.53482395,0.6055295,0.6744221,0.5873999,0.50037766,0.41335547,0.3245203,0.2374981,0.4894999,0.7433147,0.99531645,1.2473183,1.49932,1.2799516,1.0605831,0.83940166,0.6200332,0.40066472,0.34264994,0.28463513,0.22662032,0.17041849,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.9499924,1.7748904,2.5997884,3.4246864,4.249584,3.4500678,2.6505513,1.8492218,1.0497054,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,1.3506571,2.6995013,4.0501585,5.4008155,6.7496595,8.074935,9.400211,10.725487,12.050762,13.374225,11.111648,8.8508835,6.588306,4.325729,2.0631514,1.7132497,1.3633479,1.0116332,0.66173136,0.31182957,0.2991388,0.28826106,0.2755703,0.26287958,0.25018883,0.26287958,0.2755703,0.28826106,0.2991388,0.31182957,0.43692398,0.5620184,0.6871128,0.8122072,0.93730164,0.7505665,0.5620184,0.37528324,0.18673515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.17585737,0.34990177,0.52575916,0.69980353,0.87566096,0.93730164,1.0007553,1.062396,1.1258497,1.1874905,1.3869164,1.5881553,1.7875811,1.987007,2.1882458,1.8256533,1.4630609,1.1004683,0.73787576,0.37528324,0.96268314,1.550083,2.137483,2.7248828,3.3122826,4.099108,4.8877473,5.674573,6.4632115,7.250037,7.112252,6.9744673,6.836682,6.70071,6.5629244,6.836682,7.112252,7.3878226,7.663393,7.93715,7.3878226,6.836682,6.2873545,5.7380266,5.186886,6.4994707,7.8120556,9.12464,10.437225,11.74981,11.612025,11.47424,11.338268,11.200482,11.062697,12.750566,14.436621,16.124489,17.812357,19.500225,23.724428,27.950443,32.17465,36.40066,40.624866,36.1124,31.599937,27.087475,22.57501,18.062546,18.261972,18.463211,18.662638,18.862062,19.063301,19.34975,19.63801,19.92446,20.212719,20.499168,19.387821,18.274662,17.163317,16.050158,14.936998,15.488139,16.037468,16.586794,17.137936,17.687263,19.099562,20.511858,21.924156,23.338266,24.750565,23.7625,22.774435,21.788185,20.80012,19.812056,18.149569,16.487082,14.824595,13.162108,11.499621,12.60009,13.700559,14.799213,15.899682,17.00015,16.525154,16.050158,15.575162,15.100165,14.625169,13.075087,11.525003,9.97492,8.424837,6.874754,6.825804,6.775041,6.7242785,6.6753283,6.624565,8.725789,10.825199,12.92461,15.025834,17.125244,14.824595,12.525759,10.225109,7.9244595,5.6256227,4.9258194,4.2242026,3.5243993,2.8245957,2.124792,2.8499773,3.5751622,4.3003473,5.0255322,5.750717,6.2130227,6.6753283,7.137634,7.5999393,8.062244,9.400211,10.738177,12.07433,13.412297,14.750263,13.700559,12.650853,11.599335,10.549629,9.499924,9.461852,9.425592,9.38752,9.349448,9.313189,9.1500225,8.9868555,8.825501,8.662335,8.499168,9.237044,9.97492,10.712796,11.450671,12.186734,11.650098,11.111648,10.57501,10.038374,9.499924,10.600392,11.700861,12.799516,13.899984,15.000452,14.924308,14.849977,14.775645,14.699501,14.625169,12.137785,9.6504,7.1630154,4.6756306,2.1882458,3.5624714,4.936697,6.3127356,7.686961,9.063,10.962985,12.862969,14.762955,16.66294,18.562923,20.363195,22.161655,23.961926,25.762197,27.56247,27.112856,26.66324,26.211813,25.762197,25.312584,28.075539,30.836681,33.599636,36.36259,39.125546,38.612476,38.099407,37.588154,37.075085,36.562016,33.6504,30.736967,27.82535,24.911919,22.000301,22.087322,22.174345,22.26318,22.350203,22.437225,20.986855,19.538298,18.087927,16.637558,15.187187,12.174044,9.162713,6.149569,3.1382382,0.12509441,0.66173136,1.2001812,1.7368182,2.275268,2.811905,15.163619,27.511707,39.863422,52.21332,64.563225,73.80027,83.037315,92.27617,101.513214,110.75026,91.42408,72.09971,52.77353,33.44916,14.124791,11.912977,9.699349,7.4875355,5.275721,3.0620937,4.313038,5.562169,6.813113,8.062244,9.313189,9.063,8.812811,8.562622,8.312433,8.062244,6.624565,5.186886,3.7492065,2.3133402,0.87566096,1.2255627,1.5754645,1.9253663,2.275268,2.6251698,3.049403,3.4754493,3.8996825,4.325729,4.749962,5.0998635,5.4497657,5.7996674,6.149569,6.4994707,6.0244746,5.5494785,5.0744824,4.599486,4.12449,4.9620786,5.7996674,6.637256,7.474845,8.312433,8.26167,8.212721,8.161958,8.113008,8.062244,7.699652,7.3370595,6.9744673,6.6118746,6.249282,6.1749506,6.1006193,6.0244746,5.9501433,5.8758116,5.7996674,5.7253356,5.6491914,5.57486,5.5005283,5.4497657,5.4008155,5.3500524,5.2992897,5.2503395,8.036863,10.825199,13.611723,16.400059,19.188396,21.788185,24.387972,26.98776,29.58755,32.187336,32.700405,33.211662,33.72473,34.237797,34.750866,40.187943,45.625015,51.06209,56.50098,61.938053,63.575157,65.212265,66.84937,68.48829,70.12539,68.49917,66.87475,65.250336,63.624107,61.999695,61.499317,61.00075,60.500374,59.999996,59.49962,58.562317,57.625015,56.687714,55.750412,54.81311,50.423927,46.038372,41.64919,37.26182,32.87445,31.09956,29.324669,27.54978,25.774889,23.999998,22.886839,21.775494,20.662334,19.549175,18.43783,18.312735,18.187641,18.062546,17.937452,17.812357,16.749962,15.687565,14.625169,13.562773,12.500377,13.075087,13.649796,14.224504,14.799213,15.375735,14.436621,13.499319,12.562017,11.624716,10.687414,14.675932,18.662638,22.649342,26.63786,30.624563,37.613533,44.600693,51.58785,58.57501,65.562164,64.962074,64.361984,63.761894,63.161804,62.561714,59.811447,57.062996,54.312733,51.56247,48.812206,46.5877,44.363194,42.136875,39.912373,37.687866,33.43647,29.186884,24.9373,20.687716,16.438131,15.4246855,14.413053,13.399607,12.387974,11.374527,10.812509,10.25049,9.686659,9.12464,8.562622,11.874905,15.187187,18.49947,21.811752,25.125849,28.14987,31.175705,34.199726,37.22556,40.24958,34.148964,28.050158,21.949537,15.850732,9.750113,9.275117,8.80012,8.325124,7.850128,7.3751316,5.89938,4.4254417,2.94969,1.4757515,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,3.6875658,7.311678,10.937603,14.561715,18.187641,18.749659,19.311678,19.87551,20.437527,20.999546,18.20033,15.399304,12.60009,9.800876,6.9998484,5.924762,4.8496747,3.774588,2.6995013,1.6244144,1.3742256,1.1258497,0.87566096,0.62547207,0.37528324,0.2991388,0.22480737,0.15047589,0.07433146,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.11240368,0.22480737,0.33721104,0.44961473,0.5620184,0.48768693,0.41335547,0.33721104,0.26287958,0.18673515,0.51306844,0.8375887,1.162109,1.4866294,1.8129625,1.5373923,1.261822,0.9880646,0.7124943,0.43692398,0.37528324,0.31182957,0.25018883,0.18673515,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.07433146,0.099712946,0.12509441,0.15047589,0.17585737,0.8375887,1.49932,2.1628644,2.8245957,3.48814,3.7020695,3.917812,4.1317415,4.347484,4.5632267,3.972201,3.3829882,2.7919624,2.2027495,1.6117238,2.373168,3.1327994,3.8924308,4.652062,5.411693,6.492219,7.572745,8.653271,9.731983,10.812509,9.019489,7.228282,5.4352617,3.6422417,1.8492218,1.5718386,1.2944553,1.017072,0.73968875,0.46230546,0.56020546,0.65810543,0.7541924,0.8520924,0.9499924,0.8103943,0.67079616,0.5293851,0.38978696,0.25018883,0.35171473,0.4550536,0.55839247,0.65991837,0.76325727,0.61278135,0.46230546,0.31182957,0.16316663,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.04169814,0.034446288,0.027194439,0.01994259,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.09427405,0.17767033,0.25925365,0.34264994,0.42423326,0.52213323,0.6200332,0.7179332,0.81583315,0.9119202,0.91917205,0.92823684,0.9354887,0.94274056,0.9499924,1.1095331,1.2708868,1.4304274,1.5899682,1.7495089,1.4630609,1.1747998,0.8883517,0.6000906,0.31182957,0.88472575,1.4576219,2.030518,2.6016014,3.1744974,3.9051213,4.6357455,5.3645563,6.09518,6.825804,6.742408,6.6608243,6.5774283,6.495845,6.412449,6.9418335,7.473032,8.002417,8.531802,9.063,8.303369,7.5419245,6.782293,6.0226617,5.2630305,6.378002,7.4929743,8.607946,9.7229185,10.837891,10.754494,10.672911,10.589515,10.507931,10.424535,11.537694,12.64904,13.762199,14.875358,15.986704,19.387821,22.787127,26.188244,29.58755,32.986855,29.607492,26.22813,22.846954,19.467592,16.08823,16.285843,16.481644,16.679256,16.87687,17.074482,17.529535,17.984589,18.439642,18.894695,19.34975,18.136877,16.92582,15.712947,14.500074,13.287203,13.796645,14.3079,14.817343,15.326786,15.838041,16.998337,18.15682,19.317116,20.477413,21.637709,20.838192,20.036863,19.237347,18.43783,17.638313,16.36924,15.101978,13.834718,12.567456,11.300196,12.059827,12.819458,13.57909,14.340534,15.100165,14.811904,14.525456,14.237195,13.9507475,13.662486,12.3916,11.122525,9.851639,8.582565,7.311678,7.3026133,7.2917356,7.2826705,7.271793,7.262728,8.740293,10.217857,11.695421,13.172986,14.650551,13.466686,12.284635,11.102583,9.920531,8.736667,7.3950744,6.053482,4.710077,3.3666716,2.0250793,2.6306088,3.2343252,3.8398547,4.445384,5.049101,5.4044414,5.7597823,6.115123,6.4704633,6.825804,7.9842873,9.144584,10.304879,11.465176,12.625471,11.744371,10.865085,9.985798,9.104698,8.225411,8.403082,8.580752,8.756609,8.934279,9.11195,9.284182,9.458226,9.630457,9.802689,9.97492,10.342952,10.70917,11.077202,11.445232,11.813264,11.564888,11.318325,11.069949,10.823386,10.57501,11.566701,12.5602045,13.551895,14.545399,15.537089,15.343102,15.147303,14.953316,14.757515,14.561715,12.145037,9.728357,7.309865,4.893186,2.474694,3.8579843,5.239462,6.622752,8.00423,9.38752,10.694666,12.001812,13.310771,14.617917,15.925063,18.372562,20.820063,23.267561,25.715061,28.162561,27.71476,27.266956,26.819155,26.373167,25.925365,27.528025,29.130682,30.733341,32.334187,33.936848,33.13733,32.337814,31.536484,30.736967,29.93745,27.470009,25.002567,22.535126,20.067682,17.60024,17.687263,17.774284,17.863121,17.950142,18.037165,17.029158,16.022963,15.014956,14.006948,13.000754,10.680162,8.3595705,6.0407915,3.720199,1.3996071,3.5044568,5.6093063,7.7159686,9.820818,11.925668,20.905272,29.884874,38.86448,47.845894,56.8255,63.205315,69.58513,75.96494,82.34476,88.72458,73.23825,57.75555,42.269222,26.78471,11.300196,9.56519,7.8301854,6.09518,4.360175,2.6251698,3.589666,4.554162,5.520471,6.484967,7.4494634,7.250037,7.0506115,6.849373,6.6499467,6.450521,5.2992897,4.1498713,3.000453,1.8492218,0.69980353,1.0080072,1.3143979,1.6226015,1.9308052,2.2371957,2.960568,3.682127,4.405499,5.127058,5.8504305,5.7942286,5.7398396,5.6854506,5.6292486,5.57486,5.67276,5.77066,5.866747,5.964647,6.0625467,6.5230393,6.981719,7.4422116,7.902704,8.363196,8.116633,7.8718834,7.6271334,7.382384,7.137634,6.8656893,6.591932,6.319988,6.0480433,5.774286,5.8377395,5.89938,5.962834,6.0244746,6.0879283,6.189454,6.2927933,6.394319,6.497658,6.599184,7.1394467,7.6797094,8.219973,8.760235,9.300498,12.580148,15.859797,19.139446,22.420908,25.700558,26.989574,28.280403,29.56942,30.860249,32.149265,33.110134,34.06919,35.030064,35.990932,36.94999,41.085358,45.220726,49.35428,53.489647,57.625015,58.883213,60.139595,61.39779,62.654175,63.91237,62.452934,60.991688,59.532253,58.07282,56.61157,56.185524,55.757664,55.329803,54.901947,54.474087,53.442513,52.409122,51.37755,50.34416,49.312584,45.344006,41.377247,37.410484,33.441906,29.475145,27.778214,26.079466,24.382534,22.6856,20.986855,20.43934,19.891825,19.34431,18.796797,18.24928,19.500225,20.749357,22.000301,23.249432,24.500376,23.405348,22.310318,21.215288,20.120258,19.025229,19.327993,19.630758,19.933523,20.234476,20.537241,19.657953,18.776854,17.897566,17.01828,16.13718,18.852999,21.567003,24.282822,26.996826,29.712645,36.328144,42.941833,49.55733,56.172832,62.788334,63.297775,63.807217,64.31666,64.82792,65.33736,62.617916,59.89847,57.177216,54.45777,51.738327,49.736816,47.737118,45.73742,43.73772,41.738026,37.94168,34.147152,30.35262,26.558088,22.761745,21.855265,20.94697,20.04049,19.132195,18.225714,17.04185,15.859797,14.677745,13.495693,12.311829,14.752076,17.192324,19.632572,22.072819,24.513067,27.013142,29.513218,32.013294,34.511555,37.01163,32.551743,28.091856,23.631968,19.17208,14.712192,13.082338,11.452485,9.822631,8.192778,6.5629244,5.2557783,3.9468195,2.6396735,1.3325275,0.025381476,0.034446288,0.045324065,0.054388877,0.065266654,0.07433146,3.4174345,6.7605376,10.101828,13.44493,16.788034,17.074482,17.362743,17.64919,17.937452,18.225714,16.842422,15.460945,14.077655,12.694364,11.312886,10.549629,9.788185,9.024928,8.263483,7.500226,6.341743,5.185073,4.028403,2.8699198,1.7132497,1.3778516,1.0424535,0.7070554,0.37165734,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.09064813,0.1794833,0.27013144,0.36077955,0.44961473,0.38978696,0.32995918,0.27013144,0.21030366,0.15047589,0.40972954,0.67079616,0.9300498,1.1893034,1.4503701,1.2328146,1.015259,0.79770356,0.58014804,0.36259252,0.3245203,0.28826106,0.25018883,0.21211663,0.17585737,0.17223145,0.17041849,0.16679256,0.16497959,0.16316663,0.13415924,0.10696479,0.07977036,0.052575916,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.12509441,0.15047589,0.17585737,0.19942589,0.22480737,0.72518504,1.2255627,1.7241274,2.2245052,2.7248828,3.9558845,5.185073,6.414262,7.645263,8.874452,7.744976,6.6155005,5.484212,4.3547363,3.2252605,3.395679,3.5642843,3.7347028,3.9051213,4.07554,4.9095025,5.7452784,6.5792413,7.415017,8.2507925,6.92733,5.6056805,4.2822175,2.960568,1.6371052,1.4322405,1.2273756,1.0225109,0.81764615,0.61278135,0.8194591,1.0279498,1.2346275,1.4431182,1.649796,1.357909,1.064209,0.77232206,0.48043507,0.18673515,0.26831847,0.3480888,0.42785916,0.5076295,0.5873999,0.4749962,0.36259252,0.25018883,0.13778515,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.08520924,0.07070554,0.054388877,0.03988518,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.19036107,0.35534066,0.52032024,0.6852999,0.85027945,0.87022203,0.8901646,0.9101072,0.9300498,0.9499924,0.90285534,0.8557183,0.80676836,0.75963134,0.7124943,0.8321498,0.95180535,1.0732739,1.1929294,1.3125849,1.1004683,0.8883517,0.6744221,0.46230546,0.25018883,0.80676836,1.3651608,1.9217403,2.4801328,3.0367124,3.7093215,4.3819304,5.0545397,5.727149,6.399758,6.3725634,6.345369,6.3181744,6.2891674,6.261973,7.0469856,7.8319983,8.617011,9.402024,10.1870365,9.217102,8.247167,7.2772317,6.3072968,5.337362,6.2547207,7.17208,8.089439,9.006798,9.924157,9.896963,9.869768,9.842574,9.815379,9.788185,10.324821,10.863272,11.399909,11.938358,12.474996,15.049402,17.625622,20.20003,22.774435,25.350657,23.102583,20.85451,18.608248,16.360174,14.112101,14.3079,14.501887,14.697688,14.891675,15.087475,15.709321,16.33298,16.954826,17.576672,18.20033,16.887747,15.575162,14.262577,12.949992,11.637406,12.106964,12.578335,13.047892,13.517449,13.987006,14.895301,15.801782,16.710075,17.61837,18.52485,17.912071,17.29929,16.68832,16.075539,15.462758,14.590723,13.716875,12.84484,11.972805,11.10077,11.519565,11.940171,12.360779,12.779573,13.200181,13.100468,13.000754,12.899229,12.799516,12.699803,11.709926,10.720048,9.73017,8.740293,7.750415,7.7794223,7.8102427,7.83925,7.8700705,7.900891,8.754796,9.610515,10.46442,11.320138,12.175857,12.11059,12.045323,11.980057,11.91479,11.849524,9.864329,7.8809485,5.8957543,3.9105604,1.9253663,2.4094272,2.8953013,3.3793623,3.8652363,4.349297,4.597673,4.844236,5.092612,5.3391747,5.5875506,6.5701766,7.552802,8.535428,9.518054,10.500679,9.789998,9.079316,8.370448,7.6597667,6.9490857,7.3424983,7.7340984,8.127511,8.519112,8.912524,9.420154,9.927783,10.435412,10.943042,11.450671,11.447045,11.445232,11.4416065,11.439794,11.437981,11.479679,11.5231905,11.564888,11.608399,11.650098,12.534823,13.419549,14.304275,15.190813,16.075539,15.760084,15.444629,15.129172,14.81553,14.500074,12.152288,9.804502,7.456715,5.1107416,2.762955,4.1516843,5.542227,6.932769,8.323311,9.712041,10.428161,11.142468,11.856775,12.572895,13.287203,16.38193,19.476658,22.573196,25.667925,28.762651,28.316662,27.872486,27.42831,26.982323,26.538147,26.980509,27.422873,27.865234,28.307598,28.74996,27.662184,26.574406,25.486628,24.400663,23.312885,21.28962,19.268166,17.2449,15.221634,13.200181,13.287203,13.374225,13.46306,13.550082,13.637105,13.073273,12.507628,11.941984,11.378153,10.812509,9.184468,7.558241,5.9302006,4.3021603,2.6741197,6.347182,10.020245,13.693306,17.364555,21.037619,26.648737,32.25804,37.867348,43.476654,49.087776,52.610363,56.132946,59.655533,63.17812,66.70071,55.054234,43.409576,31.764917,20.120258,8.4756,7.217404,5.959208,4.702825,3.444629,2.1882458,2.8681068,3.5479677,4.227829,4.9076896,5.5875506,5.4370747,5.2865987,5.137936,4.98746,4.836984,3.975827,3.1128569,2.2498865,1.3869164,0.52575916,0.7904517,1.0551442,1.3198367,1.5845293,1.8492218,2.8699198,3.8906176,4.9095025,5.9302006,6.9508986,6.490406,6.0299134,5.569421,5.1107416,4.650249,5.319232,5.9900284,6.6608243,7.3298078,8.000604,8.082188,8.165584,8.247167,8.330563,8.412147,7.9715962,7.5328593,7.0923095,6.6517596,6.2130227,6.0299134,5.846804,5.6655083,5.482399,5.2992897,5.5005283,5.6999545,5.89938,6.1006193,6.300045,6.5792413,6.8602505,7.1394467,7.420456,7.699652,8.830941,9.960417,11.089892,12.219368,13.3506565,17.123432,20.894394,24.66717,28.439943,32.21272,32.192776,32.172832,32.152893,32.13295,32.113007,33.519867,34.926723,36.335396,37.742256,39.149113,41.982773,44.81462,47.64828,50.48013,53.311977,54.189453,55.066925,55.9444,56.821873,57.69935,56.404892,55.110435,53.814167,52.519714,51.225258,50.86992,50.514576,50.159237,49.80571,49.450367,48.322704,47.19504,46.06738,44.939716,43.812054,40.264088,36.71793,33.169964,29.621996,26.07584,24.455051,22.834263,21.215288,19.5945,17.975525,17.99184,18.00997,18.0281,18.044416,18.062546,20.687716,23.312885,25.938055,28.563225,31.188395,30.060732,28.93307,27.805407,26.677744,25.550081,25.580902,25.60991,25.64073,25.669737,25.700558,24.877472,24.054388,23.233116,22.41003,21.586945,23.030064,24.473183,25.914488,27.357605,28.800724,35.042755,41.284782,47.526814,53.770657,60.012688,61.633476,63.252453,64.87324,66.49222,68.11301,65.42257,62.732132,60.041695,57.353073,54.662636,52.887745,51.112854,49.337963,47.563072,45.78818,42.44689,39.107414,35.76794,32.426647,29.087172,28.285843,27.4827,26.679558,25.878227,25.075085,23.273,21.470917,19.667019,17.864933,16.062849,17.629248,19.19746,20.765673,22.332073,23.900286,25.874601,27.85073,29.825047,31.799364,33.775494,30.954523,28.135366,25.314396,22.49524,19.67427,16.889559,14.104849,11.320138,8.535428,5.750717,4.610364,3.4700103,2.3296568,1.1893034,0.05076295,0.058014803,0.065266654,0.072518505,0.07977036,0.0870222,3.147303,6.207584,9.267865,12.328146,15.386614,15.399304,15.411995,15.4246855,15.437376,15.4500675,15.484513,15.520773,15.555219,15.589665,15.625924,15.174497,14.724882,14.275268,13.825653,13.374225,11.30926,9.244296,7.179332,5.1143675,3.049403,2.4547513,1.8600996,1.2654479,0.67079616,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06707962,0.13415924,0.2030518,0.27013144,0.33721104,0.291887,0.24837588,0.2030518,0.15772775,0.11240368,0.30820364,0.50219065,0.6979906,0.8919776,1.0877775,0.92823684,0.7668832,0.6073425,0.44780177,0.28826106,0.2755703,0.26287958,0.25018883,0.2374981,0.22480737,0.23205921,0.23931105,0.24837588,0.25562772,0.26287958,0.21936847,0.17767033,0.13415924,0.092461094,0.05076295,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.17585737,0.19942589,0.22480737,0.25018883,0.2755703,0.61278135,0.9499924,1.2872034,1.6244144,1.9616255,4.207886,6.452334,8.696781,10.943042,13.1874895,11.517752,9.848013,8.178274,6.506723,4.836984,4.41819,3.9975824,3.576975,3.1581807,2.7375734,3.3267863,3.917812,4.507025,5.0980506,5.6872635,4.835171,3.9830787,3.1291735,2.277081,1.4249886,1.2926424,1.1602961,1.0279498,0.89560354,0.76325727,1.0805258,1.3977941,1.7150626,2.032331,2.3495996,1.9054236,1.4594349,1.015259,0.56927025,0.12509441,0.18310922,0.23931105,0.29732585,0.35534066,0.41335547,0.33721104,0.26287958,0.18673515,0.11240368,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.12690738,0.10515183,0.08339628,0.059827764,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.28463513,0.533011,0.7795739,1.0279498,1.2745126,1.2183108,1.1602961,1.1022812,1.0442665,0.9880646,0.88472575,0.78319985,0.67986095,0.57833505,0.4749962,0.55476654,0.6345369,0.71430725,0.79589057,0.87566096,0.73787576,0.6000906,0.46230546,0.3245203,0.18673515,0.7306239,1.2726997,1.8147756,2.3568513,2.9007401,3.5153344,4.1299286,4.744523,5.3591175,5.975525,6.002719,6.0299134,6.057108,6.0843024,6.11331,7.1521373,8.192778,9.233418,10.272246,11.312886,10.1326475,8.952409,7.7721705,6.591932,5.411693,6.1332526,6.8529987,7.572745,8.292491,9.012237,9.039432,9.066626,9.0956335,9.122828,9.1500225,9.11195,9.07569,9.037619,8.999546,8.963287,10.712796,12.462305,14.211814,15.963136,17.712645,16.597672,15.4827,14.367728,13.252756,12.137785,12.329959,12.522133,12.714307,12.908294,13.100468,13.889107,14.679558,15.47001,16.260462,17.050913,15.636803,14.224504,12.812206,11.399909,9.987611,10.417283,10.846955,11.276628,11.708113,12.137785,12.792264,13.446743,14.103036,14.757515,15.411995,14.9877615,14.561715,14.137483,13.713249,13.287203,12.810393,12.331772,11.854962,11.378153,10.899531,10.979301,11.060884,11.1406555,11.220426,11.300196,11.3872175,11.47424,11.563075,11.650098,11.73712,11.028252,10.31757,9.606889,8.898021,8.187339,8.258044,8.326937,8.397643,8.4683485,8.537241,8.7693,9.003172,9.235231,9.467291,9.699349,10.752681,11.804199,12.857531,13.910862,14.96238,12.335398,9.708415,7.079619,4.4526362,1.8256533,2.1900587,2.5544643,2.9206827,3.2850883,3.6494937,3.7909048,3.930503,4.070101,4.209699,4.349297,5.1542525,5.959208,6.7641635,7.570932,8.375887,7.835624,7.2953615,6.755099,6.2148356,5.674573,6.281915,6.889258,7.498413,8.105756,8.713099,9.554313,10.397341,11.240368,12.083396,12.92461,12.552953,12.179482,11.807825,11.434355,11.062697,11.39447,11.728055,12.059827,12.3916,12.725184,13.502945,14.280706,15.056654,15.834415,16.612177,16.177065,15.741954,15.306843,14.871732,14.436621,12.15954,9.882459,7.605378,5.328297,3.049403,4.4471974,5.844991,7.2427855,8.640579,10.038374,10.1598425,10.283124,10.4045925,10.527874,10.649343,14.39311,18.135065,21.87702,25.620787,29.362741,28.92038,28.478016,28.035654,27.59329,27.149115,26.432995,25.715061,24.997128,24.279196,23.563074,22.187037,20.81281,19.436771,18.062546,16.68832,15.10923,13.531953,11.954676,10.377398,8.80012,8.887142,8.974165,9.063,9.1500225,9.237044,9.115576,8.992294,8.870826,8.747544,8.624263,7.690587,6.755099,5.81961,4.8841214,3.9504454,9.189907,14.429369,19.670645,24.910107,30.149569,32.39039,34.6294,36.87022,39.10923,41.35005,42.015408,42.680763,43.34431,44.009666,44.675022,36.87022,29.065416,21.260612,13.455809,5.6491914,4.8696175,4.0900435,3.3104696,2.5308957,1.7495089,2.1447346,2.5399606,2.9351864,3.3304121,3.7256382,3.6241121,3.5243993,3.4246864,3.3249733,3.2252605,2.6505513,2.0758421,1.49932,0.9246109,0.34990177,0.5728962,0.79589057,1.017072,1.2400664,1.4630609,2.7792716,4.0972953,5.4153194,6.733343,8.049554,7.1847706,6.319988,5.4552045,4.590421,3.7256382,4.9675174,6.209397,7.453089,8.694968,9.936848,9.643148,9.347635,9.052122,8.756609,8.46291,7.8265595,7.192023,6.5574856,5.922949,5.2884116,5.1941376,5.101677,5.009216,4.9167547,4.8242936,5.163317,5.5005283,5.8377395,6.1749506,6.5121617,6.970841,7.4277077,7.8845744,8.343254,8.80012,10.520622,12.23931,13.959812,15.680313,17.400814,21.664904,25.928991,30.194891,34.460793,38.72488,37.394165,36.065266,34.73455,33.405647,32.074936,33.929596,35.784256,37.640728,39.495388,41.35005,42.88019,44.41033,45.94047,47.47061,49.00075,49.497505,49.994255,50.49282,50.989574,51.488136,50.35685,49.22737,48.097897,46.968422,45.83713,45.55431,45.2733,44.99048,44.707657,44.424835,43.2029,41.98096,40.757214,39.535275,38.31334,35.184166,32.056805,28.929443,25.802084,22.674723,21.131891,19.590874,18.048042,16.50521,14.96238,15.544341,16.128115,16.710075,17.292038,17.87581,21.875206,25.874601,29.87581,33.875206,37.8746,36.714306,35.55582,34.395527,33.23523,32.074936,31.831997,31.58906,31.347937,31.105,30.862062,30.096992,29.331923,28.56685,27.80178,27.03671,27.207129,27.377548,27.547966,27.718386,27.88699,33.757362,39.627735,45.498108,51.36848,57.23704,59.96736,62.697685,65.42801,68.158325,70.88683,68.22722,65.567604,62.90799,60.24656,57.586945,56.03686,54.48678,52.936695,51.386612,49.83834,46.952106,44.06768,41.183258,38.29702,35.412598,34.714607,34.016617,33.32044,32.622448,31.924458,29.50234,27.080221,24.658104,22.235987,19.812056,20.508232,21.202597,21.896961,22.59314,23.287504,24.737875,26.188244,27.6368,29.087172,30.537542,29.357304,28.177065,26.996826,25.8184,24.63816,20.696781,16.757214,12.817645,8.8780775,4.936697,3.9649491,2.9932013,2.0196402,1.0478923,0.07433146,0.07977036,0.08520924,0.09064813,0.09427405,0.099712946,2.8771715,5.65463,8.432089,11.209548,13.987006,13.724127,13.46306,13.200181,12.937301,12.674421,14.128417,15.580601,17.032784,18.484966,19.93715,19.799364,19.66158,19.525606,19.387821,19.250036,16.276777,13.305332,10.332074,7.360628,4.3873696,3.531651,2.6777458,1.8220274,0.968122,0.11240368,0.09064813,0.06707962,0.045324065,0.02175555,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.045324065,0.09064813,0.13415924,0.1794833,0.22480737,0.19579996,0.16497959,0.13415924,0.10515183,0.07433146,0.20486477,0.33539808,0.46411842,0.5946517,0.72518504,0.62184614,0.52032024,0.4169814,0.3154555,0.21211663,0.22480737,0.2374981,0.25018883,0.26287958,0.2755703,0.291887,0.3100166,0.32814622,0.3444629,0.36259252,0.3045777,0.24837588,0.19036107,0.13234627,0.07433146,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03988518,0.07977036,0.11965553,0.15954071,0.19942589,0.22480737,0.25018883,0.2755703,0.2991388,0.3245203,0.50037766,0.6744221,0.85027945,1.0243238,1.2001812,4.459888,7.7195945,10.979301,14.240821,17.500528,15.290526,13.080525,10.870523,8.660522,6.450521,5.4407005,4.4308805,3.4192474,2.4094272,1.3996071,1.74407,2.0903459,2.4348087,2.7792716,3.1255474,2.7430124,2.3604772,1.9779422,1.5954071,1.2128719,1.1530442,1.0932164,1.0333886,0.97174793,0.9119202,1.3397794,1.7676386,2.1954978,2.6233568,3.049403,2.4529383,1.8546607,1.258196,0.65991837,0.06164073,0.09789998,0.13234627,0.16679256,0.2030518,0.2374981,0.19942589,0.16316663,0.12509441,0.0870222,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.03988518,0.07977036,0.11965553,0.15954071,0.19942589,0.17041849,0.13959812,0.11059072,0.07977036,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.38072214,0.7106813,1.0406405,1.3705997,1.7005589,1.5645868,1.4304274,1.2944553,1.1602961,1.0243238,0.8665961,0.7106813,0.5529536,0.39522585,0.2374981,0.27738327,0.31726846,0.35715362,0.39703882,0.43692398,0.37528324,0.31182957,0.25018883,0.18673515,0.12509441,0.6526665,1.1802386,1.7078108,2.2353828,2.762955,3.3195345,3.877927,4.4345064,4.992899,5.5494785,5.632875,5.714458,5.7978544,5.8794374,5.962834,7.2572894,8.551744,9.848013,11.142468,12.436923,11.048194,9.657652,8.267109,6.87838,5.487838,6.009971,6.532104,7.0542374,7.5781837,8.100317,8.1819,8.265296,8.34688,8.430276,8.511859,7.900891,7.28811,6.6753283,6.0625467,5.4497657,6.3743763,7.2989874,8.225411,9.1500225,10.074633,10.092763,10.109079,10.127209,10.145339,10.161655,10.352016,10.542377,10.7327385,10.9230995,11.111648,12.070704,13.027949,13.985193,14.942437,15.899682,14.387671,12.87566,11.361836,9.849826,8.337815,8.727602,9.117389,9.507175,9.896963,10.28675,10.689227,11.091705,11.494183,11.896661,12.299138,12.06164,11.8241415,11.586644,11.349146,11.111648,11.030065,10.946668,10.865085,10.781689,10.700105,10.440851,10.179785,9.920531,9.659465,9.400211,9.675781,9.949538,10.225109,10.500679,10.774437,10.344765,9.915092,9.48542,9.055748,8.624263,8.734854,8.845445,8.954222,9.064813,9.175404,8.785617,8.39583,8.00423,7.614443,7.224656,9.394773,11.564888,13.735004,15.905121,18.075237,14.804652,11.535881,8.265296,4.994712,1.7241274,1.9706904,2.2154403,2.4601903,2.70494,2.94969,2.9823234,3.0149567,3.04759,3.0802233,3.1128569,3.7401419,4.367427,4.994712,5.621997,6.249282,5.8794374,5.5095935,5.139749,4.7699046,4.40006,5.223145,6.0444174,6.867502,7.690587,8.511859,9.690285,10.866898,12.045323,13.221936,14.400362,13.657047,12.915545,12.172231,11.430729,10.687414,11.30926,11.9329195,12.554766,13.178425,13.800271,14.4692545,15.140051,15.810846,16.47983,17.150625,16.59586,16.03928,15.484513,14.929747,14.37498,12.166792,9.960417,7.752228,5.5458527,3.3376641,4.74271,6.147756,7.552802,8.957849,10.362894,9.893337,9.421967,8.952409,8.482852,8.013294,12.402477,16.79166,21.182655,25.571836,29.962833,29.522284,29.081734,28.642996,28.202446,27.761896,25.885479,24.00725,22.12902,20.252605,18.374376,16.71189,15.049402,13.386916,11.724429,10.061942,8.930654,7.797552,6.6644506,5.5331616,4.40006,4.4870825,4.574105,4.6629395,4.749962,4.836984,5.1578784,5.47696,5.7978544,6.1169357,6.43783,6.1948934,5.9519563,5.710832,5.467895,5.224958,12.032633,18.840307,25.647982,32.455658,39.263332,38.132042,37.002567,35.87309,34.741802,33.612328,31.420454,29.22677,27.034899,24.843027,22.649342,18.684393,14.719443,10.754494,6.789545,2.8245957,2.521831,2.220879,1.9181144,1.6153497,1.3125849,1.4231756,1.5319533,1.6425442,1.7531348,1.8619126,1.8129625,1.7621996,1.7132497,1.6624867,1.6117238,1.3252757,1.0370146,0.7505665,0.46230546,0.17585737,0.35534066,0.53482395,0.71430725,0.89560354,1.0750868,2.6904364,4.305786,5.919323,7.5346723,9.1500225,7.8791356,6.6100616,5.3391747,4.070101,2.7992141,4.615803,6.430578,8.245354,10.060129,11.874905,11.202296,10.529687,9.857078,9.184468,8.511859,7.6833353,6.8529987,6.0226617,5.1923246,4.361988,4.360175,4.358362,4.3547363,4.3529234,4.349297,4.8242936,5.2992897,5.774286,6.249282,6.7242785,7.360628,7.995165,8.629702,9.264238,9.900589,12.210303,14.520018,16.829731,19.139446,21.44916,26.208187,30.9654,35.722614,40.479828,45.23704,42.59737,39.957695,37.318024,34.67835,32.03686,34.339325,36.64179,38.94425,41.24671,43.549175,43.777607,44.004227,44.232662,44.459282,44.687714,44.805557,44.921585,45.03943,45.157272,45.275116,44.31062,43.34431,42.379814,41.415318,40.45082,40.240517,40.030212,39.819912,39.609608,39.399303,38.08309,36.765068,35.447044,34.12902,32.81281,30.104244,27.397491,24.690737,21.982172,19.275417,17.810545,16.34567,14.880796,13.41411,11.949236,13.096842,14.244447,15.392053,16.539658,17.687263,23.062696,28.438131,33.813564,39.187187,44.562622,43.36969,42.17676,40.985645,39.792717,38.599785,38.084904,37.570023,37.05514,36.54026,36.02538,35.318325,34.609455,33.9024,33.195343,32.48829,31.384195,30.281914,29.179632,28.07735,26.97507,32.471973,37.970688,43.46759,48.964493,54.463207,58.303062,62.142918,65.98277,69.822624,73.66248,71.031876,68.403076,65.77247,63.14186,60.513065,59.18779,57.862514,56.53724,55.211964,53.88669,51.457317,49.027946,46.596764,44.167393,41.738026,41.145187,40.552345,39.959507,39.36848,38.775642,35.731678,32.68953,29.647377,26.605227,23.563074,23.385405,23.207733,23.030064,22.852394,22.674723,23.599335,24.525759,25.450369,26.374979,27.299591,27.760082,28.220575,28.679255,29.139748,29.60024,24.504002,19.409578,14.315152,9.220728,4.12449,3.3195345,2.514579,1.7096237,0.90466833,0.099712946,0.10333887,0.10515183,0.10696479,0.11059072,0.11240368,2.6070402,5.101677,7.5981264,10.092763,12.5873995,12.050762,11.512312,10.975676,10.437225,9.900589,12.770509,15.640429,18.510347,21.380268,24.250187,24.424232,24.60009,24.775948,24.949991,25.125849,21.244295,17.364555,13.484816,9.605076,5.7253356,4.610364,3.4953918,2.38042,1.2654479,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.09789998,0.08339628,0.06707962,0.052575916,0.038072214,0.10333887,0.16679256,0.23205921,0.29732585,0.36259252,0.31726846,0.27194437,0.22662032,0.18310922,0.13778515,0.17585737,0.21211663,0.25018883,0.28826106,0.3245203,0.35171473,0.38072214,0.40791658,0.43511102,0.46230546,0.38978696,0.31726846,0.24474995,0.17223145,0.099712946,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,0.2755703,0.2991388,0.3245203,0.34990177,0.37528324,0.387974,0.40066472,0.41335547,0.42423326,0.43692398,4.7118897,8.9868555,13.261822,17.536787,21.811752,19.063301,16.313038,13.562773,10.812509,8.062244,6.4632115,4.8623657,3.2633326,1.6624867,0.06164073,0.16316663,0.26287958,0.36259252,0.46230546,0.5620184,0.6508536,0.73787576,0.824898,0.9119202,1.0007553,1.0116332,1.0243238,1.0370146,1.0497054,1.062396,1.6008459,2.137483,2.6741197,3.2125697,3.7492065,3.000453,2.2498865,1.49932,0.7505665,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,0.21211663,0.17585737,0.13778515,0.099712946,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.4749962,0.8883517,1.2998942,1.7132497,2.124792,1.9126755,1.7005589,1.4866294,1.2745126,1.062396,0.85027945,0.63816285,0.42423326,0.21211663,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.5747091,1.0877775,1.6008459,2.1121013,2.6251698,3.1255474,3.6241121,4.12449,4.6248674,5.125245,5.2630305,5.4008155,5.5367875,5.674573,5.812358,7.362441,8.912524,10.462607,12.012691,13.562773,11.961927,10.362894,8.762048,7.1630154,5.562169,5.8866897,6.2130227,6.5375433,6.8620634,7.1883965,7.324369,7.462154,7.5999393,7.7377243,7.8755093,6.688019,5.5005283,4.313038,3.1255474,1.938057,2.03777,2.137483,2.2371957,2.3369088,2.4366217,3.587853,4.7372713,5.8866897,7.037921,8.187339,8.375887,8.562622,8.749357,8.937905,9.12464,10.25049,11.374527,12.500377,13.6244135,14.750263,13.136727,11.525003,9.91328,8.299743,6.688019,7.037921,7.3878226,7.7377243,8.087626,8.437528,8.588004,8.736667,8.887142,9.037619,9.188094,9.137331,9.088382,9.037619,8.9868555,8.937905,9.249735,9.563377,9.875207,10.1870365,10.500679,9.900589,9.300498,8.700407,8.100317,7.500226,7.9625316,8.424837,8.887142,9.349448,9.811753,9.663091,9.512614,9.362139,9.211663,9.063,9.211663,9.362139,9.512614,9.663091,9.811753,8.80012,7.7866745,6.775041,5.7615952,4.749962,8.036863,11.325577,14.612478,17.89938,21.188093,17.27572,13.363347,9.449161,5.5367875,1.6244144,1.7495089,1.8746033,1.9996977,2.124792,2.2498865,2.175555,2.0994108,2.0250793,1.9507477,1.8746033,2.324218,2.7756457,3.2252605,3.6748753,4.12449,3.925064,3.7256382,3.5243993,3.3249733,3.1255474,4.162562,5.199577,6.2384043,7.2754188,8.312433,9.824444,11.338268,12.850279,14.362289,15.8743,14.762955,13.649796,12.536636,11.42529,10.312131,11.225864,12.137785,13.049705,13.961625,14.875358,15.437376,15.999394,16.563227,17.125244,17.687263,17.01284,16.338419,15.662184,14.9877615,14.313339,12.174044,10.038374,7.899078,5.7615952,3.6241121,5.038223,6.450521,7.8628187,9.275117,10.687414,9.625018,8.562622,7.500226,6.43783,5.375434,10.413657,15.4500675,20.48829,25.5247,30.562923,30.124186,29.687262,29.250338,28.811602,28.374678,25.337965,22.29944,19.262728,16.224201,13.1874895,11.236742,9.287807,7.3370595,5.388125,3.437377,2.7502642,2.0631514,1.3742256,0.6871128,0.0,0.0870222,0.17585737,0.26287958,0.34990177,0.43692398,1.2001812,1.9616255,2.7248828,3.48814,4.249584,4.699199,5.1506267,5.600241,6.049856,6.4994707,14.875358,23.249432,31.625319,39.999393,48.375282,43.875507,39.375732,34.87415,30.374374,25.874601,20.8255,15.774588,10.725487,5.674573,0.62547207,0.50037766,0.37528324,0.25018883,0.12509441,0.0,0.17585737,0.34990177,0.52575916,0.69980353,0.87566096,0.69980353,0.52575916,0.34990177,0.17585737,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13778515,0.2755703,0.41335547,0.5493277,0.6871128,2.5997884,4.512464,6.4251394,8.337815,10.25049,8.575313,6.9001355,5.224958,3.5497808,1.8746033,4.262275,6.6499467,9.037619,11.42529,13.812962,12.763257,11.711739,10.662033,9.612328,8.562622,7.5382986,6.5121617,5.487838,4.461701,3.437377,3.5243993,3.6132345,3.7002566,3.787279,3.874301,4.4870825,5.0998635,5.712645,6.3254266,6.9382076,7.750415,8.562622,9.374829,10.1870365,10.999244,13.899984,16.800724,19.699652,22.600391,25.49932,30.749659,35.999996,41.25034,46.50068,51.749203,47.80057,43.850124,39.89968,35.949234,32.000603,34.750866,37.499317,40.24958,42.999847,45.75011,44.675022,43.599937,42.52485,41.449764,40.374676,40.111797,39.85073,39.587852,39.32497,39.06209,38.262577,37.46306,36.661728,35.862213,35.062695,34.92491,34.787125,34.64934,34.51337,34.375584,32.963287,31.549175,30.136877,28.724579,27.31228,25.024323,22.738176,20.450218,18.16226,15.8743,14.487384,13.100468,11.711739,10.324821,8.937905,10.649343,12.362592,14.075842,15.787278,17.500528,24.250187,30.999847,37.749508,44.50098,51.25064,50.025078,48.799515,47.575764,46.3502,45.124638,44.337814,43.549175,42.76235,41.97552,41.186886,40.53784,39.88699,39.23795,38.587097,37.938053,35.563072,33.18809,30.813112,28.438131,26.06315,31.188395,36.31183,41.437073,46.562317,51.687565,56.63695,61.58815,66.53754,71.48693,76.438126,73.836525,71.23674,68.63695,66.03716,63.437374,62.336906,61.23825,60.137783,59.037315,57.936844,55.96253,53.988213,52.012085,50.037766,48.061638,47.575764,47.088078,46.60039,46.1127,45.625015,41.962833,38.300648,34.63665,30.974466,27.31228,26.262575,25.212872,24.163166,23.11346,22.061941,22.462606,22.863272,23.262123,23.662788,24.06164,26.162863,28.262274,30.361685,32.46291,34.562317,28.311224,22.061941,15.812659,9.563377,3.3122826,2.6741197,2.03777,1.3996071,0.76325727,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,2.3369088,4.550536,6.7623506,8.974165,11.187792,10.375585,9.563377,8.749357,7.93715,7.124943,11.4126,15.700256,19.987913,24.27557,28.563225,29.050913,29.536787,30.024473,30.51216,30.999847,26.211813,21.423779,16.637558,11.849524,7.063302,5.6872635,4.313038,2.9369993,1.5627737,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.12509441,0.18673515,0.25018883,0.31182957,0.37528324,0.41335547,0.44961473,0.48768693,0.52575916,0.5620184,0.4749962,0.387974,0.2991388,0.21211663,0.12509441,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03988518,0.07977036,0.11965553,0.15954071,0.19942589,0.968122,1.7350051,2.5018883,3.2705846,4.0374675,4.8297324,5.621997,6.414262,7.208339,8.000604,10.642091,13.28539,15.926876,18.570175,21.211662,18.755098,16.29672,13.840157,11.381779,8.925215,7.230095,5.5349746,3.8398547,2.1447346,0.44961473,0.44961473,0.44961473,0.44961473,0.44961473,0.44961473,0.5728962,0.69436467,0.81764615,0.93911463,1.062396,1.020698,0.97718686,0.9354887,0.8919776,0.85027945,1.2944553,1.7404441,2.18462,2.6306088,3.0747845,2.4601903,1.845596,1.2291887,0.61459434,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.045324065,0.09064813,0.13415924,0.1794833,0.22480737,0.19217403,0.15954071,0.12690738,0.09427405,0.06164073,0.052575916,0.04169814,0.032633327,0.02175555,0.012690738,0.032633327,0.052575916,0.072518505,0.092461094,0.11240368,0.09427405,0.07795739,0.059827764,0.04169814,0.025381476,0.058014803,0.09064813,0.12328146,0.15410182,0.18673515,0.5275721,0.8665961,1.2074331,1.54827,1.887294,1.745883,1.6026589,1.4594349,1.3180238,1.1747998,0.9554313,0.73424983,0.5148814,0.2955129,0.07433146,0.51306844,0.9499924,1.3869164,1.8256533,2.2625773,1.8202144,1.3778516,0.9354887,0.49312583,0.05076295,0.61459434,1.1802386,1.745883,2.3097143,2.8753586,3.4119956,3.9504454,4.4870825,5.0255322,5.562169,5.7017674,5.8431783,5.9827766,6.1223745,6.261973,7.5419245,8.821876,10.101828,11.381779,12.661731,11.287505,9.91328,8.537241,7.1630154,5.7869763,6.3218007,6.8566246,7.3932614,7.9280853,8.46291,8.283426,8.10213,7.9226465,7.743163,7.5618668,6.4577727,5.351866,4.2477713,3.141864,2.03777,2.084907,2.132044,2.179181,2.228131,2.275268,4.006647,5.7398396,7.473032,9.2044115,10.937603,10.885027,10.832452,10.779876,10.7273,10.674724,11.256684,11.840459,12.42242,13.00438,13.588155,12.335398,11.082641,9.829884,8.577126,7.324369,7.4893484,7.654328,7.819308,7.9842873,8.149267,8.252605,8.354132,8.457471,8.560809,8.662335,8.664148,8.667774,8.669587,8.673213,8.675026,8.901647,9.130079,9.3567,9.585134,9.811753,9.547061,9.282369,9.017676,8.752983,8.488291,8.798307,9.108324,9.418341,9.728357,10.038374,9.73017,9.421967,9.115576,8.807372,8.499168,8.580752,8.660522,8.740293,8.820063,8.899834,8.549932,8.200029,7.850128,7.500226,7.1503243,9.811753,12.474996,15.138238,17.799667,20.462908,16.922194,13.383289,9.842574,6.301858,2.762955,2.8517902,2.9424384,3.0330863,3.1219215,3.2125697,2.9206827,2.6269827,2.335096,2.0432088,1.7495089,2.1592383,2.570781,2.9805105,3.39024,3.7999697,3.9123733,4.024777,4.137181,4.249584,4.361988,5.422571,6.4831543,7.5419245,8.602508,9.663091,10.80707,11.952863,13.096842,14.242634,15.386614,14.3079,13.227375,12.14685,11.068136,9.987611,10.785315,11.583018,12.380721,13.176612,13.974316,14.567154,15.159993,15.752831,16.34567,16.936697,16.367426,15.798156,15.227073,14.657803,14.0867195,12.134158,10.183411,8.23085,6.2782893,4.325729,5.351866,6.379815,7.407765,8.435715,9.461852,8.957849,8.452031,7.948028,7.4422116,6.9382076,11.298383,15.656745,20.01692,24.377094,28.73727,27.839853,26.942436,26.045021,25.147604,24.250187,21.621391,18.99441,16.367426,13.740443,11.111648,10.437225,9.762803,9.088382,8.412147,7.7377243,6.4795284,5.223145,3.9649491,2.7067533,1.4503701,3.0747845,4.699199,6.3254266,7.949841,9.576068,8.997733,8.419398,7.842876,7.264541,6.688019,7.2953615,7.902704,8.510046,9.117389,9.724731,15.522586,21.32044,27.118294,32.914337,38.71219,35.23493,31.757666,28.280403,24.80314,21.324066,18.087927,14.849977,11.612025,8.375887,5.137936,4.160749,3.1817493,2.2045624,1.2273756,0.25018883,0.38434806,0.52032024,0.6544795,0.7904517,0.9246109,0.8629702,0.7995165,0.73787576,0.6744221,0.61278135,0.5529536,0.49312583,0.43329805,0.37165734,0.31182957,0.25018883,0.18673515,0.12509441,0.06164073,0.0,0.14322405,0.28463513,0.42785916,0.56927025,0.7124943,2.222692,3.73289,5.243088,6.7532854,8.26167,6.969028,5.678199,4.3855567,3.092914,1.8002719,3.7673361,5.7344007,7.703278,9.670342,11.637406,10.912222,10.1870365,9.461852,8.736667,8.013294,7.166641,6.3218007,5.47696,4.632119,3.787279,4.15531,4.5233417,4.88956,5.2575917,5.6256227,6.5701766,7.51473,8.459284,9.40565,10.3502035,11.597522,12.84484,14.092158,15.339477,16.586794,19.54555,22.502491,25.459433,28.418188,31.37513,34.792564,38.21,41.627434,45.04487,48.462303,45.072063,41.681824,38.291584,34.903156,31.512915,33.655838,35.796947,37.93987,40.08279,42.22571,41.42257,40.619427,39.818096,39.014954,38.21181,38.494633,38.77746,39.06028,39.3431,39.62411,38.24807,36.87022,35.492367,34.114517,32.736664,32.27255,31.806616,31.342497,30.876566,30.412447,28.936695,27.462757,25.987005,24.513067,23.037315,21.019487,19.001661,16.985647,14.967819,12.949992,11.827768,10.705544,9.583321,8.459284,7.3370595,8.898021,10.457169,12.018129,13.577277,15.138238,20.834566,26.532707,32.23085,37.927177,43.62532,42.68802,41.750717,40.8116,39.8743,38.936996,38.327843,37.716873,37.10772,36.49675,35.887596,35.407158,34.926723,34.4481,33.967667,33.487232,31.891825,30.298231,28.702824,27.107416,25.512009,29.904818,34.297626,38.690434,43.083244,47.47424,52.142616,56.80918,61.477562,66.14413,70.81251,68.60794,66.401566,64.19701,61.992443,59.78788,59.204105,58.622147,58.040184,57.45822,56.87445,55.324368,53.774284,52.2242,50.674118,49.125847,49.860096,50.594345,51.33041,52.06466,52.800724,49.51745,46.235985,42.95271,39.671246,36.387974,34.738174,33.08838,31.436771,29.786976,28.137178,27.190813,26.242634,25.294455,24.348087,23.399908,25.287203,27.174496,29.06179,30.949083,32.838192,27.167244,21.49811,15.827164,10.15803,4.4870825,4.0356545,3.5824142,3.1291735,2.6777458,2.2245052,1.9344311,1.6443571,1.3542831,1.064209,0.774135,2.764768,4.7554007,6.7442207,8.734854,10.725487,10.257742,9.789998,9.322253,8.854509,8.386765,11.583018,14.777458,17.971897,21.166338,24.36259,25.002567,25.642542,26.282518,26.922495,27.56247,23.381779,19.201086,15.022208,10.843329,6.6626377,6.0879283,5.5132194,4.936697,4.361988,3.787279,3.3775494,2.9678197,2.5580902,2.1483607,1.7368182,1.5355793,1.3325275,1.1294757,0.92823684,0.72518504,0.60190356,0.48043507,0.35715362,0.23568514,0.11240368,0.09064813,0.06707962,0.045324065,0.02175555,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,0.2991388,0.32995918,0.36077955,0.38978696,0.42060733,0.44961473,0.387974,0.3245203,0.26287958,0.19942589,0.13778515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,1.6606737,3.1690586,4.6792564,6.189454,7.699652,9.273304,10.845142,12.416981,13.990632,15.56247,16.57229,17.582111,18.59193,19.601751,20.613384,18.446894,16.282217,14.117539,11.952863,9.788185,7.996978,6.207584,4.41819,2.6269827,0.8375887,0.73787576,0.63816285,0.53663695,0.43692398,0.33721104,0.4949388,0.6526665,0.8103943,0.968122,1.1258497,1.0279498,0.9300498,0.8321498,0.73424983,0.63816285,0.9898776,1.3415923,1.69512,2.0468347,2.4003625,1.9199274,1.4394923,0.96087015,0.48043507,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.03988518,0.07977036,0.11965553,0.15954071,0.19942589,0.17223145,0.14503701,0.11784257,0.09064813,0.06164073,0.054388877,0.047137026,0.03988518,0.032633327,0.025381476,0.065266654,0.10515183,0.14503701,0.18492219,0.22480737,0.19036107,0.15410182,0.11965553,0.08520924,0.05076295,0.10333887,0.15410182,0.20667773,0.25925365,0.31182957,0.58014804,0.8466535,1.114972,1.3832904,1.649796,1.5772774,1.504759,1.4322405,1.3597219,1.2872034,1.0605831,0.8321498,0.6055295,0.3770962,0.15047589,1.0243238,1.8999848,2.7756457,3.6494937,4.5251546,3.6277382,2.7303216,1.8329052,0.9354887,0.038072214,0.6544795,1.2726997,1.8909199,2.5073273,3.1255474,3.7002566,4.274966,4.8496747,5.424384,6.000906,6.1423173,6.285541,6.4269524,6.5701766,6.7134004,7.723221,8.733041,9.742861,10.752681,11.762501,10.613083,9.461852,8.312433,7.1630154,6.011784,6.7569118,7.502039,8.247167,8.992294,9.737422,9.24067,8.7421055,8.245354,7.746789,7.250037,6.2275267,5.2050157,4.1825047,3.159994,2.137483,2.132044,2.126605,2.1229792,2.1175404,2.1121013,4.4272547,6.742408,9.057561,11.372714,13.687867,13.394168,13.102281,12.810393,12.516694,12.224807,12.264692,12.304577,12.344462,12.384347,12.4242325,11.532255,10.640278,9.7483,8.854509,7.9625316,7.9425893,7.9226465,7.902704,7.8827615,7.8628187,7.9172077,7.9715962,8.027799,8.082188,8.138389,8.192778,8.247167,8.303369,8.357758,8.412147,8.55537,8.696781,8.840006,8.98323,9.12464,9.195346,9.264238,9.334945,9.40565,9.474543,9.63227,9.789998,9.947725,10.1054535,10.263181,9.79725,9.333132,8.8672,8.403082,7.93715,7.948028,7.957093,7.9679704,7.9770355,7.987913,8.299743,8.613385,8.925215,9.237044,9.550687,11.586644,13.6244135,15.662184,17.699953,19.737724,16.570478,13.403233,10.234174,7.066928,3.8996825,3.9558845,4.0102735,4.064662,4.120864,4.175253,3.6658103,3.1545548,2.6451125,2.13567,1.6244144,1.9942589,2.3641033,2.7357605,3.105605,3.4754493,3.8996825,4.325729,4.749962,5.1741953,5.600241,6.68258,7.764919,8.847258,9.929596,11.011934,11.789696,12.567456,13.345218,14.122978,14.90074,13.852847,12.804955,11.757062,10.70917,9.663091,10.344765,11.028252,11.709926,12.3916,13.075087,13.696932,14.320591,14.942437,15.564283,16.187943,15.722012,15.257894,14.791962,14.327844,13.861912,12.094274,10.328448,8.560809,6.793171,5.0255322,5.667321,6.3091097,6.9527116,7.5945,8.238102,8.290678,8.343254,8.39583,8.448405,8.499168,12.183108,15.865235,19.547363,23.22949,26.911617,25.555521,24.19761,22.839703,21.481794,20.125698,17.906631,15.689378,13.472125,11.254871,9.037619,9.637709,10.2378,10.837891,11.437981,12.038072,10.210606,8.383139,6.5556726,4.7282066,2.9007401,6.0625467,9.224354,12.387974,15.54978,18.7134,16.795286,14.877171,12.96087,11.042755,9.12464,9.88971,10.654781,11.419851,12.184921,12.949992,16.169813,19.389635,22.609457,25.829277,29.049099,26.594349,24.139597,21.684845,19.230095,16.775343,15.350354,13.925365,12.500377,11.075388,9.6504,7.819308,5.9900284,4.160749,2.3296568,0.50037766,0.5946517,0.69073874,0.7850128,0.8792868,0.97537386,1.0243238,1.0750868,1.1258497,1.1747998,1.2255627,1.1040943,0.98443866,0.86478317,0.7451276,0.62547207,0.50037766,0.37528324,0.25018883,0.12509441,0.0,0.14684997,0.2955129,0.44236287,0.58921283,0.73787576,1.845596,2.953316,4.059223,5.1669436,6.2746634,5.3645563,4.454449,3.5443418,2.6342347,1.7241274,3.2723975,4.8206677,6.3671246,7.915395,9.461852,9.063,8.662335,8.26167,7.8628187,7.462154,6.796797,6.1332526,5.467895,4.802538,4.137181,4.784408,5.431636,6.0806766,6.7279043,7.3751316,8.653271,9.929596,11.207735,12.485873,13.762199,15.444629,17.127058,18.809486,20.491917,22.174345,25.191114,28.204258,31.22103,34.235985,37.250942,38.835472,40.420002,42.00453,43.590874,45.1754,42.345367,39.51533,36.6853,33.855263,31.025229,32.560806,34.094574,35.630154,37.165733,38.6995,38.170113,37.640728,37.10953,36.580147,36.050762,36.877472,37.70418,38.532707,39.359417,40.187943,38.231754,36.27738,34.32301,32.36682,30.412447,29.620182,28.827917,28.035654,27.241575,26.44931,24.911919,23.374527,21.837133,20.299742,18.76235,17.014654,15.266958,13.519262,11.771566,10.025683,9.168152,8.31062,7.453089,6.5955577,5.7380266,7.1448855,8.551744,9.960417,11.367275,12.774135,17.420757,22.065567,26.710379,31.355188,35.999996,35.349144,34.700104,34.04925,33.40021,32.749355,32.31787,31.884573,31.453089,31.01979,30.588305,30.278288,29.968271,29.658255,29.348238,29.038221,28.22239,27.40837,26.592535,25.776703,24.962683,28.623053,32.281612,35.941982,39.602356,43.262726,47.64828,52.032024,56.417583,60.80314,65.18688,63.377544,61.56821,59.75706,57.947723,56.136574,56.07312,56.007854,55.942585,55.87732,55.812054,54.688015,53.56217,52.43813,51.31228,50.188244,52.14443,54.10243,56.06043,58.016617,59.974617,57.072063,54.16951,51.266956,48.364403,45.46185,43.211964,40.96208,38.71219,36.462303,34.212418,31.917206,29.621996,27.326784,25.033388,22.738176,24.413355,26.08672,27.761896,29.437073,31.112251,26.021452,20.932467,15.841667,10.752681,5.661882,5.3953767,5.127058,4.860553,4.592234,4.325729,3.7455807,3.1654327,2.5852847,2.0051367,1.4249886,3.1926272,4.9602656,6.7279043,8.495543,10.263181,10.139899,10.016619,9.89515,9.771869,9.6504,11.753436,13.85466,15.957697,18.060734,20.161957,20.954222,21.748299,22.540564,23.332829,24.125093,20.551744,16.980207,13.406858,9.835322,6.261973,6.48678,6.7134004,6.9382076,7.1630154,7.3878226,6.604623,5.823236,5.040036,4.256836,3.4754493,3.0693457,2.665055,2.2607644,1.8546607,1.4503701,1.2056202,0.96087015,0.71430725,0.46955732,0.22480737,0.1794833,0.13415924,0.09064813,0.045324065,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.22480737,0.24837588,0.27013144,0.291887,0.3154555,0.33721104,0.2991388,0.26287958,0.22480737,0.18673515,0.15047589,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,2.3532255,4.604925,6.8584375,9.110137,11.361836,13.715062,16.068287,18.4197,20.772924,23.124338,22.502491,21.880646,21.256987,20.63514,20.013294,18.140503,16.267714,14.394923,12.522133,10.649343,8.765674,6.880193,4.994712,3.1092308,1.2255627,1.0243238,0.824898,0.62547207,0.42423326,0.22480737,0.4169814,0.6091554,0.8031424,0.99531645,1.1874905,1.0352017,0.88291276,0.7306239,0.57833505,0.42423326,0.6852999,0.9445535,1.2056202,1.4648738,1.7241274,1.3796645,1.0352017,0.69073874,0.3444629,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.034446288,0.07070554,0.10515183,0.13959812,0.17585737,0.15228885,0.13053331,0.10696479,0.08520924,0.06164073,0.058014803,0.052575916,0.047137026,0.04169814,0.038072214,0.09789998,0.15772775,0.21755551,0.27738327,0.33721104,0.28463513,0.23205921,0.1794833,0.12690738,0.07433146,0.14684997,0.21936847,0.291887,0.36440548,0.43692398,0.6327239,0.82671094,1.0225109,1.2183108,1.4122978,1.4104849,1.4068589,1.405046,1.403233,1.3996071,1.1657349,0.9300498,0.69436467,0.4604925,0.22480737,1.5373923,2.8499773,4.162562,5.475147,6.787732,5.4352617,4.082792,2.7303216,1.3778516,0.025381476,0.69436467,1.3651608,2.034144,2.70494,3.3757362,3.9867048,4.599486,5.2122674,5.825049,6.43783,6.582867,6.7279043,6.872941,7.017978,7.1630154,7.902704,8.642392,9.382081,10.12177,10.863272,9.936848,9.012237,8.087626,7.1630154,6.2384043,7.192023,8.147454,9.102885,10.058316,11.011934,10.197914,9.382081,8.568061,7.752228,6.9382076,5.99728,5.0581656,4.117238,3.1781235,2.2371957,2.179181,2.1229792,2.0649643,2.0069497,1.9507477,4.847862,7.744976,10.642091,13.539205,16.438131,15.905121,15.372109,14.839099,14.3079,13.77489,13.272699,12.770509,12.268318,11.764315,11.262123,10.729113,10.197914,9.664904,9.131892,8.600695,8.39583,8.189152,7.9842873,7.7794223,7.574558,7.5818095,7.590874,7.5981264,7.605378,7.61263,7.7195945,7.8283725,7.935337,8.042302,8.149267,8.207282,8.265296,8.323311,8.379513,8.437528,8.841819,9.247922,9.652213,10.058316,10.462607,10.468046,10.471672,10.477111,10.48255,10.487988,9.864329,9.242483,8.620637,7.996978,7.3751316,7.315304,7.2554765,7.1956487,7.135821,7.07418,8.049554,9.024928,10.000301,10.975676,11.949236,13.363347,14.775645,16.187943,17.60024,19.012539,16.21695,13.423175,10.627586,7.8319983,5.038223,5.0581656,5.0781083,5.0980506,5.1179934,5.137936,4.409125,3.682127,2.955129,2.228131,1.49932,1.8292793,2.1592383,2.4891977,2.819157,3.149116,3.8869917,4.6248674,5.3627434,6.1006193,6.836682,7.9425893,9.046683,10.152591,11.256684,12.362592,12.772322,13.182051,13.591781,14.003323,14.413053,13.397794,12.382534,11.367275,10.352016,9.336758,9.904215,10.471672,11.039129,11.608399,12.175857,12.826711,13.479377,14.132043,14.78471,15.437376,15.076597,14.71763,14.356851,13.997884,13.637105,12.054388,10.471672,8.890768,7.308052,5.7253356,5.9827766,6.240217,6.497658,6.755099,7.0125394,7.6216946,8.232663,8.841819,9.452786,10.061942,13.067834,16.071913,19.077805,22.081884,25.087776,23.269375,21.452785,19.634384,17.817797,15.999394,14.191871,12.384347,10.576823,8.7693,6.9617763,8.838193,10.712796,12.5873995,14.462003,16.336605,13.939869,11.543133,9.144584,6.7478466,4.349297,9.050309,13.749508,18.45052,23.14972,27.85073,24.592838,21.334944,18.07705,14.819156,11.563075,12.485873,13.406858,14.329657,15.252454,16.175253,16.817041,17.460642,18.102432,18.74422,19.387821,17.955582,16.52334,15.089288,13.657047,12.224807,12.612781,13.000754,13.386916,13.77489,14.162864,11.479679,8.798307,6.115123,3.4319382,0.7505665,0.80495536,0.85934424,0.9155461,0.969935,1.0243238,1.1874905,1.3506571,1.5120108,1.6751775,1.8383441,1.6570477,1.4775645,1.2980812,1.1167849,0.93730164,0.7505665,0.5620184,0.37528324,0.18673515,0.0,0.15228885,0.3045777,0.45686656,0.6091554,0.76325727,1.4666867,2.1719291,2.8771715,3.5824142,4.2876563,3.7600844,3.2325122,2.70494,2.1773682,1.649796,2.7774587,3.9051213,5.032784,6.1604466,7.28811,7.211965,7.137634,7.063302,6.987158,6.9128265,6.4269524,5.942891,5.4570174,4.972956,4.4870825,5.4153194,6.341743,7.26998,8.198216,9.12464,10.734551,12.344462,13.954373,15.564283,17.174194,19.291735,21.409275,23.526815,25.644356,27.761896,30.834867,33.90784,36.980812,40.051968,43.124943,42.876564,42.63,42.381626,42.135063,41.88669,39.61686,37.34703,35.0772,32.80737,30.537542,31.465778,32.392204,33.32044,34.246864,35.1751,34.91766,34.660217,34.40278,34.145336,33.887897,35.26031,36.63272,38.005135,39.37755,40.74996,38.21725,35.684544,33.151833,30.619125,28.08823,26.96782,25.847408,24.726997,23.608398,22.487988,20.887142,19.288109,17.687263,16.08823,14.487384,13.009819,11.532255,10.05469,8.577126,7.0995617,6.506723,5.915697,5.3228583,4.7300196,4.137181,5.391751,6.6481338,7.902704,9.157274,10.411844,14.005136,17.596615,21.189907,24.7832,28.374678,28.012085,27.649492,27.2869,26.924307,26.561714,26.3079,26.052273,25.796644,25.54283,25.287203,25.147604,25.008005,24.868408,24.726997,24.587399,24.552952,24.516693,24.482246,24.4478,24.413355,27.339476,30.26741,33.195343,36.12328,39.0494,43.152134,47.25487,51.357605,55.46034,59.563072,58.14715,56.73304,55.317116,53.903004,52.48708,52.94032,53.391747,53.84499,54.29823,54.749657,54.049854,53.350048,52.650246,51.950443,51.25064,54.430576,57.61051,60.790447,63.970387,67.15032,64.62668,62.104847,59.583015,57.059372,54.53754,51.687565,48.837585,45.98761,43.13763,40.287655,36.645412,33.00317,29.359116,25.716875,22.074633,23.537693,25.000753,26.462002,27.925062,29.388123,24.877472,20.366821,15.857984,11.347333,6.836682,6.755099,6.6717024,6.590119,6.506723,6.4251394,5.5549173,4.6846952,3.8144734,2.9442513,2.0758421,3.6204863,5.1651306,6.7097745,8.254418,9.800876,10.022058,10.245051,10.468046,10.689227,10.912222,11.922042,12.931862,13.941682,14.953316,15.963136,16.907688,17.852243,18.796797,19.743162,20.687716,17.721708,14.757515,11.793322,8.827314,5.863121,6.887445,7.911769,8.937905,9.96223,10.988366,9.8316965,8.676839,7.5219817,6.3671246,5.2122674,4.604925,3.9975824,3.39024,2.7828975,2.175555,1.8075237,1.4394923,1.0732739,0.70524246,0.33721104,0.27013144,0.2030518,0.13415924,0.06707962,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.15047589,0.16497959,0.1794833,0.19579996,0.21030366,0.22480737,0.21211663,0.19942589,0.18673515,0.17585737,0.16316663,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,3.045777,6.0407915,9.035806,12.03082,15.025834,18.15682,21.28962,24.422419,27.555218,30.688017,28.432692,26.177366,23.92204,21.666716,19.413204,17.8323,16.25321,14.672306,13.093216,11.512312,9.5325575,7.552802,5.573047,3.5932918,1.6117238,1.3125849,1.0116332,0.7124943,0.41335547,0.11240368,0.34083697,0.56745726,0.79589057,1.0225109,1.2491312,1.0424535,0.83577573,0.62728506,0.42060733,0.21211663,0.38072214,0.5475147,0.71430725,0.88291276,1.0497054,0.83940166,0.629098,0.42060733,0.21030366,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.13234627,0.11421664,0.09789998,0.07977036,0.06164073,0.059827764,0.058014803,0.054388877,0.052575916,0.05076295,0.13053331,0.21030366,0.29007402,0.36984438,0.44961473,0.38072214,0.3100166,0.23931105,0.17041849,0.099712946,0.19217403,0.28463513,0.3770962,0.46955732,0.5620184,0.6852999,0.80676836,0.9300498,1.0533313,1.1747998,1.2418793,1.310772,1.3778516,1.4449311,1.5120108,1.2708868,1.0279498,0.7850128,0.5420758,0.2991388,2.0504606,3.7999697,5.5494785,7.3008003,9.050309,7.2427855,5.4352617,3.6277382,1.8202144,0.012690738,0.73424983,1.4576219,2.179181,2.902553,3.6241121,4.274966,4.9258194,5.57486,6.2257137,6.874754,7.021604,7.170267,7.317117,7.46578,7.61263,8.082188,8.551744,9.023115,9.492672,9.96223,9.262425,8.562622,7.8628187,7.1630154,6.4632115,7.6271334,8.792869,9.956791,11.122525,12.28826,11.155159,10.022058,8.890768,7.757667,6.624565,5.767034,4.9095025,4.0519714,3.1944401,2.3369088,2.228131,2.1175404,2.0069497,1.8981718,1.7875811,5.2666564,8.747544,12.228433,15.707508,19.188396,18.41426,17.64194,16.869617,16.097294,15.324973,14.280706,13.234627,12.19036,11.144281,10.100015,9.927783,9.755551,9.583321,9.409276,9.237044,8.847258,8.457471,8.067683,7.6778965,7.28811,7.2482243,7.208339,7.166641,7.1267557,7.0868707,7.2482243,7.407765,7.567306,7.7268467,7.8882003,7.859193,7.8319983,7.804804,7.7776093,7.750415,8.490104,9.229793,9.969481,10.70917,11.450671,11.302009,11.155159,11.008308,10.859646,10.712796,9.933222,9.151835,8.372261,7.592687,6.813113,6.68258,6.552047,6.4233265,6.2927933,6.16226,7.799365,9.438283,11.075388,12.712494,14.349599,15.138238,15.925063,16.71189,17.500528,18.287354,15.865235,13.443117,11.019187,8.597069,6.1749506,6.1604466,6.14413,6.1296263,6.115123,6.1006193,5.1542525,4.209699,3.2651455,2.3205922,1.3742256,1.6642996,1.9543737,2.2444477,2.5345216,2.8245957,3.874301,4.9258194,5.975525,7.02523,8.074935,9.202598,10.330261,11.457924,12.585587,13.713249,13.754947,13.796645,13.840157,13.881854,13.925365,12.9427395,11.9601145,10.9774885,9.994863,9.012237,9.465478,9.916905,10.370146,10.823386,11.274815,11.958302,12.639976,13.321649,14.005136,14.68681,14.432995,14.177367,13.92174,13.667925,13.412297,12.0145035,10.616709,9.220728,7.8229337,6.4251394,6.298232,6.169512,6.0426044,5.915697,5.7869763,6.9545245,8.122072,9.28962,10.457169,11.624716,13.95256,16.280403,18.608248,20.934278,23.262123,20.985043,18.70796,16.429068,14.151986,11.874905,10.477111,9.079316,7.6815224,6.285541,4.8877473,8.036863,11.187792,14.336908,17.487837,20.636953,17.669134,14.703127,11.735307,8.767487,5.7996674,12.038072,18.274662,24.513067,30.749659,36.988064,32.39039,27.792717,23.195044,10258.0,13.999697,15.080223,16.160748,17.239462,18.319986,19.400513,17.464268,15.529838,13.595407,11.6591625,9.724731,9.3150015,8.9052725,8.495543,8.0858135,7.6742706,9.875207,12.07433,14.275268,16.474392,18.675327,15.140051,11.6047735,8.069496,4.5342193,1.0007553,1.015259,1.0297627,1.0442665,1.0605831,1.0750868,1.3506571,1.6244144,1.8999848,2.175555,2.4493124,2.2100015,1.9706904,1.7295663,1.4902552,1.2491312,1.0007553,0.7505665,0.50037766,0.25018883,0.0,0.15772775,0.3154555,0.47318324,0.629098,0.7868258,1.0895905,1.3923552,1.69512,1.9978848,2.3006494,2.1556125,2.0105755,1.8655385,1.7205015,1.5754645,2.2825198,2.9895754,3.6966307,4.405499,5.1125546,5.3627434,5.612932,5.863121,6.11331,6.3616858,6.057108,5.75253,5.4479527,5.143375,4.836984,6.0444174,7.25185,8.459284,9.666717,10.874149,12.817645,14.759329,16.702824,18.644506,20.588003,23.140654,25.693306,28.245956,30.796795,33.349445,36.480434,39.609608,42.740593,45.869766,49.00075,46.91947,44.840004,42.760536,40.679253,38.599785,36.890163,35.18054,33.4691,31.759478,30.049854,30.370749,30.68983,31.010725,31.329807,31.650702,31.665205,31.679708,31.694212,31.71053,31.725033,33.643147,35.55945,37.477562,39.395676,41.311977,38.202747,35.091705,31.982473,28.873241,25.762197,24.315454,22.866898,21.420153,19.971596,18.52485,16.862366,15.199879,13.537392,11.874905,10.212419,9.004985,7.797552,6.590119,5.382686,4.175253,3.8471067,3.5207734,3.1926272,2.864481,2.5381477,3.6404288,4.74271,5.844991,6.947273,8.049554,10.589515,13.129475,15.6694355,18.209396,20.749357,20.675026,20.600695,20.52455,20.450218,20.374073,20.29793,20.219973,20.142014,20.064056,19.987913,20.01692,20.04774,20.076748,20.107569,20.136576,20.881702,21.626831,22.371958,23.117086,23.862213,26.05771,28.253208,30.446894,32.64239,34.83789,38.657803,42.477715,46.297626,50.11754,53.93745,52.91675,51.897865,50.87717,49.858284,48.837585,49.80752,50.777454,51.74739,52.717327,53.68726,53.41169,53.13793,52.862362,52.586792,52.313034,56.71491,61.116783,65.52047,69.92234,74.32421,72.183105,70.040184,67.89726,65.75615,63.61323,60.163162,56.713097,53.263027,49.81296,46.362892,41.371807,36.382534,31.393261,26.402174,21.4129,22.662033,23.912977,25.162107,26.413052,27.662184,23.73168,19.80299,15.872487,11.941984,8.013294,8.1148205,8.21816,8.319685,8.423024,8.52455,7.364254,6.205771,5.045475,3.8851788,2.7248828,4.0483456,5.369995,6.6916447,8.015107,9.336758,9.904215,10.471672,11.039129,11.606586,12.175857,12.092461,12.010877,11.927481,11.844085,11.762501,12.859344,13.957999,15.054841,16.151684,17.25034,14.891675,12.534823,10.177972,7.819308,5.462456,7.28811,9.11195,10.937603,12.763257,14.587097,13.060582,11.532255,10.00574,8.477413,6.9508986,6.1405044,5.33011,4.519716,3.7093215,2.9007401,2.4094272,1.9199274,1.4304274,0.94092757,0.44961473,0.36077955,0.27013144,0.1794833,0.09064813,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.07433146,0.08339628,0.09064813,0.09789998,0.10515183,0.11240368,0.12509441,0.13778515,0.15047589,0.16316663,0.17585737,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,3.738329,7.474845,11.213174,14.94969,18.688019,22.600391,26.512764,30.425138,34.337513,38.249886,34.362892,30.4759,26.587097,22.700104,18.813112,17.52591,16.236893,14.94969,13.662486,12.375282,10.29944,8.225411,6.149569,4.07554,1.9996977,1.6008459,1.2001812,0.7995165,0.40066472,0.0,0.26287958,0.52575916,0.7868258,1.0497054,1.3125849,1.0497054,0.7868258,0.52575916,0.26287958,0.0,0.07433146,0.15047589,0.22480737,0.2991388,0.37528324,0.2991388,0.22480737,0.15047589,0.07433146,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.16316663,0.26287958,0.36259252,0.46230546,0.5620184,0.4749962,0.387974,0.2991388,0.21211663,0.12509441,0.2374981,0.34990177,0.46230546,0.5747091,0.6871128,0.73787576,0.7868258,0.8375887,0.8883517,0.93730164,1.0750868,1.2128719,1.3506571,1.4866294,1.6244144,1.3742256,1.1258497,0.87566096,0.62547207,0.37528324,2.561716,4.749962,6.9382076,9.12464,11.312886,9.050309,6.787732,4.5251546,2.2625773,0.0,0.774135,1.550083,2.324218,3.100166,3.874301,4.5632267,5.2503395,5.9374523,6.624565,7.311678,7.462154,7.61263,7.763106,7.911769,8.062244,8.26167,8.46291,8.662335,8.861761,9.063,8.588004,8.113008,7.6380115,7.1630154,6.688019,8.062244,9.438283,10.812509,12.186734,13.562773,12.112403,10.662033,9.211663,7.763106,6.3127356,5.5367875,4.762653,3.9867048,3.2125697,2.4366217,2.275268,2.1121013,1.9507477,1.7875811,1.6244144,5.6872635,9.750113,13.812962,17.87581,21.936848,20.925215,19.911768,18.900135,17.886688,16.875055,15.2869005,13.700559,12.112403,10.524248,8.937905,9.12464,9.313189,9.499924,9.686659,9.875207,9.300498,8.725789,8.149267,7.574558,6.9998484,6.9128265,6.825804,6.736969,6.6499467,6.5629244,6.775041,6.987158,7.1992745,7.413204,7.6253204,7.512917,7.400513,7.28811,7.175706,7.063302,8.138389,9.211663,10.28675,11.361836,12.436923,12.137785,11.836833,11.537694,11.236742,10.937603,10.000301,9.063,8.125698,7.1865835,6.249282,6.049856,5.8504305,5.6491914,5.4497657,5.2503395,7.549176,9.849826,12.1504755,14.449312,16.749962,16.913128,17.074482,17.237648,17.400814,17.562168,15.511708,13.46306,11.4126,9.362139,7.311678,7.262728,7.211965,7.1630154,7.112252,7.063302,5.89938,4.7372713,3.5751622,2.4130533,1.2491312,1.49932,1.7495089,1.9996977,2.2498865,2.5000753,3.8616104,5.224958,6.588306,7.949841,9.313189,10.462607,11.612025,12.763257,13.912675,15.062093,14.737573,14.413053,14.0867195,13.762199,13.437678,12.487686,11.537694,10.587702,9.637709,8.6877165,9.024928,9.362139,9.699349,10.038374,10.375585,11.088079,11.800573,12.513068,13.225562,13.938056,13.7875805,13.637105,13.486629,13.337966,13.1874895,11.974618,10.761745,9.550687,8.337815,7.124943,6.6118746,6.1006193,5.5875506,5.0744824,4.5632267,6.2873545,8.013294,9.737422,11.463363,13.1874895,14.837286,16.487082,18.136877,19.786674,21.438282,18.700708,15.963136,13.225562,10.487988,7.750415,6.7623506,5.774286,4.788034,3.7999697,2.811905,7.2373466,11.662788,16.08823,20.511858,24.9373,21.40021,17.863121,14.324218,10.7871275,7.250037,15.025834,22.799818,30.575613,38.349598,46.125393,40.187943,34.25049,28.313036,22.375584,16.438131,17.674572,18.912827,20.149265,21.38752,22.625772,18.111496,13.600845,9.086569,4.574105,0.06164073,0.6744221,1.2872034,1.8999848,2.5127661,3.1255474,7.137634,11.14972,15.161806,19.175705,23.187792,18.800423,14.413053,10.025683,5.638314,1.2491312,1.2255627,1.2001812,1.1747998,1.1494182,1.1258497,1.5120108,1.8999848,2.2879589,2.6741197,3.0620937,2.762955,2.4620032,2.1628644,1.8619126,1.5627737,1.2491312,0.93730164,0.62547207,0.31182957,0.0,0.16316663,0.3245203,0.48768693,0.6508536,0.8122072,0.7124943,0.61278135,0.51306844,0.41335547,0.31182957,0.5493277,0.7868258,1.0243238,1.261822,1.49932,1.7875811,2.0758421,2.3622901,2.6505513,2.9369993,3.5117085,4.0882306,4.6629395,5.237649,5.812358,5.6872635,5.562169,5.4370747,5.3119802,5.186886,6.6753283,8.161958,9.6504,11.137029,12.625471,14.90074,17.174194,19.449463,21.724731,23.999998,26.98776,29.975523,32.963287,35.949234,38.936996,42.126,45.313187,48.500374,51.687565,54.874752,50.96238,47.050003,43.13763,39.225258,35.312885,34.161655,33.012238,31.862818,30.711586,29.562168,29.27572,28.98746,28.699198,28.41275,28.124489,28.41275,28.699198,28.98746,29.27572,29.562168,32.025986,34.487988,36.94999,39.411995,41.87581,38.18643,34.50068,30.813112,27.125546,23.43798,21.66309,19.888199,18.11331,16.336605,14.561715,12.837588,11.111648,9.38752,7.66158,5.9374523,5.0001507,4.062849,3.1255474,2.1882458,1.2491312,1.1874905,1.1258497,1.062396,1.0007553,0.93730164,1.887294,2.8372865,3.787279,4.7372713,5.6872635,7.175706,8.662335,10.150778,11.637406,13.125849,13.337966,13.550082,13.762199,13.974316,14.188245,14.287958,14.387671,14.487384,14.587097,14.68681,14.888049,15.087475,15.2869005,15.488139,15.687565,17.212267,18.736969,20.26167,21.788185,23.312885,24.775948,26.237194,27.700254,29.163317,30.624563,34.163467,37.700558,41.237648,44.77474,48.31183,47.688168,47.062695,46.437225,45.811752,45.18809,46.67472,48.163162,49.64979,51.138237,52.624866,52.77534,52.925816,53.07448,53.224957,53.37543,59.001053,64.62486,70.25049,75.8743,81.49992,79.73772,77.97552,76.21332,74.44931,72.68711,68.63695,64.58679,60.536633,56.48829,52.43813,46.100014,39.761894,33.42559,27.087475,20.749357,21.788185,22.8252,23.862213,24.89923,25.938055,22.5877,19.237347,15.8869915,12.538449,9.188094,9.474543,9.762803,10.049252,10.337513,10.625773,9.175404,7.7250338,6.2746634,4.8242936,3.3757362,4.4743915,5.57486,6.6753283,7.7757964,8.874452,9.788185,10.700105,11.612025,12.525759,13.437678,12.262879,11.088079,9.91328,8.736667,7.5618668,8.812811,10.061942,11.312886,12.562017,13.812962,12.06164,10.312131,8.562622,6.813113,5.0617914,7.686961,10.312131,12.937301,15.56247,18.187641,16.287657,14.387671,12.487686,10.587702,8.6877165,7.6742706,6.6626377,5.6491914,4.6375585,3.6241121,3.0131438,2.4003625,1.7875811,1.1747998,0.5620184,0.44961473,0.33721104,0.22480737,0.11240368,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,3.0856624,6.169512,9.255174,12.340837,15.4246855,18.526665,21.630457,24.732435,27.834415,30.938206,27.894243,24.85209,21.80994,18.767788,15.725637,14.764768,13.80571,12.84484,11.885782,10.924912,9.3693905,7.8156815,6.26016,4.704638,3.150929,2.6324217,2.1157274,1.5972201,1.0805258,0.5620184,0.6726091,0.78319985,0.8919776,1.0025684,1.1131591,0.9119202,0.7124943,0.51306844,0.31182957,0.11240368,0.15047589,0.18673515,0.22480737,0.26287958,0.2991388,0.23931105,0.1794833,0.11965553,0.059827764,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.09064813,0.07977036,0.07070554,0.059827764,0.05076295,0.052575916,0.054388877,0.058014803,0.059827764,0.06164073,0.15047589,0.2374981,0.3245203,0.41335547,0.50037766,0.4224203,0.3444629,0.26831847,0.19036107,0.11240368,0.19942589,0.28826106,0.37528324,0.46230546,0.5493277,0.76325727,0.97537386,1.1874905,1.3996071,1.6117238,1.5645868,1.5174497,1.4703126,1.4231756,1.3742256,1.2273756,1.0805258,0.9318628,0.7850128,0.63816285,2.3296568,4.022964,5.714458,7.407765,9.099259,7.28811,5.475147,3.6621845,1.8492218,0.038072214,0.9572442,1.8782293,2.7974012,3.7183862,4.6375585,5.3627434,6.0879283,6.813113,7.5382986,8.26167,8.009668,7.757667,7.5056653,7.25185,6.9998484,7.07418,7.1503243,7.224656,7.3008003,7.3751316,7.017978,6.6608243,6.301858,5.9447045,5.5875506,7.117691,8.647832,10.177972,11.708113,13.238253,11.9021,10.567759,9.231606,7.897265,6.5629244,5.660069,4.7572136,3.8543584,2.953316,2.0504606,2.3169663,2.5852847,2.8517902,3.1201086,3.388427,6.9019485,10.417283,13.932617,17.447952,20.963285,20.326937,19.6924,19.057863,18.423326,17.786976,15.979452,14.171928,12.364405,10.556881,8.749357,8.63514,8.519112,8.404895,8.290678,8.174648,7.6724577,7.170267,6.6680765,6.164073,5.661882,5.6074934,5.5531044,5.4969025,5.4425135,5.388125,5.7906027,6.19308,6.5955577,6.9980354,7.400513,7.304426,7.210152,7.115878,7.019791,6.925517,7.667019,8.410334,9.151835,9.89515,10.636651,10.943042,11.24762,11.552197,11.856775,12.163166,10.883214,9.603263,8.323311,7.0433598,5.7615952,5.5349746,5.3083544,5.0799212,4.853301,4.6248674,6.7297173,8.834567,10.939416,13.044266,15.149116,15.199879,15.250641,15.299591,15.350354,15.399304,13.80571,12.210303,10.614896,9.019489,7.4258947,7.502039,7.5799966,7.6579537,7.7359114,7.8120556,6.60281,5.391751,4.1825047,2.9732587,1.7621996,2.0758421,2.3876717,2.6995013,3.0131438,3.3249733,4.4798307,5.634688,6.789545,7.944402,9.099259,9.99305,10.885027,11.777005,12.670795,13.562773,13.294455,13.027949,12.75963,12.493125,12.224807,11.731681,11.240368,10.747242,10.254116,9.762803,10.032935,10.303066,10.573197,10.843329,11.111648,11.73712,12.362592,12.988064,13.611723,14.237195,13.987006,13.736817,13.486629,13.238253,12.988064,11.583018,10.177972,8.772926,7.36788,5.962834,5.8431783,5.7217097,5.6020546,5.482399,5.3627434,6.5574856,7.752228,8.94697,10.141713,11.338268,12.565643,13.793019,15.020395,16.24777,17.475147,16.492521,15.509895,14.527269,13.544643,12.562017,11.144281,9.728357,8.31062,6.892884,5.475147,8.370448,11.26575,14.159238,17.054539,19.94984,17.132496,14.315152,11.497808,8.680465,5.863121,12.228433,18.59193,24.957243,31.322554,37.687866,32.783802,27.883364,22.979301,18.07705,13.174799,14.159238,15.14549,16.129929,17.114367,18.100618,14.512766,10.924912,7.3370595,3.7492065,0.16316663,0.69073874,1.2183108,1.745883,2.2716422,2.7992141,5.9501433,9.099259,12.250188,15.399304,18.550234,15.040338,11.530442,8.020547,4.510651,1.0007553,0.9808127,0.96087015,0.93911463,0.91917205,0.89922947,1.3724127,1.845596,2.3169663,2.7901495,3.2633326,2.8608549,2.4583774,2.0540867,1.651609,1.2491312,1.0007553,0.7505665,0.50037766,0.25018883,0.0,0.13053331,0.25925365,0.38978696,0.52032024,0.6508536,0.56927025,0.4894999,0.40972954,0.32995918,0.25018883,0.4949388,0.73968875,0.98443866,1.2291887,1.4757515,1.7023718,1.9308052,2.1574254,2.3858588,2.612479,3.1654327,3.7165732,4.269527,4.8224807,5.375434,5.2630305,5.1506267,5.038223,4.9258194,4.8116026,5.964647,7.117691,8.270736,9.421967,10.57501,12.806767,15.040338,17.272095,19.505665,21.737421,24.117842,26.496449,28.876867,31.257288,33.637707,36.320892,39.002266,41.685448,44.36682,47.050003,44.406704,41.76522,39.121918,36.480434,33.837135,34.645714,35.452484,36.25925,37.067833,37.8746,36.549324,35.225864,33.90059,32.575314,31.250036,32.82006,34.390087,35.960114,37.53014,39.100163,40.789845,42.479527,44.17102,45.860703,47.55038,42.62275,37.695118,32.767487,27.839853,22.912222,20.97779,19.04336,17.107115,15.172684,13.238253,11.650098,10.061942,8.4756,6.887445,5.2992897,4.5342193,3.7691493,3.004079,2.2408218,1.4757515,1.4068589,1.3397794,1.2726997,1.2056202,1.1367276,1.8582866,2.5780327,3.2977788,4.017525,4.7372713,6.017223,7.2971745,8.577126,9.857078,11.137029,11.253058,11.367275,11.483305,11.597522,11.711739,11.999999,12.28826,12.574709,12.862969,13.149418,13.310771,13.470312,13.629852,13.789393,13.9507475,15.0421505,16.135366,17.22677,18.319986,19.413204,20.881702,22.352016,23.822329,25.29264,26.762953,30.049854,33.336758,36.62547,39.912373,43.199272,42.999847,42.80042,42.599182,42.399757,42.20033,43.772167,45.344006,46.91766,48.4895,50.06315,50.509136,50.95694,51.40474,51.852543,52.300346,57.313187,62.324215,67.33706,72.3499,77.36274,76.46713,75.57335,74.67774,73.782135,72.88835,69.663086,66.43783,63.212566,59.987305,56.762047,50.857227,44.952408,39.04759,33.14277,27.23795,27.61686,27.997581,28.378304,28.757212,29.137934,26.27164,23.40716,20.542679,17.678198,14.811904,14.14836,13.483003,12.817645,12.152288,11.486931,10.46442,9.441909,8.419398,7.3968873,6.3743763,7.112252,7.850128,8.588004,9.325879,10.061942,10.665659,11.267563,11.869466,12.473183,13.075087,11.940171,10.805257,9.670342,8.535428,7.400513,8.432089,9.465478,10.497053,11.530442,12.562017,10.872336,9.182655,7.4929743,5.803293,4.1117992,6.200332,8.287052,10.375585,12.462305,14.549025,13.274512,11.999999,10.725487,9.449161,8.174648,7.217404,6.26016,5.3029156,4.345671,3.386614,2.810092,2.231757,1.6552348,1.0768998,0.50037766,0.43692398,0.37528324,0.31182957,0.25018883,0.18673515,0.15954071,0.13234627,0.10515183,0.07795739,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,2.4329958,4.8641787,7.2971745,9.73017,12.163166,14.454751,16.748148,19.039734,21.33313,23.624716,21.427404,19.230095,17.032784,14.835473,12.638163,12.005438,11.372714,10.73999,10.107266,9.474543,8.439341,7.404139,6.3707504,5.335549,4.3003473,3.6658103,3.0294604,2.3949237,1.7603867,1.1258497,1.0823387,1.0406405,0.99712944,0.9554313,0.9119202,0.774135,0.63816285,0.50037766,0.36259252,0.22480737,0.22480737,0.22480737,0.22480737,0.22480737,0.22480737,0.1794833,0.13415924,0.09064813,0.045324065,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.06707962,0.059827764,0.052575916,0.045324065,0.038072214,0.04169814,0.047137026,0.052575916,0.058014803,0.06164073,0.13778515,0.21211663,0.28826106,0.36259252,0.43692398,0.36984438,0.30276474,0.23568514,0.16679256,0.099712946,0.16316663,0.22480737,0.28826106,0.34990177,0.41335547,0.7868258,1.162109,1.5373923,1.9126755,2.2879589,2.0558996,1.8220274,1.5899682,1.357909,1.1258497,1.0805258,1.0352017,0.9898776,0.9445535,0.89922947,2.0975976,3.294153,4.4925213,5.6908894,6.887445,5.52591,4.162562,2.7992141,1.4376793,0.07433146,1.1403534,2.2045624,3.2705846,4.3347936,5.4008155,6.16226,6.925517,7.686961,8.450218,9.211663,8.557183,7.902704,7.2482243,6.591932,5.9374523,5.8866897,5.8377395,5.7869763,5.7380266,5.6872635,5.4479527,5.2068286,4.9675174,4.7282066,4.4870825,6.1731377,7.85738,9.543435,11.227677,12.91192,11.691795,10.471672,9.253361,8.033237,6.813113,5.7833505,4.751775,3.7220123,2.6922495,1.6624867,2.3604772,3.056655,3.7546456,4.4526362,5.1506267,8.116633,11.084454,14.052273,17.020092,19.987913,19.730473,19.473032,19.21559,18.958149,18.700708,16.672005,14.645112,12.618219,10.589515,8.562622,8.145641,7.7268467,7.309865,6.892884,6.474089,6.0444174,5.614745,5.185073,4.7554007,4.325729,4.3021603,4.2804046,4.256836,4.2350807,4.213325,4.804351,5.3971896,5.9900284,6.582867,7.175706,7.0977483,7.019791,6.9418335,6.8656893,6.787732,7.1974616,7.607191,8.01692,8.42665,8.838193,9.7483,10.656594,11.566701,12.476809,13.386916,11.764315,10.141713,8.519112,6.8983226,5.275721,5.0200934,4.764466,4.510651,4.255023,3.9993954,5.910258,7.819308,9.73017,11.63922,13.550082,13.486629,13.424988,13.363347,13.299893,13.238253,12.097899,10.957546,9.817192,8.676839,7.5382986,7.743163,7.948028,8.152893,8.357758,8.562622,7.304426,6.0480433,4.7898474,3.531651,2.275268,2.6505513,3.0258346,3.3993049,3.774588,4.1498713,5.0980506,6.0444174,6.9925966,7.9407763,8.887142,9.52168,10.15803,10.792566,11.427103,12.06164,11.853149,11.642846,11.432542,11.222239,11.011934,10.9774885,10.943042,10.906783,10.872336,10.837891,11.039129,11.242181,11.445232,11.648285,11.849524,12.387974,12.92461,13.46306,13.999697,14.538147,14.188245,13.838344,13.486629,13.136727,12.786825,11.189605,9.592385,7.995165,6.397945,4.800725,5.0726695,5.3446136,5.618371,5.8903155,6.16226,6.827617,7.4929743,8.158332,8.821876,9.487233,10.292189,11.097144,11.9021,12.707055,13.512011,14.284332,15.056654,15.83079,16.603111,17.375433,15.528025,13.680615,11.833207,9.985798,8.138389,9.501737,10.866898,12.232059,13.597219,14.96238,12.864782,10.767185,8.669587,6.5719895,4.4743915,9.431031,14.384046,19.340685,24.295511,29.250338,25.381475,21.514427,17.647377,13.780329,9.91328,10.645717,11.378153,12.11059,12.843027,13.575464,10.912222,8.2507925,5.5875506,2.9243085,0.26287958,0.70524246,1.1476053,1.5899682,2.032331,2.474694,4.762653,7.0506115,9.336758,11.624716,13.912675,11.280253,8.647832,6.01541,3.3829882,0.7505665,0.73424983,0.7197462,0.70524246,0.69073874,0.6744221,1.2328146,1.789394,2.3477864,2.904366,3.4627585,2.956942,2.4529383,1.9471219,1.4431182,0.93730164,0.7505665,0.5620184,0.37528324,0.18673515,0.0,0.09789998,0.19579996,0.291887,0.38978696,0.48768693,0.42785916,0.3680314,0.30820364,0.24837588,0.18673515,0.4405499,0.69255173,0.9445535,1.1983683,1.4503701,1.6171626,1.7857682,1.9525607,2.1193533,2.2879589,2.817344,3.346729,3.877927,4.407312,4.936697,4.836984,4.7372713,4.6375585,4.537845,4.4381323,5.2557783,6.071612,6.889258,7.706904,8.52455,10.714609,12.904668,15.094727,17.284784,19.474844,21.247921,23.019186,24.792263,26.56534,28.336605,30.515787,32.693153,34.87052,37.04789,39.225258,37.852844,36.480434,35.10802,33.735607,32.363194,35.127964,37.89273,40.657497,43.422268,46.187035,43.824745,41.462456,39.100163,36.737873,34.375584,37.227375,40.079163,42.932766,45.784557,48.63816,49.55552,50.472878,51.390236,52.3076,53.224957,47.05726,40.889557,34.72186,28.554161,22.388275,20.29249,18.196705,16.102734,14.006948,11.912977,10.462607,9.012237,7.5618668,6.11331,4.6629395,4.070101,3.4772623,2.8844235,2.2933977,1.7005589,1.6280404,1.5555218,1.4830034,1.4104849,1.3379664,1.8274662,2.3169663,2.808279,3.2977788,3.787279,4.860553,5.9320135,7.0052876,8.076748,9.1500225,9.168152,9.184468,9.202598,9.220728,9.237044,9.712041,10.1870365,10.662033,11.137029,11.612025,11.731681,11.853149,11.972805,12.092461,12.212116,12.872034,13.531953,14.191871,14.851789,15.511708,16.989273,18.466837,19.9444,21.421967,22.89953,25.938055,28.974768,32.013294,35.050007,38.08672,38.31334,38.538147,38.762955,38.98776,39.212566,40.869614,42.526665,44.185524,45.84257,47.49962,48.244747,48.989876,49.735004,50.48013,51.225258,55.625317,60.02538,64.42544,68.8255,73.225555,73.198364,73.16936,73.142166,73.11497,73.087776,70.68741,68.28705,65.88669,63.488136,61.087772,55.61444,50.142918,44.669586,39.198063,33.72473,33.447346,33.169964,32.892582,32.615196,32.337814,29.957394,27.576973,25.198366,22.817947,20.437527,18.820364,17.203201,15.584227,13.967064,12.349901,11.755249,11.160598,10.564133,9.969481,9.374829,9.750113,10.125396,10.500679,10.874149,11.249433,11.543133,11.83502,12.126906,12.420607,12.712494,11.617464,10.522435,9.427405,8.3323765,7.2373466,8.05318,8.8672,9.683033,10.497053,11.312886,9.683033,8.05318,6.4233265,4.7934732,3.1618068,4.7118897,6.261973,7.8120556,9.362139,10.912222,10.263181,9.612328,8.963287,8.312433,7.663393,6.7605376,5.857682,4.954827,4.0519714,3.149116,2.6070402,2.0649643,1.5228885,0.9808127,0.43692398,0.42423326,0.41335547,0.40066472,0.387974,0.37528324,0.3208944,0.26469254,0.21030366,0.15410182,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,1.7803292,3.5606585,5.3391747,7.119504,8.899834,10.382836,11.86584,13.347031,14.830034,16.313038,14.960567,13.608097,12.255627,10.903157,9.550687,9.244296,8.939718,8.63514,8.330563,8.024173,7.509291,6.9944096,6.4795284,5.964647,5.4497657,4.6973863,3.9450066,3.1926272,2.4402475,1.6878681,1.4920682,1.2980812,1.1022812,0.90829426,0.7124943,0.63816285,0.5620184,0.48768693,0.41335547,0.33721104,0.2991388,0.26287958,0.22480737,0.18673515,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.045324065,0.03988518,0.034446288,0.030820364,0.025381476,0.032633327,0.03988518,0.047137026,0.054388877,0.06164073,0.12509441,0.18673515,0.25018883,0.31182957,0.37528324,0.31726846,0.25925365,0.2030518,0.14503701,0.0870222,0.12509441,0.16316663,0.19942589,0.2374981,0.2755703,0.8122072,1.3506571,1.887294,2.4257438,2.962381,2.5453994,2.126605,1.7096237,1.2926424,0.87566096,0.9318628,0.9898776,1.0478923,1.1040943,1.162109,1.8655385,2.5671551,3.2705846,3.972201,4.6756306,3.7618973,2.8499773,1.938057,1.0243238,0.11240368,1.3216497,2.5327086,3.7419548,4.953014,6.16226,6.9617763,7.763106,8.562622,9.362139,10.161655,9.104698,8.047741,6.9907837,5.9320135,4.8750563,4.699199,4.5251546,4.349297,4.175253,3.9993954,3.877927,3.7546456,3.633177,3.5098956,3.386614,5.2267714,7.066928,8.907085,10.747242,12.5873995,11.483305,10.377398,9.273304,8.167397,7.063302,5.904819,4.748149,3.589666,2.4329958,1.2745126,2.4021754,3.529838,4.6575007,5.7851634,6.9128265,9.333132,11.751623,14.171928,16.592234,19.012539,19.132195,19.25185,19.373318,19.492973,19.612629,17.364555,15.118295,12.870221,10.622148,8.375887,7.654328,6.9345818,6.2148356,5.4950895,4.7753434,4.41819,4.059223,3.7020695,3.3449159,2.9877625,2.9968271,3.007705,3.0167696,3.0276475,3.0367124,3.8199122,4.603112,5.384499,6.167699,6.9508986,6.889258,6.82943,6.7696023,6.7097745,6.6499467,6.7279043,6.8058615,6.882006,6.9599633,7.037921,8.551744,10.067381,11.583018,13.096842,14.612478,12.647227,10.681975,8.716724,6.7532854,4.788034,4.505212,4.2223897,3.9395678,3.6567454,3.3757362,5.090799,6.8058615,8.520925,10.234174,11.949236,11.775192,11.599335,11.42529,11.249433,11.075388,10.390089,9.704789,9.019489,8.334189,7.650702,7.9824743,8.314246,8.647832,8.979604,9.313189,8.007855,6.7025228,5.3971896,4.0918565,2.7883365,3.2252605,3.6621845,4.099108,4.537845,4.974769,5.714458,6.454147,7.1956487,7.935337,8.675026,9.052122,9.429218,9.808127,10.185224,10.56232,10.410031,10.257742,10.1054535,9.953164,9.800876,10.223296,10.645717,11.068136,11.490557,11.912977,12.047136,12.183108,12.317267,12.45324,12.5873995,13.037014,13.486629,13.938056,14.387671,14.837286,14.387671,13.938056,13.486629,13.037014,12.5873995,10.798005,9.006798,7.217404,5.42801,3.636803,4.3021603,4.9675174,5.632875,6.298232,6.9617763,7.0977483,7.231908,7.36788,7.502039,7.6380115,8.020547,8.403082,8.785617,9.168152,9.550687,12.077957,14.6052265,17.132496,19.659767,22.187037,19.909956,17.632874,15.355793,13.0769,10.799818,10.634838,10.469859,10.304879,10.139899,9.97492,8.597069,7.219217,5.8431783,4.465327,3.0874753,6.6336303,10.177972,13.722314,17.268469,20.81281,17.97915,15.147303,12.3154545,9.481794,6.6499467,7.130382,7.610817,8.089439,8.569874,9.050309,7.311678,5.57486,3.8380418,2.0994108,0.36259252,0.7197462,1.0768998,1.4358664,1.79302,2.1501737,3.5751622,5.0001507,6.4251394,7.850128,9.275117,7.520169,5.765221,4.0102735,2.2553256,0.50037766,0.4894999,0.48043507,0.46955732,0.4604925,0.44961473,1.0932164,1.7350051,2.3767939,3.0203958,3.6621845,3.054842,2.4474995,1.840157,1.2328146,0.62547207,0.50037766,0.37528324,0.25018883,0.12509441,0.0,0.065266654,0.13053331,0.19579996,0.25925365,0.3245203,0.28463513,0.24474995,0.20486477,0.16497959,0.12509441,0.38434806,0.64541465,0.90466833,1.1657349,1.4249886,1.5319533,1.6407311,1.7476959,1.8546607,1.9616255,2.469255,2.9768846,3.484514,3.9921436,4.499773,4.4127507,4.325729,4.2368937,4.1498713,4.062849,4.5450974,5.027345,5.5095935,5.9918413,6.4759026,8.62245,10.770811,12.917358,15.065719,17.212267,18.378002,19.541924,20.707659,21.873394,23.037315,24.71068,26.38223,28.055595,29.727148,31.400513,31.297173,31.195646,31.092308,30.990782,30.887444,35.61021,40.332977,45.055748,49.7767,54.49947,51.100163,47.70086,44.29974,40.900436,37.499317,41.634686,45.770054,49.905422,54.04079,58.174343,58.31938,58.464417,58.609455,58.75449,58.89953,51.491764,44.08581,36.678047,29.27028,21.862516,19.607191,17.351866,15.0965395,12.843027,10.587702,9.275117,7.9625316,6.6499467,5.337362,4.024777,3.6041696,3.1853752,2.764768,2.3441606,1.9253663,1.8474089,1.7694515,1.693307,1.6153497,1.5373923,1.7966459,2.0577126,2.3169663,2.5780327,2.8372865,3.7020695,4.5668526,5.431636,6.298232,7.1630154,7.083245,7.0016613,6.921891,6.8421206,6.7623506,7.4258947,8.087626,8.749357,9.412902,10.074633,10.154404,10.234174,10.315757,10.395528,10.475298,10.701918,10.930351,11.156972,11.385405,11.612025,13.096842,14.581658,16.068287,17.553104,19.03792,21.824444,24.61278,27.399303,30.18764,32.974163,33.625015,34.27587,34.92491,35.575764,36.224804,37.967064,39.70932,41.45339,43.19565,44.937904,45.98036,47.02281,48.065266,49.107716,50.15017,53.93745,57.724728,61.51201,65.299286,69.08838,69.92778,70.76718,71.6084,72.4478,73.2872,71.71174,70.138084,68.56262,66.98715,65.41169,60.371655,55.33343,50.29158,45.25336,40.21332,39.277836,38.342346,37.406857,36.473183,35.537693,33.643147,31.746788,29.852242,27.957697,26.06315,23.492369,20.9234,18.352621,15.781839,13.212872,13.044266,12.877473,12.710681,12.542075,12.375282,12.387974,12.400664,12.413355,12.4242325,12.436923,12.420607,12.402477,12.384347,12.368031,12.349901,11.294757,10.239613,9.184468,8.129324,7.07418,7.6724577,8.270736,8.8672,9.465478,10.061942,8.491917,6.921891,5.351866,3.7818398,2.2118144,3.2252605,4.2368937,5.2503395,6.261973,7.2754188,7.250037,7.224656,7.1992745,7.175706,7.1503243,6.301858,5.4552045,4.606738,3.7600844,2.911618,2.4058013,1.8981718,1.3905423,0.88291276,0.37528324,0.41335547,0.44961473,0.48768693,0.52575916,0.5620184,0.48043507,0.39703882,0.3154555,0.23205921,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.07433146,0.07433146,0.07433146,0.07433146,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,1.1276628,2.2553256,3.3829882,4.510651,5.638314,6.3091097,6.981719,7.654328,8.326937,8.999546,8.491917,7.9842873,7.476658,6.969028,6.4632115,6.484967,6.506723,6.530291,6.552047,6.5756154,6.5792413,6.58468,6.590119,6.5955577,6.599184,5.730775,4.860553,3.9903307,3.1201086,2.2498865,1.9017978,1.5555218,1.2074331,0.85934424,0.51306844,0.50037766,0.48768693,0.4749962,0.46230546,0.44961473,0.37528324,0.2991388,0.22480737,0.15047589,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.02175555,0.01994259,0.018129626,0.014503701,0.012690738,0.02175555,0.032633327,0.04169814,0.052575916,0.06164073,0.11240368,0.16316663,0.21211663,0.26287958,0.31182957,0.26469254,0.21755551,0.17041849,0.12328146,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.13778515,0.8375887,1.5373923,2.2371957,2.9369993,3.636803,3.0348995,2.4329958,1.8292793,1.2273756,0.62547207,0.7850128,0.9445535,1.1059072,1.2654479,1.4249886,1.6316663,1.840157,2.0468347,2.2553256,2.4620032,1.9996977,1.5373923,1.0750868,0.61278135,0.15047589,1.504759,2.8608549,4.215138,5.569421,6.925517,7.763106,8.600695,9.438283,10.275872,11.111648,9.652213,8.192778,6.733343,5.272095,3.8126602,3.5117085,3.2125697,2.911618,2.612479,2.3133402,2.3079014,2.3024626,2.2970235,2.2915847,2.2879589,4.2822175,6.2782893,8.272549,10.266808,12.262879,11.273002,10.283124,9.293246,8.303369,7.311678,6.0281005,4.74271,3.4573197,2.1719291,0.8883517,2.4456866,4.0030212,5.560356,7.117691,8.675026,10.547816,12.420607,14.293397,16.164375,18.037165,18.53573,19.03248,19.529232,20.027798,20.52455,18.057108,15.589665,13.122223,10.654781,8.187339,7.1648283,6.1423173,5.1198063,4.0972953,3.0747845,2.7901495,2.5055144,2.2190661,1.9344311,1.649796,1.693307,1.7350051,1.7767034,1.8202144,1.8619126,2.8354735,3.8072214,4.780782,5.75253,6.7242785,6.68258,6.640882,6.5973706,6.5556726,6.5121617,6.258347,6.002719,5.7470913,5.4932766,5.237649,7.3570023,9.4781685,11.597522,13.716875,15.838041,13.53014,11.222239,8.914337,6.6082487,4.3003473,3.9903307,3.680314,3.3702974,3.0602808,2.7502642,4.269527,5.7906027,7.309865,8.829127,10.3502035,10.061942,9.775495,9.487233,9.200785,8.912524,8.682278,8.452031,8.221786,7.993352,7.763106,8.221786,8.682278,9.142771,9.603263,10.061942,8.709473,7.3570023,6.004532,4.652062,3.299592,3.7999697,4.3003473,4.800725,5.2992897,5.7996674,6.3326783,6.8656893,7.3968873,7.9298983,8.46291,8.582565,8.70222,8.821876,8.943344,9.063,8.966913,8.872639,8.778365,8.682278,8.588004,9.467291,10.346578,11.227677,12.106964,12.988064,13.055143,13.122223,13.189302,13.258195,13.325275,13.687867,14.05046,14.413053,14.775645,15.138238,14.587097,14.037769,13.486629,12.937301,12.387974,10.4045925,8.423024,6.439643,4.458075,2.474694,3.531651,4.590421,5.6473784,6.7043357,7.763106,7.36788,6.972654,6.5774283,6.1822023,5.7869763,5.7470913,5.7072062,5.667321,5.6274357,5.5875506,9.869768,14.151986,18.436016,22.718235,27.000452,24.291885,21.585133,18.876566,16.169813,13.46306,11.7679405,10.07282,8.3777,6.68258,4.98746,4.329355,3.673062,3.0149567,2.3568513,1.7005589,3.834416,5.9700856,8.105756,10.239613,12.375282,10.576823,8.780178,6.981719,5.185073,3.386614,3.6150475,3.8416677,4.070101,4.2967215,4.5251546,3.7129474,2.9007401,2.08672,1.2745126,0.46230546,0.73424983,1.0080072,1.2799516,1.551896,1.8256533,2.3876717,2.94969,3.5117085,4.07554,4.6375585,3.7600844,2.8826106,2.0051367,1.1276628,0.25018883,0.24474995,0.23931105,0.23568514,0.23024625,0.22480737,0.95180535,1.6806163,2.4076142,3.1346123,3.8616104,3.152742,2.4420607,1.7331922,1.0225109,0.31182957,0.25018883,0.18673515,0.12509441,0.06164073,0.0,0.032633327,0.065266654,0.09789998,0.13053331,0.16316663,0.14322405,0.12328146,0.10333887,0.08339628,0.06164073,0.32995918,0.5982776,0.86478317,1.1331016,1.3996071,1.4467441,1.4956942,1.5428312,1.5899682,1.6371052,2.1229792,2.6070402,3.092914,3.576975,4.062849,3.9867048,3.9123733,3.8380418,3.7618973,3.6875658,3.834416,3.9830787,4.1299286,4.2767787,4.4254417,6.530291,8.63514,10.73999,12.84484,14.94969,15.508082,16.064661,16.623055,17.179634,17.738026,18.905573,20.073122,21.24067,22.408218,23.575766,24.743313,25.909048,27.076595,28.244144,29.411692,36.09246,42.773228,49.45218,56.132946,62.8119,58.375584,53.93745,49.499317,45.063,40.624866,46.041996,51.45913,56.878075,62.295208,67.71234,67.08505,66.45777,65.83048,65.2032,64.57591,55.92627,47.28025,38.63242,29.984589,21.336756,18.92189,16.507025,14.092158,11.677292,9.262425,8.087626,6.9128265,5.7380266,4.5632267,3.386614,3.1400511,2.8916752,2.6451125,2.3967366,2.1501737,2.0667772,1.9851941,1.9017978,1.8202144,1.7368182,1.7676386,1.7966459,1.8274662,1.8582866,1.887294,2.5453994,3.2016919,3.8597972,4.517903,5.1741953,4.9983377,4.8206677,4.6429973,4.465327,4.2876563,5.137936,5.9882154,6.836682,7.686961,8.537241,8.577126,8.617011,8.656897,8.696781,8.736667,8.531802,8.326937,8.122072,7.9172077,7.7123427,9.2044115,10.698292,12.19036,13.682428,15.174497,17.712645,20.24898,22.787127,25.325274,27.861609,28.936695,30.011782,31.08687,32.161957,33.23704,35.06451,36.891975,38.71944,40.54691,42.374374,43.714153,45.055748,46.395527,47.735306,49.075085,52.24958,55.42408,58.60039,61.774887,64.94939,66.657196,68.365005,70.072815,71.780624,73.486626,72.73787,71.987305,71.23674,70.48798,69.73742,65.130684,60.52213,55.915394,51.308655,46.700104,45.108322,43.51473,41.922947,40.329353,38.73757,37.327087,35.918415,34.50793,33.097446,31.68696,28.164373,24.641787,21.119202,17.598429,14.075842,14.335095,14.594349,14.855415,15.114669,15.375735,15.025834,14.675932,14.324218,13.974316,13.6244135,13.29808,12.969934,12.6417885,12.3154545,11.9873085,10.97205,9.956791,8.943344,7.9280853,6.9128265,7.2917356,7.6724577,8.05318,8.432089,8.812811,7.3026133,5.7924156,4.2822175,2.7720199,1.261822,1.7368182,2.2118144,2.6868105,3.1618068,3.636803,4.2368937,4.836984,5.4370747,6.037165,6.637256,5.844991,5.0527267,4.2604623,3.4681973,2.6741197,2.2027495,1.7295663,1.258196,0.7850128,0.31182957,0.40066472,0.48768693,0.5747091,0.66173136,0.7505665,0.6399758,0.5293851,0.42060733,0.3100166,0.19942589,0.15954071,0.11965553,0.07977036,0.03988518,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.099712946,0.099712946,0.099712946,0.099712946,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06164073,0.12509441,0.18673515,0.25018883,0.31182957,0.25018883,0.18673515,0.12509441,0.06164073,0.0,0.4749962,0.9499924,1.4249886,1.8999848,2.374981,2.2371957,2.0994108,1.9616255,1.8256533,1.6878681,2.0250793,2.3622901,2.6995013,3.0367124,3.3757362,3.7256382,4.07554,4.4254417,4.7753434,5.125245,5.6491914,6.1749506,6.70071,7.224656,7.750415,6.7623506,5.774286,4.788034,3.7999697,2.811905,2.3133402,1.8129625,1.3125849,0.8122072,0.31182957,0.36259252,0.41335547,0.46230546,0.51306844,0.5620184,0.44961473,0.33721104,0.22480737,0.11240368,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.099712946,0.13778515,0.17585737,0.21211663,0.25018883,0.21211663,0.17585737,0.13778515,0.099712946,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.8629702,1.7241274,2.5870976,3.4500678,4.313038,3.5243993,2.7375734,1.9507477,1.162109,0.37528324,0.63816285,0.89922947,1.162109,1.4249886,1.6878681,1.3996071,1.1131591,0.824898,0.53663695,0.25018883,0.2374981,0.22480737,0.21211663,0.19942589,0.18673515,1.6878681,3.1871881,4.688321,6.187641,7.686961,8.562622,9.438283,10.312131,11.187792,12.06164,10.199727,8.337815,6.474089,4.612177,2.7502642,2.324218,1.8999848,1.4757515,1.0497054,0.62547207,0.73787576,0.85027945,0.96268314,1.0750868,1.1874905,3.3376641,5.487838,7.6380115,9.788185,11.938358,11.062697,10.1870365,9.313189,8.437528,7.5618668,6.149569,4.7372713,3.3249733,1.9126755,0.50037766,2.4873846,4.4743915,6.4632115,8.450218,10.437225,11.762501,13.087777,14.413053,15.738328,17.06179,17.937452,18.813112,19.68696,20.562622,21.438282,18.749659,16.062849,13.374225,10.687414,8.000604,6.6753283,5.3500524,4.024777,2.6995013,1.3742256,1.162109,0.9499924,0.73787576,0.52575916,0.31182957,0.387974,0.46230546,0.53663695,0.61278135,0.6871128,1.8492218,3.0131438,4.175253,5.337362,6.4994707,6.4759026,6.450521,6.4251394,6.399758,6.3743763,5.7869763,5.199577,4.612177,4.024777,3.437377,6.16226,8.887142,11.612025,14.336908,17.06179,14.413053,11.762501,9.11195,6.4632115,3.8126602,3.4754493,3.1382382,2.7992141,2.4620032,2.124792,3.4500678,4.7753434,6.1006193,7.4258947,8.749357,8.350506,7.949841,7.549176,7.1503243,6.7496595,6.9744673,7.1992745,7.4258947,7.650702,7.8755093,8.46291,9.050309,9.637709,10.225109,10.812509,9.412902,8.013294,6.6118746,5.2122674,3.8126602,4.3746786,4.936697,5.5005283,6.0625467,6.624565,6.9508986,7.2754188,7.5999393,7.9244595,8.2507925,8.113008,7.9752226,7.837437,7.699652,7.5618668,7.5256076,7.4875355,7.4494634,7.413204,7.3751316,8.713099,10.049252,11.3872175,12.725184,14.06315,14.06315,14.06315,14.06315,14.06315,14.06315,14.336908,14.612478,14.888049,15.161806,15.437376,14.788336,14.137483,13.486629,12.837588,12.186734,10.012992,7.837437,5.661882,3.48814,1.3125849,2.762955,4.213325,5.661882,7.112252,8.562622,7.6380115,6.7134004,5.7869763,4.8623657,3.9377546,3.4754493,3.0131438,2.5508385,2.08672,1.6244144,7.663393,13.700559,19.737724,25.774889,31.812054,28.675629,25.537392,22.399153,19.262728,16.124489,12.899229,9.675781,6.450521,3.2252605,0.0,0.06164073,0.12509441,0.18673515,0.25018883,0.31182957,1.0370146,1.7621996,2.4873846,3.2125697,3.9377546,3.1744974,2.4130533,1.649796,0.8883517,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.11240368,0.22480737,0.33721104,0.44961473,0.5620184,0.7505665,0.93730164,1.1258497,1.3125849,1.49932,1.2001812,0.89922947,0.6000906,0.2991388,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.8122072,1.6244144,2.4366217,3.2506418,4.062849,3.2506418,2.4366217,1.6244144,0.8122072,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.2755703,0.5493277,0.824898,1.1004683,1.3742256,1.3633479,1.3506571,1.3379664,1.3252757,1.3125849,1.7748904,2.2371957,2.6995013,3.1618068,3.6241121,3.5624714,3.5008307,3.437377,3.3757362,3.3122826,3.1255474,2.9369993,2.7502642,2.561716,2.374981,4.4381323,6.4994707,8.562622,10.625773,12.687112,12.638163,12.5873995,12.536636,12.487686,12.436923,13.100468,13.762199,14.425743,15.087475,15.749206,18.187641,20.624262,23.062696,25.49932,27.937754,36.574707,45.211662,53.850426,62.48738,71.12434,65.649185,60.175854,54.700706,49.22556,43.750412,50.451122,57.15002,63.85073,70.54963,77.250336,75.85073,74.44931,73.0497,71.65009,70.25049,60.36259,50.47469,40.586792,30.700708,20.81281,18.236591,15.662184,13.087777,10.511557,7.93715,6.9001355,5.863121,4.8242936,3.787279,2.7502642,2.6741197,2.5997884,2.525457,2.4493124,2.374981,2.2879589,2.1991236,2.1121013,2.0250793,1.938057,1.7368182,1.5373923,1.3379664,1.1367276,0.93730164,1.3869164,1.8383441,2.2879589,2.7375734,3.1871881,2.911618,2.6378605,2.3622901,2.08672,1.8129625,2.8499773,3.8869917,4.9258194,5.962834,6.9998484,6.9998484,6.9998484,6.9998484,6.9998484,6.9998484,6.3616858,5.7253356,5.087173,4.4508233,3.8126602,5.3119802,6.813113,8.312433,9.811753,11.312886,13.600845,15.8869915,18.17495,20.462908,22.750868,24.250187,25.749508,27.25064,28.74996,30.24928,32.161957,34.07463,35.98731,37.899982,39.812656,41.449764,43.08687,44.72579,46.362892,47.999996,50.563526,53.125244,55.68696,58.25049,60.812202,63.388424,65.96283,68.53724,71.11164,73.68787,73.7622,73.83834,73.912674,73.987,74.06315,69.88789,65.71264,61.537388,57.362137,53.186882,50.936996,48.68711,46.437225,44.187336,41.93745,41.01284,40.08823,39.161804,38.237194,37.312584,32.83638,28.361986,23.887594,19.413204,14.936998,15.625924,16.313038,17.00015,17.687263,18.374376,17.661882,16.949387,16.236893,15.524399,14.811904,14.175554,13.537392,12.899229,12.262879,11.624716,10.649343,9.675781,8.700407,7.7250338,6.7496595,6.9128265,7.07418,7.2373466,7.400513,7.5618668,6.11331,4.6629395,3.2125697,1.7621996,0.31182957,0.25018883,0.18673515,0.12509441,0.06164073,0.0,1.2255627,2.4493124,3.6748753,4.900438,6.1241875,5.388125,4.650249,3.9123733,3.1744974,2.4366217,1.9996977,1.5627737,1.1258497,0.6871128,0.25018883,0.387974,0.52575916,0.66173136,0.7995165,0.93730164,0.7995165,0.66173136,0.52575916,0.387974,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.38072214,0.75963134,1.1403534,1.5192627,1.8999848,2.3604772,2.819157,3.2796493,3.7401419,4.2006345,4.795286,5.389938,5.9845896,6.5792413,7.175706,6.717026,6.26016,5.803293,5.3446136,4.8877473,5.1596913,5.431636,5.7053933,5.977338,6.249282,5.8431783,5.4352617,5.027345,4.6194286,4.213325,3.437377,2.663242,1.887294,1.1131591,0.33721104,0.42967212,0.52213323,0.61459434,0.7070554,0.7995165,0.6417888,0.48587397,0.32814622,0.17041849,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.04169814,0.034446288,0.027194439,0.01994259,0.012690738,0.06164073,0.11240368,0.16316663,0.21211663,0.26287958,0.3825351,0.50219065,0.62184614,0.7433147,0.8629702,0.70524246,0.5475147,0.38978696,0.23205921,0.07433146,0.099712946,0.12509441,0.15047589,0.17585737,0.19942589,0.3100166,0.42060733,0.5293851,0.6399758,0.7505665,0.61822027,0.48587397,0.35171473,0.21936847,0.0870222,0.78319985,1.4775645,2.1719291,2.8681068,3.5624714,3.002266,2.4420607,1.8818551,1.3216497,0.76325727,0.9880646,1.2128719,1.4376793,1.6624867,1.887294,1.9217403,1.9579996,1.9924458,2.0268922,2.0631514,2.561716,3.0620937,3.5624714,4.062849,4.5632267,5.863121,7.1630154,8.46291,9.762803,11.062697,10.832452,10.602205,10.371959,10.141713,9.91328,8.568061,7.2228427,5.8776245,4.5324063,3.1871881,2.6523643,2.1175404,1.5827163,1.0478923,0.51306844,0.60190356,0.69255173,0.78319985,0.872035,0.96268314,2.6868105,4.4127507,6.1368785,7.8628187,9.5869465,8.917963,8.247167,7.5781837,6.9073873,6.2365913,5.1143675,3.9921436,2.8699198,1.7476959,0.62547207,2.2897718,3.9540713,5.620184,7.2844834,8.950596,10.098202,11.245807,12.3916,13.539205,14.68681,15.459132,16.233267,17.005589,17.77791,18.550234,16.34567,14.139296,11.934732,9.73017,7.5256076,6.354434,5.185073,4.0157123,2.8445382,1.6751775,1.5446441,1.4141108,1.2853905,1.1548572,1.0243238,1.1004683,1.1747998,1.2491312,1.3252757,1.3996071,2.1592383,2.9206827,3.680314,4.439945,5.199577,5.18326,5.1651306,5.147001,5.130684,5.1125546,4.6429973,4.171627,3.7020695,3.2325122,2.762955,4.942136,7.12313,9.302311,11.483305,13.662486,11.5503845,9.438283,7.324369,5.2122674,3.100166,2.8499773,2.5997884,2.3495996,2.0994108,1.8492218,2.907992,3.9649491,5.0219064,6.0806766,7.137634,6.796797,6.4577727,6.1169357,5.7779117,5.4370747,5.638314,5.8377395,6.037165,6.2365913,6.43783,7.2355337,8.033237,8.829127,9.626831,10.424535,9.242483,8.0604315,6.876567,5.6945157,4.512464,4.9095025,5.3083544,5.7053933,6.1024323,6.4994707,6.53573,6.5701766,6.604623,6.639069,6.6753283,6.644508,6.6155005,6.58468,6.5556726,6.5248523,6.414262,6.305484,6.1948934,6.0843024,5.975525,7.230095,8.484665,9.739235,10.995618,12.250188,12.130532,12.009064,11.889409,11.769753,11.650098,11.949236,12.250188,12.549327,12.850279,13.149418,12.565643,11.980057,11.39447,10.810696,10.225109,8.417585,6.6100616,4.802538,2.9950142,1.1874905,2.4003625,3.6132345,4.8242936,6.037165,7.250037,6.836682,6.4251394,6.011784,5.600241,5.186886,4.95664,4.7282066,4.49796,4.267714,4.0374675,8.560809,13.082338,17.60568,22.127209,26.65055,23.900286,21.15002,18.399757,15.649493,12.899229,10.319383,7.7395372,5.1596913,2.5798457,0.0,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,0.83033687,1.4104849,1.9906329,2.570781,3.149116,2.5399606,1.9308052,1.3198367,0.7106813,0.099712946,0.0870222,0.07433146,0.06164073,0.05076295,0.038072214,0.11965553,0.2030518,0.28463513,0.3680314,0.44961473,0.6000906,0.7505665,0.89922947,1.0497054,1.2001812,0.9644961,0.7306239,0.4949388,0.25925365,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.6653573,1.3180238,1.9706904,2.6233568,3.2742105,2.619731,1.9652514,1.310772,0.6544795,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.21936847,0.4405499,0.65991837,0.8792868,1.1004683,1.0895905,1.0805258,1.0696479,1.0605831,1.0497054,1.502946,1.9543737,2.4076142,2.8608549,3.3122826,3.2270734,3.141864,3.056655,2.9732587,2.8880494,2.7031271,2.518205,2.333283,2.1483607,1.9616255,3.6059825,5.2467136,6.889258,8.531802,10.174346,10.462607,10.749055,11.037316,11.325577,11.612025,13.189302,14.766581,16.34567,17.922949,19.500225,22.627586,25.754946,28.882307,32.009666,35.137028,41.680008,48.222992,54.765972,61.307144,67.85013,63.23432,58.62033,54.004528,49.39054,44.77474,52.933067,61.08959,69.24792,77.404434,85.56277,81.71022,77.85768,74.005135,70.15259,66.30004,56.602505,46.90497,37.20743,27.509893,17.812357,15.683939,13.557334,11.430729,9.302311,7.175706,6.1803894,5.185073,4.1897564,3.1944401,2.1991236,2.1392958,2.079468,2.0196402,1.9598125,1.8999848,1.8329052,1.7658255,1.696933,1.6298534,1.5627737,1.5754645,1.5881553,1.6008459,1.6117238,1.6244144,2.039583,2.4547513,2.8699198,3.2850883,3.7002566,3.5497808,3.3993049,3.2506418,3.100166,2.94969,3.7256382,4.499773,5.275721,6.049856,6.825804,6.8058615,6.784106,6.7641635,6.7442207,6.7242785,6.2873545,5.8504305,5.411693,4.974769,4.537845,5.8377395,7.137634,8.437528,9.737422,11.037316,12.810393,14.581658,16.354736,18.127813,19.899076,21.374828,22.85058,24.324518,25.80027,27.27421,28.936695,30.599182,32.26167,33.924156,35.586643,36.93186,38.27708,39.622295,40.967514,42.312733,44.30518,46.297626,48.29007,50.282516,52.274963,54.465023,56.65508,58.84514,61.0352,63.225258,64.590416,65.95558,67.32074,68.68409,70.04925,66.93276,63.81447,60.697987,57.579693,54.463207,53.587547,52.711887,51.83804,50.96238,50.08853,48.152287,46.217854,44.283424,42.34718,40.41275,36.152287,31.891825,27.633175,23.372713,19.112251,20.366821,21.623205,22.877775,24.132345,25.386915,23.33464,21.282368,19.230095,17.17782,15.125546,14.5508375,13.974316,13.399607,12.824898,12.250188,11.057259,9.864329,8.673213,7.4802837,6.2873545,6.4070096,6.526665,6.6481338,6.7677894,6.887445,5.8304877,4.7717175,3.7147603,2.657803,1.6008459,1.5392052,1.4793775,1.4195497,1.3597219,1.2998942,2.2879589,3.2760234,4.262275,5.2503395,6.2384043,5.567608,4.896812,4.227829,3.5570326,2.8880494,2.3532255,1.8165885,1.2817645,0.7469406,0.21211663,0.3208944,0.42785916,0.53482395,0.6417888,0.7505665,0.72337204,0.69436467,0.6671702,0.6399758,0.61278135,0.83940166,1.067835,1.2944553,1.5228885,1.7495089,1.938057,2.124792,2.3133402,2.5000753,2.6868105,2.324218,1.9616255,1.6008459,1.2382535,0.87566096,0.7179332,0.56020546,0.40247768,0.24474995,0.0870222,0.07070554,0.052575916,0.034446288,0.018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.28463513,0.56927025,0.8557183,1.1403534,1.4249886,2.4819458,3.540716,4.597673,5.65463,6.7134004,7.5654926,8.417585,9.269678,10.12177,10.975676,9.710228,8.444779,7.179332,5.915697,4.650249,4.670192,4.690134,4.710077,4.7300196,4.749962,4.9221935,5.0944247,5.2666564,5.4407005,5.612932,4.5632267,3.5117085,2.4620032,1.4122978,0.36259252,0.49675176,0.6327239,0.7668832,0.90285534,1.0370146,0.83577573,0.6327239,0.42967212,0.22662032,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.034446288,0.032633327,0.030820364,0.027194439,0.025381476,0.12509441,0.22480737,0.3245203,0.42423326,0.52575916,0.7650702,1.0043813,1.2455053,1.4848163,1.7241274,1.3977941,1.0696479,0.7433147,0.41516843,0.0870222,0.099712946,0.11240368,0.12509441,0.13778515,0.15047589,0.40791658,0.6653573,0.922798,1.1802386,1.4376793,1.1856775,0.9318628,0.67986095,0.42785916,0.17585737,0.7016165,1.2291887,1.7567607,2.2843328,2.811905,2.4801328,2.1483607,1.8147756,1.4830034,1.1494182,1.3379664,1.5247015,1.7132497,1.8999848,2.08672,2.4456866,2.8028402,3.159994,3.5171473,3.874301,4.8877473,5.89938,6.9128265,7.9244595,8.937905,10.038374,11.137029,12.237497,13.337966,14.436621,13.102281,11.7679405,10.431787,9.097446,7.763106,6.9345818,6.107871,5.279347,4.4526362,3.6241121,2.9805105,2.335096,1.6896812,1.0442665,0.40066472,0.46774435,0.53482395,0.60190356,0.67079616,0.73787576,2.03777,3.3376641,4.6375585,5.9374523,7.2373466,6.773228,6.3072968,5.8431783,5.377247,4.9131284,4.079166,3.247016,2.4148662,1.5827163,0.7505665,2.0921588,3.435564,4.7771564,6.1205616,7.462154,8.432089,9.402024,10.371959,11.341894,12.311829,12.982625,13.651608,14.322405,14.9932,15.662184,13.939869,12.217555,10.49524,8.772926,7.0506115,6.035352,5.0200934,4.004834,2.9895754,1.9743162,1.9271792,1.8800422,1.8329052,1.7857682,1.7368182,1.8129625,1.887294,1.9616255,2.03777,2.1121013,2.469255,2.8282216,3.1853752,3.5425289,3.8996825,3.8906176,3.87974,3.870675,3.8597972,3.8507326,3.4972048,3.1454902,2.7919624,2.4402475,2.08672,3.7220123,5.3573046,6.9925966,8.627889,10.263181,8.6877165,7.112252,5.5367875,3.9631362,2.3876717,2.2245052,2.0631514,1.8999848,1.7368182,1.5754645,2.3641033,3.1545548,3.9450066,4.7354584,5.524097,5.2449007,4.9657044,4.6846952,4.405499,4.12449,4.3003473,4.4743915,4.650249,4.8242936,5.0001507,6.008158,7.0143523,8.02236,9.030367,10.038374,9.072064,8.107569,7.1430726,6.1767635,5.2122674,5.4443264,5.678199,5.910258,6.1423173,6.3743763,6.1205616,5.864934,5.6093063,5.3554916,5.0998635,5.177821,5.2557783,5.331923,5.40988,5.487838,5.3047285,5.121619,4.940323,4.7572136,4.574105,5.7470913,6.9200783,8.093065,9.264238,10.437225,10.197914,9.956791,9.71748,9.4781685,9.237044,9.563377,9.8878975,10.212419,10.536939,10.863272,10.342952,9.822631,9.302311,8.781991,8.26167,6.8221784,5.382686,3.9431937,2.5018883,1.062396,2.03777,3.0131438,3.9867048,4.9620786,5.9374523,6.037165,6.1368785,6.2384043,6.338117,6.43783,6.439643,6.4432693,6.445082,6.446895,6.450521,9.458226,12.464118,15.471823,18.479528,21.487232,19.124943,16.762651,14.400362,12.038072,9.675781,7.7395372,5.805106,3.870675,1.9344311,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.62184614,1.0569572,1.4920682,1.9271792,2.3622901,1.9054236,1.4467441,0.9898776,0.533011,0.07433146,0.07433146,0.07433146,0.07433146,0.07433146,0.07433146,0.12690738,0.1794833,0.23205921,0.28463513,0.33721104,0.44961473,0.5620184,0.6744221,0.7868258,0.89922947,0.7306239,0.56020546,0.38978696,0.21936847,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.5166943,1.0098201,1.502946,1.9942589,2.4873846,1.9906329,1.4920682,0.99531645,0.49675176,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.16497959,0.32995918,0.4949388,0.65991837,0.824898,0.81764615,0.8103943,0.8031424,0.79589057,0.7868258,1.2291887,1.6733645,2.1157274,2.5580902,3.000453,2.8916752,2.7847104,2.6777458,2.570781,2.4620032,2.280707,2.0975976,1.9144884,1.7331922,1.550083,2.7720199,3.9957695,5.217706,6.439643,7.66158,8.287052,8.912524,9.537996,10.161655,10.7871275,13.279951,15.772775,18.265598,20.75842,23.249432,27.067532,30.88563,34.701916,38.520016,42.338116,46.785313,51.23251,55.679707,60.126904,64.574104,60.819454,57.06481,53.310165,49.55552,45.800873,55.415016,65.02915,74.64511,84.26106,93.875206,87.56972,81.266045,74.96056,68.65508,62.349598,52.84242,43.335243,33.828068,24.31908,14.811904,13.1331005,11.452485,9.771869,8.093065,6.412449,5.4606433,4.507025,3.5552197,2.6016014,1.649796,1.6044719,1.5591478,1.5156367,1.4703126,1.4249886,1.3778516,1.3307146,1.2817645,1.2346275,1.1874905,1.4122978,1.6371052,1.8619126,2.08672,2.3133402,2.6922495,3.0729716,3.4518807,3.832603,4.213325,4.1879435,4.162562,4.137181,4.1117992,4.0882306,4.599486,5.1125546,5.6256227,6.1368785,6.6499467,6.6100616,6.5701766,6.530291,6.490406,6.450521,6.2130227,5.975525,5.7380266,5.5005283,5.2630305,6.3616858,7.462154,8.562622,9.663091,10.761745,12.019942,13.278138,14.534521,15.792717,17.0491,18.49947,19.94984,21.40021,22.85058,24.299137,25.71325,27.125546,28.537844,29.950142,31.36244,32.41577,33.46729,34.520622,35.57214,36.62547,38.046833,39.47001,40.893185,42.31455,43.73772,45.543434,47.347332,49.15304,50.95694,52.76265,55.41683,58.07282,60.726994,63.382984,66.03716,63.97764,61.91811,59.856773,57.79725,55.73772,56.2381,56.736664,57.23704,57.73742,58.237797,55.291733,52.34748,49.40323,46.457165,43.512917,39.46638,35.423477,31.376944,27.332224,23.287504,25.109531,26.933372,28.7554,30.577427,32.399456,29.0074,25.615349,22.223295,18.82943,15.437376,14.924308,14.413053,13.899984,13.386916,12.87566,11.465176,10.05469,8.644206,7.2355337,5.825049,5.903006,5.979151,6.057108,6.1350656,6.2130227,5.5476656,4.882308,4.216951,3.5534067,2.8880494,2.8300345,2.7720199,2.715818,2.657803,2.5997884,3.350355,4.100921,4.8496747,5.600241,6.350808,5.7470913,5.145188,4.5432844,3.9395678,3.3376641,2.70494,2.0722163,1.4394923,0.80676836,0.17585737,0.2520018,0.32995918,0.40791658,0.48587397,0.5620184,0.64541465,0.726998,0.8103943,0.8919776,0.97537386,1.4793775,1.9851941,2.4891977,2.9950142,3.5008307,3.8507326,4.2006345,4.550536,4.900438,5.2503395,4.5251546,3.7999697,3.0747845,2.3495996,1.6244144,1.3343405,1.0442665,0.7541924,0.46411842,0.17585737,0.13959812,0.10515183,0.07070554,0.034446288,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.19036107,0.38072214,0.56927025,0.75963134,0.9499924,2.6052272,4.2604623,5.915697,7.569119,9.224354,10.3357,11.445232,12.554766,13.664299,14.775645,12.701616,10.629399,8.557183,6.484967,4.4127507,4.1806917,3.9468195,3.7147603,3.482701,3.2506418,4.0030212,4.7554007,5.5077806,6.26016,7.0125394,5.6872635,4.361988,3.0367124,1.7132497,0.387974,0.5656443,0.7433147,0.91917205,1.0968424,1.2745126,1.0279498,0.7795739,0.533011,0.28463513,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.027194439,0.030820364,0.032633327,0.034446288,0.038072214,0.18673515,0.33721104,0.48768693,0.63816285,0.7868258,1.1476053,1.5083848,1.8673514,2.228131,2.5870976,2.0903459,1.5917811,1.0950294,0.5982776,0.099712946,0.099712946,0.099712946,0.099712946,0.099712946,0.099712946,0.5058166,0.9101072,1.3143979,1.7205015,2.124792,1.7531348,1.3796645,1.0080072,0.6345369,0.26287958,0.62184614,0.9826257,1.3434052,1.7023718,2.0631514,1.9579996,1.8528478,1.7476959,1.6425442,1.5373923,1.6878681,1.8383441,1.987007,2.137483,2.2879589,2.9678197,3.6476808,4.327542,5.0074024,5.6872635,7.211965,8.736667,10.263181,11.787883,13.312584,14.211814,15.112856,16.012085,16.913128,17.812357,15.372109,12.931862,10.491614,8.05318,5.612932,5.3029156,4.992899,4.6828823,4.3728657,4.062849,3.3068438,2.5526514,1.7966459,1.0424535,0.28826106,0.33177215,0.3770962,0.4224203,0.46774435,0.51306844,1.3869164,2.2625773,3.1382382,4.0120864,4.8877473,4.6266804,4.367427,4.1081734,3.8471067,3.587853,3.045777,2.5018883,1.9598125,1.4177368,0.87566096,1.8945459,2.9152439,3.9359417,4.954827,5.975525,6.7677894,7.560054,8.352319,9.144584,9.936848,10.504305,11.071762,11.63922,12.206677,12.774135,11.535881,10.2958145,9.055748,7.8156815,6.5756154,5.714458,4.855114,3.9957695,3.1346123,2.275268,2.3097143,2.3441606,2.38042,2.4148662,2.4493124,2.525457,2.5997884,2.6741197,2.7502642,2.8245957,2.7792716,2.7357605,2.6904364,2.6451125,2.5997884,2.5979755,2.5943494,2.5925364,2.5907235,2.5870976,2.3532255,2.1175404,1.8818551,1.647983,1.4122978,2.5018883,3.5932918,4.6828823,5.772473,6.8620634,5.825049,4.788034,3.7492065,2.712192,1.6751775,1.6008459,1.5247015,1.4503701,1.3742256,1.2998942,1.8220274,2.3441606,2.8681068,3.39024,3.9123733,3.6930048,3.4718235,3.2524548,3.0330863,2.811905,2.962381,3.1128569,3.2633326,3.4119956,3.5624714,4.780782,5.99728,7.215591,8.432089,9.6504,8.901647,8.154706,7.407765,6.6608243,5.9120708,5.979151,6.0480433,6.115123,6.1822023,6.249282,5.7053933,5.1596913,4.615803,4.070101,3.5243993,3.7093215,3.8942437,4.079166,4.265901,4.4508233,4.195195,3.9395678,3.6857529,3.4301252,3.1744974,4.265901,5.3554916,6.445082,7.5346723,8.624263,8.265296,7.9045167,7.5455503,7.1847706,6.825804,7.175706,7.5256076,7.8755093,8.225411,8.575313,8.120259,7.665206,7.210152,6.755099,6.300045,5.2267714,4.15531,3.0820365,2.0105755,0.93730164,1.6751775,2.4130533,3.150929,3.8869917,4.6248674,5.237649,5.8504305,6.4632115,7.07418,7.686961,7.9226465,8.158332,8.392203,8.627889,8.861761,10.355642,11.847711,13.339779,14.831847,16.325727,14.349599,12.375282,10.399154,8.424837,6.450521,5.1596913,3.870675,2.5798457,1.2908293,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.41516843,0.70524246,0.99531645,1.2853905,1.5754645,1.2708868,0.9644961,0.65991837,0.35534066,0.05076295,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.13415924,0.15772775,0.1794833,0.2030518,0.22480737,0.2991388,0.37528324,0.44961473,0.52575916,0.6000906,0.4949388,0.38978696,0.28463513,0.1794833,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.36984438,0.7016165,1.0352017,1.3669738,1.7005589,1.3597219,1.020698,0.67986095,0.34083697,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.11059072,0.21936847,0.32995918,0.4405499,0.5493277,0.54570174,0.5402629,0.53482395,0.5293851,0.52575916,0.9572442,1.3905423,1.8220274,2.2553256,2.6868105,2.5580902,2.427557,2.2970235,2.1683033,2.03777,1.8582866,1.6769904,1.4975071,1.3180238,1.1367276,1.93987,2.7430124,3.5443418,4.347484,5.1506267,6.11331,7.07418,8.036863,8.999546,9.96223,13.370599,16.777155,20.185526,23.592083,27.000452,31.507477,36.014503,40.52334,45.030365,49.537388,51.890614,54.242027,56.595253,58.946667,61.299892,58.40459,55.50929,52.6158,49.720497,46.8252,57.898773,68.970535,80.0423,91.115875,102.18764,93.429214,84.67261,75.914185,67.15757,58.39915,49.082336,39.765522,30.446894,21.13008,11.813264,10.58045,9.347635,8.1148205,6.882006,5.6491914,4.7390842,3.83079,2.9206827,2.0105755,1.1004683,1.0696479,1.0406405,1.0098201,0.9808127,0.9499924,0.922798,0.89560354,0.8665961,0.83940166,0.8122072,1.2491312,1.6878681,2.124792,2.561716,3.000453,3.3449159,3.6893787,4.0356545,4.3801174,4.7245803,4.8242936,4.9258194,5.0255322,5.125245,5.224958,5.475147,5.7253356,5.975525,6.2257137,6.4759026,6.414262,6.354434,6.294606,6.2347784,6.1749506,6.1368785,6.1006193,6.0625467,6.0244746,5.9882154,6.887445,7.7866745,8.6877165,9.5869465,10.487988,11.22949,11.972805,12.714307,13.457622,14.199123,15.625924,17.0491,18.475903,19.90089,21.325878,22.487988,23.650097,24.812206,25.974316,27.138237,27.89787,28.6575,29.417131,30.176762,30.938206,31.790298,32.64239,33.494484,34.34839,35.20048,36.62003,38.03958,39.460945,40.880493,42.30004,46.24505,50.190056,54.135063,58.08007,62.025074,61.022507,60.01994,59.017372,58.0148,57.012234,58.886837,60.763252,62.637856,64.51246,66.38706,62.43299,58.477108,54.523037,50.567154,46.61308,42.78229,38.953316,35.122524,31.293547,27.462757,29.852242,32.241726,34.633022,37.02251,39.411995,34.68016,29.948328,25.214684,20.482851,15.749206,15.299591,14.849977,14.400362,13.9507475,13.499319,11.873092,10.245051,8.617011,6.9907837,5.3627434,5.3971896,5.431636,5.467895,5.5023413,5.5367875,5.2648435,4.992899,4.7191415,4.4471974,4.175253,4.120864,4.064662,4.0102735,3.9558845,3.8996825,4.4127507,4.9258194,5.4370747,5.9501433,6.4632115,5.9265747,5.391751,4.856927,4.322103,3.787279,3.056655,2.327844,1.5972201,0.8684091,0.13778515,0.18492219,0.23205921,0.27919623,0.32814622,0.37528324,0.56745726,0.75963134,0.95180535,1.1457924,1.3379664,2.1193533,2.902553,3.6857529,4.4671397,5.2503395,5.763408,6.2746634,6.787732,7.3008003,7.8120556,6.7242785,5.636501,4.550536,3.4627585,2.374981,1.9525607,1.5301404,1.1077201,0.6852999,0.26287958,0.21030366,0.15772775,0.10515183,0.052575916,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.09427405,0.19036107,0.28463513,0.38072214,0.4749962,2.7266958,4.9802084,7.231908,9.48542,11.73712,13.1059065,14.47288,15.839854,17.206827,18.575615,15.694818,12.815832,9.935035,7.0542374,4.175253,3.6893787,3.2053177,2.7194438,2.2353828,1.7495089,3.0820365,4.4145637,5.7470913,7.079619,8.412147,6.813113,5.2122674,3.6132345,2.0123885,0.41335547,0.6327239,0.8520924,1.0732739,1.2926424,1.5120108,1.2201238,0.92823684,0.6345369,0.34264994,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.01994259,0.027194439,0.034446288,0.04169814,0.05076295,0.25018883,0.44961473,0.6508536,0.85027945,1.0497054,1.5301404,2.0105755,2.4891977,2.9696326,3.4500678,2.7828975,2.1157274,1.4467441,0.7795739,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.05076295,0.60190356,1.1548572,1.7078108,2.2607644,2.811905,2.3205922,1.8274662,1.3343405,0.8430276,0.34990177,0.5420758,0.73424983,0.92823684,1.1204109,1.3125849,1.4358664,1.5573349,1.6806163,1.8020848,1.9253663,2.03777,2.1501737,2.2625773,2.374981,2.4873846,3.489953,4.4925213,5.4950895,6.497658,7.500226,9.537996,11.575767,13.611723,15.649493,17.687263,18.387066,19.08687,19.786674,20.48829,21.188093,17.64194,14.097597,10.553255,7.0071006,3.4627585,3.6694362,3.877927,4.0846047,4.2930956,4.499773,3.63499,2.770207,1.9054236,1.0406405,0.17585737,0.19761293,0.21936847,0.24293698,0.26469254,0.28826106,0.73787576,1.1874905,1.6371052,2.08672,2.5381477,2.4819458,2.427557,2.373168,2.3169663,2.2625773,2.0105755,1.7567607,1.504759,1.2527572,1.0007553,1.696933,2.3949237,3.092914,3.7890918,4.4870825,5.101677,5.718084,6.3326783,6.947273,7.5618668,8.027799,8.491917,8.957849,9.421967,9.8878975,9.130079,8.372261,7.614443,6.8566246,6.1006193,5.3953767,4.690134,3.9848917,3.2796493,2.5744069,2.6922495,2.810092,2.9279346,3.045777,3.1618068,3.2379513,3.3122826,3.386614,3.4627585,3.53709,3.0892882,2.6432993,2.1954978,1.7476959,1.2998942,1.305333,1.310772,1.3143979,1.3198367,1.3252757,1.2074331,1.0895905,0.97174793,0.8557183,0.73787576,1.2817645,1.8274662,2.373168,2.9170568,3.4627585,2.962381,2.4620032,1.9616255,1.4630609,0.96268314,0.97537386,0.9880646,1.0007553,1.0116332,1.0243238,1.2799516,1.5355793,1.789394,2.0450218,2.3006494,2.1392958,1.9797552,1.8202144,1.6606737,1.49932,1.6244144,1.7495089,1.8746033,1.9996977,2.124792,3.5515938,4.9802084,6.4070096,7.835624,9.262425,8.733041,8.201842,7.6724577,7.1430726,6.6118746,6.5157876,6.4178877,6.319988,6.2220874,6.1241875,5.290225,4.454449,3.6204863,2.7847104,1.9507477,2.2426348,2.5345216,2.8282216,3.1201086,3.4119956,3.0856624,2.7575161,2.42937,2.1030366,1.7748904,2.7828975,3.7890918,4.797099,5.805106,6.813113,6.3326783,5.8522434,5.371808,4.893186,4.4127507,4.788034,5.163317,5.5367875,5.9120708,6.2873545,5.8975673,5.5077806,5.1179934,4.7282066,4.3366065,3.633177,2.9279346,2.222692,1.5174497,0.8122072,1.3125849,1.8129625,2.3133402,2.811905,3.3122826,4.4381323,5.562169,6.688019,7.8120556,8.937905,9.40565,9.873394,10.339326,10.80707,11.274815,11.253058,11.22949,11.207735,11.184166,11.162411,9.574255,7.987913,6.399758,4.8116026,3.2252605,2.5798457,1.9344311,1.2908293,0.64541465,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.20667773,0.35171473,0.49675176,0.6417888,0.7868258,0.6345369,0.48224804,0.32995918,0.17767033,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.15047589,0.14322405,0.13415924,0.12690738,0.11965553,0.11240368,0.15047589,0.18673515,0.22480737,0.26287958,0.2991388,0.25925365,0.21936847,0.1794833,0.13959812,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.2229944,0.39522585,0.56745726,0.73968875,0.9119202,0.7306239,0.5475147,0.36440548,0.18310922,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.054388877,0.11059072,0.16497959,0.21936847,0.2755703,0.27194437,0.27013144,0.26831847,0.26469254,0.26287958,0.6852999,1.1077201,1.5301404,1.9525607,2.374981,2.222692,2.0704033,1.9181144,1.7658255,1.6117238,1.4358664,1.258196,1.0805258,0.90285534,0.72518504,1.1077201,1.4902552,1.8727903,2.2553256,2.6378605,3.9377546,5.237649,6.5375433,7.837437,9.137331,13.4594345,17.781536,22.105453,26.427555,30.749659,35.947422,41.145187,46.34295,51.540714,56.738476,56.99592,57.253357,57.5108,57.768238,58.02568,55.989723,53.955578,51.919624,49.88548,47.84952,60.38072,72.9101,85.4413,97.97069,110.50007,99.28871,88.08097,76.86961,65.660065,54.45052,45.32225,36.195797,27.067532,17.939264,8.812811,8.027799,7.2427855,6.4577727,5.67276,4.8877473,4.019338,3.152742,2.2843328,1.4177368,0.5493277,0.53482395,0.52032024,0.5058166,0.4894999,0.4749962,0.46774435,0.4604925,0.45324063,0.44417584,0.43692398,1.0877775,1.7368182,2.3876717,3.0367124,3.6875658,3.9975824,4.307599,4.6176157,4.9276323,5.237649,5.462456,5.6872635,5.9120708,6.1368785,6.3616858,6.350808,6.338117,6.3254266,6.3127356,6.300045,6.2202744,6.1405044,6.060734,5.979151,5.89938,6.0625467,6.2257137,6.3870673,6.550234,6.7134004,7.413204,8.113008,8.812811,9.512614,10.212419,10.440851,10.667472,10.894093,11.122525,11.349146,12.750566,14.150173,15.54978,16.949387,18.350807,19.262728,20.174648,21.086567,22.000301,22.912222,23.379965,23.84771,24.315454,24.7832,25.24913,25.531952,25.814774,26.097597,26.380419,26.66324,27.696629,28.73183,29.767033,30.802235,31.837437,37.073273,42.307293,47.54313,52.777153,58.01299,58.06738,58.12177,58.17797,58.232357,58.286747,61.537388,64.78803,68.03686,71.2875,74.53815,69.57244,64.60855,59.64284,54.67714,49.713245,46.098198,42.48315,38.868103,35.253056,31.63801,34.59495,37.551895,40.51065,43.46759,46.424534,40.35292,34.279495,28.207886,22.136272,16.062849,15.674874,15.2869005,14.90074,14.512766,14.124791,12.279196,10.435412,8.589817,6.7442207,4.900438,4.893186,4.8841214,4.876869,4.8696175,4.8623657,4.9820213,5.101677,5.223145,5.3428006,5.462456,5.40988,5.3573046,5.3047285,5.2521524,5.199577,5.475147,5.750717,6.0244746,6.300045,6.5756154,6.107871,5.6401267,5.1723824,4.704638,4.2368937,3.4101827,2.5816586,1.7549478,0.92823684,0.099712946,0.11784257,0.13415924,0.15228885,0.17041849,0.18673515,0.4894999,0.79226464,1.0950294,1.3977941,1.7005589,2.759329,3.8199122,4.880495,5.9392653,6.9998484,7.6742706,8.350506,9.024928,9.699349,10.375585,8.925215,7.474845,6.0244746,4.5759177,3.1255474,2.570781,2.0142014,1.4594349,0.90466833,0.34990177,0.27919623,0.21030366,0.13959812,0.07070554,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.8499773,5.6999545,8.549932,11.399909,14.249886,15.8743,17.500528,19.124943,20.749357,22.375584,18.688019,15.000452,11.312886,7.6253204,3.9377546,3.199879,2.4620032,1.7241274,0.9880646,0.25018883,2.1628644,4.07554,5.9882154,7.900891,9.811753,7.93715,6.0625467,4.1879435,2.3133402,0.43692398,0.69980353,0.96268314,1.2255627,1.4866294,1.7495089,1.4122978,1.0750868,0.73787576,0.40066472,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.31182957,0.5620184,0.8122072,1.062396,1.3125849,1.9126755,2.5127661,3.1128569,3.7129474,4.313038,3.4754493,2.6378605,1.8002719,0.96268314,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.69980353,1.3996071,2.0994108,2.7992141,3.5008307,2.8880494,2.275268,1.6624867,1.0497054,0.43692398,0.46230546,0.48768693,0.51306844,0.53663695,0.5620184,0.9119202,1.261822,1.6117238,1.9616255,2.3133402,2.3876717,2.4620032,2.5381477,2.612479,2.6868105,4.0120864,5.337362,6.6626377,7.987913,9.313189,11.862214,14.413053,16.962078,19.512917,22.061941,22.562319,23.062696,23.563074,24.06164,24.562017,19.911768,15.263332,10.613083,5.962834,1.3125849,2.03777,2.762955,3.48814,4.213325,4.936697,3.9631362,2.9877625,2.0123885,1.0370146,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.0870222,0.11240368,0.13778515,0.16316663,0.18673515,0.33721104,0.48768693,0.63816285,0.7868258,0.93730164,0.97537386,1.0116332,1.0497054,1.0877775,1.1258497,1.49932,1.8746033,2.2498865,2.6251698,3.000453,3.437377,3.874301,4.313038,4.749962,5.186886,5.5494785,5.9120708,6.2746634,6.637256,6.9998484,6.7242785,6.450521,6.1749506,5.89938,5.6256227,5.0744824,4.5251546,3.975827,3.4246864,2.8753586,3.0747845,3.2742105,3.4754493,3.6748753,3.874301,3.9504454,4.024777,4.099108,4.175253,4.249584,3.3993049,2.5508385,1.7005589,0.85027945,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.099712946,0.13778515,0.17585737,0.21211663,0.25018883,0.34990177,0.44961473,0.5493277,0.6508536,0.7505665,0.73787576,0.72518504,0.7124943,0.69980353,0.6871128,0.5873999,0.48768693,0.387974,0.28826106,0.18673515,0.28826106,0.387974,0.48768693,0.5873999,0.6871128,2.324218,3.9631362,5.600241,7.2373466,8.874452,8.562622,8.2507925,7.93715,7.6253204,7.311678,7.0506115,6.787732,6.5248523,6.261973,6.000906,4.8750563,3.7492065,2.6251698,1.49932,0.37528324,0.774135,1.1747998,1.5754645,1.9743162,2.374981,1.9743162,1.5754645,1.1747998,0.774135,0.37528324,1.2998942,2.2245052,3.150929,4.07554,5.0001507,4.40006,3.7999697,3.199879,2.5997884,1.9996977,2.4003625,2.7992141,3.199879,3.6005437,3.9993954,3.6748753,3.350355,3.0258346,2.6995013,2.374981,2.03777,1.7005589,1.3633479,1.0243238,0.6871128,0.9499924,1.2128719,1.4757515,1.7368182,1.9996977,3.636803,5.275721,6.9128265,8.549932,10.1870365,10.88684,11.586644,12.28826,12.988064,13.687867,12.1504755,10.613083,9.07569,7.5382986,6.000906,4.800725,3.6005437,2.4003625,1.2001812,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.41335547,0.824898,1.2382535,1.649796,2.0631514,1.887294,1.7132497,1.5373923,1.3633479,1.1874905,1.0116332,0.8375887,0.66173136,0.48768693,0.31182957,0.2755703,0.2374981,0.19942589,0.16316663,0.12509441,1.7621996,3.3993049,5.038223,6.6753283,8.312433,13.550082,18.787731,24.025381,29.26303,34.50068,40.387367,46.274055,52.16256,58.049248,63.93775,62.099407,60.262875,58.424534,56.588,54.749657,53.574856,52.40006,51.225258,50.050457,48.87566,62.862663,76.84967,90.83849,104.82549,65535.0,105.15002,91.48753,77.82504,64.16256,50.500072,41.56217,32.626076,23.686356,14.750263,5.812358,5.475147,5.137936,4.800725,4.461701,4.12449,3.299592,2.474694,1.649796,0.824898,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.9246109,1.7875811,2.6505513,3.5117085,4.3746786,4.650249,4.9258194,5.199577,5.475147,5.750717,6.1006193,6.450521,6.8004227,7.1503243,7.500226,7.224656,6.9508986,6.6753283,6.399758,6.1241875,6.0244746,5.924762,5.825049,5.7253356,5.6256227,5.9882154,6.350808,6.7134004,7.07418,7.4367723,7.93715,8.437528,8.937905,9.438283,9.936848,9.6504,9.362139,9.07569,8.78743,8.499168,9.875207,11.249433,12.625471,13.999697,15.375735,16.037468,16.699198,17.362743,18.024473,18.688019,18.862062,19.03792,19.211964,19.387821,19.561867,19.275417,18.987158,18.700708,18.412449,18.124187,18.77504,19.424082,20.074934,20.725788,21.374828,27.899681,34.424534,40.949387,47.47424,54.000904,55.11225,56.22541,57.336754,58.449913,59.563072,64.18794,68.812805,73.437675,78.062546,82.68741,76.71188,70.738174,64.76265,58.787125,52.8116,49.412296,46.01299,42.611874,39.212566,35.813263,39.33766,42.86206,46.388275,49.912674,53.437073,46.02387,38.612476,31.199272,23.787882,16.374678,16.050158,15.725637,15.399304,15.074784,14.750263,12.687112,10.625773,8.562622,6.4994707,4.4381323,4.3873696,4.3366065,4.2876563,4.2368937,4.1879435,4.699199,5.2122674,5.7253356,6.2365913,6.7496595,6.70071,6.6499467,6.599184,6.550234,6.4994707,6.5375433,6.5756154,6.6118746,6.6499467,6.688019,6.2873545,5.8866897,5.487838,5.087173,4.688321,3.7618973,2.8372865,1.9126755,0.9880646,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.41335547,0.824898,1.2382535,1.649796,2.0631514,3.3993049,4.7372713,6.0752378,7.413204,8.749357,9.5869465,10.424535,11.262123,12.099712,12.937301,11.124338,9.311376,7.500226,5.6872635,3.874301,3.1871881,2.5000753,1.8129625,1.1258497,0.43692398,0.34990177,0.26287958,0.17585737,0.0870222,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.11421664,0.23024625,0.3444629,0.4604925,0.5747091,0.54570174,0.5148814,0.48587397,0.4550536,0.42423326,0.36077955,0.2955129,0.23024625,0.16497959,0.099712946,2.373168,4.64481,6.9182653,9.189907,11.46155,12.852092,14.242634,15.633177,17.021906,18.412449,15.656745,12.902855,10.147152,7.3932614,4.6375585,3.8180993,2.9968271,2.1773682,1.357909,0.53663695,2.3949237,4.25321,6.109684,7.9679704,9.824444,7.9734097,6.1205616,4.267714,2.4148662,0.5620184,0.7469406,0.9318628,1.1167849,1.3017071,1.4866294,1.2201238,0.95180535,0.6852999,0.4169814,0.15047589,0.12328146,0.09427405,0.06707962,0.03988518,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.27194437,0.48224804,0.69255173,0.90285534,1.1131591,1.5917811,2.0722163,2.5526514,3.0330863,3.5117085,2.8354735,2.1574254,1.4793775,0.8031424,0.12509441,0.15954071,0.19579996,0.23024625,0.26469254,0.2991388,0.87566096,1.4503701,2.0250793,2.5997884,3.1744974,3.0149567,2.855416,2.6958754,2.5345216,2.374981,2.0921588,1.8093367,1.5283275,1.2455053,0.96268314,1.3669738,1.7730774,2.1773682,2.5816586,2.9877625,3.2633326,3.53709,3.8126602,4.0882306,4.361988,5.772473,7.1829576,8.593443,10.002114,11.4126,14.3079,17.203201,20.098503,22.991991,25.887293,25.406858,24.928236,24.4478,23.967365,23.48693,19.188396,14.888049,10.587702,6.2873545,1.987007,2.6016014,3.2180085,3.832603,4.4471974,5.0617914,4.269527,3.4772623,2.6849976,1.892733,1.1004683,1.2291887,1.3597219,1.4902552,1.6207886,1.7495089,1.6117238,1.4757515,1.3379664,1.2001812,1.062396,1.0968424,1.1331016,1.167548,1.2019942,1.2382535,1.1947423,1.1530442,1.1095331,1.067835,1.0243238,1.3125849,1.6008459,1.887294,2.175555,2.4620032,2.8481643,3.2325122,3.6168604,4.0030212,4.3873696,4.708264,5.027345,5.3482394,5.667321,5.9882154,5.7017674,5.4171324,5.132497,4.847862,4.5632267,4.1099863,3.6567454,3.2053177,2.752077,2.3006494,2.4620032,2.6251698,2.7883365,2.94969,3.1128569,3.1726844,3.2325122,3.29234,3.3521678,3.4119956,2.7321346,2.0522738,1.3724127,0.69255173,0.012690738,0.01994259,0.027194439,0.034446288,0.04169814,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.07977036,0.11059072,0.13959812,0.17041849,0.19942589,0.27919623,0.36077955,0.4405499,0.52032024,0.6000906,0.59283876,0.5855869,0.57833505,0.56927025,0.5620184,0.48587397,0.40791658,0.32995918,0.2520018,0.17585737,0.2520018,0.32995918,0.40791658,0.48587397,0.5620184,1.8746033,3.1871881,4.499773,5.812358,7.124943,6.965402,6.8058615,6.644508,6.484967,6.3254266,6.069799,5.814171,5.560356,5.3047285,5.049101,4.269527,3.489953,2.7103791,1.9308052,1.1494182,1.6226015,2.0957847,2.5671551,3.0403383,3.5117085,3.007705,2.5018883,1.9978848,1.4920682,0.9880646,1.6207886,2.2516994,2.8844235,3.5171473,4.1498713,3.7673361,3.3848011,3.002266,2.619731,2.2371957,2.5381477,2.8372865,3.1382382,3.437377,3.738329,3.4047437,3.0729716,2.7393866,2.4076142,2.0758421,2.1392958,2.2045624,2.269829,2.335096,2.4003625,2.6958754,2.9895754,3.2850883,3.5806012,3.874301,4.7554007,5.634688,6.5157876,7.3950744,8.274362,9.015862,9.755551,10.49524,11.234929,11.974618,10.765372,9.554313,8.345067,7.135821,5.924762,4.7390842,3.5552197,2.3695421,1.1856775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.15228885,0.3045777,0.45686656,0.6091554,0.76325727,0.6091554,0.45686656,0.3045777,0.15228885,0.0,0.058014803,0.11421664,0.17223145,0.23024625,0.28826106,0.25018883,0.21211663,0.17585737,0.13778515,0.099712946,0.08520924,0.07070554,0.054388877,0.03988518,0.025381476,0.030820364,0.034446288,0.03988518,0.045324065,0.05076295,0.17041849,0.29007402,0.40972954,0.5293851,0.6508536,0.52575916,0.40066472,0.2755703,0.15047589,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.15047589,0.13234627,0.11421664,0.09789998,0.07977036,0.06164073,0.052575916,0.04169814,0.032633327,0.02175555,0.012690738,0.032633327,0.052575916,0.072518505,0.092461094,0.11240368,0.09064813,0.06707962,0.045324065,0.02175555,0.0,0.33721104,0.6744221,1.0116332,1.3506571,1.6878681,1.6080978,1.5283275,1.4467441,1.3669738,1.2872034,1.1548572,1.0225109,0.8901646,0.75781834,0.62547207,0.52213323,0.42060733,0.31726846,0.21574254,0.11240368,1.5446441,2.9768846,4.409125,5.8431783,7.2754188,11.644659,16.013899,20.38495,24.75419,29.125244,33.780933,38.434807,43.090496,47.74437,52.40006,51.79634,51.19444,50.592533,49.99063,49.386913,50.73757,52.088226,53.437073,54.787727,56.138386,66.379814,76.62305,86.86448,97.10771,107.349144,94.40821,81.47091,68.52998,55.589058,42.649944,35.178726,27.70932,20.239914,12.770509,5.2992897,5.0001507,4.699199,4.40006,4.099108,3.7999697,3.147303,2.4946365,1.84197,1.1893034,0.53663695,0.4749962,0.41335547,0.34990177,0.28826106,0.22480737,0.2374981,0.25018883,0.26287958,0.2755703,0.28826106,1.0533313,1.8165885,2.5816586,3.346729,4.1117992,4.360175,4.606738,4.855114,5.101677,5.3500524,5.667321,5.9845896,6.301858,6.6191263,6.9382076,6.8004227,6.6626377,6.5248523,6.3870673,6.249282,6.155008,6.060734,5.964647,5.870373,5.774286,6.0824895,6.390693,6.697084,7.0052876,7.311678,7.7268467,8.1420145,8.557183,8.972352,9.38752,8.887142,8.386765,7.8882003,7.3878226,6.887445,8.045928,9.202598,10.359268,11.517752,12.674421,13.41411,14.155612,14.895301,15.63499,16.374678,16.38737,16.400059,16.41275,16.425442,16.438131,16.262274,16.08823,15.912373,15.738328,15.56247,16.184317,16.807976,17.429823,18.051668,18.675327,24.28826,29.89938,35.51231,41.125244,46.738174,48.009064,49.28176,50.554462,51.82716,53.09986,57.079315,61.06058,65.04003,69.019485,72.99894,69.68665,66.374374,63.06209,59.74981,56.437527,53.92657,51.41743,48.90829,46.39734,43.8882,45.276928,46.66747,48.058014,49.446743,50.837284,45.440094,40.042904,34.645714,29.248526,23.849524,24.077955,24.304577,24.53301,24.75963,24.988064,22.205166,19.422268,16.63937,13.858286,11.075388,10.460794,9.844387,9.229793,8.615198,8.000604,7.9280853,7.855567,7.783048,7.71053,7.6380115,7.473032,7.308052,7.1430726,6.978093,6.813113,6.9128265,7.0125394,7.112252,7.211965,7.311678,6.688019,6.0625467,5.4370747,4.8134155,4.1879435,3.8180993,3.4482548,3.0784104,2.7067533,2.3369088,1.983381,1.6280404,1.2726997,0.91735905,0.5620184,1.1548572,1.7476959,2.3405347,2.9333735,3.5243993,4.441758,5.3609304,6.2782893,7.1956487,8.113008,8.696781,9.282369,9.867955,10.451729,11.037316,9.547061,8.056806,6.5665503,5.0781083,3.587853,2.9424384,2.2970235,1.651609,1.0080072,0.36259252,0.30276474,0.24293698,0.18310922,0.12328146,0.06164073,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.23024625,0.4604925,0.69073874,0.91917205,1.1494182,1.0895905,1.0297627,0.969935,0.9101072,0.85027945,0.7197462,0.58921283,0.4604925,0.32995918,0.19942589,1.8945459,3.589666,5.2847857,6.979906,8.675026,9.829884,10.98474,12.139598,13.294455,14.449312,12.627284,10.805257,8.98323,7.159389,5.337362,4.4345064,3.531651,2.6306088,1.7277533,0.824898,2.6269827,4.4290676,6.2329655,8.03505,9.837135,8.007855,6.1767635,4.347484,2.518205,0.6871128,0.79589057,0.90285534,1.0098201,1.1167849,1.2255627,1.0279498,0.83033687,0.6327239,0.43511102,0.2374981,0.19579996,0.15228885,0.11059072,0.06707962,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.23205921,0.40247768,0.5728962,0.7433147,0.9119202,1.2726997,1.6316663,1.9924458,2.3532255,2.712192,2.1954978,1.6769904,1.1602961,0.6417888,0.12509441,0.21936847,0.3154555,0.40972954,0.5058166,0.6000906,1.0497054,1.49932,1.9507477,2.4003625,2.8499773,3.141864,3.435564,3.727451,4.019338,4.313038,3.7220123,3.1327994,2.5417736,1.9525607,1.3633479,1.8220274,2.2825198,2.7430124,3.2016919,3.6621845,4.137181,4.612177,5.087173,5.562169,6.037165,7.5328593,9.026741,10.522435,12.018129,13.512011,16.751774,19.991539,23.233116,26.47288,29.712645,28.253208,26.791962,25.332525,23.87309,22.411844,18.463211,14.512766,10.56232,6.6118746,2.663242,3.1672456,3.673062,4.177066,4.6828823,5.186886,4.5777307,3.966762,3.3576066,2.7466383,2.137483,2.3967366,2.657803,2.9170568,3.1781235,3.437377,3.1382382,2.8372865,2.5381477,2.2371957,1.938057,1.8582866,1.7767034,1.696933,1.6171626,1.5373923,1.4141108,1.2926424,1.1693609,1.0478923,0.9246109,1.1258497,1.3252757,1.5247015,1.7241274,1.9253663,2.2571385,2.5907235,2.9224956,3.254268,3.587853,3.8652363,4.1426196,4.420003,4.6973863,4.974769,4.6792564,4.3855567,4.0900435,3.7945306,3.5008307,3.1454902,2.7901495,2.4348087,2.079468,1.7241274,1.8492218,1.9743162,2.0994108,2.2245052,2.3495996,2.3949237,2.4402475,2.4855716,2.5308957,2.5744069,2.0649643,1.5555218,1.0442665,0.53482395,0.025381476,0.027194439,0.030820364,0.032633327,0.034446288,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.059827764,0.08339628,0.10515183,0.12690738,0.15047589,0.21030366,0.27013144,0.32995918,0.38978696,0.44961473,0.44780177,0.44417584,0.44236287,0.4405499,0.43692398,0.3825351,0.32814622,0.27194437,0.21755551,0.16316663,0.21755551,0.27194437,0.32814622,0.3825351,0.43692398,1.4249886,2.4130533,3.3993049,4.3873696,5.375434,5.368182,5.3591175,5.351866,5.3446136,5.337362,5.090799,4.842423,4.59586,4.347484,4.099108,3.6658103,3.2306993,2.7955883,2.3604772,1.9253663,2.469255,3.0149567,3.5606585,4.1045475,4.650249,4.0392804,3.4301252,2.819157,2.2100015,1.6008459,1.93987,2.280707,2.619731,2.960568,3.299592,3.1346123,2.9696326,2.8046532,2.6396735,2.474694,2.6741197,2.8753586,3.0747845,3.2742105,3.4754493,3.1346123,2.7955883,2.4547513,2.1157274,1.7748904,2.2426348,2.7103791,3.1781235,3.6458678,4.1117992,4.439945,4.7680917,5.0944247,5.422571,5.750717,5.8721857,5.995467,6.1169357,6.240217,6.3616858,7.1430726,7.9226465,8.70222,9.481794,10.263181,9.380268,8.497355,7.614443,6.733343,5.8504305,4.6792564,3.5098956,2.3405347,1.1693609,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.26831847,0.53482395,0.8031424,1.0696479,1.3379664,1.0696479,0.8031424,0.53482395,0.26831847,0.0,0.11421664,0.23024625,0.3444629,0.4604925,0.5747091,0.4749962,0.37528324,0.2755703,0.17585737,0.07433146,0.07070554,0.065266654,0.059827764,0.054388877,0.05076295,0.047137026,0.045324065,0.04169814,0.03988518,0.038072214,0.26469254,0.49312583,0.7197462,0.9481794,1.1747998,0.9499924,0.72518504,0.50037766,0.2755703,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,0.2991388,0.26469254,0.23024625,0.19579996,0.15954071,0.12509441,0.10515183,0.08520924,0.065266654,0.045324065,0.025381476,0.065266654,0.10515183,0.14503701,0.18492219,0.22480737,0.1794833,0.13415924,0.09064813,0.045324065,0.0,0.26287958,0.52575916,0.7868258,1.0497054,1.3125849,1.3270886,1.3415923,1.357909,1.3724127,1.3869164,1.2980812,1.2074331,1.1167849,1.0279498,0.93730164,0.7705091,0.60190356,0.43511102,0.26831847,0.099712946,1.3270886,2.5544643,3.7818398,5.009216,6.2365913,9.741048,13.2418785,16.744522,20.247166,23.74981,27.172684,30.595556,34.01843,37.43949,40.862362,41.495087,42.12781,42.760536,43.39326,44.02417,47.900284,51.774586,55.6507,59.525,63.3993,69.89877,76.394615,82.89227,89.38993,95.88759,83.67004,71.452484,59.23493,47.017372,34.799816,28.797098,22.794378,16.79166,10.790753,4.788034,4.5251546,4.262275,3.9993954,3.738329,3.4754493,2.9950142,2.514579,2.034144,1.5555218,1.0750868,0.9499924,0.824898,0.69980353,0.5747091,0.44961473,0.46230546,0.4749962,0.48768693,0.50037766,0.51306844,1.1802386,1.8474089,2.514579,3.1817493,3.8507326,4.070101,4.2894692,4.510651,4.7300196,4.949388,5.235836,5.520471,5.805106,6.089741,6.3743763,6.3743763,6.3743763,6.3743763,6.3743763,6.3743763,6.285541,6.1948934,6.104245,6.01541,5.924762,6.1767635,6.430578,6.68258,6.9345818,7.1883965,7.518356,7.8483152,8.178274,8.508233,8.838193,8.125698,7.413204,6.70071,5.9882154,5.275721,6.2148356,7.155763,8.094878,9.035806,9.97492,10.792566,11.610212,12.427858,13.245504,14.06315,13.912675,13.762199,13.611723,13.46306,13.312584,13.24913,13.1874895,13.125849,13.062395,13.000754,13.595407,14.190058,14.78471,15.379361,15.975826,20.675026,25.374224,30.075235,34.774437,39.47545,40.90769,42.339928,43.772167,45.20441,46.63665,49.9725,53.306538,56.64239,59.97643,63.31228,62.66324,62.012386,61.363346,60.71249,60.061638,58.44266,56.821873,55.202896,53.582108,51.963135,51.218006,50.472878,49.72775,48.982624,48.237495,44.854507,41.47333,38.090343,34.707355,31.324368,32.105755,32.885326,33.6649,34.444477,35.225864,31.723219,28.220575,24.717932,21.215288,17.712645,16.532406,15.352167,14.171928,12.993503,11.813264,11.155159,10.497053,9.840761,9.182655,8.52455,8.245354,7.9643445,7.6851482,7.404139,7.124943,7.28811,7.4494634,7.61263,7.7757964,7.93715,7.0868707,6.2365913,5.388125,4.537845,3.6875658,3.872488,4.0574102,4.2423325,4.4272547,4.612177,3.9141862,3.2180085,2.520018,1.8220274,1.1258497,1.8981718,2.6704938,3.442816,4.215138,4.98746,5.484212,5.9827766,6.4795284,6.978093,7.474845,7.806617,8.140202,8.471974,8.805559,9.137331,7.9697833,6.8022356,5.634688,4.4671397,3.299592,2.6976883,2.0957847,1.4920682,0.8901646,0.28826106,0.25562772,0.2229944,0.19036107,0.15772775,0.12509441,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.3444629,0.69073874,1.0352017,1.3796645,1.7241274,1.6352923,1.5446441,1.455809,1.3651608,1.2745126,1.0805258,0.88472575,0.69073874,0.4949388,0.2991388,1.4177368,2.5345216,3.6531196,4.7699046,5.8866897,6.8076744,7.7268467,8.647832,9.567003,10.487988,9.597824,8.70766,7.817495,6.92733,6.037165,5.0527267,4.068288,3.0820365,2.0975976,1.1131591,2.8608549,4.606738,6.354434,8.10213,9.849826,8.042302,6.2347784,4.4272547,2.619731,0.8122072,0.8430276,0.872035,0.90285534,0.9318628,0.96268314,0.83577573,0.7070554,0.58014804,0.45324063,0.3245203,0.26831847,0.21030366,0.15228885,0.09427405,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.19217403,0.32270733,0.45324063,0.581961,0.7124943,0.95180535,1.1929294,1.4322405,1.6733645,1.9126755,1.5555218,1.1983683,0.83940166,0.48224804,0.12509441,0.27919623,0.43511102,0.58921283,0.7451276,0.89922947,1.2255627,1.550083,1.8746033,2.1991236,2.525457,3.2705846,4.0157123,4.76084,5.504154,6.249282,5.351866,4.454449,3.5570326,2.659616,1.7621996,2.277081,2.7919624,3.3068438,3.8217251,4.3366065,5.0128417,5.6872635,6.3616858,7.037921,7.7123427,9.293246,10.872336,12.45324,14.0323305,15.613234,19.19746,22.781689,26.367727,29.951954,33.537994,31.097748,28.6575,26.217253,23.777004,21.336756,17.738026,14.137483,10.536939,6.9382076,3.3376641,3.73289,4.1281157,4.5233417,4.9167547,5.3119802,4.8841214,4.458075,4.0302157,3.6023567,3.1744974,3.5642843,3.9558845,4.345671,4.7354584,5.125245,4.6629395,4.2006345,3.738329,3.2742105,2.811905,2.617918,2.422118,2.228131,2.032331,1.8383441,1.6352923,1.4322405,1.2291887,1.0279498,0.824898,0.93730164,1.0497054,1.162109,1.2745126,1.3869164,1.6679256,1.9471219,2.228131,2.5073273,2.7883365,3.0222087,3.2578938,3.491766,3.727451,3.9631362,3.6567454,3.3521678,3.04759,2.7430124,2.4366217,2.179181,1.9217403,1.6642996,1.4068589,1.1494182,1.2382535,1.3252757,1.4122978,1.49932,1.5881553,1.6171626,1.647983,1.6769904,1.7078108,1.7368182,1.3977941,1.0569572,0.7179332,0.3770962,0.038072214,0.034446288,0.032633327,0.030820364,0.027194439,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.03988518,0.054388877,0.07070554,0.08520924,0.099712946,0.13959812,0.1794833,0.21936847,0.25925365,0.2991388,0.30276474,0.3045777,0.30820364,0.3100166,0.31182957,0.27919623,0.24837588,0.21574254,0.18310922,0.15047589,0.18310922,0.21574254,0.24837588,0.27919623,0.31182957,0.97537386,1.6371052,2.3006494,2.962381,3.6241121,3.7691493,3.9141862,4.059223,4.2042603,4.349297,4.1099863,3.870675,3.6295512,3.39024,3.149116,3.0602808,2.9696326,2.8807976,2.7901495,2.6995013,3.3177216,3.9341288,4.552349,5.1705694,5.7869763,5.0726695,4.358362,3.6422417,2.9279346,2.2118144,2.2607644,2.3079014,2.3550384,2.4021754,2.4493124,2.5018883,2.5544643,2.6070402,2.659616,2.712192,2.811905,2.911618,3.0131438,3.1128569,3.2125697,2.864481,2.518205,2.1701162,1.8220274,1.4757515,2.3441606,3.2143826,4.0846047,4.954827,5.825049,6.185828,6.544795,6.9055743,7.264541,7.6253204,6.9907837,6.354434,5.719897,5.08536,4.4508233,5.2702823,6.089741,6.9092,7.7304726,8.549932,7.995165,7.440398,6.885632,6.3308654,5.774286,4.6194286,3.4645715,2.3097143,1.1548572,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.3825351,0.7650702,1.1476053,1.5301404,1.9126755,1.5301404,1.1476053,0.7650702,0.3825351,0.0,0.17223145,0.3444629,0.5166943,0.69073874,0.8629702,0.69980353,0.53663695,0.37528324,0.21211663,0.05076295,0.054388877,0.059827764,0.065266654,0.07070554,0.07433146,0.065266654,0.054388877,0.045324065,0.034446288,0.025381476,0.36077955,0.69436467,1.0297627,1.3651608,1.7005589,1.3742256,1.0497054,0.72518504,0.40066472,0.07433146,0.15047589,0.22480737,0.2991388,0.37528324,0.44961473,0.39703882,0.3444629,0.291887,0.23931105,0.18673515,0.15772775,0.12690738,0.09789998,0.06707962,0.038072214,0.09789998,0.15772775,0.21755551,0.27738327,0.33721104,0.27013144,0.2030518,0.13415924,0.06707962,0.0,0.18673515,0.37528324,0.5620184,0.7505665,0.93730164,1.0478923,1.1566701,1.2672608,1.3778516,1.4866294,1.4394923,1.3923552,1.3452182,1.2980812,1.2491312,1.017072,0.7850128,0.5529536,0.3208944,0.0870222,1.1095331,2.132044,3.1545548,4.177066,5.199577,7.835624,10.469859,13.1059065,15.740141,18.374376,20.564434,22.754494,24.944551,27.134611,29.324669,31.19202,33.059372,34.926723,36.795887,38.66324,45.063,51.462757,57.862514,64.26227,70.66203,73.41592,76.168,78.920074,81.67215,84.424225,72.930046,61.435863,49.93987,38.445686,26.949688,22.41547,17.879436,13.345218,8.809185,4.274966,4.0501585,3.825351,3.6005437,3.3757362,3.149116,2.8427253,2.5345216,2.228131,1.9199274,1.6117238,1.4249886,1.2382535,1.0497054,0.8629702,0.6744221,0.6871128,0.69980353,0.7124943,0.72518504,0.73787576,1.3071461,1.8782293,2.4474995,3.0167696,3.587853,3.780027,3.972201,4.164375,4.358362,4.550536,4.802538,5.0545397,5.3083544,5.560356,5.812358,5.9501433,6.0879283,6.2257137,6.3616858,6.4994707,6.414262,6.3308654,6.245656,6.1604466,6.0752378,6.2728505,6.4704633,6.6680765,6.8656893,7.063302,7.308052,7.552802,7.797552,8.042302,8.287052,7.362441,6.43783,5.5132194,4.5867953,3.6621845,4.3855567,5.1071157,5.8304877,6.552047,7.2754188,8.1692095,9.064813,9.960417,10.854207,11.74981,11.437981,11.124338,10.812509,10.500679,10.1870365,10.2378,10.28675,10.337513,10.388275,10.437225,11.004683,11.57214,12.139598,12.707055,13.274512,17.063604,20.84907,24.63816,28.42544,32.21272,33.8045,35.398094,36.989876,38.581657,40.17525,42.86569,45.55431,48.244747,50.935184,53.62562,55.63801,57.6504,59.662785,61.675175,63.68756,62.95694,62.228127,61.497505,60.76688,60.03807,57.157272,54.278286,51.397488,48.518505,45.637707,44.270733,42.901947,41.534973,40.168,38.799213,40.13174,41.464268,42.796795,44.129322,45.46185,41.23946,37.01707,32.79468,28.57229,24.349901,22.604017,20.859947,19.114065,17.369995,15.624111,14.382232,13.140353,11.896661,10.654781,9.412902,9.017676,8.62245,8.227224,7.8319983,7.4367723,7.663393,7.8882003,8.113008,8.337815,8.562622,7.4875355,6.412449,5.337362,4.262275,3.1871881,3.926877,4.668379,5.408067,6.147756,6.887445,5.846804,4.8079767,3.7673361,2.7266958,1.6878681,2.6396735,3.5932918,4.5450974,5.4969025,6.450521,6.526665,6.604623,6.68258,6.7605376,6.836682,6.9182653,6.9980354,7.077806,7.157576,7.2373466,6.392506,5.5476656,4.702825,3.8579843,3.0131438,2.4529383,1.892733,1.3325275,0.77232206,0.21211663,0.20667773,0.2030518,0.19761293,0.19217403,0.18673515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.4604925,0.91917205,1.3796645,1.840157,2.3006494,2.179181,2.0595255,1.93987,1.8202144,1.7005589,1.4394923,1.1802386,0.91917205,0.65991837,0.40066472,0.93911463,1.4793775,2.0196402,2.5599031,3.100166,3.785466,4.4707656,5.1542525,5.8395524,6.5248523,6.5665503,6.6100616,6.6517596,6.695271,6.736969,5.669134,4.603112,3.5352771,2.467442,1.3996071,3.092914,4.784408,6.4777155,8.1692095,9.862516,8.076748,6.2927933,4.507025,2.72307,0.93730164,0.8901646,0.8430276,0.79589057,0.7469406,0.69980353,0.6417888,0.5855869,0.5275721,0.46955732,0.41335547,0.34083697,0.26831847,0.19579996,0.12328146,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.15228885,0.24293698,0.33177215,0.4224203,0.51306844,0.6327239,0.7523795,0.872035,0.9916905,1.1131591,0.9155461,0.7179332,0.52032024,0.32270733,0.12509441,0.34083697,0.55476654,0.7705091,0.98443866,1.2001812,1.3996071,1.6008459,1.8002719,1.9996977,2.1991236,3.397492,4.59586,5.7924156,6.9907837,8.187339,6.981719,5.7779117,4.572292,3.3666716,2.1628644,2.7321346,3.303218,3.872488,4.441758,5.0128417,5.8866897,6.7623506,7.6380115,8.511859,9.38752,11.05182,12.717933,14.382232,16.048346,17.712645,21.643147,25.571836,29.50234,33.432842,37.363346,33.942284,30.523039,27.101978,23.68273,20.26167,17.01284,13.762199,10.511557,7.262728,4.0120864,4.2967215,4.5831695,4.8678045,5.1524396,5.4370747,5.1923246,4.947575,4.702825,4.458075,4.213325,4.7318325,5.2521524,5.772473,6.2927933,6.813113,6.187641,5.562169,4.936697,4.313038,3.6875658,3.3775494,3.0675328,2.7575161,2.4474995,2.137483,1.8546607,1.5718386,1.2908293,1.0080072,0.72518504,0.7505665,0.774135,0.7995165,0.824898,0.85027945,1.0768998,1.305333,1.5319533,1.7603867,1.987007,2.179181,2.373168,2.565342,2.7575161,2.94969,2.6342347,2.3205922,2.0051367,1.6896812,1.3742256,1.214685,1.0551442,0.89560354,0.73424983,0.5747091,0.62547207,0.6744221,0.72518504,0.774135,0.824898,0.83940166,0.8557183,0.87022203,0.88472575,0.89922947,0.7306239,0.56020546,0.38978696,0.21936847,0.05076295,0.04169814,0.034446288,0.027194439,0.01994259,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.01994259,0.027194439,0.034446288,0.04169814,0.05076295,0.07070554,0.09064813,0.11059072,0.13053331,0.15047589,0.15772775,0.16497959,0.17223145,0.1794833,0.18673515,0.17767033,0.16679256,0.15772775,0.14684997,0.13778515,0.14684997,0.15772775,0.16679256,0.17767033,0.18673515,0.52575916,0.8629702,1.2001812,1.5373923,1.8746033,2.1719291,2.469255,2.7683938,3.0657198,3.3630457,3.1291735,2.8971143,2.665055,2.4329958,2.1991236,2.4547513,2.7103791,2.9641938,3.2198215,3.4754493,4.164375,4.855114,5.5458527,6.2347784,6.925517,6.104245,5.2847857,4.465327,3.6458678,2.8245957,2.5798457,2.335096,2.0903459,1.845596,1.6008459,1.8691645,2.1392958,2.4094272,2.6795588,2.94969,2.94969,2.94969,2.94969,2.94969,2.94969,2.5943494,2.2408218,1.8854811,1.5301404,1.1747998,2.4474995,3.720199,4.992899,6.265599,7.5382986,7.9298983,8.323311,8.714911,9.108324,9.499924,8.107569,6.7152133,5.3228583,3.930503,2.5381477,3.397492,4.256836,5.1179934,5.977338,6.836682,6.6100616,6.3816285,6.155008,5.9283876,5.6999545,4.559601,3.4192474,2.280707,1.1403534,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.49675176,0.99531645,1.4920682,1.9906329,2.4873846,1.9906329,1.4920682,0.99531645,0.49675176,0.0,0.23024625,0.4604925,0.69073874,0.91917205,1.1494182,0.9246109,0.69980353,0.4749962,0.25018883,0.025381476,0.03988518,0.054388877,0.07070554,0.08520924,0.099712946,0.08339628,0.065266654,0.047137026,0.030820364,0.012690738,0.4550536,0.8974165,1.3397794,1.7821422,2.2245052,1.8002719,1.3742256,0.9499924,0.52575916,0.099712946,0.19942589,0.2991388,0.40066472,0.50037766,0.6000906,0.5293851,0.4604925,0.38978696,0.3208944,0.25018883,0.21030366,0.17041849,0.13053331,0.09064813,0.05076295,0.13053331,0.21030366,0.29007402,0.36984438,0.44961473,0.36077955,0.27013144,0.1794833,0.09064813,0.0,0.11240368,0.22480737,0.33721104,0.44961473,0.5620184,0.7668832,0.97174793,1.1766127,1.3832904,1.5881553,1.5827163,1.5772774,1.5718386,1.5682126,1.5627737,1.2654479,0.968122,0.67079616,0.37165734,0.07433146,0.8919776,1.7096237,2.5272698,3.3449159,4.162562,5.9302006,7.6978393,9.465478,11.233116,13.000754,13.957999,14.915243,15.872487,16.829731,17.786976,20.890768,23.992746,27.094727,30.196705,33.300495,42.22571,51.149113,60.07614,68.99954,77.92476,76.93307,75.93956,74.947876,73.95437,72.96268,62.190056,51.41743,40.64481,29.872185,19.099562,16.032028,12.964496,9.896963,6.82943,3.7618973,3.5751622,3.386614,3.199879,3.0131438,2.8245957,2.6904364,2.5544643,2.420305,2.2843328,2.1501737,1.8999848,1.649796,1.3996071,1.1494182,0.89922947,0.9119202,0.9246109,0.93730164,0.9499924,0.96268314,1.4358664,1.9072367,2.38042,2.8517902,3.3249733,3.489953,3.6549325,3.8199122,3.9848917,4.1498713,4.36924,4.590421,4.8097897,5.029158,5.2503395,5.52591,5.7996674,6.0752378,6.350808,6.624565,6.544795,6.4650245,6.3852544,6.305484,6.2257137,6.3671246,6.510349,6.6517596,6.794984,6.9382076,7.0977483,7.2572894,7.41683,7.5781837,7.7377243,6.599184,5.462456,4.325729,3.1871881,2.0504606,2.5544643,3.0602808,3.5642843,4.070101,4.574105,5.5476656,6.5194135,7.4929743,8.464723,9.438283,8.963287,8.488291,8.013294,7.5382986,7.063302,7.224656,7.3878226,7.549176,7.7123427,7.8755093,8.415772,8.954222,9.494485,10.034748,10.57501,13.45037,16.325727,19.199274,22.074633,24.949991,26.703125,28.454447,30.207582,31.958904,33.71204,35.75706,37.802082,39.847103,41.892128,43.93715,48.612778,53.286594,57.962227,62.637856,67.311676,67.47303,67.63257,67.79211,67.95346,68.11301,63.09654,58.081882,53.067226,48.052574,43.037918,43.685146,44.332375,44.979603,45.62683,46.27587,48.15954,50.045017,51.9305,53.814167,55.69965,50.757515,45.815376,40.87324,35.931107,30.987156,28.677443,26.367727,24.058014,21.748299,19.436771,17.609306,15.781839,13.954373,12.126906,10.29944,9.789998,9.280556,8.7693,8.259857,7.750415,8.036863,8.325124,8.613385,8.899834,9.188094,7.8882003,6.586493,5.2865987,3.9867048,2.6868105,3.9830787,5.277534,6.5719895,7.8682575,9.162713,7.7794223,6.397945,5.0146546,3.633177,2.2498865,3.3829882,4.514277,5.6473784,6.78048,7.911769,7.569119,7.228282,6.885632,6.542982,6.200332,6.0281005,5.8540564,5.6818247,5.5095935,5.337362,4.8152285,4.2930956,3.7691493,3.247016,2.7248828,2.2081885,1.6896812,1.1729867,0.6544795,0.13778515,0.15954071,0.18310922,0.20486477,0.22662032,0.25018883,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.5747091,1.1494182,1.7241274,2.3006494,2.8753586,2.7248828,2.5744069,2.4257438,2.275268,2.124792,1.8002719,1.4757515,1.1494182,0.824898,0.50037766,0.46230546,0.42423326,0.387974,0.34990177,0.31182957,0.76325727,1.2128719,1.6624867,2.1121013,2.561716,3.53709,4.512464,5.487838,6.4632115,7.4367723,6.2873545,5.137936,3.9867048,2.8372865,1.6878681,3.3249733,4.9620786,6.599184,8.238102,9.875207,8.113008,6.350808,4.5867953,2.8245957,1.062396,0.93730164,0.8122072,0.6871128,0.5620184,0.43692398,0.44961473,0.46230546,0.4749962,0.48768693,0.50037766,0.41335547,0.3245203,0.2374981,0.15047589,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.11240368,0.16316663,0.21211663,0.26287958,0.31182957,0.31182957,0.31182957,0.31182957,0.31182957,0.31182957,0.2755703,0.2374981,0.19942589,0.16316663,0.12509441,0.40066472,0.6744221,0.9499924,1.2255627,1.49932,1.5754645,1.649796,1.7241274,1.8002719,1.8746033,3.5243993,5.1741953,6.825804,8.4756,10.125396,8.613385,7.0995617,5.5875506,4.07554,2.561716,3.1871881,3.8126602,4.4381323,5.0617914,5.6872635,6.7623506,7.837437,8.912524,9.987611,11.062697,12.812206,14.561715,16.313038,18.062546,19.812056,24.08702,28.361986,32.63695,36.91192,41.186886,36.786823,32.386765,27.986704,23.586643,19.188396,16.287657,13.386916,10.487988,7.5872483,4.688321,4.8623657,5.038223,5.2122674,5.388125,5.562169,5.5005283,5.4370747,5.375434,5.3119802,5.2503395,5.89938,6.550234,7.1992745,7.850128,8.499168,7.7123427,6.925517,6.1368785,5.3500524,4.5632267,4.137181,3.7129474,3.2869012,2.8626678,2.4366217,2.0758421,1.7132497,1.3506571,0.9880646,0.62547207,0.5620184,0.50037766,0.43692398,0.37528324,0.31182957,0.48768693,0.66173136,0.8375887,1.0116332,1.1874905,1.3379664,1.4866294,1.6371052,1.7875811,1.938057,1.6117238,1.2872034,0.96268314,0.63816285,0.31182957,0.25018883,0.18673515,0.12509441,0.06164073,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.5747091,1.0243238,1.4757515,1.9253663,2.374981,2.1501737,1.9253663,1.7005589,1.4757515,1.2491312,1.8492218,2.4493124,3.049403,3.6494937,4.249584,5.0128417,5.774286,6.5375433,7.3008003,8.062244,7.137634,6.2130227,5.2865987,4.361988,3.437377,2.9007401,2.3622901,1.8256533,1.2872034,0.7505665,1.2382535,1.7241274,2.2118144,2.6995013,3.1871881,3.0874753,2.9877625,2.8880494,2.7883365,2.6868105,2.324218,1.9616255,1.6008459,1.2382535,0.87566096,2.5508385,4.2242026,5.89938,7.574558,9.249735,9.675781,10.100015,10.524248,10.950294,11.374527,9.224354,7.07418,4.9258194,2.7756457,0.62547207,1.5247015,2.4257438,3.3249733,4.2242026,5.125245,5.224958,5.3246713,5.424384,5.524097,5.6256227,4.499773,3.3757362,2.2498865,1.1258497,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.61278135,1.2255627,1.8383441,2.4493124,3.0620937,2.4493124,1.8383441,1.2255627,0.61278135,0.0,0.28826106,0.5747091,0.8629702,1.1494182,1.4376793,1.1494182,0.8629702,0.5747091,0.28826106,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.5493277,1.1004683,1.649796,2.1991236,2.7502642,2.2245052,1.7005589,1.1747998,0.6508536,0.12509441,0.25018883,0.37528324,0.50037766,0.62547207,0.7505665,0.66173136,0.5747091,0.48768693,0.40066472,0.31182957,0.26287958,0.21211663,0.16316663,0.11240368,0.06164073,0.16316663,0.26287958,0.36259252,0.46230546,0.5620184,0.44961473,0.33721104,0.22480737,0.11240368,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.48768693,0.7868258,1.0877775,1.3869164,1.6878681,1.7241274,1.7621996,1.8002719,1.8383441,1.8746033,1.5120108,1.1494182,0.7868258,0.42423326,0.06164073,0.6744221,1.2872034,1.8999848,2.5127661,3.1255474,4.024777,4.9258194,5.825049,6.7242785,7.6253204,7.3497505,7.07418,6.8004227,6.5248523,6.249282,10.587702,14.924308,19.262728,23.599335,27.937754,39.388424,50.837284,62.287956,73.73682,85.187485,80.45022,75.712944,70.97567,66.23659,61.499317,51.450066,41.400814,31.349749,21.300497,11.249433,9.6504,8.049554,6.450521,4.8496747,3.2506418,3.100166,2.94969,2.7992141,2.6505513,2.5000753,2.5381477,2.5744069,2.612479,2.6505513,2.6868105,2.374981,2.0631514,1.7495089,1.4376793,1.1258497,1.1367276,1.1494182,1.162109,1.1747998,1.1874905,1.5627737,1.938057,2.3133402,2.6868105,3.0620937,3.199879,3.3376641,3.4754493,3.6132345,3.7492065,3.9377546,4.12449,4.313038,4.499773,4.688321,5.0998635,5.5132194,5.924762,6.338117,6.7496595,6.6753283,6.599184,6.5248523,6.450521,6.3743763,6.4632115,6.550234,6.637256,6.7242785,6.813113,6.887445,6.9617763,7.037921,7.112252,7.1883965,5.8377395,4.4870825,3.1382382,1.7875811,0.43692398,0.72518504,1.0116332,1.2998942,1.5881553,1.8746033,2.9243085,3.975827,5.0255322,6.0752378,7.124943,6.48678,5.8504305,5.2122674,4.574105,3.9377546,4.213325,4.4870825,4.762653,5.038223,5.3119802,5.825049,6.338117,6.849373,7.362441,7.8755093,9.837135,11.800573,13.762199,15.725637,17.687263,19.59994,21.512613,23.42529,25.337965,27.25064,28.650248,30.049854,31.449461,32.849068,34.25049,41.587547,48.92461,56.26348,63.59873,70.9376,71.987305,73.03701,74.086716,75.13824,76.18794,69.03761,61.88729,54.736965,47.588455,40.43813,43.09956,45.762802,48.42423,51.08747,53.750713,56.187336,58.62577,61.062393,63.499016,65.93745,60.273754,54.611874,48.94999,43.28811,37.624413,34.749054,31.875507,29.000149,26.12479,23.249432,20.838192,18.425138,16.012085,13.600845,11.187792,10.56232,9.936848,9.313189,8.6877165,8.062244,8.412147,8.762048,9.11195,9.461852,9.811753,8.287052,6.7623506,5.237649,3.7129474,2.1882458,4.0374675,5.8885026,7.7377243,9.5869465,11.437981,9.712041,7.987913,6.261973,4.537845,2.811905,4.12449,5.4370747,6.7496595,8.062244,9.374829,8.611572,7.850128,7.0868707,6.3254266,5.562169,5.137936,4.7118897,4.2876563,3.8634233,3.437377,3.2379513,3.0367124,2.8372865,2.6378605,2.4366217,1.9616255,1.4866294,1.0116332,0.53663695,0.06164073,0.11240368,0.16316663,0.21211663,0.26287958,0.31182957,0.0,0.0,0.0,0.0,0.0,0.0,0.17223145,0.3444629,0.5166943,0.69073874,0.8629702,0.69980353,0.53663695,0.37528324,0.21211663,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.4604925,0.91917205,1.3796645,1.840157,2.3006494,2.179181,2.0595255,1.93987,1.8202144,1.7005589,1.4394923,1.1802386,0.91917205,0.65991837,0.40066472,0.37165734,0.3444629,0.31726846,0.29007402,0.26287958,0.62184614,0.9826257,1.3434052,1.7023718,2.0631514,3.5243993,4.98746,6.450521,7.911769,9.374829,8.040489,6.7043357,5.369995,4.0356545,2.6995013,3.872488,5.045475,6.2166486,7.3896356,8.562622,7.0524244,5.542227,4.0320287,2.521831,1.0116332,0.90829426,0.8031424,0.6979906,0.59283876,0.48768693,0.49675176,0.5076295,0.5166943,0.5275721,0.53663695,0.45324063,0.3680314,0.28282216,0.19761293,0.11240368,0.09064813,0.06707962,0.045324065,0.02175555,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.027194439,0.04169814,0.058014803,0.072518505,0.0870222,0.15410182,0.2229944,0.29007402,0.35715362,0.42423326,0.44417584,0.46411842,0.48587397,0.5058166,0.52575916,0.533011,0.5402629,0.5475147,0.55476654,0.5620184,0.8031424,1.0424535,1.2817645,1.5228885,1.7621996,1.8220274,1.8818551,1.9416829,2.0033236,2.0631514,3.343103,4.6230545,5.903006,7.1829576,8.46291,7.3497505,6.2384043,5.125245,4.0120864,2.9007401,3.4319382,3.9649491,4.49796,5.029158,5.562169,7.262728,8.963287,10.662033,12.362592,14.06315,17.4407,20.818249,24.195799,27.573347,30.950897,32.919773,34.890465,36.85934,38.830032,40.800724,35.822327,30.845745,25.86735,20.890768,15.912373,13.54283,11.173288,8.801933,6.432391,4.062849,4.2804046,4.49796,4.7155156,4.933071,5.1506267,5.1905117,5.230397,5.2702823,5.3101673,5.3500524,5.7978544,6.245656,6.6916447,7.1394467,7.5872483,6.8403077,6.093367,5.3446136,4.597673,3.8507326,3.6096084,3.3702974,3.1291735,2.8898623,2.6505513,2.3495996,2.0504606,1.7495089,1.4503701,1.1494182,0.99531645,0.83940166,0.6852999,0.5293851,0.37528324,0.4949388,0.61459434,0.73424983,0.8557183,0.97537386,1.0950294,1.214685,1.3343405,1.455809,1.5754645,1.3143979,1.0551442,0.79589057,0.53482395,0.2755703,0.22662032,0.1794833,0.13234627,0.08520924,0.038072214,0.03988518,0.04169814,0.045324065,0.047137026,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.059827764,0.07070554,0.07977036,0.09064813,0.099712946,0.09064813,0.07977036,0.07070554,0.059827764,0.05076295,0.11421664,0.1794833,0.24474995,0.3100166,0.37528324,0.8665961,1.3597219,1.8528478,2.3441606,2.8372865,2.5526514,2.268016,1.983381,1.696933,1.4122978,1.8129625,2.2118144,2.612479,3.0131438,3.4119956,4.7245803,6.037165,7.3497505,8.662335,9.97492,8.54268,7.1104393,5.678199,4.2441454,2.811905,2.8318477,2.8517902,2.8717327,2.8916752,2.913431,2.8427253,2.7720199,2.7031271,2.6324217,2.561716,2.9243085,3.2869012,3.6494937,4.0120864,4.3746786,3.6549325,2.9351864,2.2154403,1.4956942,0.774135,2.1574254,3.540716,4.9221935,6.305484,7.686961,8.352319,9.017676,9.683033,10.348391,11.011934,9.333132,7.652515,5.9718986,4.2930956,2.612479,3.0820365,3.5534067,4.022964,4.4925213,4.9620786,4.8696175,4.7771564,4.6846952,4.592234,4.499773,3.6005437,2.6995013,1.8002719,0.89922947,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.5166943,1.0098201,1.502946,1.9942589,2.4873846,1.9906329,1.4920682,0.99531645,0.49675176,0.0,0.23024625,0.4604925,0.69073874,0.91917205,1.1494182,1.0551442,0.96087015,0.86478317,0.7705091,0.6744221,0.56020546,0.44417584,0.32995918,0.21574254,0.099712946,0.09427405,0.09064813,0.08520924,0.07977036,0.07433146,0.50219065,0.9300498,1.357909,1.7857682,2.2118144,1.8691645,1.5283275,1.1856775,0.8430276,0.50037766,0.52032024,0.5402629,0.56020546,0.58014804,0.6000906,0.5293851,0.4604925,0.38978696,0.3208944,0.25018883,0.2374981,0.22480737,0.21211663,0.19942589,0.18673515,0.26469254,0.34264994,0.42060733,0.49675176,0.5747091,0.4604925,0.3444629,0.23024625,0.11421664,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.40066472,0.6508536,0.89922947,1.1494182,1.3996071,1.452183,1.504759,1.5573349,1.6099107,1.6624867,1.3669738,1.0732739,0.7777609,0.48224804,0.18673515,0.66173136,1.1367276,1.6117238,2.08672,2.561716,3.3666716,4.171627,4.9783955,5.7833505,6.588306,6.4233265,6.258347,6.093367,5.9283876,5.7615952,9.131892,12.50219,15.872487,19.242785,22.613083,31.942587,41.272095,50.603413,59.93292,69.26242,65.33373,61.406857,57.47998,53.55129,49.624413,42.07161,34.520622,26.96782,19.415016,11.862214,10.442664,9.023115,7.6017523,6.1822023,4.762653,4.421816,4.082792,3.7419548,3.4029307,3.0620937,2.9442513,2.8282216,2.7103791,2.5925364,2.474694,2.1628644,1.8492218,1.5373923,1.2255627,0.9119202,1.1167849,1.3216497,1.5283275,1.7331922,1.938057,2.2045624,2.472881,2.7393866,3.007705,3.2742105,3.3666716,3.4591327,3.5534067,3.6458678,3.738329,3.917812,4.0972953,4.2767787,4.458075,4.6375585,5.1143675,5.5929894,6.069799,6.546608,7.02523,6.849373,6.6753283,6.4994707,6.3254266,6.149569,6.1241875,6.1006193,6.0752378,6.049856,6.0244746,6.1278133,6.2293396,6.3326783,6.434204,6.5375433,5.33011,4.122677,2.9152439,1.7078108,0.50037766,0.79226464,1.0841516,1.3778516,1.6697385,1.9616255,2.7774587,3.5932918,4.407312,5.223145,6.037165,5.4896507,4.942136,4.3946214,3.8471067,3.299592,3.5352771,3.7691493,4.004834,4.2405195,4.4743915,5.038223,5.600241,6.16226,6.7242785,7.28811,8.812811,10.337513,11.862214,13.386916,14.911617,16.557787,18.202145,19.848314,21.492672,23.137028,24.910107,26.683184,28.454447,30.227526,32.000603,38.22269,44.44478,50.666866,56.888954,63.112854,64.41819,65.72171,67.02704,68.332375,69.6377,64.53422,59.43254,54.32905,49.22737,44.125698,45.342194,46.560505,47.777004,48.995316,50.21181,51.542526,52.87143,54.20214,55.532856,56.86176,52.40187,47.941982,43.482094,39.022205,34.562317,32.314243,30.067984,27.81991,25.571836,23.325577,21.842573,20.35957,18.87838,17.395376,15.912373,14.777458,13.642544,12.507628,11.372714,10.2378,10.388275,10.536939,10.687414,10.837891,10.988366,10.477111,9.967669,9.458226,8.94697,8.437528,9.782746,11.127964,12.473183,13.8184,15.161806,13.272699,11.381779,9.492672,7.603565,5.712645,6.3145485,6.9182653,7.520169,8.122072,8.725789,8.002417,7.2790446,6.5574856,5.8359265,5.1125546,4.652062,4.1915693,3.73289,3.2723975,2.811905,2.6523643,2.4928236,2.333283,2.1719291,2.0123885,1.6207886,1.2273756,0.83577573,0.44236287,0.05076295,0.09064813,0.13053331,0.17041849,0.21030366,0.25018883,0.0,0.0,0.0,0.0,0.0,0.0,0.3444629,0.69073874,1.0352017,1.3796645,1.7241274,1.3996071,1.0750868,0.7505665,0.42423326,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.3444629,0.69073874,1.0352017,1.3796645,1.7241274,1.6352923,1.5446441,1.455809,1.3651608,1.2745126,1.0805258,0.88472575,0.69073874,0.4949388,0.2991388,0.28282216,0.26469254,0.24837588,0.23024625,0.21211663,0.48224804,0.7523795,1.0225109,1.2926424,1.5627737,3.5117085,5.462456,7.413204,9.362139,11.312886,9.791811,8.272549,6.7532854,5.23221,3.7129474,4.420003,5.127058,5.8341136,6.542982,7.250037,5.9918413,4.7354584,3.4772623,2.220879,0.96268314,0.8774739,0.79226464,0.7070554,0.62184614,0.53663695,0.54570174,0.5529536,0.56020546,0.56745726,0.5747091,0.49312583,0.40972954,0.32814622,0.24474995,0.16316663,0.13053331,0.09789998,0.065266654,0.032633327,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.04169814,0.059827764,0.07795739,0.09427405,0.11240368,0.19761293,0.28282216,0.3680314,0.45324063,0.53663695,0.57833505,0.61822027,0.65810543,0.6979906,0.73787576,0.7904517,0.8430276,0.89560354,0.9481794,1.0007553,1.2056202,1.4104849,1.6153497,1.8202144,2.0250793,2.0704033,2.1157274,2.1592383,2.2045624,2.2498865,3.159994,4.070101,4.9802084,5.8903155,6.8004227,6.0879283,5.375434,4.6629395,3.9504454,3.2379513,3.6766882,4.117238,4.557788,4.9983377,5.4370747,7.763106,10.087324,12.413355,14.737573,17.06179,22.06738,27.07297,32.07856,37.082336,42.087925,41.75253,41.41713,41.081734,40.748146,40.41275,34.85783,29.302914,23.747997,18.193079,12.638163,10.798005,8.957849,7.117691,5.277534,3.437377,3.6966307,3.9576974,4.216951,4.478018,4.7372713,4.880495,5.0219064,5.1651306,5.3083544,5.4497657,5.6945157,5.9392653,6.185828,6.430578,6.6753283,5.9682727,5.2594047,4.552349,3.8452935,3.1382382,3.0820365,3.0276475,2.9732587,2.9170568,2.8626678,2.6251698,2.3876717,2.1501737,1.9126755,1.6751775,1.4268016,1.1802386,0.9318628,0.6852999,0.43692398,0.50219065,0.56745726,0.6327239,0.6979906,0.76325727,0.8520924,0.94274056,1.0333886,1.1222239,1.2128719,1.017072,0.823085,0.62728506,0.43329805,0.2374981,0.20486477,0.17223145,0.13959812,0.10696479,0.07433146,0.06707962,0.059827764,0.052575916,0.045324065,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.045324065,0.052575916,0.059827764,0.06707962,0.07433146,0.06707962,0.059827764,0.052575916,0.045324065,0.038072214,0.15410182,0.27194437,0.38978696,0.5076295,0.62547207,1.1602961,1.69512,2.229944,2.764768,3.299592,2.955129,2.610666,2.2643902,1.9199274,1.5754645,1.7748904,1.9743162,2.175555,2.374981,2.5744069,4.4381323,6.300045,8.161958,10.025683,11.887595,9.947725,8.007855,6.0679855,4.1281157,2.1882458,2.764768,3.343103,3.919625,4.49796,5.0744824,4.4471974,3.8199122,3.1926272,2.565342,1.938057,2.762955,3.587853,4.4127507,5.237649,6.0625467,4.985647,3.9069343,2.8300345,1.7531348,0.6744221,1.7658255,2.855416,3.9450066,5.034597,6.1241875,7.0306687,7.935337,8.840006,9.744674,10.649343,9.440096,8.23085,7.019791,5.810545,4.599486,4.6393714,4.6792564,4.7191415,4.76084,4.800725,4.514277,4.229642,3.9450066,3.6603715,3.3757362,2.6995013,2.0250793,1.3506571,0.6744221,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.4224203,0.79589057,1.167548,1.5392052,1.9126755,1.5301404,1.1476053,0.7650702,0.3825351,0.0,0.17223145,0.3444629,0.5166943,0.69073874,0.8629702,0.96087015,1.0569572,1.1548572,1.2527572,1.3506571,1.0950294,0.83940166,0.5855869,0.32995918,0.07433146,0.09064813,0.10515183,0.11965553,0.13415924,0.15047589,0.4550536,0.75963134,1.064209,1.3705997,1.6751775,1.5156367,1.3542831,1.1947423,1.0352017,0.87566096,0.7904517,0.70524246,0.6200332,0.53482395,0.44961473,0.39703882,0.3444629,0.291887,0.23931105,0.18673515,0.21211663,0.2374981,0.26287958,0.28826106,0.31182957,0.3680314,0.4224203,0.47680917,0.533011,0.5873999,0.46955732,0.35171473,0.23568514,0.11784257,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.31182957,0.51306844,0.7124943,0.9119202,1.1131591,1.1802386,1.2473183,1.3143979,1.3832904,1.4503701,1.2219368,0.99531645,0.7668832,0.5402629,0.31182957,0.6508536,0.9880646,1.3252757,1.6624867,1.9996977,2.7103791,3.4192474,4.1299286,4.84061,5.5494785,5.4950895,5.4407005,5.384499,5.33011,5.275721,7.6778965,10.080072,12.482247,14.884423,17.286598,24.498564,31.706903,38.917053,46.12721,53.33736,50.219063,47.10258,43.984283,40.8678,37.749508,32.694965,27.640427,22.584074,17.529535,12.474996,11.234929,9.994863,8.754796,7.51473,6.2746634,5.7452784,5.2158933,4.6846952,4.15531,3.6241121,3.3521678,3.0802233,2.808279,2.5345216,2.2625773,1.9507477,1.6371052,1.3252757,1.0116332,0.69980353,1.0968424,1.4956942,1.892733,2.2897718,2.6868105,2.8481643,3.007705,3.1672456,3.3267863,3.48814,3.5352771,3.5824142,3.6295512,3.6766882,3.7256382,3.8978696,4.070101,4.2423325,4.4145637,4.5867953,5.130684,5.67276,6.2148356,6.7569118,7.3008003,7.02523,6.7496595,6.474089,6.200332,5.924762,5.7869763,5.6491914,5.5132194,5.375434,5.237649,5.368182,5.4969025,5.6274357,5.7579694,5.8866897,4.8224807,3.7582715,2.6922495,1.6280404,0.5620184,0.85934424,1.1566701,1.455809,1.7531348,2.0504606,2.6306088,3.2107568,3.7909048,4.36924,4.949388,4.4925213,4.0356545,3.576975,3.1201086,2.663242,2.857229,3.053029,3.247016,3.442816,3.636803,4.249584,4.8623657,5.475147,6.0879283,6.70071,7.7866745,8.874452,9.96223,11.050007,12.137785,13.515636,14.891675,16.269526,17.647377,19.025229,21.169964,23.3147,25.459433,27.604168,29.750715,34.85783,39.964947,45.072063,50.17918,55.288105,56.847256,58.408215,59.96736,61.526512,63.08747,60.03263,56.977787,53.922947,50.868103,47.813263,47.584827,47.358208,47.129776,46.903156,46.67472,46.897717,47.120712,47.341892,47.564888,47.78788,44.529987,41.272095,38.0142,34.758118,31.500225,29.879436,28.26046,26.639671,25.020697,23.399908,22.846954,22.295815,21.74286,21.189907,20.636953,18.992596,17.346426,15.702069,14.057712,12.413355,12.362592,12.311829,12.262879,12.212116,12.163166,12.66717,13.172986,13.67699,14.182806,14.68681,15.528025,16.367426,17.206827,18.048042,18.887444,16.831545,14.777458,12.721559,10.667472,8.613385,8.504607,8.397643,8.290678,8.1819,8.074935,7.3932614,6.7097745,6.0281005,5.3446136,4.6629395,4.168001,3.673062,3.1781235,2.6831846,2.1882458,2.0667772,1.9471219,1.8274662,1.7078108,1.5881553,1.2781386,0.968122,0.65810543,0.3480888,0.038072214,0.06707962,0.09789998,0.12690738,0.15772775,0.18673515,0.0,0.0,0.0,0.0,0.0,0.0,0.5166943,1.0352017,1.551896,2.0704033,2.5870976,2.0994108,1.6117238,1.1258497,0.63816285,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.23024625,0.4604925,0.69073874,0.91917205,1.1494182,1.0895905,1.0297627,0.969935,0.9101072,0.85027945,0.7197462,0.58921283,0.4604925,0.32995918,0.19942589,0.19217403,0.18492219,0.17767033,0.17041849,0.16316663,0.34264994,0.52213323,0.7016165,0.88291276,1.062396,3.5008307,5.9374523,8.375887,10.812509,13.24913,11.544946,9.840761,8.134763,6.430578,4.7245803,4.9675174,5.2104545,5.4533916,5.6945157,5.9374523,4.933071,3.926877,2.9224956,1.9181144,0.9119202,0.8466535,0.78319985,0.7179332,0.6526665,0.5873999,0.59283876,0.5982776,0.60190356,0.6073425,0.61278135,0.533011,0.45324063,0.37165734,0.291887,0.21211663,0.17041849,0.12690738,0.08520924,0.04169814,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.058014803,0.07795739,0.09789998,0.11784257,0.13778515,0.23931105,0.34264994,0.44417584,0.5475147,0.6508536,0.7106813,0.7705091,0.83033687,0.8901646,0.9499924,1.0478923,1.1457924,1.2418793,1.3397794,1.4376793,1.6080978,1.7767034,1.9471219,2.1175404,2.2879589,2.3169663,2.3477864,2.3767939,2.4076142,2.4366217,2.9768846,3.5171473,4.0574102,4.597673,5.137936,4.8242936,4.512464,4.2006345,3.8869917,3.5751622,3.923251,4.269527,4.6176157,4.9657044,5.3119802,8.26167,11.213174,14.162864,17.112555,20.062244,26.694061,33.32769,39.959507,46.59314,53.224957,50.58528,47.94561,45.304123,42.664448,40.024776,33.893337,27.760082,21.626831,15.495391,9.362139,8.05318,6.742408,5.431636,4.122677,2.811905,3.1146698,3.4174345,3.720199,4.022964,4.325729,4.5704784,4.8152285,5.0599785,5.3047285,5.5494785,5.5929894,5.634688,5.678199,5.719897,5.763408,5.0944247,4.4272547,3.7600844,3.092914,2.4257438,2.5544643,2.6849976,2.8155308,2.9442513,3.0747845,2.9007401,2.7248828,2.5508385,2.374981,2.1991236,1.8600996,1.5192627,1.1802386,0.83940166,0.50037766,0.5094425,0.52032024,0.5293851,0.5402629,0.5493277,0.6091554,0.67079616,0.7306239,0.7904517,0.85027945,0.7197462,0.58921283,0.4604925,0.32995918,0.19942589,0.18310922,0.16497959,0.14684997,0.13053331,0.11240368,0.09427405,0.07795739,0.059827764,0.04169814,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.030820364,0.034446288,0.03988518,0.045324065,0.05076295,0.045324065,0.03988518,0.034446288,0.030820364,0.025381476,0.19579996,0.36440548,0.53482395,0.70524246,0.87566096,1.452183,2.030518,2.6070402,3.1853752,3.7618973,3.3576066,2.953316,2.5472124,2.1429217,1.7368182,1.7368182,1.7368182,1.7368182,1.7368182,1.7368182,4.1498713,6.5629244,8.974165,11.3872175,13.800271,11.352772,8.9052725,6.4577727,4.0102735,1.5627737,2.6976883,3.832603,4.9675174,6.1024323,7.2373466,6.051669,4.8678045,3.682127,2.4982624,1.3125849,2.5997884,3.8869917,5.1741953,6.4632115,7.750415,6.3145485,4.880495,3.444629,2.0105755,0.5747091,1.3724127,2.1701162,2.9678197,3.7655232,4.5632267,5.7072062,6.8529987,7.996978,9.142771,10.28675,9.547061,8.807372,8.067683,7.327995,6.588306,6.1967063,5.806919,5.4171324,5.027345,4.6375585,4.160749,3.682127,3.2053177,2.7266958,2.2498865,1.8002719,1.3506571,0.89922947,0.44961473,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.32814622,0.58014804,0.8321498,1.0841516,1.3379664,1.0696479,0.8031424,0.53482395,0.26831847,0.0,0.11421664,0.23024625,0.3444629,0.4604925,0.5747091,0.86478317,1.1548572,1.4449311,1.7350051,2.0250793,1.6298534,1.2346275,0.83940166,0.44417584,0.05076295,0.08520924,0.11965553,0.15410182,0.19036107,0.22480737,0.40791658,0.58921283,0.77232206,0.9554313,1.1367276,1.1602961,1.1820517,1.2056202,1.2273756,1.2491312,1.0605831,0.87022203,0.67986095,0.4894999,0.2991388,0.26469254,0.23024625,0.19579996,0.15954071,0.12509441,0.18673515,0.25018883,0.31182957,0.37528324,0.43692398,0.46955732,0.50219065,0.53482395,0.56745726,0.6000906,0.48043507,0.36077955,0.23931105,0.11965553,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.22480737,0.37528324,0.52575916,0.6744221,0.824898,0.90829426,0.9898776,1.0732739,1.1548572,1.2382535,1.0768998,0.91735905,0.75781834,0.5982776,0.43692398,0.63816285,0.8375887,1.0370146,1.2382535,1.4376793,2.0522738,2.666868,3.2832751,3.8978696,4.512464,4.5668526,4.6230545,4.6774435,4.7318325,4.788034,6.2220874,7.6579537,9.092008,10.527874,11.961927,17.052727,22.141712,27.232512,32.32331,37.412296,35.104393,32.798306,30.490404,28.182503,25.874601,23.316511,20.760235,18.202145,15.645867,13.087777,12.027194,10.968424,9.907841,8.847258,7.7866745,7.066928,6.347182,5.6274357,4.9076896,4.1879435,3.7600844,3.3322253,2.904366,2.47832,2.0504606,1.7368182,1.4249886,1.1131591,0.7995165,0.48768693,1.0768998,1.6679256,2.2571385,2.8481643,3.437377,3.489953,3.5425289,3.5951047,3.6476808,3.7002566,3.7020695,3.7056956,3.7075086,3.7093215,3.7129474,3.877927,4.0429068,4.207886,4.3728657,4.537845,5.145188,5.75253,6.359873,6.967215,7.574558,7.1992745,6.825804,6.450521,6.0752378,5.6999545,5.4497657,5.199577,4.949388,4.699199,4.4508233,4.606738,4.764466,4.9221935,5.0799212,5.237649,4.314851,3.392053,2.469255,1.54827,0.62547207,0.92823684,1.2291887,1.5319533,1.8347181,2.137483,2.4819458,2.8282216,3.1726844,3.5171473,3.8616104,3.4953918,3.1273603,2.759329,2.3931105,2.0250793,2.179181,2.335096,2.4891977,2.6451125,2.7992141,3.4627585,4.12449,4.788034,5.4497657,6.11331,6.7623506,7.413204,8.062244,8.713099,9.362139,10.473485,11.583018,12.692551,13.802084,14.91343,17.429823,19.948027,22.464418,24.982624,27.50083,31.492973,35.485115,39.47726,43.469402,47.46336,49.278137,51.09291,52.90769,54.72246,56.53724,55.529232,54.523037,53.51503,52.507023,51.500828,49.827465,48.15591,46.482548,44.810997,43.13763,42.252907,41.36818,40.48164,39.596916,38.71219,36.658104,34.602203,32.54812,30.492218,28.438131,27.444628,26.452936,25.459433,24.467743,23.47424,23.85315,24.230246,24.607342,24.984438,25.363346,23.207733,21.052122,18.89651,16.74271,14.587097,14.336908,14.0867195,13.838344,13.588155,13.337966,14.857228,16.378304,17.897566,19.41683,20.937904,21.273302,21.606888,21.942286,22.277683,22.613083,20.392202,18.171324,15.952258,13.7331915,11.512312,10.694666,9.87702,9.059374,8.241728,7.4258947,6.782293,6.1405044,5.4969025,4.855114,4.213325,3.682127,3.152742,2.6233568,2.0921588,1.5627737,1.4830034,1.403233,1.3216497,1.2418793,1.162109,0.9354887,0.7070554,0.48043507,0.2520018,0.025381476,0.045324065,0.065266654,0.08520924,0.10515183,0.12509441,0.0,0.0,0.0,0.0,0.0,0.0,0.69073874,1.3796645,2.0704033,2.759329,3.4500678,2.7992141,2.1501737,1.49932,0.85027945,0.19942589,0.15954071,0.11965553,0.07977036,0.03988518,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.11421664,0.23024625,0.3444629,0.4604925,0.5747091,0.54570174,0.5148814,0.48587397,0.4550536,0.42423326,0.36077955,0.2955129,0.23024625,0.16497959,0.099712946,0.10333887,0.10515183,0.10696479,0.11059072,0.11240368,0.2030518,0.291887,0.3825351,0.47318324,0.5620184,3.48814,6.412449,9.336758,12.262879,15.187187,13.29808,11.407161,9.518054,7.6271334,5.7380266,5.5150323,5.292038,5.0708566,4.847862,4.6248674,3.872488,3.1201086,2.3677292,1.6153497,0.8629702,0.81764615,0.77232206,0.726998,0.68167394,0.63816285,0.6399758,0.6417888,0.64541465,0.64722764,0.6508536,0.5728962,0.4949388,0.4169814,0.34083697,0.26287958,0.21030366,0.15772775,0.10515183,0.052575916,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.072518505,0.09427405,0.11784257,0.13959812,0.16316663,0.28282216,0.40247768,0.52213323,0.6417888,0.76325727,0.8430276,0.922798,1.0025684,1.0823387,1.162109,1.305333,1.4467441,1.5899682,1.7331922,1.8746033,2.0105755,2.1447346,2.280707,2.4148662,2.5508385,2.565342,2.5798457,2.5943494,2.610666,2.6251698,2.7955883,2.9641938,3.1346123,3.3050308,3.4754493,3.5624714,3.6494937,3.738329,3.825351,3.9123733,4.168001,4.421816,4.6774435,4.933071,5.186886,8.762048,12.337211,15.912373,19.487535,23.062696,31.322554,39.582413,47.84227,56.102127,64.361984,59.418037,54.472275,49.526512,44.58256,39.636803,32.927025,26.217253,19.507477,12.797703,6.0879283,5.3083544,4.5269675,3.7473936,2.9678197,2.1882458,2.5327086,2.8771715,3.2216346,3.5679104,3.9123733,4.2604623,4.606738,4.954827,5.3029156,5.6491914,5.4896507,5.33011,5.1705694,5.009216,4.8496747,4.2223897,3.5951047,2.9678197,2.3405347,1.7132497,2.0268922,2.3423476,2.657803,2.9732587,3.2869012,3.1744974,3.0620937,2.94969,2.8372865,2.7248828,2.2933977,1.8600996,1.4268016,0.99531645,0.5620184,0.5166943,0.47318324,0.42785916,0.3825351,0.33721104,0.3680314,0.39703882,0.42785916,0.45686656,0.48768693,0.4224203,0.35715362,0.291887,0.22662032,0.16316663,0.15954071,0.15772775,0.15410182,0.15228885,0.15047589,0.12328146,0.09427405,0.06707962,0.03988518,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.014503701,0.018129626,0.01994259,0.02175555,0.025381476,0.02175555,0.01994259,0.018129626,0.014503701,0.012690738,0.23568514,0.45686656,0.67986095,0.90285534,1.1258497,1.745883,2.3641033,2.9841363,3.6041696,4.2242026,3.7600844,3.294153,2.8300345,2.3641033,1.8999848,1.7005589,1.49932,1.2998942,1.1004683,0.89922947,3.8616104,6.825804,9.788185,12.750566,15.712947,12.757817,9.802689,6.8475595,3.8924308,0.93730164,2.6306088,4.322103,6.01541,7.706904,9.400211,7.6579537,5.915697,4.171627,2.42937,0.6871128,2.4384346,4.1879435,5.9374523,7.686961,9.438283,7.645263,5.8522434,4.059223,2.268016,0.4749962,0.9808127,1.4848163,1.9906329,2.4946365,3.000453,4.3855567,5.77066,7.155763,8.540867,9.924157,9.655839,9.385707,9.115576,8.845445,8.575313,7.755854,6.9345818,6.115123,5.295664,4.4743915,3.8054085,3.1346123,2.465629,1.794833,1.1258497,0.89922947,0.6744221,0.44961473,0.22480737,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.23205921,0.36440548,0.49675176,0.629098,0.76325727,0.6091554,0.45686656,0.3045777,0.15228885,0.0,0.058014803,0.11421664,0.17223145,0.23024625,0.28826106,0.7705091,1.2527572,1.7350051,2.2172532,2.6995013,2.1646774,1.6298534,1.0950294,0.56020546,0.025381476,0.07977036,0.13415924,0.19036107,0.24474995,0.2991388,0.36077955,0.42060733,0.48043507,0.5402629,0.6000906,0.80495536,1.0098201,1.214685,1.4195497,1.6244144,1.3307146,1.0352017,0.73968875,0.44417584,0.15047589,0.13234627,0.11421664,0.09789998,0.07977036,0.06164073,0.16316663,0.26287958,0.36259252,0.46230546,0.5620184,0.5728962,0.581961,0.59283876,0.60190356,0.61278135,0.4894999,0.3680314,0.24474995,0.12328146,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.13778515,0.2374981,0.33721104,0.43692398,0.53663695,0.6345369,0.7324369,0.83033687,0.92823684,1.0243238,0.9318628,0.83940166,0.7469406,0.6544795,0.5620184,0.62547207,0.6871128,0.7505665,0.8122072,0.87566096,1.3941683,1.9144884,2.4348087,2.955129,3.4754493,3.6404288,3.8054085,3.9703882,4.135368,4.3003473,4.7680917,5.235836,5.7017674,6.169512,6.637256,9.606889,12.576522,15.547967,18.5176,21.487232,19.989725,18.492218,16.99471,15.497204,13.999697,13.939869,13.880041,13.820213,13.760386,13.700559,12.819458,11.940171,11.060884,10.179785,9.300498,8.39039,7.4802837,6.5701766,5.660069,4.749962,4.168001,3.584227,3.002266,2.420305,1.8383441,1.5247015,1.2128719,0.89922947,0.5873999,0.2755703,1.0569572,1.840157,2.6233568,3.4047437,4.1879435,4.1317415,4.077353,4.022964,3.966762,3.9123733,3.870675,3.827164,3.785466,3.7419548,3.7002566,3.8579843,4.0157123,4.171627,4.329355,4.4870825,5.1596913,5.8323007,6.5049095,7.177519,7.850128,7.3751316,6.9001355,6.4251394,5.9501433,5.475147,5.1125546,4.749962,4.3873696,4.024777,3.6621845,3.8471067,4.0320287,4.216951,4.401873,4.5867953,3.8072214,3.0276475,2.2480736,1.4666867,0.6871128,0.99531645,1.3017071,1.6099107,1.9181144,2.2245052,2.335096,2.4456866,2.5544643,2.665055,2.7756457,2.4982624,2.220879,1.9416829,1.6642996,1.3869164,1.502946,1.6171626,1.7331922,1.8474089,1.9616255,2.675933,3.386614,4.099108,4.8116026,5.524097,5.7380266,5.9501433,6.16226,6.3743763,6.588306,7.4295206,8.272549,9.115576,9.956791,10.799818,13.68968,16.579542,19.469404,22.359268,25.24913,28.128115,31.005285,33.882458,36.75963,39.636803,41.707203,43.777607,45.84801,47.9166,49.987003,51.027645,52.068287,53.107113,54.147755,55.188393,52.0701,48.9518,45.83532,42.717026,39.60054,37.608097,35.61565,33.623203,31.630758,29.6365,28.784407,27.932314,27.080221,26.22813,25.374224,25.009819,24.645412,24.279196,23.91479,23.550385,24.85753,26.164677,27.471823,28.78078,30.087927,27.422873,24.757816,22.092762,19.427708,16.762651,16.313038,15.861609,15.411995,14.96238,14.512766,17.047287,19.583622,22.118143,24.652666,27.187187,27.016768,26.848164,26.677744,26.507326,26.336908,23.952862,21.567003,19.182957,16.797098,14.413053,12.884725,11.358211,9.829884,8.303369,6.775041,6.1731377,5.569421,4.9675174,4.365614,3.7618973,3.198066,2.6324217,2.0667772,1.502946,0.93730164,0.8974165,0.8575313,0.81764615,0.7777609,0.73787576,0.59283876,0.44780177,0.30276474,0.15772775,0.012690738,0.02175555,0.032633327,0.04169814,0.052575916,0.06164073,0.0,0.0,0.0,0.0,0.0,0.0,0.8629702,1.7241274,2.5870976,3.4500678,4.313038,3.5008307,2.6868105,1.8746033,1.062396,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,3.4754493,6.887445,10.29944,13.713249,17.125244,15.049402,12.975373,10.899531,8.825501,6.7496595,6.0625467,5.375434,4.688321,3.9993954,3.3122826,2.811905,2.3133402,1.8129625,1.3125849,0.8122072,0.7868258,0.76325727,0.73787576,0.7124943,0.6871128,0.6871128,0.6871128,0.6871128,0.6871128,0.6871128,0.61278135,0.53663695,0.46230546,0.387974,0.31182957,0.25018883,0.18673515,0.12509441,0.06164073,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.0870222,0.11240368,0.13778515,0.16316663,0.18673515,0.3245203,0.46230546,0.6000906,0.73787576,0.87566096,0.97537386,1.0750868,1.1747998,1.2745126,1.3742256,1.5627737,1.7495089,1.938057,2.124792,2.3133402,2.4130533,2.5127661,2.612479,2.712192,2.811905,2.811905,2.811905,2.811905,2.811905,2.811905,2.612479,2.4130533,2.2118144,2.0123885,1.8129625,2.3006494,2.7883365,3.2742105,3.7618973,4.249584,4.4127507,4.574105,4.7372713,4.900438,5.0617914,9.262425,13.46306,17.661882,21.862516,26.06315,35.949234,45.83713,55.72503,65.61293,75.500824,68.250786,61.00075,53.7489,46.50068,39.25064,31.96253,24.674421,17.388124,10.100015,2.811905,2.561716,2.3133402,2.0631514,1.8129625,1.5627737,1.9507477,2.3369088,2.7248828,3.1128569,3.5008307,3.9504454,4.40006,4.8496747,5.2992897,5.750717,5.388125,5.0255322,4.6629395,4.3003473,3.9377546,3.350355,2.762955,2.175555,1.5881553,1.0007553,1.49932,1.9996977,2.5000753,3.000453,3.5008307,3.4500678,3.3993049,3.350355,3.299592,3.2506418,2.7248828,2.1991236,1.6751775,1.1494182,0.62547207,0.52575916,0.42423326,0.3245203,0.22480737,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.13778515,0.15047589,0.16316663,0.17585737,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.2755703,0.5493277,0.824898,1.1004683,1.3742256,2.03777,2.6995013,3.3630457,4.024777,4.688321,4.162562,3.636803,3.1128569,2.5870976,2.0631514,1.6624867,1.261822,0.8629702,0.46230546,0.06164073,3.5751622,7.0868707,10.600392,14.112101,17.625622,14.162864,10.700105,7.2373466,3.774588,0.31182957,2.561716,4.8116026,7.063302,9.313189,11.563075,9.262425,6.9617763,4.6629395,2.3622901,0.06164073,2.275268,4.4870825,6.70071,8.912524,11.124338,8.974165,6.825804,4.6756306,2.525457,0.37528324,0.5873999,0.7995165,1.0116332,1.2255627,1.4376793,3.0620937,4.688321,6.3127356,7.93715,9.563377,9.762803,9.96223,10.161655,10.362894,10.56232,9.313189,8.062244,6.813113,5.562169,4.313038,3.4500678,2.5870976,1.7241274,0.8629702,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.13778515,0.15047589,0.16316663,0.17585737,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.0,0.0,0.0,0.0,0.0,0.6744221,1.3506571,2.0250793,2.6995013,3.3757362,2.6995013,2.0250793,1.3506571,0.6744221,0.0,0.07433146,0.15047589,0.22480737,0.2991388,0.37528324,0.31182957,0.25018883,0.18673515,0.12509441,0.06164073,0.44961473,0.8375887,1.2255627,1.6117238,1.9996977,1.6008459,1.2001812,0.7995165,0.40066472,0.0,0.0,0.0,0.0,0.0,0.0,0.13778515,0.2755703,0.41335547,0.5493277,0.6871128,0.6744221,0.66173136,0.6508536,0.63816285,0.62547207,0.50037766,0.37528324,0.25018883,0.12509441,0.0,0.0,0.0,0.0,0.0,0.0,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,0.36259252,0.4749962,0.5873999,0.69980353,0.8122072,0.7868258,0.76325727,0.73787576,0.7124943,0.6871128,0.61278135,0.53663695,0.46230546,0.387974,0.31182957,0.73787576,1.162109,1.5881553,2.0123885,2.4366217,2.712192,2.9877625,3.2633326,3.53709,3.8126602,3.3122826,2.811905,2.3133402,1.8129625,1.3125849,2.1628644,3.0131438,3.8634233,4.7118897,5.562169,4.8750563,4.1879435,3.5008307,2.811905,2.124792,4.5632267,6.9998484,9.438283,11.874905,14.313339,13.611723,12.91192,12.212116,11.512312,10.812509,9.712041,8.613385,7.512917,6.412449,5.3119802,4.574105,3.8380418,3.100166,2.3622901,1.6244144,1.3125849,1.0007553,0.6871128,0.37528324,0.06164073,1.0370146,2.0123885,2.9877625,3.9631362,4.936697,4.7753434,4.612177,4.4508233,4.2876563,4.12449,4.0374675,3.9504454,3.8616104,3.774588,3.6875658,3.8380418,3.9867048,4.137181,4.2876563,4.4381323,5.1741953,5.9120708,6.6499467,7.3878226,8.125698,7.549176,6.9744673,6.399758,5.825049,5.2503395,4.7753434,4.3003473,3.825351,3.350355,2.8753586,3.0874753,3.299592,3.5117085,3.7256382,3.9377546,3.299592,2.663242,2.0250793,1.3869164,0.7505665,1.062396,1.3742256,1.6878681,1.9996977,2.3133402,2.1882458,2.0631514,1.938057,1.8129625,1.6878681,1.49932,1.3125849,1.1258497,0.93730164,0.7505665,0.824898,0.89922947,0.97537386,1.0497054,1.1258497,1.887294,2.6505513,3.4119956,4.175253,4.936697,4.7118897,4.4870825,4.262275,4.0374675,3.8126602,4.3873696,4.9620786,5.5367875,6.11331,6.688019,9.949538,13.212872,16.474392,19.737724,22.999243,24.763256,26.525455,28.287655,30.049854,31.812054,34.138084,36.462303,38.788334,41.112553,43.43677,46.52606,49.61172,52.699196,55.78667,58.874146,54.312733,49.749508,45.18809,40.624866,36.061638,32.96147,29.86312,26.762953,23.662788,20.562622,20.912523,21.262424,21.612328,21.962229,22.31213,22.57501,22.837889,23.100769,23.361835,23.624716,25.861912,28.10092,30.338116,32.575314,34.812508,31.63801,28.4617,25.287203,22.112705,18.938208,18.287354,17.638313,16.98746,16.338419,15.687565,19.237347,22.787127,26.336908,29.886688,33.438282,32.762047,32.087624,31.413202,30.736967,30.062546,27.511707,24.962683,22.411844,19.862818,17.31198,15.074784,12.837588,10.600392,8.363196,6.1241875,5.562169,5.0001507,4.4381323,3.874301,3.3122826,2.712192,2.1121013,1.5120108,0.9119202,0.31182957,0.31182957,0.31182957,0.31182957,0.31182957,0.31182957,0.25018883,0.18673515,0.12509441,0.06164073,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.69255173,1.3851035,2.077655,2.770207,3.4627585,2.8155308,2.1683033,1.5192627,0.872035,0.22480737,0.1794833,0.13415924,0.09064813,0.045324065,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.0870222,0.16316663,0.2374981,0.31182957,0.387974,0.31182957,0.2374981,0.16316663,0.0870222,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,0.24474995,0.23931105,0.23568514,0.23024625,0.22480737,2.9406252,5.65463,8.370448,11.084454,13.800271,12.335398,10.870523,9.40565,7.9407763,6.474089,5.870373,5.2648435,4.6593137,4.0555973,3.4500678,2.9351864,2.420305,1.9054236,1.3905423,0.87566096,0.83940166,0.80495536,0.7705091,0.73424983,0.69980353,0.67986095,0.65991837,0.6399758,0.6200332,0.6000906,0.54570174,0.4894999,0.43511102,0.38072214,0.3245203,0.35534066,0.38434806,0.41516843,0.44417584,0.4749962,0.40066472,0.3245203,0.25018883,0.17585737,0.099712946,0.14322405,0.18492219,0.22662032,0.27013144,0.31182957,0.43692398,0.5620184,0.6871128,0.8122072,0.93730164,1.1331016,1.3270886,1.5228885,1.7168756,1.9126755,1.9181144,1.9217403,1.9271792,1.9326181,1.938057,2.0250793,2.1121013,2.1991236,2.2879589,2.374981,2.4891977,2.6052272,2.7194438,2.8354735,2.94969,3.056655,3.1654327,3.2723975,3.3793623,3.48814,3.9069343,4.327542,4.748149,5.1669436,5.5875506,5.6274357,5.667321,5.7072062,5.7470913,5.7869763,9.202598,12.618219,16.032028,19.447649,22.863272,30.807673,38.752075,46.69829,54.642693,62.587093,56.578938,50.57259,44.564434,38.558086,32.54993,26.715816,20.87989,15.043963,9.20985,3.3757362,3.2506418,3.1255474,3.000453,2.8753586,2.7502642,3.2723975,3.7945306,4.3166637,4.84061,5.3627434,5.52591,5.6872635,5.8504305,6.011784,6.1749506,5.7344007,5.295664,4.855114,4.4145637,3.975827,3.4192474,2.864481,2.3097143,1.7549478,1.2001812,1.6117238,2.0250793,2.4366217,2.8499773,3.2633326,4.0030212,4.74271,5.482399,6.2220874,6.9617763,6.3743763,5.7869763,5.199577,4.612177,4.024777,3.388427,2.7502642,2.1121013,1.4757515,0.8375887,0.69073874,0.5420758,0.39522585,0.24837588,0.099712946,0.099712946,0.099712946,0.099712946,0.099712946,0.099712946,0.11059072,0.11965553,0.13053331,0.13959812,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.09427405,0.07795739,0.059827764,0.04169814,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.24837588,0.4949388,0.7433147,0.9898776,1.2382535,1.9199274,2.6016014,3.2850883,3.966762,4.650249,4.552349,4.454449,4.358362,4.2604623,4.162562,3.339477,2.518205,1.69512,0.872035,0.05076295,2.859042,5.669134,8.479226,11.289318,14.09941,11.332829,8.564435,5.7978544,3.0294604,0.26287958,2.1501737,4.0374675,5.924762,7.8120556,9.699349,7.7921133,5.8848767,3.97764,2.0704033,0.16316663,2.675933,5.186886,7.699652,10.212419,12.725184,10.417283,8.109382,5.803293,3.4953918,1.1874905,1.4503701,1.7132497,1.9743162,2.2371957,2.5000753,3.53709,4.574105,5.612932,6.6499467,7.686961,8.272549,8.858135,9.441909,10.027496,10.613083,9.179029,7.746789,6.3145485,4.882308,3.4500678,2.759329,2.0704033,1.3796645,0.69073874,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.11059072,0.11965553,0.13053331,0.13959812,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.0,0.0,0.0,0.0,0.0,0.5402629,1.0805258,1.6207886,2.1592383,2.6995013,2.1592383,1.6207886,1.0805258,0.5402629,0.0,0.06707962,0.13415924,0.2030518,0.27013144,0.33721104,0.28826106,0.2374981,0.18673515,0.13778515,0.0870222,0.40791658,0.726998,1.0478923,1.3669738,1.6878681,1.4376793,1.1874905,0.93730164,0.6871128,0.43692398,0.40791658,0.3770962,0.3480888,0.31726846,0.28826106,0.6345369,0.9826257,1.3307146,1.6769904,2.0250793,1.7205015,1.4159238,1.1095331,0.80495536,0.50037766,0.40066472,0.2991388,0.19942589,0.099712946,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.13053331,0.24837588,0.36440548,0.48224804,0.6000906,0.7016165,0.80495536,0.90829426,1.0098201,1.1131591,1.1059072,1.0968424,1.0895905,1.0823387,1.0750868,0.9101072,0.7451276,0.58014804,0.41516843,0.25018883,0.6345369,1.020698,1.405046,1.789394,2.175555,2.3495996,2.525457,2.6995013,2.8753586,3.049403,2.6505513,2.2498865,1.8492218,1.4503701,1.0497054,1.7295663,2.4094272,3.0892882,3.7691493,4.4508233,3.8996825,3.350355,2.7992141,2.2498865,1.7005589,3.6494937,5.600241,7.549176,9.499924,11.450671,11.519565,11.59027,11.6591625,11.729868,11.800573,10.3502035,8.899834,7.4494634,5.999093,4.550536,4.1408067,3.729264,3.3195345,2.909805,2.5000753,2.7974012,3.094727,3.392053,3.6893787,3.9867048,4.3909955,4.7916603,5.195951,5.5984282,6.000906,5.6528172,5.3047285,4.95664,4.610364,4.262275,4.249584,4.2368937,4.2242026,4.213325,4.2006345,4.459888,4.7191415,4.9802084,5.239462,5.5005283,6.4033837,7.304426,8.207282,9.110137,10.012992,9.402024,8.792869,8.1819,7.572745,6.9617763,6.294606,5.6274357,4.9602656,4.2930956,3.6241121,3.584227,3.5443418,3.5044568,3.4645715,3.4246864,3.0693457,2.715818,2.3604772,2.0051367,1.649796,1.7241274,1.8002719,1.8746033,1.9507477,2.0250793,1.9108626,1.794833,1.6806163,1.5645868,1.4503701,1.3270886,1.2056202,1.0823387,0.96087015,0.8375887,0.8520924,0.8665961,0.88291276,0.8974165,0.9119202,1.5192627,2.126605,2.7357605,3.343103,3.9504454,3.7727752,3.5951047,3.4174345,3.2397642,3.0620937,3.6241121,4.1879435,4.749962,5.3119802,5.8758116,8.582565,11.289318,13.997884,16.704638,19.413204,21.402023,23.392656,25.38329,27.372108,29.362741,31.492973,33.623203,35.75162,37.881855,40.012085,42.588303,45.162712,47.737118,50.311523,52.887745,49.584526,46.283123,42.979904,39.678497,36.375282,33.74286,31.110437,28.478016,25.845594,23.213173,23.002869,22.792566,22.582262,22.371958,22.161655,22.23236,22.303066,22.371958,22.442663,22.513369,24.112402,25.71325,27.31228,28.913128,30.51216,27.959509,25.406858,22.854206,20.303368,17.750717,17.357304,16.965704,16.57229,16.18069,15.787278,18.709774,21.632269,24.554766,27.47726,30.399757,29.754341,29.11074,28.465326,27.81991,27.174496,25.602657,24.029007,22.457167,20.885328,19.311678,17.059978,14.806465,12.554766,10.303066,8.049554,6.972654,5.8957543,4.8170414,3.7401419,2.663242,2.1918716,1.7223145,1.2527572,0.78319985,0.31182957,0.2991388,0.28826106,0.2755703,0.26287958,0.25018883,0.20486477,0.15954071,0.11421664,0.07070554,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.52213323,1.0442665,1.5682126,2.0903459,2.612479,2.1302311,1.647983,1.1657349,0.68167394,0.19942589,0.15954071,0.11965553,0.07977036,0.03988518,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.17585737,0.3245203,0.4749962,0.62547207,0.774135,0.62547207,0.4749962,0.3245203,0.17585737,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0870222,0.17585737,0.26287958,0.34990177,0.43692398,0.42785916,0.4169814,0.40791658,0.39703882,0.387974,2.4058013,4.421816,6.439643,8.457471,10.475298,9.619579,8.765674,7.909956,7.0542374,6.200332,5.678199,5.1542525,4.632119,4.1099863,3.587853,3.056655,2.5272698,1.9978848,1.4666867,0.93730164,0.8919776,0.8466535,0.8031424,0.75781834,0.7124943,0.6726091,0.6327239,0.59283876,0.5529536,0.51306844,0.47680917,0.44236287,0.40791658,0.37165734,0.33721104,0.4604925,0.581961,0.70524246,0.82671094,0.9499924,0.7868258,0.62547207,0.46230546,0.2991388,0.13778515,0.19761293,0.2574407,0.31726846,0.3770962,0.43692398,0.5493277,0.66173136,0.774135,0.8883517,1.0007553,1.2908293,1.5790904,1.8691645,2.1592383,2.4493124,2.2716422,2.0957847,1.9181144,1.7404441,1.5627737,1.6371052,1.7132497,1.7875811,1.8619126,1.938057,2.1683033,2.3967366,2.6269827,2.857229,3.0874753,3.5026438,3.917812,4.3329806,4.748149,5.163317,5.5150323,5.866747,6.2202744,6.5719895,6.925517,6.8421206,6.7605376,6.677141,6.5955577,6.5121617,9.142771,11.771566,14.402175,17.032784,19.66158,25.664299,31.667017,37.669735,43.672455,49.675175,44.91071,40.144432,35.379963,30.6155,25.84922,21.46729,17.08536,12.701616,8.319685,3.9377546,3.9377546,3.9377546,3.9377546,3.9377546,3.9377546,4.59586,5.2521524,5.910258,6.5683637,7.224656,7.0995617,6.9744673,6.849373,6.7242785,6.599184,6.0824895,5.565795,5.047288,4.5305934,4.0120864,3.489953,2.9678197,2.4456866,1.9217403,1.3996071,1.7241274,2.0504606,2.374981,2.6995013,3.0258346,4.554162,6.0843024,7.614443,9.144584,10.674724,10.025683,9.374829,8.725789,8.074935,7.4258947,6.249282,5.0744824,3.8996825,2.7248828,1.550083,1.2545701,0.96087015,0.6653573,0.36984438,0.07433146,0.07433146,0.07433146,0.07433146,0.07433146,0.07433146,0.08339628,0.09064813,0.09789998,0.10515183,0.11240368,0.09064813,0.06707962,0.045324065,0.02175555,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.045324065,0.09064813,0.13415924,0.1794833,0.22480737,0.19036107,0.15410182,0.11965553,0.08520924,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.21936847,0.4405499,0.65991837,0.8792868,1.1004683,1.8020848,2.5055144,3.207131,3.9105604,4.612177,4.942136,5.272095,5.6020546,5.9320135,6.261973,5.0182805,3.7727752,2.5272698,1.2817645,0.038072214,2.1447346,4.25321,6.359873,8.4683485,10.57501,8.502794,6.430578,4.3565493,2.2843328,0.21211663,1.7368182,3.2633326,4.788034,6.3127356,7.837437,6.3218007,4.8079767,3.29234,1.7767034,0.26287958,3.0747845,5.8866897,8.700407,11.512312,14.324218,11.860401,9.394773,6.929143,4.465327,1.9996977,2.3133402,2.6251698,2.9369993,3.2506418,3.5624714,4.0120864,4.461701,4.9131284,5.3627434,5.812358,6.782293,7.752228,8.722163,9.692098,10.662033,9.046683,7.4331465,5.8177967,4.2024474,2.5870976,2.0704033,1.551896,1.0352017,0.5166943,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.08339628,0.09064813,0.09789998,0.10515183,0.11240368,0.09064813,0.06707962,0.045324065,0.02175555,0.0,0.0,0.0,0.0,0.0,0.0,0.40429065,0.8103943,1.214685,1.6207886,2.0250793,1.6207886,1.214685,0.8103943,0.40429065,0.0,0.059827764,0.11965553,0.1794833,0.23931105,0.2991388,0.26287958,0.22480737,0.18673515,0.15047589,0.11240368,0.36440548,0.61822027,0.87022203,1.1222239,1.3742256,1.2745126,1.1747998,1.0750868,0.97537386,0.87566096,0.81583315,0.7541924,0.69436467,0.6345369,0.5747091,1.1331016,1.6896812,2.2480736,2.8046532,3.3630457,2.764768,2.1683033,1.5700256,0.97174793,0.37528324,0.2991388,0.22480737,0.15047589,0.07433146,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.21030366,0.39522585,0.58014804,0.7650702,0.9499924,1.0424535,1.1349145,1.2273756,1.3198367,1.4122978,1.4231756,1.4322405,1.4431182,1.452183,1.4630609,1.2074331,0.95180535,0.6979906,0.44236287,0.18673515,0.533011,0.8774739,1.2219368,1.5682126,1.9126755,1.987007,2.0631514,2.137483,2.2118144,2.2879589,1.987007,1.6878681,1.3869164,1.0877775,0.7868258,1.2980812,1.8075237,2.3169663,2.8282216,3.3376641,2.9243085,2.5127661,2.0994108,1.6878681,1.2745126,2.7375734,4.2006345,5.661882,7.124943,8.588004,9.427405,10.266808,11.108022,11.947423,12.786825,10.986553,9.188094,7.3878226,5.5875506,3.787279,3.7056956,3.6222992,3.540716,3.4573197,3.3757362,4.2822175,5.1905117,6.096993,7.0052876,7.911769,7.743163,7.572745,7.402326,7.231908,7.063302,6.530291,5.99728,5.464269,4.933071,4.40006,4.461701,4.5251546,4.5867953,4.650249,4.7118897,5.081734,5.4533916,5.823236,6.19308,6.5629244,7.6307597,8.696781,9.764616,10.832452,11.900287,11.254871,10.609457,9.965856,9.32044,8.675026,7.8156815,6.9545245,6.09518,5.235836,4.3746786,4.082792,3.7909048,3.4972048,3.2053177,2.911618,2.8390994,2.7683938,2.6958754,2.6233568,2.5508385,2.3876717,2.2245052,2.0631514,1.8999848,1.7368182,1.6316663,1.5283275,1.4231756,1.3180238,1.2128719,1.1548572,1.0968424,1.0406405,0.9826257,0.9246109,0.8792868,0.83577573,0.7904517,0.7451276,0.69980353,1.1530442,1.6044719,2.0577126,2.5091403,2.962381,2.8318477,2.7031271,2.572594,2.4420607,2.3133402,2.8626678,3.4119956,3.9631362,4.512464,5.0617914,7.215591,9.367578,11.519565,13.671551,15.825351,18.042604,20.259857,22.47711,24.694363,26.911617,28.84786,30.782291,32.716724,34.652966,36.5874,38.65055,40.711887,42.77504,44.838192,46.89953,44.85813,42.814926,40.771717,38.73032,36.68711,34.522434,32.357758,30.193079,28.028402,25.861912,25.093216,24.322706,23.552197,22.781689,22.01299,21.88971,21.768242,21.64496,21.521679,21.40021,22.362894,23.325577,24.28826,25.24913,26.211813,24.282822,22.352016,20.423023,18.492218,16.563227,16.427254,16.293095,16.157122,16.022963,15.8869915,18.182201,20.477413,22.772623,25.067833,27.363045,26.746637,26.132042,25.517448,24.902855,24.28826,23.691795,23.097143,22.502491,21.90784,21.313189,19.045172,16.777155,14.50914,12.242936,9.97492,8.383139,6.789545,5.197764,3.6059825,2.0123885,1.6733645,1.3325275,0.9916905,0.6526665,0.31182957,0.28826106,0.26287958,0.2374981,0.21211663,0.18673515,0.15954071,0.13234627,0.10515183,0.07795739,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.35171473,0.70524246,1.0569572,1.4104849,1.7621996,1.4449311,1.1276628,0.8103943,0.49312583,0.17585737,0.13959812,0.10515183,0.07070554,0.034446288,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.26287958,0.48768693,0.7124943,0.93730164,1.162109,0.93730164,0.7124943,0.48768693,0.26287958,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.12509441,0.25018883,0.37528324,0.50037766,0.62547207,0.6091554,0.5946517,0.58014804,0.5656443,0.5493277,1.8691645,3.1908143,4.510651,5.8304877,7.1503243,6.9055743,6.6608243,6.414262,6.169512,5.924762,5.484212,5.045475,4.604925,4.164375,3.7256382,3.1799364,2.6342347,2.0903459,1.5446441,1.0007553,0.9445535,0.8901646,0.83577573,0.7795739,0.72518504,0.6653573,0.6055295,0.54570174,0.48587397,0.42423326,0.40972954,0.39522585,0.38072214,0.36440548,0.34990177,0.5656443,0.7795739,0.99531645,1.209246,1.4249886,1.1747998,0.9246109,0.6744221,0.42423326,0.17585737,0.2520018,0.32995918,0.40791658,0.48587397,0.5620184,0.66173136,0.76325727,0.8629702,0.96268314,1.062396,1.4467441,1.8329052,2.2172532,2.6016014,2.9877625,2.6269827,2.268016,1.9072367,1.54827,1.1874905,1.2491312,1.3125849,1.3742256,1.4376793,1.49932,1.845596,2.1900587,2.5345216,2.8807976,3.2252605,3.9468195,4.670192,5.391751,6.115123,6.836682,7.12313,7.407765,7.6924005,7.9770355,8.26167,8.056806,7.851941,7.647076,7.4422116,7.2373466,9.082943,10.926725,12.772322,14.617917,16.4617,20.522736,24.581959,28.642996,32.70222,36.763256,33.24067,29.718082,26.195496,22.67291,19.150324,16.220575,13.290829,10.359268,7.4295206,4.499773,4.6248674,4.749962,4.8750563,5.0001507,5.125245,5.91751,6.7097745,7.502039,8.294304,9.088382,8.675026,8.26167,7.850128,7.4367723,7.02523,6.430578,5.8341136,5.239462,4.64481,4.0501585,3.5606585,3.0693457,2.5798457,2.0903459,1.6008459,1.8383441,2.0758421,2.3133402,2.5508385,2.7883365,5.1071157,7.4277077,9.7483,12.067079,14.387671,13.675177,12.962683,12.250188,11.537694,10.825199,9.11195,7.400513,5.6872635,3.975827,2.2625773,1.8202144,1.3778516,0.9354887,0.49312583,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.054388877,0.059827764,0.065266654,0.07070554,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06707962,0.13415924,0.2030518,0.27013144,0.33721104,0.28463513,0.23205921,0.1794833,0.12690738,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.19217403,0.38434806,0.57833505,0.7705091,0.96268314,1.6842422,2.4076142,3.1291735,3.8525455,4.574105,5.331923,6.089741,6.8475595,7.605378,8.363196,6.695271,5.027345,3.3594196,1.693307,0.025381476,1.4304274,2.8354735,4.2405195,5.6455655,7.0506115,5.67276,4.2949085,2.9170568,1.5392052,0.16316663,1.3252757,2.4873846,3.6494937,4.8134155,5.975525,4.853301,3.729264,2.6070402,1.4848163,0.36259252,3.4754493,6.588306,9.699349,12.812206,15.925063,13.301706,10.680162,8.056806,5.4352617,2.811905,3.1744974,3.53709,3.8996825,4.262275,4.6248674,4.4870825,4.349297,4.213325,4.07554,3.9377546,5.292038,6.6481338,8.002417,9.3567,10.712796,8.914337,7.117691,5.319232,3.5225863,1.7241274,1.3796645,1.0352017,0.69073874,0.3444629,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.054388877,0.059827764,0.065266654,0.07070554,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.27013144,0.5402629,0.8103943,1.0805258,1.3506571,1.0805258,0.8103943,0.5402629,0.27013144,0.0,0.052575916,0.10515183,0.15772775,0.21030366,0.26287958,0.2374981,0.21211663,0.18673515,0.16316663,0.13778515,0.32270733,0.5076295,0.69255173,0.8774739,1.062396,1.1131591,1.162109,1.2128719,1.261822,1.3125849,1.2219368,1.1331016,1.0424535,0.95180535,0.8629702,1.6298534,2.3967366,3.1654327,3.9323158,4.699199,3.8090343,2.9206827,2.030518,1.1403534,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.29007402,0.5420758,0.79589057,1.0478923,1.2998942,1.3832904,1.4648738,1.54827,1.6298534,1.7132497,1.7404441,1.7676386,1.794833,1.8220274,1.8492218,1.504759,1.1602961,0.81583315,0.46955732,0.12509441,0.42967212,0.73424983,1.0406405,1.3452182,1.649796,1.6244144,1.6008459,1.5754645,1.550083,1.5247015,1.3252757,1.1258497,0.9246109,0.72518504,0.52575916,0.86478317,1.2056202,1.5446441,1.8854811,2.2245052,1.9507477,1.6751775,1.3996071,1.1258497,0.85027945,1.8256533,2.7992141,3.774588,4.749962,5.7253356,7.3352466,8.945157,10.555068,12.164979,13.77489,11.624716,9.474543,7.324369,5.1741953,3.0258346,3.2705846,3.5153344,3.7600844,4.004834,4.249584,5.767034,7.2844834,8.801933,10.319383,11.836833,11.095331,10.352016,9.610515,8.8672,8.125698,7.407765,6.6898317,5.9718986,5.2557783,4.537845,4.6756306,4.8116026,4.949388,5.087173,5.224958,5.7053933,6.185828,6.6644506,7.1448855,7.6253204,8.858135,10.089137,11.321951,12.554766,13.7875805,13.107719,12.427858,11.747997,11.068136,10.388275,9.334945,8.283426,7.230095,6.1767635,5.125245,4.5795436,4.0356545,3.489953,2.9442513,2.4003625,2.610666,2.819157,3.0294604,3.2397642,3.4500678,3.049403,2.6505513,2.2498865,1.8492218,1.4503701,1.3542831,1.260009,1.1657349,1.0696479,0.97537386,0.9826257,0.9898776,0.99712944,1.0043813,1.0116332,0.90829426,0.8031424,0.6979906,0.59283876,0.48768693,0.7850128,1.0823387,1.3796645,1.6769904,1.9743162,1.892733,1.8093367,1.7277533,1.6443571,1.5627737,2.0994108,2.6378605,3.1744974,3.7129474,4.249584,5.846804,7.4458375,9.043057,10.640278,12.237497,14.683184,17.127058,19.572744,22.016617,24.462305,26.202747,27.943192,29.681824,31.422268,33.162712,34.712795,36.26288,37.81296,39.363045,40.913128,40.12993,39.346725,38.565342,37.78214,37.00075,35.302006,33.605076,31.908142,30.209396,28.512463,27.181747,25.852846,24.522131,23.19323,21.862516,21.54706,21.233418,20.917963,20.602507,20.287052,20.613384,20.937904,21.262424,21.586945,21.913279,20.60432,19.297174,17.990028,16.682882,15.375735,15.497204,15.620485,15.741954,15.865235,15.986704,17.654629,19.322556,20.99048,22.656593,24.324518,23.740746,23.155159,22.56957,21.985798,21.40021,21.782745,22.165281,22.547815,22.930351,23.312885,21.030367,18.747847,16.465326,14.182806,11.900287,9.791811,7.6851482,5.576673,3.4700103,1.3633479,1.1530442,0.94274056,0.7324369,0.52213323,0.31182957,0.2755703,0.2374981,0.19942589,0.16316663,0.12509441,0.11421664,0.10515183,0.09427405,0.08520924,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.18310922,0.36440548,0.5475147,0.7306239,0.9119202,0.75963134,0.6073425,0.4550536,0.30276474,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.34990177,0.6508536,0.9499924,1.2491312,1.550083,1.2491312,0.9499924,0.6508536,0.34990177,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.16316663,0.3245203,0.48768693,0.6508536,0.8122072,0.79226464,0.77232206,0.7523795,0.7324369,0.7124943,1.3343405,1.9579996,2.5798457,3.2016919,3.825351,4.1897564,4.554162,4.9203806,5.2847857,5.6491914,5.292038,4.934884,4.5777307,4.220577,3.8616104,3.303218,2.7430124,2.182807,1.6226015,1.062396,0.99712944,0.9318628,0.8665961,0.8031424,0.73787576,0.65810543,0.57833505,0.49675176,0.4169814,0.33721104,0.34264994,0.3480888,0.35171473,0.35715362,0.36259252,0.67079616,0.97718686,1.2853905,1.5917811,1.8999848,1.5627737,1.2255627,0.8883517,0.5493277,0.21211663,0.30820364,0.40247768,0.49675176,0.59283876,0.6871128,0.774135,0.8629702,0.9499924,1.0370146,1.1258497,1.6044719,2.084907,2.565342,3.045777,3.5243993,2.9823234,2.4402475,1.8981718,1.3542831,0.8122072,0.8629702,0.9119202,0.96268314,1.0116332,1.062396,1.5228885,1.983381,2.4420607,2.902553,3.3630457,4.3928084,5.422571,6.452334,7.4820967,8.511859,8.729415,8.94697,9.164526,9.382081,9.599637,9.273304,8.945157,8.617011,8.290678,7.9625316,9.023115,10.081885,11.142468,12.203052,13.261822,15.379361,17.496902,19.614443,21.731983,23.849524,21.57063,19.289923,17.009214,14.730321,12.449615,10.97205,9.494485,8.01692,6.539356,5.0617914,5.3119802,5.562169,5.812358,6.0625467,6.3127356,7.2391596,8.167397,9.0956335,10.022058,10.950294,10.25049,9.550687,8.8508835,8.149267,7.4494634,6.776854,6.104245,5.431636,4.76084,4.0882306,3.6295512,3.1726844,2.715818,2.2571385,1.8002719,1.9507477,2.0994108,2.2498865,2.4003625,2.5508385,5.660069,8.7693,11.880343,14.989574,18.100618,17.32467,16.550535,15.774588,15.000452,14.224504,11.974618,9.724731,7.474845,5.224958,2.9750717,2.3858588,1.794833,1.2056202,0.61459434,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.027194439,0.030820364,0.032633327,0.034446288,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.09064813,0.1794833,0.27013144,0.36077955,0.44961473,0.38072214,0.3100166,0.23931105,0.17041849,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.16497959,0.32995918,0.4949388,0.65991837,0.824898,1.5682126,2.3097143,3.053029,3.7945306,4.537845,5.7217097,6.9073873,8.093065,9.27693,10.462607,8.372261,6.281915,4.1915693,2.1030366,0.012690738,0.71430725,1.4177368,2.1193533,2.8227828,3.5243993,2.8427253,2.1592383,1.4775645,0.79407763,0.11240368,0.9119202,1.7132497,2.5127661,3.3122826,4.1117992,3.3829882,2.6523643,1.9217403,1.1929294,0.46230546,3.876114,7.28811,10.700105,14.112101,17.52591,14.744824,11.965553,9.184468,6.4051967,3.6241121,4.0374675,4.4508233,4.8623657,5.275721,5.6872635,4.9620786,4.2368937,3.5117085,2.7883365,2.0631514,3.8017826,5.542227,7.2826705,9.023115,10.761745,8.781991,6.8022356,4.8224807,2.8427253,0.8629702,0.69073874,0.5166943,0.3444629,0.17223145,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.027194439,0.030820364,0.032633327,0.034446288,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.13415924,0.27013144,0.40429065,0.5402629,0.6744221,0.5402629,0.40429065,0.27013144,0.13415924,0.0,0.045324065,0.09064813,0.13415924,0.1794833,0.22480737,0.21211663,0.19942589,0.18673515,0.17585737,0.16316663,0.27919623,0.39703882,0.5148814,0.6327239,0.7505665,0.9499924,1.1494182,1.3506571,1.550083,1.7495089,1.6298534,1.5101979,1.3905423,1.2708868,1.1494182,2.128418,3.105605,4.082792,5.0599785,6.037165,4.855114,3.673062,2.4891977,1.3071461,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.36984438,0.69073874,1.0098201,1.3307146,1.649796,1.7223145,1.794833,1.8673514,1.93987,2.0123885,2.0577126,2.1030366,2.1483607,2.1918716,2.2371957,1.8020848,1.3669738,0.9318628,0.49675176,0.06164073,0.32814622,0.59283876,0.8575313,1.1222239,1.3869164,1.261822,1.1367276,1.0116332,0.8883517,0.76325727,0.66173136,0.5620184,0.46230546,0.36259252,0.26287958,0.43329805,0.60190356,0.77232206,0.94274056,1.1131591,0.97537386,0.8375887,0.69980353,0.5620184,0.42423326,0.9119202,1.3996071,1.887294,2.374981,2.8626678,5.243088,7.6216946,10.002114,12.382534,14.762955,12.262879,9.762803,7.262728,4.762653,2.2625773,2.8354735,3.4083695,3.9794528,4.552349,5.125245,7.25185,9.380268,11.506873,13.635292,15.761897,14.447499,13.1331005,11.81689,10.502492,9.188094,8.285239,7.382384,6.4795284,5.576673,4.6756306,4.8877473,5.0998635,5.3119802,5.52591,5.7380266,6.3272395,6.9182653,7.507478,8.096691,8.6877165,10.085511,11.483305,12.879286,14.277081,15.674874,14.960567,14.244447,13.53014,12.815832,12.099712,10.854207,9.610515,8.365009,7.119504,5.8758116,5.0781083,4.2804046,3.482701,2.6849976,1.887294,2.38042,2.8717327,3.3648586,3.8579843,4.349297,3.7129474,3.0747845,2.4366217,1.8002719,1.162109,1.0768998,0.9916905,0.90829426,0.823085,0.73787576,0.8103943,0.88291276,0.9554313,1.0279498,1.1004683,0.9354887,0.7705091,0.6055295,0.4405499,0.2755703,0.4169814,0.56020546,0.7016165,0.8448406,0.9880646,0.95180535,0.91735905,0.88291276,0.8466535,0.8122072,1.3379664,1.8619126,2.3876717,2.911618,3.437377,4.4798307,5.522284,6.5647373,7.607191,8.649645,11.321951,13.994258,16.668379,19.340685,22.01299,23.557636,25.10228,26.646925,28.191568,29.738026,30.77504,31.812054,32.849068,33.887897,34.92491,35.401722,35.88034,36.35715,36.835773,37.312584,36.08158,34.852394,33.623203,32.392204,31.163013,29.272095,27.382986,25.492067,23.60296,21.71204,21.20441,20.696781,20.189152,19.683334,19.175705,18.862062,18.550234,18.236591,17.92476,17.612932,16.927631,16.242332,15.557032,14.871732,14.188245,14.567154,14.947877,15.326786,15.707508,16.08823,17.127058,18.167698,19.208338,20.247166,21.287807,20.73304,20.178274,19.621695,19.066927,18.512161,19.871883,21.233418,22.59314,23.952862,25.312584,23.01556,20.716722,18.4197,16.122677,13.825653,11.202296,8.5789385,5.957395,3.3358512,0.7124943,0.6327239,0.5529536,0.47318324,0.39159992,0.31182957,0.26287958,0.21211663,0.16316663,0.11240368,0.06164073,0.07070554,0.07795739,0.08520924,0.092461094,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.43692398,0.8122072,1.1874905,1.5627737,1.938057,1.5627737,1.1874905,0.8122072,0.43692398,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.19942589,0.40066472,0.6000906,0.7995165,1.0007553,0.97537386,0.9499924,0.9246109,0.89922947,0.87566096,0.7995165,0.72518504,0.6508536,0.5747091,0.50037766,1.4757515,2.4493124,3.4246864,4.40006,5.375434,5.0998635,4.8242936,4.550536,4.274966,3.9993954,3.4246864,2.8499773,2.275268,1.7005589,1.1258497,1.0497054,0.97537386,0.89922947,0.824898,0.7505665,0.6508536,0.5493277,0.44961473,0.34990177,0.25018883,0.2755703,0.2991388,0.3245203,0.34990177,0.37528324,0.774135,1.1747998,1.5754645,1.9743162,2.374981,1.9507477,1.5247015,1.1004683,0.6744221,0.25018883,0.36259252,0.4749962,0.5873999,0.69980353,0.8122072,0.8883517,0.96268314,1.0370146,1.1131591,1.1874905,1.7621996,2.3369088,2.911618,3.48814,4.062849,3.3376641,2.612479,1.887294,1.162109,0.43692398,0.4749962,0.51306844,0.5493277,0.5873999,0.62547207,1.2001812,1.7748904,2.3495996,2.9243085,3.5008307,4.836984,6.1749506,7.512917,8.8508835,10.1870365,10.337513,10.487988,10.636651,10.7871275,10.937603,10.487988,10.038374,9.5869465,9.137331,8.6877165,8.963287,9.237044,9.512614,9.788185,10.061942,10.2378,10.411844,10.587702,10.761745,10.937603,9.900589,8.861761,7.8247466,6.787732,5.750717,5.7253356,5.6999545,5.674573,5.6491914,5.6256227,5.999093,6.3743763,6.7496595,7.124943,7.500226,8.562622,9.625018,10.687414,11.74981,12.812206,11.8241415,10.837891,9.849826,8.861761,7.8755093,7.124943,6.3743763,5.6256227,4.8750563,4.12449,3.7002566,3.2742105,2.8499773,2.4257438,1.9996977,2.0631514,2.124792,2.1882458,2.2498865,2.3133402,6.2130227,10.112705,14.012388,17.912071,21.811752,20.974165,20.138388,19.3008,18.463211,17.625622,14.837286,12.050762,9.262425,6.474089,3.6875658,2.94969,2.2118144,1.4757515,0.73787576,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.11240368,0.22480737,0.33721104,0.44961473,0.5620184,0.4749962,0.387974,0.2991388,0.21211663,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13778515,0.2755703,0.41335547,0.5493277,0.6871128,1.4503701,2.2118144,2.9750717,3.738329,4.499773,6.11331,7.7250338,9.336758,10.950294,12.562017,10.049252,7.5382986,5.0255322,2.5127661,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.50037766,0.93730164,1.3742256,1.8129625,2.2498865,1.9126755,1.5754645,1.2382535,0.89922947,0.5620184,4.274966,7.987913,11.700861,15.411995,19.124943,16.187943,13.250943,10.312131,7.3751316,4.4381323,4.900438,5.3627434,5.825049,6.2873545,6.7496595,5.4370747,4.12449,2.811905,1.49932,0.18673515,2.3133402,4.4381323,6.5629244,8.6877165,10.812509,8.649645,6.48678,4.325729,2.1628644,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.18673515,0.18673515,0.18673515,0.18673515,0.18673515,0.2374981,0.28826106,0.33721104,0.387974,0.43692398,0.7868258,1.1367276,1.4866294,1.8383441,2.1882458,2.03777,1.887294,1.7368182,1.5881553,1.4376793,2.6251698,3.8126602,5.0001507,6.187641,7.3751316,5.89938,4.4254417,2.94969,1.4757515,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.44961473,0.8375887,1.2255627,1.6117238,1.9996977,2.0631514,2.124792,2.1882458,2.2498865,2.3133402,2.374981,2.4366217,2.5000753,2.561716,2.6251698,2.0994108,1.5754645,1.0497054,0.52575916,0.0,0.22480737,0.44961473,0.6744221,0.89922947,1.1258497,0.89922947,0.6744221,0.44961473,0.22480737,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,3.150929,6.300045,9.4509735,12.60009,15.749206,12.899229,10.049252,7.1992745,4.349297,1.49932,2.4003625,3.299592,4.2006345,5.0998635,6.000906,8.73848,11.47424,14.211814,16.949387,19.68696,17.799667,15.912373,14.025079,12.137785,10.25049,9.162713,8.074935,6.987158,5.89938,4.8116026,5.0998635,5.388125,5.674573,5.962834,6.249282,6.9508986,7.650702,8.350506,9.050309,9.750113,11.312886,12.87566,14.438434,15.999394,17.562168,16.811602,16.062849,15.312282,14.561715,13.812962,12.375282,10.937603,9.499924,8.062244,6.624565,5.57486,4.5251546,3.4754493,2.4257438,1.3742256,2.1501737,2.9243085,3.7002566,4.4743915,5.2503395,4.3746786,3.5008307,2.6251698,1.7495089,0.87566096,0.7995165,0.72518504,0.6508536,0.5747091,0.50037766,0.63816285,0.774135,0.9119202,1.0497054,1.1874905,0.96268314,0.73787576,0.51306844,0.28826106,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.5747091,1.0877775,1.6008459,2.1121013,2.6251698,3.1128569,3.6005437,4.0882306,4.574105,5.0617914,7.9625316,10.863272,13.762199,16.66294,19.561867,20.912523,22.26318,23.612024,24.962683,26.31334,26.837286,27.363045,27.88699,28.41275,28.936695,30.675327,32.412144,34.150776,35.887596,37.624413,36.86297,36.099712,35.33827,34.57501,33.811752,31.36244,28.913128,26.462002,24.01269,21.563377,20.861761,20.161957,19.462152,18.76235,18.062546,17.112555,16.162561,15.212569,14.262577,13.312584,13.24913,13.1874895,13.125849,13.062395,13.000754,13.637105,14.275268,14.911617,15.54978,16.187943,16.599485,17.01284,17.424383,17.837738,18.24928,17.725336,17.199575,16.67563,16.14987,15.624111,17.962833,20.299742,22.638464,24.975372,27.31228,25.000753,22.687414,20.374073,18.062546,15.749206,12.612781,9.474543,6.338117,3.199879,0.06164073,0.11240368,0.16316663,0.21211663,0.26287958,0.31182957,0.25018883,0.18673515,0.12509441,0.06164073,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.059827764,0.07070554,0.07977036,0.09064813,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.35171473,0.6544795,0.9572442,1.260009,1.5627737,1.2926424,1.0225109,0.7523795,0.48224804,0.21211663,0.17041849,0.12690738,0.08520924,0.04169814,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.19036107,0.34264994,0.4949388,0.64722764,0.7995165,0.8575313,0.9155461,0.97174793,1.0297627,1.0877775,0.9880646,0.8883517,0.7868258,0.6871128,0.5873999,1.3542831,2.1229792,2.8898623,3.6567454,4.4254417,4.274966,4.12449,3.975827,3.825351,3.6748753,3.4301252,3.1853752,2.9406252,2.6958754,2.4493124,2.0975976,1.745883,1.3923552,1.0406405,0.6871128,0.58921283,0.49312583,0.39522585,0.29732585,0.19942589,0.21936847,0.23931105,0.25925365,0.27919623,0.2991388,0.62728506,0.9554313,1.2817645,1.6099107,1.938057,1.6008459,1.261822,0.9246109,0.5873999,0.25018883,0.36077955,0.46955732,0.58014804,0.69073874,0.7995165,0.83033687,0.85934424,0.8901646,0.91917205,0.9499924,1.4104849,1.8691645,2.3296568,2.7901495,3.2506418,2.6704938,2.0903459,1.5101979,0.9300498,0.34990177,0.45324063,0.55476654,0.65810543,0.75963134,0.8629702,1.4431182,2.0232663,2.6034143,3.1817493,3.7618973,4.7390842,5.718084,6.695271,7.6724577,8.649645,8.999546,9.349448,9.699349,10.049252,10.399154,10.038374,9.675781,9.313189,8.950596,8.588004,8.680465,8.772926,8.865387,8.957849,9.050309,9.267865,9.48542,9.702975,9.920531,10.138086,9.360326,8.582565,7.804804,7.027043,6.249282,6.1405044,6.0299134,5.919323,5.810545,5.6999545,5.9447045,6.189454,6.434204,6.680767,6.925517,8.417585,9.909654,11.401722,12.895603,14.387671,13.062395,11.73712,10.411844,9.088382,7.763106,7.0506115,6.338117,5.6256227,4.9131284,4.2006345,3.6875658,3.1744974,2.663242,2.1501737,1.6371052,1.693307,1.7476959,1.8020848,1.8582866,1.9126755,5.2575917,8.602508,11.947423,15.292339,18.637255,18.33993,18.042604,17.745277,17.447952,17.150625,14.382232,11.615651,8.847258,6.0806766,3.3122826,2.6541772,1.9978848,1.3397794,0.68167394,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.09064813,0.1794833,0.27013144,0.36077955,0.44961473,0.3825351,0.3154555,0.24837588,0.1794833,0.11240368,0.09427405,0.07795739,0.059827764,0.04169814,0.025381476,0.02175555,0.01994259,0.018129626,0.014503701,0.012690738,0.014503701,0.018129626,0.01994259,0.02175555,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.034446288,0.045324065,0.054388877,0.065266654,0.07433146,0.17041849,0.26469254,0.36077955,0.4550536,0.5493277,1.1602961,1.7694515,2.38042,2.9895754,3.6005437,4.893186,6.185828,7.476658,8.7693,10.061942,8.2779875,6.492219,4.708264,2.9224956,1.1367276,1.1403534,1.1421664,1.1457924,1.1476053,1.1494182,1.1403534,1.1294757,1.1204109,1.1095331,1.1004683,1.2400664,1.3796645,1.5192627,1.6606737,1.8002719,1.5301404,1.260009,0.9898776,0.7197462,0.44961473,3.4246864,6.399758,9.374829,12.349901,15.324973,13.172986,11.019187,8.8672,6.7152133,4.5632267,4.7300196,4.896812,5.0654173,5.23221,5.4008155,4.349297,3.299592,2.2498865,1.2001812,0.15047589,1.8492218,3.5497808,5.2503395,6.9490857,8.649645,6.9200783,5.1905117,3.4591327,1.7295663,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.15772775,0.16497959,0.17223145,0.1794833,0.18673515,0.40972954,0.6327239,0.8557183,1.0768998,1.2998942,1.5319533,1.7658255,1.9978848,2.229944,2.4620032,2.2045624,1.9471219,1.6896812,1.4322405,1.1747998,2.1193533,3.0657198,4.0102735,4.954827,5.89938,4.7191415,3.540716,2.3604772,1.1802386,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.36077955,0.67079616,0.9808127,1.2908293,1.6008459,1.649796,1.7005589,1.7495089,1.8002719,1.8492218,1.9072367,1.9652514,2.0232663,2.079468,2.137483,1.7223145,1.3071461,0.8919776,0.47680917,0.06164073,0.23024625,0.39703882,0.5656443,0.7324369,0.89922947,0.7197462,0.5402629,0.36077955,0.1794833,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.521831,5.045475,7.567306,10.089137,12.612781,10.825199,9.037619,7.250037,5.462456,3.6748753,3.8996825,4.12449,4.349297,4.574105,4.800725,7.6325727,10.46442,13.29808,16.129929,18.961775,17.034595,15.107417,13.180238,11.253058,9.325879,8.326937,7.3298078,6.3326783,5.335549,4.3366065,4.6756306,5.0128417,5.3500524,5.6872635,6.0244746,6.677141,7.3298078,7.9824743,8.63514,9.287807,11.182353,13.0769,14.973258,16.867804,18.76235,17.76522,16.768091,15.769149,14.772019,13.77489,12.469557,11.164224,9.860703,8.55537,7.250037,6.742408,6.2347784,5.727149,5.219519,4.7118897,4.748149,4.782595,4.8170414,4.853301,4.8877473,4.64481,4.401873,4.160749,3.917812,3.6748753,3.0403383,2.4058013,1.7694515,1.1349145,0.50037766,0.7433147,0.98443866,1.2273756,1.4703126,1.7132497,1.3941683,1.0768998,0.75963134,0.44236287,0.12509441,0.10333887,0.07977036,0.058014803,0.034446288,0.012690738,0.01994259,0.027194439,0.034446288,0.04169814,0.05076295,0.72337204,1.3941683,2.0667772,2.7393866,3.4119956,3.6132345,3.8126602,4.0120864,4.213325,4.4127507,6.6608243,8.907085,11.155159,13.40142,15.649493,16.769903,17.890314,19.010725,20.129324,21.249735,22.15259,23.055445,23.9583,24.859343,25.762197,27.471823,29.183258,30.892883,32.602505,34.31213,34.437225,34.562317,34.687412,34.812508,34.937603,33.32769,31.717781,30.10787,28.49796,26.888048,25.925365,24.962683,23.999998,23.037315,22.074633,20.89258,19.71053,18.526665,17.344612,16.162561,15.825351,15.488139,15.1509285,14.811904,14.474693,14.871732,15.270584,15.667623,16.064661,16.4617,16.914942,17.368181,17.819609,18.27285,18.724277,17.620184,16.514277,15.410182,14.304275,13.200181,15.404743,17.609306,19.815681,22.020243,24.224806,23.18054,22.13446,21.090193,20.045927,18.999847,15.241576,11.485118,7.7268467,3.9703882,0.21211663,0.3825351,0.5529536,0.72337204,0.8919776,1.062396,0.8557183,0.64722764,0.4405499,0.23205921,0.025381476,0.06164073,0.099712946,0.13778515,0.17585737,0.21211663,0.19942589,0.18673515,0.17585737,0.16316663,0.15047589,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.045324065,0.052575916,0.059827764,0.06707962,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.26831847,0.49675176,0.726998,0.9572442,1.1874905,1.0225109,0.8575313,0.69255173,0.5275721,0.36259252,0.29007402,0.21755551,0.14503701,0.072518505,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.1794833,0.28463513,0.38978696,0.4949388,0.6000906,0.73968875,0.8792868,1.020698,1.1602961,1.2998942,1.1747998,1.0497054,0.9246109,0.7995165,0.6744221,1.2346275,1.794833,2.3550384,2.9152439,3.4754493,3.4500678,3.4246864,3.3993049,3.3757362,3.350355,3.435564,3.5207734,3.6041696,3.6893787,3.774588,3.1454902,2.514579,1.8854811,1.2545701,0.62547207,0.5293851,0.43511102,0.34083697,0.24474995,0.15047589,0.16497959,0.1794833,0.19579996,0.21030366,0.22480737,0.48043507,0.73424983,0.9898776,1.2455053,1.49932,1.2491312,1.0007553,0.7505665,0.50037766,0.25018883,0.35715362,0.46411842,0.5728962,0.67986095,0.7868258,0.77232206,0.75781834,0.7433147,0.726998,0.7124943,1.0569572,1.403233,1.7476959,2.0921588,2.4366217,2.0033236,1.5682126,1.1331016,0.6979906,0.26287958,0.42967212,0.5982776,0.7650702,0.9318628,1.1004683,1.6842422,2.269829,2.855416,3.43919,4.024777,4.6429973,5.2594047,5.8776245,6.495845,7.112252,7.66158,8.212721,8.762048,9.313189,9.862516,9.5869465,9.313189,9.037619,8.762048,8.488291,8.397643,8.306994,8.21816,8.127511,8.036863,8.29793,8.557183,8.81825,9.077503,9.336758,8.820063,8.303369,7.7848616,7.268167,6.7496595,6.5556726,6.359873,6.165886,5.9700856,5.774286,5.8903155,6.004532,6.1205616,6.2347784,6.350808,8.272549,10.194288,12.117842,14.039582,15.963136,14.300649,12.638163,10.975676,9.313189,7.650702,6.9744673,6.300045,5.6256227,4.949388,4.274966,3.6748753,3.0747845,2.474694,1.8746033,1.2745126,1.3216497,1.3705997,1.4177368,1.4648738,1.5120108,4.3021603,7.0923095,9.882459,12.672608,15.462758,15.705695,15.946819,16.189756,16.432693,16.67563,13.927178,11.18054,8.432089,5.6854506,2.9369993,2.3604772,1.7821422,1.2056202,0.62728506,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06707962,0.13415924,0.2030518,0.27013144,0.33721104,0.29007402,0.24293698,0.19579996,0.14684997,0.099712946,0.09064813,0.07977036,0.07070554,0.059827764,0.05076295,0.045324065,0.03988518,0.034446288,0.030820364,0.025381476,0.030820364,0.034446288,0.03988518,0.045324065,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.07070554,0.09064813,0.11059072,0.13053331,0.15047589,0.2030518,0.25562772,0.30820364,0.36077955,0.41335547,0.87022203,1.3270886,1.7857682,2.2426348,2.6995013,3.673062,4.64481,5.618371,6.590119,7.5618668,6.5049095,5.4479527,4.3891826,3.3322253,2.275268,2.280707,2.2843328,2.2897718,2.2952106,2.3006494,2.268016,2.2353828,2.2027495,2.1701162,2.137483,1.9797552,1.8220274,1.6642996,1.5083848,1.3506571,1.1476053,0.9445535,0.7433147,0.5402629,0.33721104,2.5744069,4.8116026,7.0506115,9.287807,11.525003,10.15803,8.789243,7.422269,6.055295,4.688321,4.559601,4.4326935,4.305786,4.177066,4.0501585,3.2633326,2.474694,1.6878681,0.89922947,0.11240368,1.3869164,2.663242,3.9377546,5.2122674,6.48678,5.1905117,3.8924308,2.5943494,1.2980812,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.12690738,0.14322405,0.15772775,0.17223145,0.18673515,0.581961,0.97718686,1.3724127,1.7676386,2.1628644,2.277081,2.3931105,2.5073273,2.6233568,2.7375734,2.373168,2.0069497,1.6425442,1.2781386,0.9119202,1.6153497,2.3169663,3.0203958,3.7220123,4.4254417,3.540716,2.6541772,1.7694515,0.88472575,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.27013144,0.50219065,0.73424983,0.968122,1.2001812,1.2382535,1.2745126,1.3125849,1.3506571,1.3869164,1.4394923,1.4920682,1.5446441,1.5972201,1.649796,1.3452182,1.0406405,0.73424983,0.42967212,0.12509441,0.23568514,0.3444629,0.4550536,0.5656443,0.6744221,0.5402629,0.40429065,0.27013144,0.13415924,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.8945459,3.7890918,5.6854506,7.5799966,9.474543,8.749357,8.024173,7.3008003,6.5756154,5.8504305,5.4008155,4.949388,4.499773,4.0501585,3.6005437,6.528478,9.4546,12.382534,15.310469,18.236591,16.269526,14.302462,12.335398,10.368333,8.399456,7.4929743,6.58468,5.678199,4.7699046,3.8616104,4.249584,4.6375585,5.0255322,5.411693,5.7996674,6.4051967,7.0107265,7.614443,8.219973,8.825501,11.05182,13.279951,15.508082,17.7344,19.96253,18.717026,17.473333,16.227829,14.982323,13.736817,12.565643,11.392657,10.21967,9.046683,7.8755093,7.909956,7.944402,7.9806614,8.015107,8.049554,7.344311,6.640882,5.9356394,5.230397,4.5251546,4.914942,5.3047285,5.6945157,6.0843024,6.4759026,5.279347,4.0846047,2.8898623,1.69512,0.50037766,0.8466535,1.1947423,1.5428312,1.889107,2.2371957,1.8274662,1.4177368,1.0080072,0.5982776,0.18673515,0.15410182,0.12328146,0.09064813,0.058014803,0.025381476,0.027194439,0.030820364,0.032633327,0.034446288,0.038072214,0.87022203,1.7023718,2.5345216,3.3666716,4.2006345,4.1117992,4.024777,3.9377546,3.8507326,3.7618973,5.3573046,6.9527116,8.548119,10.141713,11.73712,12.627284,13.517449,14.407614,15.297778,16.187943,17.467894,18.747847,20.027798,21.307749,22.5877,24.27013,25.952559,27.634989,29.317417,30.999847,32.013294,33.024925,34.038372,35.050007,36.061638,35.292942,34.522434,33.751923,32.983227,32.21272,30.987156,29.763407,28.537844,27.31228,26.08672,24.672607,23.256683,21.842573,20.428463,19.012539,18.399757,17.786976,17.174194,16.563227,15.950445,16.108173,16.2659,16.421816,16.579542,16.73727,17.230396,17.721708,18.214834,18.70796,19.199274,17.515032,15.828977,14.144734,12.460492,10.774437,12.848466,14.920682,16.992899,19.065115,21.137331,21.360325,21.583319,21.8045,22.027494,22.25049,17.872185,13.49388,9.117389,4.740897,0.36259252,0.6526665,0.94274056,1.2328146,1.5228885,1.8129625,1.4594349,1.1077201,0.7541924,0.40247768,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,0.2991388,0.2991388,0.2991388,0.2991388,0.2991388,0.2991388,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.030820364,0.034446288,0.03988518,0.045324065,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.18310922,0.34083697,0.49675176,0.6544795,0.8122072,0.7523795,0.69255173,0.6327239,0.5728962,0.51306844,0.40972954,0.30820364,0.20486477,0.10333887,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.17041849,0.22662032,0.28463513,0.34264994,0.40066472,0.62184614,0.8448406,1.067835,1.2908293,1.5120108,1.3633479,1.2128719,1.062396,0.9119202,0.76325727,1.114972,1.4666867,1.8202144,2.1719291,2.525457,2.6251698,2.7248828,2.8245957,2.9243085,3.0258346,3.43919,3.8543584,4.269527,4.6846952,5.0998635,4.1933823,3.2850883,2.3767939,1.4703126,0.5620184,0.46955732,0.3770962,0.28463513,0.19217403,0.099712946,0.11059072,0.11965553,0.13053331,0.13959812,0.15047589,0.33177215,0.5148814,0.6979906,0.8792868,1.062396,0.89922947,0.73787576,0.5747091,0.41335547,0.25018883,0.35534066,0.4604925,0.5656443,0.67079616,0.774135,0.71430725,0.6544795,0.5946517,0.53482395,0.4749962,0.70524246,0.9354887,1.1657349,1.3941683,1.6244144,1.3343405,1.0442665,0.7541924,0.46411842,0.17585737,0.40791658,0.6399758,0.872035,1.1059072,1.3379664,1.9271792,2.518205,3.1074178,3.6966307,4.2876563,4.5450974,4.802538,5.0599785,5.317419,5.57486,6.3254266,7.07418,7.8247466,8.575313,9.325879,9.137331,8.950596,8.762048,8.575313,8.386765,8.1148205,7.842876,7.569119,7.2971745,7.02523,7.327995,7.6307597,7.931711,8.234476,8.537241,8.2798,8.02236,7.764919,7.507478,7.250037,6.970841,6.6898317,6.4106355,6.1296263,5.8504305,5.8341136,5.81961,5.805106,5.7906027,5.774286,8.127511,10.480737,12.8321495,15.185374,17.536787,15.537089,13.537392,11.537694,9.537996,7.5382986,6.9001355,6.261973,5.6256227,4.98746,4.349297,3.6621845,2.9750717,2.2879589,1.6008459,0.9119202,0.95180535,0.9916905,1.0333886,1.0732739,1.1131591,3.346729,5.582112,7.817495,10.052877,12.28826,13.069647,13.852847,14.634234,15.417434,16.200634,13.472125,10.745429,8.01692,5.290225,2.561716,2.0649643,1.5682126,1.0696479,0.5728962,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.045324065,0.09064813,0.13415924,0.1794833,0.22480737,0.19761293,0.17041849,0.14322405,0.11421664,0.0870222,0.08520924,0.08339628,0.07977036,0.07795739,0.07433146,0.06707962,0.059827764,0.052575916,0.045324065,0.038072214,0.045324065,0.052575916,0.059827764,0.06707962,0.07433146,0.07433146,0.07433146,0.07433146,0.07433146,0.07433146,0.10515183,0.13415924,0.16497959,0.19579996,0.22480737,0.23568514,0.24474995,0.25562772,0.26469254,0.2755703,0.58014804,0.88472575,1.1893034,1.4956942,1.8002719,2.4529383,3.105605,3.7582715,4.409125,5.0617914,4.7318325,4.401873,4.071914,3.7419548,3.4119956,3.4192474,3.4283123,3.435564,3.442816,3.4500678,3.395679,3.339477,3.2850883,3.2306993,3.1744974,2.7194438,2.2643902,1.8093367,1.3542831,0.89922947,0.7650702,0.630911,0.4949388,0.36077955,0.22480737,1.7259403,3.2252605,4.7245803,6.2257137,7.7250338,7.1430726,6.5592985,5.977338,5.3953767,4.8116026,4.3891826,3.966762,3.5443418,3.1219215,2.6995013,2.175555,1.649796,1.1258497,0.6000906,0.07433146,0.9246109,1.7748904,2.6251698,3.4754493,4.325729,3.4591327,2.5943494,1.7295663,0.86478317,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.09789998,0.11965553,0.14322405,0.16497959,0.18673515,0.7541924,1.3216497,1.889107,2.4583774,3.0258346,3.0222087,3.0203958,3.0167696,3.0149567,3.0131438,2.5399606,2.0667772,1.5954071,1.1222239,0.6508536,1.1095331,1.5700256,2.030518,2.4891977,2.94969,2.3604772,1.7694515,1.1802386,0.58921283,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.1794833,0.33539808,0.4894999,0.64541465,0.7995165,0.824898,0.85027945,0.87566096,0.89922947,0.9246109,0.97174793,1.020698,1.067835,1.114972,1.162109,0.968122,0.77232206,0.57833505,0.3825351,0.18673515,0.23931105,0.291887,0.3444629,0.39703882,0.44961473,0.36077955,0.27013144,0.1794833,0.09064813,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.2672608,2.5345216,3.8017826,5.0708566,6.338117,6.6753283,7.0125394,7.3497505,7.686961,8.024173,6.9001355,5.774286,4.650249,3.5243993,2.4003625,5.422571,8.444779,11.466989,14.489197,17.513218,15.504456,13.497506,11.490557,9.481794,7.474845,6.6571984,5.8395524,5.0219064,4.2042603,3.386614,3.825351,4.262275,4.699199,5.137936,5.57486,6.1332526,6.6898317,7.2482243,7.804804,8.363196,10.9230995,13.483003,16.042906,18.60281,21.162712,19.670645,18.176764,16.684694,15.192626,13.700559,12.659918,11.619277,10.58045,9.539809,8.499168,9.077503,9.655839,10.232361,10.810696,11.3872175,9.9422865,8.497355,7.0524244,5.6074934,4.162562,5.185073,6.207584,7.230095,8.252605,9.275117,7.520169,5.765221,4.0102735,2.2553256,0.50037766,0.95180535,1.405046,1.8582866,2.3097143,2.762955,2.2607644,1.7567607,1.2545701,0.7523795,0.25018883,0.20667773,0.16497959,0.12328146,0.07977036,0.038072214,0.034446288,0.032633327,0.030820364,0.027194439,0.025381476,1.017072,2.0105755,3.002266,3.9957695,4.98746,4.612177,4.2368937,3.8616104,3.48814,3.1128569,4.0555973,4.9983377,5.9392653,6.882006,7.8247466,8.484665,9.144584,9.804502,10.46442,11.124338,12.783199,14.440247,16.097294,17.754343,19.413204,21.068438,22.72186,24.377094,26.03233,27.687565,29.58755,31.487534,33.38752,35.287502,37.18749,37.258194,37.327087,37.397793,37.466686,37.53739,36.050762,34.562317,33.07569,31.587248,30.100618,28.452635,26.804651,25.15667,23.510498,21.862516,20.974165,20.087626,19.199274,18.312735,17.424383,17.3428,17.259403,17.17782,17.094423,17.01284,17.545853,18.07705,18.610062,19.143072,19.67427,17.40988,15.14549,12.879286,10.614896,8.350506,10.290376,12.230246,14.170115,16.109985,18.049856,19.540112,21.030367,22.52062,24.009064,25.49932,20.502794,15.504456,10.507931,5.5095935,0.51306844,0.922798,1.3325275,1.742257,2.1519866,2.561716,2.0649643,1.5682126,1.0696479,0.5728962,0.07433146,0.13778515,0.19942589,0.26287958,0.3245203,0.387974,0.40066472,0.41335547,0.42423326,0.43692398,0.44961473,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.014503701,0.018129626,0.01994259,0.02175555,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.09789998,0.18310922,0.26831847,0.35171473,0.43692398,0.48224804,0.5275721,0.5728962,0.61822027,0.66173136,0.5293851,0.39703882,0.26469254,0.13234627,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.15954071,0.17041849,0.1794833,0.19036107,0.19942589,0.5058166,0.8103943,1.114972,1.4195497,1.7241274,1.550083,1.3742256,1.2001812,1.0243238,0.85027945,0.99531645,1.1403534,1.2853905,1.4304274,1.5754645,1.8002719,2.0250793,2.2498865,2.474694,2.6995013,3.444629,4.1897564,4.934884,5.6800117,6.4251394,5.239462,4.0555973,2.8699198,1.6842422,0.50037766,0.40972954,0.3208944,0.23024625,0.13959812,0.05076295,0.054388877,0.059827764,0.065266654,0.07070554,0.07433146,0.18492219,0.2955129,0.40429065,0.5148814,0.62547207,0.5493277,0.4749962,0.40066472,0.3245203,0.25018883,0.35171473,0.4550536,0.55839247,0.65991837,0.76325727,0.65810543,0.5529536,0.44780177,0.34264994,0.2374981,0.35171473,0.46774435,0.581961,0.6979906,0.8122072,0.6671702,0.52213323,0.3770962,0.23205921,0.0870222,0.38434806,0.68167394,0.9808127,1.2781386,1.5754645,2.1701162,2.764768,3.3594196,3.9558845,4.550536,4.4471974,4.345671,4.2423325,4.1408067,4.0374675,4.98746,5.9374523,6.887445,7.837437,8.78743,8.6877165,8.588004,8.488291,8.386765,8.287052,7.8319983,7.3769445,6.921891,6.4668374,6.011784,6.35806,6.7025228,7.0469856,7.3932614,7.7377243,7.7395372,7.743163,7.744976,7.746789,7.750415,7.3841968,7.019791,6.6553855,6.2891674,5.924762,5.7797246,5.634688,5.4896507,5.3446136,5.199577,7.9824743,10.765372,13.548269,16.329353,19.112251,16.775343,14.438434,12.099712,9.762803,7.4258947,6.825804,6.2257137,5.6256227,5.0255322,4.4254417,3.6494937,2.8753586,2.0994108,1.3252757,0.5493277,0.581961,0.61459434,0.64722764,0.67986095,0.7124943,2.3931105,4.071914,5.75253,7.4331465,9.11195,10.435412,11.757062,13.080525,14.402175,15.725637,13.017072,10.310318,7.6017523,4.894999,2.1882458,1.7694515,1.35247,0.9354887,0.5166943,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.10515183,0.09789998,0.09064813,0.08339628,0.07433146,0.07977036,0.08520924,0.09064813,0.09427405,0.099712946,0.09064813,0.07977036,0.07070554,0.059827764,0.05076295,0.059827764,0.07070554,0.07977036,0.09064813,0.099712946,0.099712946,0.099712946,0.099712946,0.099712946,0.099712946,0.13959812,0.1794833,0.21936847,0.25925365,0.2991388,0.26831847,0.23568514,0.2030518,0.17041849,0.13778515,0.29007402,0.44236287,0.5946517,0.7469406,0.89922947,1.2328146,1.5645868,1.8981718,2.229944,2.561716,2.960568,3.3576066,3.7546456,4.1516843,4.550536,4.559601,4.5704784,4.5795436,4.590421,4.599486,4.5233417,4.445384,4.367427,4.2894692,4.213325,3.4591327,2.7067533,1.9543737,1.2019942,0.44961473,0.3825351,0.3154555,0.24837588,0.1794833,0.11240368,0.87566096,1.6371052,2.4003625,3.1618068,3.925064,4.1281157,4.329355,4.5324063,4.7354584,4.936697,4.220577,3.5026438,2.7847104,2.0667772,1.3506571,1.0877775,0.824898,0.5620184,0.2991388,0.038072214,0.46230546,0.8883517,1.3125849,1.7368182,2.1628644,1.7295663,1.2980812,0.86478317,0.43329805,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.06707962,0.09789998,0.12690738,0.15772775,0.18673515,0.92823684,1.6679256,2.4076142,3.147303,3.8869917,3.7673361,3.6476808,3.5280252,3.4083695,3.2869012,2.7067533,2.128418,1.54827,0.968122,0.387974,0.6055295,0.823085,1.0406405,1.258196,1.4757515,1.1802386,0.88472575,0.58921283,0.2955129,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.09064813,0.16679256,0.24474995,0.32270733,0.40066472,0.41335547,0.42423326,0.43692398,0.44961473,0.46230546,0.5058166,0.5475147,0.58921283,0.6327239,0.6744221,0.58921283,0.5058166,0.42060733,0.33539808,0.25018883,0.24474995,0.23931105,0.23568514,0.23024625,0.22480737,0.1794833,0.13415924,0.09064813,0.045324065,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.6399758,1.2799516,1.9199274,2.5599031,3.199879,4.599486,5.999093,7.400513,8.80012,10.199727,8.399456,6.599184,4.800725,3.000453,1.2001812,4.3184767,7.4349594,10.553255,13.669738,16.788034,14.739386,12.692551,10.645717,8.597069,6.550234,5.823236,5.0944247,4.367427,3.6404288,2.911618,3.3993049,3.8869917,4.3746786,4.8623657,5.3500524,5.859495,6.3707504,6.880193,7.3896356,7.900891,10.792566,13.684241,16.57773,19.469404,22.362894,20.62245,18.882006,17.141562,15.40293,13.662486,12.754191,11.847711,10.939416,10.032935,9.12464,10.245051,11.365462,12.485873,13.604471,14.724882,12.540262,10.355642,8.1692095,5.9845896,3.7999697,5.4552045,7.1104393,8.765674,10.420909,12.07433,9.759177,7.4458375,5.130684,2.8155308,0.50037766,1.0569572,1.6153497,2.1719291,2.7303216,3.2869012,2.6922495,2.0975976,1.502946,0.90829426,0.31182957,0.25925365,0.20667773,0.15410182,0.10333887,0.05076295,0.04169814,0.034446288,0.027194439,0.01994259,0.012690738,1.1657349,2.3169663,3.4700103,4.6230545,5.774286,5.1125546,4.4508233,3.787279,3.1255474,2.4620032,2.752077,3.0421512,3.3322253,3.6222992,3.9123733,4.3420453,4.7717175,5.2032027,5.632875,6.0625467,8.096691,10.1326475,12.166792,14.202749,16.236893,17.864933,19.492973,21.119202,22.747242,24.375282,27.161806,29.950142,32.73848,35.525,38.31334,39.223446,40.13174,41.041847,41.951954,42.86206,41.112553,39.363045,37.61172,35.862213,34.112705,32.232662,30.35262,28.472578,26.592535,24.712494,23.550385,22.388275,21.224354,20.062244,18.900135,18.577427,18.25472,17.932013,17.609306,17.288412,17.859495,18.43239,19.005287,19.578182,20.149265,17.304728,14.46019,11.615651,8.7693,5.924762,7.7322855,9.539809,11.347333,13.154857,14.96238,17.719896,20.477413,23.234928,25.992445,28.74996,23.13159,17.515032,11.896661,6.2801023,0.66173136,1.1929294,1.7223145,2.2516994,2.7828975,3.3122826,2.6704938,2.0268922,1.3851035,0.7433147,0.099712946,0.17585737,0.25018883,0.3245203,0.40066472,0.4749962,0.50037766,0.52575916,0.5493277,0.5747091,0.6000906,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.21211663,0.36259252,0.51306844,0.66173136,0.8122072,0.6508536,0.48768693,0.3245203,0.16316663,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.387974,0.774135,1.162109,1.550083,1.938057,1.7368182,1.5373923,1.3379664,1.1367276,0.93730164,0.87566096,0.8122072,0.7505665,0.6871128,0.62547207,0.97537386,1.3252757,1.6751775,2.0250793,2.374981,3.4500678,4.5251546,5.600241,6.6753283,7.750415,6.2873545,4.8242936,3.3630457,1.8999848,0.43692398,0.34990177,0.26287958,0.17585737,0.0870222,0.0,0.0,0.0,0.0,0.0,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.19942589,0.21211663,0.22480737,0.2374981,0.25018883,0.34990177,0.44961473,0.5493277,0.6508536,0.7505665,0.6000906,0.44961473,0.2991388,0.15047589,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.36259252,0.72518504,1.0877775,1.4503701,1.8129625,2.4130533,3.0131438,3.6132345,4.213325,4.8116026,4.349297,3.8869917,3.4246864,2.962381,2.5000753,3.6494937,4.800725,5.9501433,7.0995617,8.2507925,8.238102,8.225411,8.212721,8.200029,8.187339,7.549176,6.9128265,6.2746634,5.638314,5.0001507,5.388125,5.774286,6.16226,6.550234,6.9382076,7.1992745,7.462154,7.7250338,7.987913,8.2507925,7.799365,7.3497505,6.9001355,6.450521,6.000906,5.7253356,5.4497657,5.1741953,4.900438,4.6248674,7.837437,11.050007,14.262577,17.475147,20.687716,18.011784,15.337664,12.661731,9.987611,7.311678,6.7496595,6.187641,5.6256227,5.0617914,4.499773,3.636803,2.7756457,1.9126755,1.0497054,0.18673515,0.21211663,0.2374981,0.26287958,0.28826106,0.31182957,1.4376793,2.561716,3.6875658,4.8134155,5.9374523,7.799365,9.663091,11.525003,13.386916,15.250641,12.562017,9.875207,7.1865835,4.499773,1.8129625,1.4757515,1.1367276,0.7995165,0.46230546,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.17585737,0.22480737,0.2755703,0.3245203,0.37528324,0.2991388,0.22480737,0.15047589,0.07433146,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,1.1874905,2.3133402,3.437377,4.5632267,5.6872635,5.6999545,5.712645,5.7253356,5.7380266,5.750717,5.6491914,5.5494785,5.4497657,5.3500524,5.2503395,4.2006345,3.150929,2.0994108,1.0497054,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,1.1131591,2.0994108,3.0874753,4.07554,5.0617914,4.0501585,3.0367124,2.0250793,1.0116332,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,1.1004683,2.0123885,2.9243085,3.8380418,4.749962,4.512464,4.274966,4.0374675,3.7999697,3.5624714,2.8753586,2.1882458,1.49932,0.8122072,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.21211663,0.2374981,0.26287958,0.28826106,0.31182957,0.25018883,0.18673515,0.12509441,0.06164073,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,2.525457,4.98746,7.4494634,9.91328,12.375282,9.900589,7.4258947,4.949388,2.474694,0.0,3.2125697,6.4251394,9.637709,12.850279,16.062849,13.974316,11.887595,9.799063,7.7123427,5.6256227,4.98746,4.349297,3.7129474,3.0747845,2.4366217,2.9750717,3.5117085,4.0501585,4.5867953,5.125245,5.5875506,6.049856,6.5121617,6.9744673,7.4367723,10.662033,13.887294,17.112555,20.337814,23.563074,21.574255,19.587248,17.60024,15.613234,13.6244135,12.850279,12.07433,11.300196,10.524248,9.750113,11.4126,13.075087,14.737573,16.400059,18.062546,15.136425,12.212116,9.287807,6.3616858,3.437377,5.7253356,8.013294,10.29944,12.5873995,14.875358,11.999999,9.12464,6.249282,3.3757362,0.50037766,1.162109,1.8256533,2.4873846,3.149116,3.8126602,3.1255474,2.4366217,1.7495089,1.062396,0.37528324,0.31182957,0.25018883,0.18673515,0.12509441,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,1.3125849,2.6251698,3.9377546,5.2503395,6.5629244,5.612932,4.6629395,3.7129474,2.762955,1.8129625,1.4503701,1.0877775,0.72518504,0.36259252,0.0,0.19942589,0.40066472,0.6000906,0.7995165,1.0007553,3.4119956,5.825049,8.238102,10.649343,13.062395,14.663241,16.262274,17.863121,19.462152,21.063,24.737875,28.41275,32.087624,35.7625,39.437374,41.186886,42.938206,44.687714,46.437225,48.186733,46.174343,44.161957,42.149567,40.13718,38.12479,36.012688,33.90059,31.786673,29.674572,27.56247,26.12479,24.68711,23.249432,21.811752,20.375887,19.812056,19.250036,18.688019,18.124187,17.562168,18.17495,18.787731,19.400513,20.013294,20.624262,17.199575,13.77489,10.3502035,6.925517,3.5008307,5.176008,6.849373,8.52455,10.199727,11.874905,15.899682,19.926271,23.949236,27.974012,32.000603,25.762197,19.523794,13.287203,7.0506115,0.8122072,1.4630609,2.1121013,2.762955,3.4119956,4.062849,3.2742105,2.4873846,1.7005589,0.9119202,0.12509441,0.21211663,0.2991388,0.387974,0.4749962,0.5620184,0.6000906,0.63816285,0.6744221,0.7124943,0.7505665,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.17223145,0.2955129,0.4169814,0.5402629,0.66173136,0.5656443,0.46774435,0.36984438,0.27194437,0.17585737,0.25925365,0.3444629,0.42967212,0.5148814,0.6000906,0.48224804,0.36440548,0.24837588,0.13053331,0.012690738,0.40791658,0.8031424,1.1983683,1.5917811,1.987007,1.9072367,1.8274662,1.7476959,1.6679256,1.5881553,1.4431182,1.2980812,1.1530442,1.0080072,0.8629702,1.0950294,1.3270886,1.5591478,1.79302,2.0250793,2.907992,3.7890918,4.6720047,5.5549173,6.43783,5.282973,4.1281157,2.9732587,1.8165885,0.66173136,0.5293851,0.39703882,0.26469254,0.13234627,0.0,0.0,0.0,0.0,0.0,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.15954071,0.17041849,0.1794833,0.19036107,0.19942589,0.27919623,0.36077955,0.4405499,0.52032024,0.6000906,0.48043507,0.36077955,0.23931105,0.11965553,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.29007402,0.58014804,0.87022203,1.1602961,1.4503701,1.9308052,2.4094272,2.8898623,3.3702974,3.8507326,3.482701,3.1146698,2.7466383,2.38042,2.0123885,2.9351864,3.8579843,4.780782,5.7017674,6.624565,6.695271,6.7641635,6.834869,6.9055743,6.9744673,7.0125394,7.0506115,7.0868707,7.124943,7.1630154,7.217404,7.271793,7.327995,7.382384,7.4367723,7.7359114,8.033237,8.330563,8.627889,8.925215,8.653271,8.379513,8.107569,7.835624,7.5618668,6.9182653,6.2728505,5.6274357,4.9820213,4.3366065,6.8620634,9.38752,11.912977,14.436621,16.962078,14.817343,12.672608,10.527874,8.383139,6.2365913,5.732588,5.2267714,4.7227674,4.216951,3.7129474,3.002266,2.2933977,1.5827163,0.872035,0.16316663,0.18492219,0.20667773,0.23024625,0.2520018,0.2755703,1.1874905,2.0994108,3.0131438,3.925064,4.836984,6.3218007,7.806617,9.293246,10.778063,12.262879,10.101828,7.9425893,5.7815375,3.6222992,1.4630609,1.1893034,0.91735905,0.64541465,0.37165734,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.065266654,0.07977036,0.09427405,0.11059072,0.12509441,0.40247768,0.67986095,0.9572442,1.2346275,1.5120108,1.2817645,1.0533313,0.823085,0.59283876,0.36259252,0.3770962,0.39159992,0.40791658,0.4224203,0.43692398,0.41335547,0.387974,0.36259252,0.33721104,0.31182957,0.28826106,0.26287958,0.2374981,0.21211663,0.18673515,0.19217403,0.19761293,0.2030518,0.20667773,0.21211663,0.2520018,0.291887,0.33177215,0.37165734,0.41335547,1.2400664,2.0667772,2.8953013,3.7220123,4.550536,4.615803,4.6792564,4.744523,4.8097897,4.8750563,4.7898474,4.704638,4.6194286,4.5342193,4.4508233,3.6222992,2.7955883,1.9670644,1.1403534,0.31182957,0.67079616,1.0279498,1.3851035,1.742257,2.0994108,1.8202144,1.5392052,1.260009,0.9808127,0.69980353,1.6026589,2.5055144,3.4083695,4.309412,5.2122674,4.3565493,3.5026438,2.6469254,1.79302,0.93730164,0.78319985,0.62728506,0.47318324,0.31726846,0.16316663,0.15047589,0.13778515,0.12509441,0.11240368,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.8792868,1.6099107,2.3405347,3.0693457,3.7999697,3.6966307,3.5951047,3.491766,3.39024,3.2869012,2.6505513,2.0123885,1.3742256,0.73787576,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.17041849,0.19036107,0.21030366,0.23024625,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,2.0504606,4.0501585,6.049856,8.049554,10.049252,8.0604315,6.069799,4.079166,2.0903459,0.099712946,2.657803,5.2140803,7.7721705,10.330261,12.8865385,12.092461,11.298383,10.502492,9.708415,8.912524,8.093065,7.271793,6.452334,5.632875,4.8134155,5.045475,5.277534,5.5095935,5.7416525,5.975525,5.977338,5.979151,5.9827766,5.9845896,5.9882154,8.560809,11.13159,13.704185,16.276777,18.849373,17.694515,16.539658,15.384801,14.229943,13.075087,12.754191,12.43511,12.114216,11.795135,11.47424,12.63091,13.785768,14.940624,16.095482,17.25034,15.129172,13.009819,10.890467,8.7693,6.6499467,8.234476,9.820818,11.405348,12.989877,14.574407,11.954676,9.334945,6.7152133,4.0954823,1.4757515,1.9851941,2.4946365,3.005892,3.5153344,4.024777,3.8507326,3.6748753,3.5008307,3.3249733,3.150929,2.5345216,1.9199274,1.305333,0.69073874,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,1.0497054,2.0994108,3.149116,4.2006345,5.2503395,4.4907084,3.729264,2.9696326,2.2100015,1.4503701,1.162109,0.87566096,0.5873999,0.2991388,0.012690738,0.19942589,0.387974,0.5747091,0.76325727,0.9499924,2.8699198,4.7898474,6.7097745,8.629702,10.549629,11.947423,13.345218,14.743011,16.138992,17.536787,20.655083,23.771564,26.88986,30.006344,33.124638,35.02825,36.930046,38.831844,40.735455,42.637253,41.694515,40.751774,39.809032,38.868103,37.925365,36.69255,35.459736,34.22692,32.99592,31.763105,30.265598,28.768091,27.270584,25.773077,24.27557,23.14972,22.025682,20.899832,19.775795,18.649946,18.958149,19.26454,19.572744,19.879135,20.187338,17.491463,14.7974,12.103338,9.407463,6.7134004,8.109382,9.507175,10.90497,12.302764,13.700559,16.14987,18.600996,21.050308,23.49962,25.950747,21.27149,16.594046,11.916603,7.2409725,2.561716,3.0348995,3.5080826,3.9794528,4.4526362,4.9258194,4.478018,4.0302157,3.5824142,3.1346123,2.6868105,3.0856624,3.482701,3.87974,4.2767787,4.6756306,4.604925,4.5342193,4.465327,4.3946214,4.325729,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.13234627,0.22662032,0.32270733,0.4169814,0.51306844,0.48043507,0.44780177,0.41516843,0.3825351,0.34990177,0.48224804,0.61459434,0.7469406,0.8792868,1.0116332,0.81583315,0.61822027,0.42060733,0.2229944,0.025381476,0.42785916,0.83033687,1.2328146,1.6352923,2.03777,2.077655,2.1175404,2.1574254,2.1973107,2.2371957,2.0105755,1.7821422,1.5555218,1.3270886,1.1004683,1.214685,1.3307146,1.4449311,1.5591478,1.6751775,2.3641033,3.054842,3.7455807,4.4345064,5.125245,4.2767787,3.4301252,2.5816586,1.7350051,0.8883517,0.7106813,0.533011,0.35534066,0.17767033,0.0,0.0,0.0,0.0,0.0,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.11965553,0.12690738,0.13415924,0.14322405,0.15047589,0.21030366,0.27013144,0.32995918,0.38978696,0.44961473,0.36077955,0.27013144,0.1794833,0.09064813,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.21755551,0.43511102,0.6526665,0.87022203,1.0877775,1.4467441,1.8075237,2.1683033,2.5272698,2.8880494,2.6142921,2.3423476,2.0704033,1.7966459,1.5247015,2.220879,2.9152439,3.6096084,4.305786,5.0001507,5.1524396,5.3047285,5.4570174,5.6093063,5.7615952,6.474089,7.1865835,7.900891,8.613385,9.325879,9.046683,8.7693,8.491917,8.214534,7.93715,8.270736,8.602508,8.934279,9.267865,9.599637,9.5053625,9.409276,9.3150015,9.220728,9.12464,8.109382,7.0959353,6.0806766,5.0654173,4.0501585,5.8866897,7.7250338,9.563377,11.399909,13.238253,11.622903,10.007553,8.392203,6.776854,5.163317,4.7155156,4.267714,3.8199122,3.3721104,2.9243085,2.3677292,1.8093367,1.2527572,0.69436467,0.13778515,0.15772775,0.17767033,0.19761293,0.21755551,0.2374981,0.93730164,1.6371052,2.3369088,3.0367124,3.738329,4.844236,5.9519563,7.059676,8.167397,9.275117,7.6416373,6.009971,4.3783045,2.7448254,1.1131591,0.90466833,0.6979906,0.4894999,0.28282216,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.054388877,0.072518505,0.09064813,0.10696479,0.12509441,0.69255173,1.260009,1.8274662,2.3949237,2.962381,2.4891977,2.0178273,1.5446441,1.0732739,0.6000906,0.629098,0.65991837,0.69073874,0.7197462,0.7505665,0.6508536,0.5493277,0.44961473,0.34990177,0.25018883,0.2755703,0.2991388,0.3245203,0.34990177,0.37528324,0.38434806,0.39522585,0.40429065,0.41516843,0.42423326,0.49312583,0.56020546,0.62728506,0.69436467,0.76325727,1.2926424,1.8220274,2.3532255,2.8826106,3.4119956,3.529838,3.6476808,3.7655232,3.8833659,3.9993954,3.930503,3.8597972,3.7890918,3.720199,3.6494937,3.045777,2.4402475,1.8347181,1.2291887,0.62547207,1.3397794,2.0540867,2.770207,3.484514,4.2006345,3.6150475,3.0294604,2.4456866,1.8600996,1.2745126,2.0921588,2.909805,3.727451,4.5450974,5.3627434,4.664753,3.966762,3.2705846,2.572594,1.8746033,1.5645868,1.2545701,0.9445535,0.6345369,0.3245203,0.2991388,0.2755703,0.25018883,0.22480737,0.19942589,0.15954071,0.11965553,0.07977036,0.03988518,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.65991837,1.2074331,1.7549478,2.3024626,2.8499773,2.8826106,2.9152439,2.9478772,2.9805105,3.0131438,2.4257438,1.8383441,1.2491312,0.66173136,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.12690738,0.14322405,0.15772775,0.17223145,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,1.5754645,3.1128569,4.650249,6.187641,7.7250338,6.2202744,4.7155156,3.2107568,1.7041848,0.19942589,2.1030366,4.004834,5.908445,7.8102427,9.712041,10.210606,10.707357,11.205922,11.702674,12.199425,11.1968565,10.194288,9.19172,8.189152,7.1883965,7.115878,7.0433598,6.970841,6.8983226,6.825804,6.3671246,5.910258,5.4515786,4.994712,4.537845,6.4577727,8.3777,10.297627,12.217555,14.137483,13.8147745,13.492067,13.16936,12.846653,12.525759,12.659918,12.79589,12.930049,13.064208,13.200181,13.847408,14.494636,15.141864,15.790904,16.438131,15.121921,13.807523,12.493125,11.176914,9.862516,10.745429,11.628342,12.509441,13.392355,14.275268,11.909351,9.545248,7.179332,4.8152285,2.4493124,2.808279,3.1654327,3.5225863,3.87974,4.2368937,4.5759177,4.9131284,5.2503395,5.5875506,5.924762,4.7572136,3.589666,2.422118,1.2545701,0.0870222,0.07070554,0.052575916,0.034446288,0.018129626,0.0,0.7868258,1.5754645,2.3622901,3.149116,3.9377546,3.3666716,2.7974012,2.228131,1.6570477,1.0877775,0.87566096,0.66173136,0.44961473,0.2374981,0.025381476,0.19942589,0.37528324,0.5493277,0.72518504,0.89922947,2.327844,3.7546456,5.18326,6.6100616,8.036863,9.233418,10.428161,11.622903,12.817645,14.012388,16.57229,19.132195,21.692097,24.252,26.811903,28.867804,30.92189,32.97779,35.031876,37.087776,37.214684,37.34159,37.47031,37.597218,37.724125,37.37241,37.020695,36.667168,36.315453,35.961926,34.40459,32.847256,31.28992,29.732586,28.175251,26.487383,24.799515,23.111647,21.425592,19.737724,19.739536,19.743162,19.744976,19.746788,19.750414,17.785164,15.819912,13.85466,11.889409,9.924157,11.044568,12.164979,13.28539,14.405801,15.524399,16.400059,17.27572,18.149569,19.025229,19.899076,16.782595,13.664299,10.547816,7.4295206,4.313038,4.606738,4.902251,5.197764,5.4932766,5.7869763,5.6800117,5.573047,5.464269,5.3573046,5.2503395,5.957395,6.6644506,7.3733187,8.080374,8.78743,8.609759,8.432089,8.254418,8.076748,7.900891,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.092461094,0.15954071,0.22662032,0.2955129,0.36259252,0.39522585,0.42785916,0.4604925,0.49312583,0.52575916,0.70524246,0.88472575,1.064209,1.2455053,1.4249886,1.1476053,0.87022203,0.59283876,0.3154555,0.038072214,0.44780177,0.8575313,1.2672608,1.6769904,2.08672,2.2480736,2.4076142,2.5671551,2.7266958,2.8880494,2.5780327,2.268016,1.9579996,1.647983,1.3379664,1.3343405,1.3325275,1.3307146,1.3270886,1.3252757,1.8220274,2.3205922,2.817344,3.3159087,3.8126602,3.2723975,2.7321346,2.1918716,1.651609,1.1131591,0.8901646,0.6671702,0.44417584,0.2229944,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.07977036,0.08520924,0.09064813,0.09427405,0.099712946,0.13959812,0.1794833,0.21936847,0.25925365,0.2991388,0.23931105,0.1794833,0.11965553,0.059827764,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14503701,0.29007402,0.43511102,0.58014804,0.72518504,0.9644961,1.2056202,1.4449311,1.6842422,1.9253663,1.7476959,1.5700256,1.3923552,1.214685,1.0370146,1.504759,1.9725033,2.4402475,2.907992,3.3757362,3.6096084,3.8452935,4.079166,4.314851,4.550536,5.9374523,7.324369,8.713099,10.100015,11.486931,10.877775,10.266808,9.657652,9.046683,8.437528,8.805559,9.171778,9.539809,9.907841,10.275872,10.357455,10.440851,10.522435,10.605831,10.687414,9.302311,7.9172077,6.532104,5.147001,3.7618973,4.9131284,6.0625467,7.211965,8.363196,9.512614,8.42665,7.3424983,6.258347,5.1723824,4.0882306,3.6966307,3.3068438,2.9170568,2.5272698,2.137483,1.7331922,1.3270886,0.922798,0.5166943,0.11240368,0.13053331,0.14684997,0.16497959,0.18310922,0.19942589,0.6871128,1.1747998,1.6624867,2.1501737,2.6378605,3.3666716,4.0972953,4.8279195,5.5567303,6.2873545,5.18326,4.077353,2.9732587,1.8673514,0.76325727,0.6200332,0.47680917,0.33539808,0.19217403,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.045324065,0.065266654,0.08520924,0.10515183,0.12509441,0.9826257,1.840157,2.6976883,3.5552197,4.4127507,3.6966307,2.9823234,2.268016,1.551896,0.8375887,0.88291276,0.92823684,0.97174793,1.017072,1.062396,0.8883517,0.7124943,0.53663695,0.36259252,0.18673515,0.26287958,0.33721104,0.41335547,0.48768693,0.5620184,0.57833505,0.59283876,0.6073425,0.62184614,0.63816285,0.7324369,0.82671094,0.922798,1.017072,1.1131591,1.3452182,1.5772774,1.8093367,2.0432088,2.275268,2.4456866,2.6142921,2.7847104,2.955129,3.1255474,3.0693457,3.0149567,2.960568,2.904366,2.8499773,2.467442,2.084907,1.7023718,1.3198367,0.93730164,2.0105755,3.0820365,4.15531,5.2267714,6.300045,5.40988,4.519716,3.6295512,2.7393866,1.8492218,2.5816586,3.3140955,4.0483456,4.780782,5.5132194,4.972956,4.4326935,3.8924308,3.3521678,2.811905,2.3477864,1.8818551,1.4177368,0.95180535,0.48768693,0.44961473,0.41335547,0.37528324,0.33721104,0.2991388,0.23931105,0.1794833,0.11965553,0.059827764,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.4405499,0.80495536,1.1693609,1.5355793,1.8999848,2.0667772,2.2353828,2.4021754,2.570781,2.7375734,2.1991236,1.6624867,1.1258497,0.5873999,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.08520924,0.09427405,0.10515183,0.11421664,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,1.1004683,2.175555,3.2506418,4.325729,5.4008155,4.3801174,3.3594196,2.3405347,1.3198367,0.2991388,1.54827,2.7955883,4.0429068,5.290225,6.5375433,8.326937,10.118144,11.907538,13.696932,15.488139,14.302462,13.116784,11.9329195,10.747242,9.563377,9.184468,8.807372,8.430276,8.05318,7.6742706,6.7569118,5.8395524,4.9221935,4.004834,3.0874753,4.3547363,5.621997,6.889258,8.158332,9.425592,9.935035,10.444477,10.955733,11.465176,11.974618,12.565643,13.154857,13.745882,14.335095,14.924308,15.065719,15.2053175,15.344915,15.484513,15.624111,15.114669,14.6052265,14.095784,13.584529,13.075087,13.254569,13.435865,13.615349,13.794832,13.974316,11.864027,9.755551,7.645263,5.5349746,3.4246864,3.6295512,3.834416,4.0392804,4.2441454,4.4508233,5.2992897,6.149569,6.9998484,7.850128,8.700407,6.979906,5.2594047,3.540716,1.8202144,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.52575916,1.0497054,1.5754645,2.0994108,2.6251698,2.2444477,1.8655385,1.4848163,1.1059072,0.72518504,0.5873999,0.44961473,0.31182957,0.17585737,0.038072214,0.19942589,0.36259252,0.52575916,0.6871128,0.85027945,1.7857682,2.7194438,3.6549325,4.590421,5.52591,6.5176005,7.509291,8.502794,9.494485,10.487988,12.489499,14.492823,16.494333,18.497658,20.499168,22.707355,24.915545,27.12192,29.330109,31.538298,32.73485,33.93322,35.129776,36.328144,37.5247,38.052273,38.579845,39.107414,39.634987,40.16256,38.5454,36.926422,35.309258,33.692097,32.074936,29.825047,27.575161,25.325274,23.075388,20.8255,20.522736,20.219973,19.917208,19.614443,19.311678,18.07705,16.842422,15.607795,14.373167,13.136727,13.979754,14.8227825,15.66581,16.507025,17.350052,16.650248,15.950445,15.250641,14.5508375,13.849221,12.291886,10.734551,9.177217,7.6198816,6.0625467,6.1803894,6.298232,6.414262,6.532104,6.6499467,6.882006,7.115878,7.3479376,7.5799966,7.8120556,8.830941,9.848013,10.865085,11.882156,12.899229,12.6145935,12.329959,12.045323,11.760688,11.47424,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.052575916,0.092461094,0.13234627,0.17223145,0.21211663,0.3100166,0.40791658,0.5058166,0.60190356,0.69980353,0.92823684,1.1548572,1.3832904,1.6099107,1.8383441,1.4793775,1.1222239,0.7650702,0.40791658,0.05076295,0.46774435,0.88472575,1.3017071,1.7205015,2.137483,2.4166791,2.6976883,2.9768846,3.2578938,3.53709,3.1454902,2.752077,2.3604772,1.9670644,1.5754645,1.455809,1.3343405,1.214685,1.0950294,0.97537386,1.2799516,1.5845293,1.889107,2.1954978,2.5000753,2.268016,2.034144,1.8020848,1.5700256,1.3379664,1.0696479,0.8031424,0.53482395,0.26831847,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.03988518,0.04169814,0.045324065,0.047137026,0.05076295,0.07070554,0.09064813,0.11059072,0.13053331,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.072518505,0.14503701,0.21755551,0.29007402,0.36259252,0.48224804,0.60190356,0.72337204,0.8430276,0.96268314,0.8792868,0.79770356,0.71430725,0.6327239,0.5493277,0.7904517,1.0297627,1.2708868,1.5101979,1.7495089,2.0667772,2.3858588,2.7031271,3.0203958,3.3376641,5.4008155,7.462154,9.525306,11.588457,13.649796,12.707055,11.764315,10.823386,9.880646,8.937905,9.340384,9.742861,10.145339,10.547816,10.950294,11.209548,11.470614,11.729868,11.989121,12.250188,10.49524,8.740293,6.985345,5.230397,3.4754493,3.9377546,4.40006,4.8623657,5.3246713,5.7869763,5.23221,4.6774435,4.122677,3.5679104,3.0131438,2.6795588,2.3477864,2.0142014,1.6824293,1.3506571,1.0968424,0.8448406,0.59283876,0.34083697,0.0870222,0.10333887,0.11784257,0.13234627,0.14684997,0.16316663,0.43692398,0.7124943,0.9880646,1.261822,1.5373923,1.889107,2.2426348,2.5943494,2.9478772,3.299592,2.72307,2.1447346,1.5682126,0.9898776,0.41335547,0.33539808,0.2574407,0.1794833,0.10333887,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.034446288,0.058014803,0.07977036,0.10333887,0.12509441,1.2726997,2.420305,3.5679104,4.7155156,5.863121,4.9058766,3.9468195,2.9895754,2.032331,1.0750868,1.1349145,1.1947423,1.2545701,1.3143979,1.3742256,1.1258497,0.87566096,0.62547207,0.37528324,0.12509441,0.25018883,0.37528324,0.50037766,0.62547207,0.7505665,0.7705091,0.7904517,0.8103943,0.83033687,0.85027945,0.97174793,1.0950294,1.2183108,1.3397794,1.4630609,1.3977941,1.3325275,1.2672608,1.2019942,1.1367276,1.3597219,1.5827163,1.8057107,2.0268922,2.2498865,2.2100015,2.1701162,2.1302311,2.0903459,2.0504606,1.889107,1.7295663,1.5700256,1.4104849,1.2491312,2.6795588,4.1099863,5.540414,6.970841,8.399456,7.2047133,6.009971,4.8152285,3.6204863,2.4257438,3.0729716,3.720199,4.367427,5.0146546,5.661882,5.279347,4.896812,4.514277,4.1317415,3.7492065,3.1291735,2.5091403,1.889107,1.2708868,0.6508536,0.6000906,0.5493277,0.50037766,0.44961473,0.40066472,0.3208944,0.23931105,0.15954071,0.07977036,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.21936847,0.40247768,0.5855869,0.7668832,0.9499924,1.2527572,1.5555218,1.8582866,2.1592383,2.4620032,1.9743162,1.4866294,1.0007553,0.51306844,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.04169814,0.047137026,0.052575916,0.058014803,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.62547207,1.2382535,1.8492218,2.4620032,3.0747845,2.5399606,2.0051367,1.4703126,0.9354887,0.40066472,0.9916905,1.5845293,2.1773682,2.770207,3.3630457,6.445082,9.527119,12.610968,15.693004,18.77504,17.408066,16.03928,14.672306,13.305332,11.938358,11.254871,10.573197,9.88971,9.208037,8.52455,7.1466985,5.77066,4.3928084,3.0149567,1.6371052,2.2516994,2.8681068,3.482701,4.0972953,4.7118897,6.055295,7.3968873,8.740293,10.081885,11.42529,12.469557,13.515636,14.559902,15.604169,16.650248,16.282217,15.914186,15.547967,15.179935,14.811904,15.107417,15.40293,15.6966305,15.992143,16.287657,15.765523,15.243389,14.719443,14.19731,13.675177,11.820516,9.965856,8.109382,6.2547207,4.40006,4.4526362,4.505212,4.557788,4.610364,4.6629395,6.0244746,7.3878226,8.749357,10.112705,11.47424,9.202598,6.930956,4.6575007,2.3858588,0.11240368,0.09064813,0.06707962,0.045324065,0.02175555,0.0,0.26287958,0.52575916,0.7868258,1.0497054,1.3125849,1.1222239,0.9318628,0.7433147,0.5529536,0.36259252,0.2991388,0.2374981,0.17585737,0.11240368,0.05076295,0.19942589,0.34990177,0.50037766,0.6508536,0.7995165,1.2418793,1.6842422,2.126605,2.570781,3.0131438,3.8017826,4.592234,5.382686,6.1731377,6.9617763,8.406708,9.851639,11.29657,12.741501,14.188245,16.54691,18.907387,21.267864,23.626528,25.987005,28.255022,30.523039,32.78924,35.05726,37.325275,38.732132,40.140804,41.547665,42.95452,44.363194,42.68439,41.0074,39.33041,37.65342,35.974617,33.162712,30.348993,27.537088,24.725183,21.913279,21.304123,20.696781,20.089437,19.482096,18.874754,18.37075,17.864933,17.359118,16.855114,16.349297,16.914942,17.480585,18.044416,18.610062,19.175705,16.900436,14.625169,12.349901,10.074633,7.799365,7.802991,7.804804,7.806617,7.8102427,7.8120556,7.752228,7.6924005,7.6325727,7.572745,7.512917,8.0858135,8.656897,9.229793,9.802689,10.375585,11.702674,13.029762,14.356851,15.685752,17.01284,16.619429,16.227829,15.834415,15.442815,15.049402,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.22480737,0.387974,0.5493277,0.7124943,0.87566096,1.1494182,1.4249886,1.7005589,1.9743162,2.2498865,1.8129625,1.3742256,0.93730164,0.50037766,0.06164073,0.48768693,0.9119202,1.3379664,1.7621996,2.1882458,2.5870976,2.9877625,3.386614,3.787279,4.1879435,3.7129474,3.2379513,2.762955,2.2879589,1.8129625,1.5754645,1.3379664,1.1004683,0.8629702,0.62547207,0.73787576,0.85027945,0.96268314,1.0750868,1.1874905,1.261822,1.3379664,1.4122978,1.4866294,1.5627737,1.2491312,0.93730164,0.62547207,0.31182957,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.52575916,0.9246109,1.3252757,1.7241274,2.124792,4.8623657,7.5999393,10.337513,13.075087,15.812659,14.538147,13.261822,11.9873085,10.712796,9.438283,9.875207,10.312131,10.750868,11.187792,11.624716,12.06164,12.500377,12.937301,13.374225,13.812962,11.6881695,9.563377,7.4367723,5.3119802,3.1871881,2.962381,2.7375734,2.5127661,2.2879589,2.0631514,2.03777,2.0123885,1.987007,1.9616255,1.938057,1.6624867,1.3869164,1.1131591,0.8375887,0.5620184,0.46230546,0.36259252,0.26287958,0.16316663,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.18673515,0.25018883,0.31182957,0.37528324,0.43692398,0.41335547,0.387974,0.36259252,0.33721104,0.31182957,0.26287958,0.21211663,0.16316663,0.11240368,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,1.5627737,3.000453,4.4381323,5.8758116,7.311678,6.11331,4.9131284,3.7129474,2.5127661,1.3125849,1.3869164,1.4630609,1.5373923,1.6117238,1.6878681,1.3633479,1.0370146,0.7124943,0.387974,0.06164073,0.2374981,0.41335547,0.5873999,0.76325727,0.93730164,0.96268314,0.9880646,1.0116332,1.0370146,1.062396,1.2128719,1.3633479,1.5120108,1.6624867,1.8129625,1.4503701,1.0877775,0.72518504,0.36259252,0.0,0.2755703,0.5493277,0.824898,1.1004683,1.3742256,1.3506571,1.3252757,1.2998942,1.2745126,1.2491312,1.3125849,1.3742256,1.4376793,1.49932,1.5627737,3.350355,5.137936,6.925517,8.713099,10.500679,8.999546,7.500226,5.999093,4.499773,3.000453,3.5624714,4.12449,4.688321,5.2503395,5.812358,5.5875506,5.3627434,5.137936,4.9131284,4.688321,3.9123733,3.1382382,2.3622901,1.5881553,0.8122072,0.7505665,0.6871128,0.62547207,0.5620184,0.50037766,0.40066472,0.2991388,0.19942589,0.099712946,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.43692398,0.87566096,1.3125849,1.7495089,2.1882458,1.7495089,1.3125849,0.87566096,0.43692398,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.15047589,0.2991388,0.44961473,0.6000906,0.7505665,0.69980353,0.6508536,0.6000906,0.5493277,0.50037766,0.43692398,0.37528324,0.31182957,0.25018883,0.18673515,4.5632267,8.937905,13.312584,17.687263,22.061941,20.511858,18.961775,17.411694,15.861609,14.313339,13.325275,12.337211,11.349146,10.362894,9.374829,7.5364857,5.6999545,3.8616104,2.0250793,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,2.175555,4.349297,6.5248523,8.700407,10.874149,12.375282,13.874602,15.375735,16.875055,18.374376,17.500528,16.624866,15.749206,14.875358,13.999697,15.100165,16.200634,17.29929,18.399757,19.500225,18.274662,17.050913,15.825351,14.599788,13.374225,11.775192,10.174346,8.575313,6.9744673,5.375434,5.275721,5.1741953,5.0744824,4.974769,4.8750563,6.7496595,8.624263,10.500679,12.375282,14.249886,11.42529,8.600695,5.774286,2.94969,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.19942589,0.33721104,0.4749962,0.61278135,0.7505665,0.69980353,0.6508536,0.6000906,0.5493277,0.50037766,1.0877775,1.6751775,2.2625773,2.8499773,3.437377,4.325729,5.2122674,6.1006193,6.987158,7.8755093,10.388275,12.899229,15.411995,17.92476,20.437527,23.77519,27.112856,30.45052,33.788185,37.125847,39.411995,41.69995,43.98791,46.274055,48.562016,46.8252,45.086567,43.349747,41.61293,39.8743,36.500374,33.124638,29.750715,26.374979,22.999243,22.087322,21.175404,20.26167,19.34975,18.43783,18.662638,18.887444,19.112251,19.337059,19.561867,19.850128,20.138388,20.424837,20.713097,20.999546,17.150625,13.299893,9.449161,5.600241,1.7495089,3.3122826,4.8750563,6.43783,8.000604,9.563377,9.325879,9.086569,8.8508835,8.613385,8.375887,9.287807,10.199727,11.111648,12.025381,12.937301,14.574407,16.213324,17.85043,19.487535,21.12464,20.624262,20.125698,19.62532,19.124943,18.624565,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.26469254,0.4169814,0.56927025,0.72337204,0.87566096,1.1004683,1.3252757,1.550083,1.7748904,1.9996977,1.7803292,1.5591478,1.3397794,1.1204109,0.89922947,1.1566701,1.4141108,1.6733645,1.9308052,2.1882458,2.6505513,3.1128569,3.5751622,4.0374675,4.499773,4.100921,3.7002566,3.299592,2.9007401,2.5000753,2.1193533,1.7404441,1.3597219,0.9808127,0.6000906,0.6979906,0.79589057,0.8919776,0.9898776,1.0877775,1.1222239,1.1566701,1.1929294,1.2273756,1.261822,1.0098201,0.75781834,0.5058166,0.2520018,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.059827764,0.07070554,0.07977036,0.09064813,0.099712946,0.42423326,0.7505665,1.0750868,1.3996071,1.7241274,4.02659,6.3290524,8.6333275,10.93579,13.238253,12.130532,11.022813,9.915092,8.807372,7.699652,8.201842,8.705847,9.208037,9.710228,10.212419,10.741803,11.273002,11.802386,12.331772,12.862969,11.091705,9.322253,7.552802,5.7833505,4.0120864,3.7220123,3.4319382,3.141864,2.8517902,2.561716,2.6868105,2.811905,2.9369993,3.0620937,3.1871881,2.8028402,2.4166791,2.032331,1.647983,1.261822,1.0279498,0.79226464,0.55839247,0.32270733,0.0870222,0.09064813,0.092461094,0.09427405,0.09789998,0.099712946,0.15228885,0.20486477,0.2574407,0.3100166,0.36259252,0.34264994,0.32270733,0.30276474,0.28282216,0.26287958,0.21936847,0.17767033,0.13415924,0.092461094,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,1.3996071,2.6995013,3.9993954,5.2992897,6.599184,5.5929894,4.5849824,3.576975,2.570781,1.5627737,1.6624867,1.7621996,1.8619126,1.9616255,2.0631514,2.0450218,2.0268922,2.0105755,1.9924458,1.9743162,1.8147756,1.6552348,1.4956942,1.3343405,1.1747998,1.167548,1.1602961,1.1530442,1.1457924,1.1367276,1.2726997,1.4068589,1.5428312,1.6769904,1.8129625,1.6606737,1.5083848,1.3542831,1.2019942,1.0497054,1.3905423,1.7295663,2.0704033,2.4094272,2.7502642,3.0892882,3.4301252,3.7709622,4.1099863,4.4508233,4.2876563,4.12449,3.9631362,3.7999697,3.636803,5.5095935,7.382384,9.255174,11.127964,13.000754,11.144281,9.28962,7.4349594,5.580299,3.7256382,3.9105604,4.0954823,4.2804046,4.465327,4.650249,4.4707656,4.2894692,4.1099863,3.930503,3.7492065,3.1291735,2.5091403,1.889107,1.2708868,0.6508536,0.6000906,0.5493277,0.50037766,0.44961473,0.40066472,0.3208944,0.23931105,0.15954071,0.07977036,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.052575916,0.054388877,0.058014803,0.059827764,0.06164073,0.07070554,0.07795739,0.08520924,0.092461094,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.34990177,0.69980353,1.0497054,1.3996071,1.7495089,1.3996071,1.0497054,0.69980353,0.34990177,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.11965553,0.23931105,0.36077955,0.48043507,0.6000906,0.56020546,0.52032024,0.48043507,0.4405499,0.40066472,0.34990177,0.2991388,0.25018883,0.19942589,0.15047589,3.7546456,7.360628,10.964798,14.57078,18.17495,16.856926,15.540715,14.222692,12.904668,11.586644,10.772624,9.956791,9.142771,8.326937,7.512917,6.0389786,4.5668526,3.094727,1.6226015,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,1.7404441,3.4790752,5.219519,6.9599633,8.700407,9.953164,11.204109,12.456866,13.709623,14.96238,14.743011,14.521831,14.302462,14.083094,13.861912,15.214382,16.566853,17.919323,19.271791,20.624262,18.92733,17.230396,15.531651,13.834718,12.137785,11.677292,11.2168,10.75812,10.297627,9.837135,9.935035,10.032935,10.130835,10.226922,10.324821,10.64753,10.970237,11.292944,11.615651,11.936545,9.683033,7.4277077,5.1723824,2.9170568,0.66173136,0.53663695,0.41335547,0.28826106,0.16316663,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.15954071,0.27013144,0.38072214,0.4894999,0.6000906,0.56020546,0.52032024,0.48043507,0.4405499,0.40066472,0.89560354,1.3905423,1.8854811,2.38042,2.8753586,3.7473936,4.6194286,5.4932766,6.3653116,7.2373466,9.224354,11.213174,13.200181,15.187187,17.174194,19.877321,22.580448,25.281763,27.98489,30.688017,33.066624,35.447044,37.827465,40.207886,42.58649,41.957394,41.32648,40.697384,40.068287,39.437374,36.614594,33.79181,30.97084,28.148058,25.325274,24.422419,23.519564,22.616709,21.715666,20.81281,20.669586,20.528175,20.38495,20.241728,20.100317,19.882761,19.665205,19.447649,19.230095,19.012539,15.754644,12.496751,9.24067,5.9827766,2.7248828,3.97764,5.230397,6.4831543,7.7340984,8.9868555,8.714911,8.442966,8.1692095,7.897265,7.6253204,8.239915,8.854509,9.469104,10.085511,10.700105,12.170418,13.640731,15.10923,16.579542,18.049856,17.553104,17.054539,16.557787,16.059223,15.56247,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.032633327,0.065266654,0.09789998,0.13053331,0.16316663,0.3045777,0.44780177,0.58921283,0.7324369,0.87566096,1.0497054,1.2255627,1.3996071,1.5754645,1.7495089,1.7476959,1.745883,1.742257,1.7404441,1.7368182,1.8274662,1.9181144,2.0069497,2.0975976,2.1882458,2.712192,3.2379513,3.7618973,4.2876563,4.8116026,4.4870825,4.162562,3.8380418,3.5117085,3.1871881,2.665055,2.1429217,1.6207886,1.0968424,0.5747091,0.65810543,0.73968875,0.823085,0.90466833,0.9880646,0.9826257,0.97718686,0.97174793,0.968122,0.96268314,0.7705091,0.57833505,0.38434806,0.19217403,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.045324065,0.052575916,0.059827764,0.06707962,0.07433146,0.3245203,0.5747091,0.824898,1.0750868,1.3252757,3.1926272,5.0599785,6.92733,8.794682,10.662033,9.7229185,8.781991,7.842876,6.9019485,5.962834,6.530291,7.0977483,7.665206,8.232663,8.80012,9.421967,10.045626,10.667472,11.289318,11.912977,10.497053,9.082943,7.667019,6.2529078,4.836984,4.4816437,4.1281157,3.7727752,3.4174345,3.0620937,3.3376641,3.6132345,3.8869917,4.162562,4.4381323,3.9431937,3.4482548,2.953316,2.4583774,1.9616255,1.5917811,1.2219368,0.8520924,0.48224804,0.11240368,0.10515183,0.09789998,0.09064813,0.08339628,0.07433146,0.11784257,0.15954071,0.2030518,0.24474995,0.28826106,0.27194437,0.2574407,0.24293698,0.22662032,0.21211663,0.17767033,0.14322405,0.10696479,0.072518505,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,1.2382535,2.4003625,3.5624714,4.7245803,5.8866897,5.0726695,4.256836,3.442816,2.6269827,1.8129625,1.938057,2.0631514,2.1882458,2.3133402,2.4366217,2.7266958,3.0167696,3.3068438,3.5969179,3.8869917,3.392053,2.8971143,2.4021754,1.9072367,1.4122978,1.3724127,1.3325275,1.2926424,1.2527572,1.2128719,1.3325275,1.452183,1.5718386,1.693307,1.8129625,1.8691645,1.9271792,1.9851941,2.0432088,2.0994108,2.5055144,2.909805,3.3159087,3.720199,4.12449,4.8297324,5.5349746,6.240217,6.94546,7.650702,7.262728,6.874754,6.48678,6.1006193,5.712645,7.6706448,9.626831,11.584831,13.54283,15.50083,13.289016,11.080828,8.870826,6.6608243,4.4508233,4.256836,4.064662,3.872488,3.680314,3.48814,3.3521678,3.2180085,3.0820365,2.9478772,2.811905,2.3477864,1.8818551,1.4177368,0.95180535,0.48768693,0.44961473,0.41335547,0.37528324,0.33721104,0.2991388,0.23931105,0.1794833,0.11965553,0.059827764,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.10515183,0.11059072,0.11421664,0.11965553,0.12509441,0.11421664,0.10515183,0.09427405,0.08520924,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.26287958,0.52575916,0.7868258,1.0497054,1.3125849,1.0497054,0.7868258,0.52575916,0.26287958,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.09064813,0.1794833,0.27013144,0.36077955,0.44961473,0.42060733,0.38978696,0.36077955,0.32995918,0.2991388,0.26287958,0.22480737,0.18673515,0.15047589,0.11240368,2.9478772,5.7815375,8.617011,11.452485,14.287958,13.201994,12.117842,11.0318775,9.947725,8.861761,8.219973,7.5781837,6.9345818,6.2927933,5.6491914,4.5432844,3.435564,2.327844,1.2201238,0.11240368,0.09064813,0.06707962,0.045324065,0.02175555,0.0,1.305333,2.610666,3.9141862,5.219519,6.5248523,7.5292335,8.535428,9.539809,10.54419,11.5503845,11.985496,12.420607,12.855718,13.290829,13.724127,15.330412,16.934883,18.539356,20.14564,21.750113,19.579996,17.40988,15.239763,13.069647,10.899531,11.579392,12.259253,12.940927,13.620788,14.300649,14.594349,14.889862,15.185374,15.480887,15.774588,14.545399,13.314397,12.085209,10.854207,9.625018,7.9407763,6.2547207,4.5704784,2.8844235,1.2001812,0.97537386,0.7505665,0.52575916,0.2991388,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.11965553,0.2030518,0.28463513,0.3680314,0.44961473,0.42060733,0.38978696,0.36077955,0.32995918,0.2991388,0.70342946,1.1040943,1.5083848,1.9108626,2.3133402,3.1708715,4.02659,4.8841214,5.7416525,6.599184,8.062244,9.525306,10.988366,12.449615,13.912675,15.979452,18.048042,20.11482,22.181597,24.250187,26.723068,29.19595,31.667017,34.1399,36.612778,37.08959,37.56821,38.04502,38.521828,39.00045,36.73062,34.45898,32.18915,29.919321,27.649492,26.757515,25.865538,24.971746,24.07977,23.187792,22.678349,22.167093,21.657652,21.148209,20.636953,19.915394,19.192022,18.470463,17.747091,17.025532,14.3604765,11.695421,9.030367,6.3653116,3.7002566,4.6429973,5.5857377,6.526665,7.4694057,8.412147,8.105756,7.797552,7.4893484,7.1829576,6.874754,7.192023,7.509291,7.8283725,8.145641,8.46291,9.764616,11.068136,12.3698435,13.671551,14.975071,14.480132,13.985193,13.490254,12.995316,12.500377,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.04169814,0.08520924,0.12690738,0.17041849,0.21211663,0.3444629,0.47680917,0.6091554,0.7433147,0.87566096,1.0007553,1.1258497,1.2491312,1.3742256,1.49932,1.7150626,1.9308052,2.1447346,2.3604772,2.5744069,2.4982624,2.420305,2.3423476,2.2643902,2.1882458,2.7756457,3.3630457,3.9504454,4.537845,5.125245,4.8750563,4.6248674,4.3746786,4.12449,3.874301,3.2107568,2.5453994,1.8800422,1.214685,0.5493277,0.61822027,0.6852999,0.7523795,0.8194591,0.8883517,0.8430276,0.79770356,0.7523795,0.7070554,0.66173136,0.5293851,0.39703882,0.26469254,0.13234627,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.030820364,0.034446288,0.03988518,0.045324065,0.05076295,0.22480737,0.40066472,0.5747091,0.7505665,0.9246109,2.3568513,3.7890918,5.223145,6.6553855,8.087626,7.315304,6.542982,5.77066,4.9983377,4.2242026,4.856927,5.4896507,6.1223745,6.755099,7.3878226,8.10213,8.81825,9.5325575,10.246864,10.962985,9.902402,8.841819,7.783048,6.722465,5.661882,5.243088,4.8224807,4.401873,3.9830787,3.5624714,3.9867048,4.4127507,4.836984,5.2630305,5.6872635,5.081734,4.478018,3.872488,3.2669585,2.663242,2.1574254,1.651609,1.1476053,0.6417888,0.13778515,0.11965553,0.10333887,0.08520924,0.06707962,0.05076295,0.08339628,0.11421664,0.14684997,0.1794833,0.21211663,0.2030518,0.19217403,0.18310922,0.17223145,0.16316663,0.13415924,0.10696479,0.07977036,0.052575916,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,1.0750868,2.0994108,3.1255474,4.1498713,5.1741953,4.552349,3.930503,3.3068438,2.6849976,2.0631514,2.2118144,2.3622901,2.5127661,2.663242,2.811905,3.4101827,4.006647,4.604925,5.2032027,5.7996674,4.9693303,4.1408067,3.3104696,2.4801328,1.649796,1.5772774,1.504759,1.4322405,1.3597219,1.2872034,1.3923552,1.4975071,1.6026589,1.7078108,1.8129625,2.079468,2.3477864,2.6142921,2.8826106,3.149116,3.6204863,4.0900435,4.559601,5.029158,5.5005283,6.5701766,7.6398244,8.709473,9.77912,10.850581,10.2378,9.625018,9.012237,8.399456,7.7866745,9.829884,11.873092,13.914488,15.957697,17.999092,15.435563,12.870221,10.304879,7.7395372,5.1741953,4.604925,4.0356545,3.4645715,2.8953013,2.324218,2.2353828,2.1447346,2.0558996,1.9652514,1.8746033,1.5645868,1.2545701,0.9445535,0.6345369,0.3245203,0.2991388,0.2755703,0.25018883,0.22480737,0.19942589,0.15954071,0.11965553,0.07977036,0.03988518,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.15772775,0.16497959,0.17223145,0.1794833,0.18673515,0.15954071,0.13234627,0.10515183,0.07795739,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.17585737,0.34990177,0.52575916,0.69980353,0.87566096,0.69980353,0.52575916,0.34990177,0.17585737,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.059827764,0.11965553,0.1794833,0.23931105,0.2991388,0.27919623,0.25925365,0.23931105,0.21936847,0.19942589,0.17585737,0.15047589,0.12509441,0.099712946,0.07433146,2.1392958,4.2042603,6.2692246,8.334189,10.399154,9.547061,8.694968,7.842876,6.9907837,6.1368785,5.667321,5.197764,4.7282066,4.256836,3.787279,3.045777,2.3024626,1.5591478,0.81764615,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.87022203,1.7404441,2.610666,3.4808881,4.349297,5.1071157,5.864934,6.622752,7.380571,8.138389,9.22798,10.31757,11.407161,12.496751,13.588155,15.444629,17.302916,19.15939,21.017675,22.87415,20.232662,17.589363,14.947877,12.304577,9.663091,11.483305,13.301706,15.121921,16.942135,18.76235,19.255476,19.746788,20.239914,20.73304,21.224354,18.441456,15.660371,12.877473,10.094576,7.311678,6.1967063,5.081734,3.966762,2.8517902,1.7368182,1.4122978,1.0877775,0.76325727,0.43692398,0.11240368,0.09064813,0.06707962,0.045324065,0.02175555,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.07977036,0.13415924,0.19036107,0.24474995,0.2991388,0.27919623,0.25925365,0.23931105,0.21936847,0.19942589,0.5094425,0.8194591,1.1294757,1.4394923,1.7495089,2.5925364,3.435564,4.2767787,5.1198063,5.962834,6.9001355,7.837437,8.774739,9.712041,10.649343,12.083396,13.515636,14.947877,16.380117,17.812357,20.377699,22.94304,25.508383,28.071913,30.637255,32.221783,33.808125,35.392654,36.977184,38.561714,36.844837,35.127964,33.409275,31.692398,29.975523,29.092611,28.209698,27.326784,26.445684,25.562773,24.685299,23.807825,22.930351,22.052877,21.175404,19.948027,18.720652,17.493277,16.2659,15.036712,12.964496,10.89228,8.820063,6.7478466,4.6756306,5.3083544,5.9392653,6.5719895,7.2047133,7.837437,7.494787,7.1521373,6.8094873,6.4668374,6.1241875,6.14413,6.165886,6.185828,6.205771,6.2257137,7.360628,8.495543,9.630457,10.765372,11.900287,11.407161,10.915848,10.422722,9.929596,9.438283,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.052575916,0.10515183,0.15772775,0.21030366,0.26287958,0.38434806,0.5076295,0.629098,0.7523795,0.87566096,0.9499924,1.0243238,1.1004683,1.1747998,1.2491312,1.6824293,2.1157274,2.5472124,2.9805105,3.4119956,3.1672456,2.9224956,2.6777458,2.4329958,2.1882458,2.8372865,3.48814,4.137181,4.788034,5.4370747,5.2630305,5.087173,4.9131284,4.7372713,4.5632267,3.7546456,2.9478772,2.1392958,1.3325275,0.52575916,0.57833505,0.629098,0.68167394,0.73424983,0.7868258,0.7016165,0.61822027,0.533011,0.44780177,0.36259252,0.29007402,0.21755551,0.14503701,0.072518505,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.014503701,0.018129626,0.01994259,0.02175555,0.025381476,0.12509441,0.22480737,0.3245203,0.42423326,0.52575916,1.5228885,2.520018,3.5171473,4.514277,5.5132194,4.9076896,4.3021603,3.6966307,3.092914,2.4873846,3.1853752,3.881553,4.5795436,5.277534,5.975525,6.782293,7.5890613,8.397643,9.2044115,10.012992,9.30775,8.602508,7.897265,7.192023,6.48678,6.002719,5.516845,5.032784,4.5469103,4.062849,4.6375585,5.2122674,5.7869763,6.3616858,6.9382076,6.2220874,5.5077806,4.7916603,4.077353,3.3630457,2.72307,2.0830941,1.4431182,0.8031424,0.16316663,0.13415924,0.10696479,0.07977036,0.052575916,0.025381476,0.047137026,0.07070554,0.092461094,0.11421664,0.13778515,0.13234627,0.12690738,0.12328146,0.11784257,0.11240368,0.092461094,0.072518505,0.052575916,0.032633327,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.9119202,1.8002719,2.6868105,3.5751622,4.461701,4.0320287,3.6023567,3.1726844,2.7430124,2.3133402,2.4873846,2.663242,2.8372865,3.0131438,3.1871881,4.0918565,4.9983377,5.903006,6.8076744,7.7123427,6.548421,5.382686,4.216951,3.053029,1.887294,1.7821422,1.6769904,1.5718386,1.4666867,1.3633479,1.452183,1.5428312,1.6316663,1.7223145,1.8129625,2.2897718,2.7683938,3.245203,3.7220123,4.2006345,4.7354584,5.2702823,5.805106,6.33993,6.874754,8.31062,9.744674,11.18054,12.6145935,14.05046,13.212872,12.375282,11.537694,10.700105,9.862516,11.989121,14.117539,16.245958,18.372562,20.499168,17.580297,14.6596155,11.740746,8.820063,5.89938,4.953014,4.004834,3.056655,2.1102884,1.162109,1.1167849,1.0732739,1.0279498,0.9826257,0.93730164,0.78319985,0.62728506,0.47318324,0.31726846,0.16316663,0.15047589,0.13778515,0.12509441,0.11240368,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03988518,0.07977036,0.11965553,0.15954071,0.19942589,0.21030366,0.21936847,0.23024625,0.23931105,0.25018883,0.20486477,0.15954071,0.11421664,0.07070554,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0870222,0.17585737,0.26287958,0.34990177,0.43692398,0.34990177,0.26287958,0.17585737,0.0870222,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.13959812,0.13053331,0.11965553,0.11059072,0.099712946,0.0870222,0.07433146,0.06164073,0.05076295,0.038072214,1.3325275,2.6269827,3.923251,5.217706,6.5121617,5.8921285,5.272095,4.652062,4.0320287,3.4119956,3.1146698,2.817344,2.520018,2.222692,1.9253663,1.54827,1.1693609,0.79226464,0.41516843,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.43511102,0.87022203,1.305333,1.7404441,2.175555,2.6849976,3.1944401,3.7056956,4.215138,4.7245803,6.4704633,8.214534,9.960417,11.704487,13.45037,15.5606575,17.669134,19.77942,21.88971,23.999998,20.885328,17.770658,14.654177,11.539507,8.424837,11.385405,14.34416,17.304728,20.265295,23.225864,23.91479,24.605528,25.294455,25.985193,26.675932,22.339325,18.004532,13.669738,9.334945,5.0001507,4.454449,3.9105604,3.3648586,2.819157,2.275268,1.8492218,1.4249886,1.0007553,0.5747091,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.03988518,0.06707962,0.09427405,0.12328146,0.15047589,0.13959812,0.13053331,0.11965553,0.11059072,0.099712946,0.31726846,0.53482395,0.7523795,0.969935,1.1874905,2.0142014,2.8427253,3.6694362,4.49796,5.3246713,5.7380266,6.149569,6.5629244,6.9744673,7.3878226,8.185526,8.98323,9.77912,10.576823,11.374527,14.0323305,16.690134,19.347937,22.003927,24.66173,27.355793,30.048042,32.74029,35.43254,38.12479,36.959057,35.79513,34.6294,33.465477,32.29974,31.427706,30.555672,29.681824,28.809788,27.937754,26.692247,25.446743,24.20305,22.957544,21.71204,19.980661,18.247469,16.514277,14.782897,13.049705,11.570327,10.089137,8.609759,7.130382,5.6491914,5.9718986,6.294606,6.6173134,6.9400206,7.262728,6.885632,6.506723,6.1296263,5.75253,5.375434,5.0980506,4.8206677,4.5432844,4.264088,3.9867048,4.954827,5.922949,6.889258,7.85738,8.825501,8.334189,7.844689,7.3551893,6.8656893,6.3743763,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06164073,0.12509441,0.18673515,0.25018883,0.31182957,0.42423326,0.53663695,0.6508536,0.76325727,0.87566096,0.89922947,0.9246109,0.9499924,0.97537386,1.0007553,1.649796,2.3006494,2.94969,3.6005437,4.249584,3.8380418,3.4246864,3.0131438,2.5997884,2.1882458,2.9007401,3.6132345,4.325729,5.038223,5.750717,5.6491914,5.5494785,5.4497657,5.3500524,5.2503395,4.3003473,3.350355,2.4003625,1.4503701,0.50037766,0.53663695,0.5747091,0.61278135,0.6508536,0.6871128,0.5620184,0.43692398,0.31182957,0.18673515,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.6871128,1.2491312,1.8129625,2.374981,2.9369993,2.5000753,2.0631514,1.6244144,1.1874905,0.7505665,1.5120108,2.275268,3.0367124,3.7999697,4.5632267,5.462456,6.3616858,7.262728,8.161958,9.063,8.713099,8.363196,8.013294,7.663393,7.311678,6.7623506,6.2130227,5.661882,5.1125546,4.5632267,5.2865987,6.011784,6.736969,7.462154,8.187339,7.362441,6.5375433,5.712645,4.8877473,4.062849,3.2869012,2.5127661,1.7368182,0.96268314,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.7505665,1.49932,2.2498865,3.000453,3.7492065,3.5117085,3.2742105,3.0367124,2.7992141,2.561716,2.762955,2.962381,3.1618068,3.3630457,3.5624714,4.7753434,5.9882154,7.1992745,8.412147,9.625018,8.125698,6.624565,5.125245,3.6241121,2.124792,1.987007,1.8492218,1.7132497,1.5754645,1.4376793,1.5120108,1.5881553,1.6624867,1.7368182,1.8129625,2.5000753,3.1871881,3.874301,4.5632267,5.2503395,5.8504305,6.450521,7.0506115,7.650702,8.2507925,10.049252,11.849524,13.649796,15.4500675,17.25034,16.187943,15.125546,14.06315,13.000754,11.938358,14.150173,16.361988,18.575615,20.78743,22.999243,19.725033,16.450823,13.174799,9.900589,6.624565,5.2992897,3.975827,2.6505513,1.3252757,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,0.26287958,0.2755703,0.28826106,0.2991388,0.31182957,0.25018883,0.18673515,0.12509441,0.06164073,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.52575916,1.0497054,1.5754645,2.0994108,2.6251698,2.2371957,1.8492218,1.4630609,1.0750868,0.6871128,0.5620184,0.43692398,0.31182957,0.18673515,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.26287958,0.52575916,0.7868258,1.0497054,1.3125849,3.7129474,6.11331,8.511859,10.912222,13.312584,15.674874,18.037165,20.399454,22.761745,25.125849,21.537996,17.950142,14.362289,10.774437,7.1883965,11.287505,15.386614,19.487535,23.588457,27.687565,28.575916,29.462456,30.350807,31.237345,32.125698,26.237194,20.350506,14.462003,8.575313,2.6868105,2.712192,2.7375734,2.762955,2.7883365,2.811905,2.2879589,1.7621996,1.2382535,0.7124943,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.12509441,0.25018883,0.37528324,0.50037766,0.62547207,1.4376793,2.2498865,3.0620937,3.874301,4.688321,4.574105,4.461701,4.349297,4.2368937,4.12449,4.2876563,4.4508233,4.612177,4.7753434,4.936697,7.686961,10.437225,13.1874895,15.937754,18.688019,22.487988,26.287958,30.087927,33.887897,37.687866,37.075085,36.462303,35.84952,35.23674,34.62577,33.762802,32.899834,32.03686,31.175705,30.312735,28.699198,27.087475,25.47575,23.862213,22.25049,20.01148,17.774284,15.537089,13.299893,11.062697,10.174346,9.287807,8.399456,7.512917,6.624565,6.637256,6.6499467,6.6626377,6.6753283,6.688019,6.2746634,5.863121,5.4497657,5.038223,4.6248674,4.0501585,3.4754493,2.9007401,2.324218,1.7495089,2.5508385,3.350355,4.1498713,4.949388,5.750717,5.2630305,4.7753434,4.2876563,3.7999697,3.3122826,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,0.34264994,0.43511102,0.5275721,0.6200332,0.7124943,0.73787576,0.76325727,0.7868258,0.8122072,0.8375887,1.3669738,1.8981718,2.427557,2.956942,3.48814,3.3068438,3.1273603,2.9478772,2.7683938,2.5870976,3.0276475,3.4681973,3.9069343,4.347484,4.788034,4.670192,4.552349,4.4345064,4.3166637,4.2006345,3.43919,2.6795588,1.9199274,1.1602961,0.40066472,0.4405499,0.48043507,0.52032024,0.56020546,0.6000906,0.4949388,0.38978696,0.28463513,0.1794833,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.5493277,1.0007553,1.4503701,1.8999848,2.3495996,1.9996977,1.649796,1.2998942,0.9499924,0.6000906,1.209246,1.8202144,2.42937,3.0403383,3.6494937,4.3946214,5.139749,5.8848767,6.630004,7.3751316,7.5455503,7.7141557,7.8845744,8.054993,8.225411,8.517298,8.809185,9.102885,9.394773,9.688472,9.683033,9.677594,9.672155,9.666717,9.663091,8.517298,7.3733187,6.2275267,5.081734,3.9377546,3.1853752,2.4329958,1.6806163,0.92823684,0.17585737,0.13959812,0.10515183,0.07070554,0.034446288,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.36440548,0.7306239,1.0950294,1.4594349,1.8256533,1.4721256,1.1204109,0.7668832,0.41516843,0.06164073,1.2328146,2.4021754,3.5733492,4.74271,5.9120708,5.18326,4.4526362,3.7220123,2.9932013,2.2625773,2.4076142,2.5526514,2.6976883,2.8427253,2.9877625,3.9341288,4.882308,5.8304877,6.776854,7.7250338,6.733343,5.7398396,4.748149,3.7546456,2.762955,2.9170568,3.0729716,3.2270734,3.3829882,3.53709,3.2796493,3.0222087,2.764768,2.5073273,2.2498865,3.2723975,4.2949085,5.317419,6.33993,7.362441,7.3841968,7.407765,7.4295206,7.453089,7.474845,9.775495,12.07433,14.37498,16.67563,18.974466,17.420757,15.865235,14.309713,12.754191,11.200482,12.639976,14.079468,15.520773,16.960264,18.399757,15.780026,13.1602955,10.540565,7.9190207,5.2992897,4.2477713,3.1944401,2.1429217,1.0895905,0.038072214,0.032633327,0.027194439,0.02175555,0.018129626,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03988518,0.07977036,0.11965553,0.15954071,0.19942589,0.21030366,0.21936847,0.23024625,0.23931105,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.42060733,0.83940166,1.260009,1.6806163,2.0994108,1.789394,1.4793775,1.1693609,0.85934424,0.5493277,0.44961473,0.34990177,0.25018883,0.15047589,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.21030366,0.42060733,0.629098,0.83940166,1.0497054,2.9823234,4.914942,6.8475595,8.780178,10.712796,12.650853,14.587097,16.525154,18.463211,20.399454,17.772472,15.14549,12.516694,9.88971,7.262728,12.217555,17.172382,22.127209,27.082035,32.03686,31.106812,30.176762,29.246712,28.316662,27.386612,22.34295,17.297476,12.252001,7.208339,2.1628644,2.179181,2.1973107,2.2154403,2.231757,2.2498865,1.8292793,1.4104849,0.9898776,0.56927025,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.21936847,0.42785916,0.6345369,0.8430276,1.0497054,1.7223145,2.3949237,3.0675328,3.7401419,4.4127507,4.401873,4.3928084,4.3819304,4.3728657,4.361988,4.41819,4.4725785,4.5269675,4.5831695,4.6375585,6.9146395,9.193533,11.470614,13.747695,16.024776,19.230095,22.435411,25.64073,28.844234,32.049553,31.915394,31.77942,31.645262,31.509289,31.37513,31.039732,30.704334,30.370749,30.03535,29.699953,28.372864,27.043962,25.716875,24.389786,23.062696,21.050308,19.03792,17.025532,15.013144,13.000754,12.284635,11.570327,10.854207,10.139899,9.425592,9.164526,8.9052725,8.644206,8.384952,8.125698,7.8845744,7.645263,7.404139,7.1648283,6.925517,6.548421,6.169512,5.7924156,5.4153194,5.038223,5.433449,5.826862,6.2220874,6.6173134,7.0125394,6.156821,5.3029156,4.4471974,3.5932918,2.7375734,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.25925365,0.33177215,0.40429065,0.47680917,0.5493277,0.5747091,0.6000906,0.62547207,0.6508536,0.6744221,1.0841516,1.4956942,1.9054236,2.3151531,2.7248828,2.7774587,2.8300345,2.8826106,2.9351864,2.9877625,3.1545548,3.3231604,3.489953,3.6567454,3.825351,3.6893787,3.5552197,3.4192474,3.2850883,3.149116,2.5798457,2.0105755,1.4394923,0.87022203,0.2991388,0.34264994,0.38434806,0.42785916,0.46955732,0.51306844,0.42785916,0.34264994,0.2574407,0.17223145,0.0870222,0.07070554,0.052575916,0.034446288,0.018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.41335547,0.7505665,1.0877775,1.4249886,1.7621996,1.49932,1.2382535,0.97537386,0.7124943,0.44961473,0.90829426,1.3651608,1.8220274,2.280707,2.7375734,3.3267863,3.917812,4.507025,5.0980506,5.6872635,6.378002,7.066928,7.757667,8.448405,9.137331,10.272246,11.407161,12.542075,13.67699,14.811904,14.077655,13.343405,12.607342,11.873092,11.137029,9.672155,8.207282,6.742408,5.277534,3.8126602,3.0820365,2.3532255,1.6226015,0.8919776,0.16316663,0.13053331,0.09789998,0.065266654,0.032633327,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.7306239,1.4594349,2.1900587,2.9206827,3.6494937,2.9442513,2.2408218,1.5355793,0.83033687,0.12509441,1.7150626,3.3050308,4.894999,6.484967,8.074935,6.8529987,5.6292486,4.407312,3.1853752,1.9616255,2.0522738,2.1429217,2.231757,2.322405,2.4130533,3.094727,3.778214,4.459888,5.143375,5.825049,5.3391747,4.855114,4.36924,3.8851788,3.3993049,3.8471067,4.2949085,4.74271,5.1905117,5.638314,5.047288,4.458075,3.8670492,3.2778363,2.6868105,4.0447197,5.4026284,6.7605376,8.116633,9.474543,8.919776,8.365009,7.8102427,7.2554765,6.70071,9.499924,12.299138,15.100165,17.89938,20.700407,18.651758,16.604925,14.558089,12.509441,10.462607,11.129777,11.7969475,12.464118,13.1331005,13.800271,11.83502,9.869768,7.9045167,5.9392653,3.975827,3.1944401,2.4148662,1.6352923,0.8557183,0.07433146,0.065266654,0.054388877,0.045324065,0.034446288,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.15772775,0.16497959,0.17223145,0.1794833,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.3154555,0.629098,0.9445535,1.260009,1.5754645,1.3415923,1.1095331,0.8774739,0.64541465,0.41335547,0.33721104,0.26287958,0.18673515,0.11240368,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.15772775,0.3154555,0.47318324,0.629098,0.7868258,2.2516994,3.7165732,5.18326,6.6481338,8.113008,9.625018,11.137029,12.650853,14.162864,15.674874,14.006948,12.340837,10.672911,9.004985,7.3370595,13.147605,18.958149,24.766882,30.577427,36.387974,33.639523,30.892883,28.144432,25.397793,22.649342,18.446894,14.244447,10.042,5.8395524,1.6371052,1.647983,1.6570477,1.6679256,1.6769904,1.6878681,1.3724127,1.0569572,0.7433147,0.42785916,0.11240368,0.09064813,0.06707962,0.045324065,0.02175555,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.3154555,0.6055295,0.89560354,1.1856775,1.4757515,2.0069497,2.5399606,3.0729716,3.6041696,4.137181,4.229642,4.322103,4.4145637,4.507025,4.599486,4.5469103,4.494334,4.441758,4.3891826,4.3366065,6.1423173,7.948028,9.751925,11.557636,13.363347,15.9722,18.582867,21.19172,23.802385,26.413052,26.755701,27.098352,27.439188,27.78184,28.124489,28.316662,28.510649,28.702824,28.894999,29.087172,28.044718,27.002264,25.959812,24.917358,23.874905,22.087322,20.299742,18.512161,16.72458,14.936998,14.394923,13.852847,13.310771,12.766883,12.224807,11.691795,11.160598,10.627586,10.094576,9.563377,9.494485,9.427405,9.360326,9.293246,9.224354,9.04487,8.865387,8.685904,8.504607,8.325124,8.314246,8.3051815,8.294304,8.285239,8.274362,7.0524244,5.8304877,4.606738,3.3848011,2.1628644,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.17767033,0.23024625,0.28282216,0.33539808,0.387974,0.41335547,0.43692398,0.46230546,0.48768693,0.51306844,0.8031424,1.0932164,1.3832904,1.6733645,1.9616255,2.2480736,2.5327086,2.817344,3.101979,3.386614,3.2832751,3.1781235,3.0729716,2.9678197,2.8626678,2.7103791,2.5580902,2.4058013,2.2516994,2.0994108,1.7205015,1.3397794,0.96087015,0.58014804,0.19942589,0.24474995,0.29007402,0.33539808,0.38072214,0.42423326,0.36077955,0.2955129,0.23024625,0.16497959,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.2755703,0.50037766,0.72518504,0.9499924,1.1747998,1.0007553,0.824898,0.6508536,0.4749962,0.2991388,0.6055295,0.9101072,1.214685,1.5192627,1.8256533,2.2607644,2.6958754,3.1291735,3.5642843,3.9993954,5.2104545,6.4197006,7.6307597,8.840006,10.049252,12.027194,14.005136,15.983078,17.959208,19.93715,18.472277,17.007402,15.542528,14.077655,12.612781,10.827013,9.043057,7.2572894,5.473334,3.6875658,2.9805105,2.2716422,1.5645868,0.8575313,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.0950294,2.1900587,3.2850883,4.3801174,5.475147,4.41819,3.3594196,2.3024626,1.2455053,0.18673515,2.1973107,4.207886,6.2166486,8.227224,10.2378,8.5227375,6.8076744,5.092612,3.3775494,1.6624867,1.696933,1.7331922,1.7676386,1.8020848,1.8383441,2.2553256,2.6723068,3.0892882,3.5080826,3.925064,3.9468195,3.9703882,3.9921436,4.0157123,4.0374675,4.7771564,5.516845,6.258347,6.9980354,7.7377243,6.814926,5.8921285,4.9693303,4.0483456,3.1255474,4.8170414,6.510349,8.201842,9.89515,11.586644,10.455356,9.322253,8.189152,7.057863,5.924762,9.224354,12.525759,15.825351,19.124943,22.424534,19.884573,17.344612,14.804652,12.264692,9.724731,9.619579,9.514427,9.409276,9.304124,9.200785,7.890013,6.5792413,5.2702823,3.9595103,2.6505513,2.1429217,1.6352923,1.1276628,0.6200332,0.11240368,0.09789998,0.08339628,0.06707962,0.052575916,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.10515183,0.11059072,0.11421664,0.11965553,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.21030366,0.42060733,0.630911,0.83940166,1.0497054,0.89560354,0.73968875,0.5855869,0.42967212,0.2755703,0.22480737,0.17585737,0.12509441,0.07433146,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.10515183,0.21030366,0.3154555,0.42060733,0.52575916,1.5228885,2.520018,3.5171473,4.514277,5.5132194,6.599184,7.686961,8.774739,9.862516,10.950294,10.243238,9.53437,8.827314,8.120259,7.413204,14.077655,20.742105,27.40837,34.07282,40.73727,36.17223,31.60719,27.04215,22.47711,17.912071,14.55265,11.193231,7.8319983,4.4725785,1.1131591,1.114972,1.1167849,1.1204109,1.1222239,1.1258497,0.9155461,0.70524246,0.4949388,0.28463513,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.40972954,0.78319985,1.1548572,1.5283275,1.8999848,2.2933977,2.6849976,3.0784104,3.4700103,3.8616104,4.0574102,4.25321,4.4471974,4.6429973,4.836984,4.6774435,4.517903,4.358362,4.1970086,4.0374675,5.369995,6.7025228,8.03505,9.367578,10.700105,12.714307,14.730321,16.744522,18.760536,20.774738,21.594198,22.41547,23.234928,24.054388,24.87566,25.595406,26.315151,27.034899,27.754644,28.47439,27.716572,26.960567,26.202747,25.44493,24.68711,23.124338,21.561563,20.000603,18.43783,16.875055,16.50521,16.135366,15.765523,15.3956785,15.025834,14.219066,13.41411,12.609155,11.804199,10.999244,11.104396,11.209548,11.314699,11.419851,11.525003,11.543133,11.559449,11.5775795,11.595709,11.612025,11.1968565,10.781689,10.368333,9.953164,9.537996,7.948028,6.35806,4.7680917,3.1781235,1.5881553,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.09427405,0.12690738,0.15954071,0.19217403,0.22480737,0.25018883,0.2755703,0.2991388,0.3245203,0.34990177,0.52032024,0.69073874,0.85934424,1.0297627,1.2001812,1.7168756,2.2353828,2.752077,3.2705846,3.787279,3.4101827,3.0330863,2.6541772,2.277081,1.8999848,1.7295663,1.5591478,1.3905423,1.2201238,1.0497054,0.85934424,0.67079616,0.48043507,0.29007402,0.099712946,0.14684997,0.19579996,0.24293698,0.29007402,0.33721104,0.291887,0.24837588,0.2030518,0.15772775,0.11240368,0.09064813,0.06707962,0.045324065,0.02175555,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.13778515,0.25018883,0.36259252,0.4749962,0.5873999,0.50037766,0.41335547,0.3245203,0.2374981,0.15047589,0.30276474,0.4550536,0.6073425,0.75963134,0.9119202,1.1929294,1.4721256,1.7531348,2.032331,2.3133402,4.0429068,5.772473,7.502039,9.233418,10.962985,13.782142,16.603111,19.422268,22.243238,25.062395,22.866898,20.673212,18.477715,16.282217,14.0867195,11.98187,9.87702,7.7721705,5.667321,3.5624714,2.8771715,2.1918716,1.5065719,0.823085,0.13778515,0.11059072,0.08339628,0.054388877,0.027194439,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.4594349,2.9206827,4.3801174,5.8395524,7.3008003,5.8903155,4.4798307,3.0693457,1.6606737,0.25018883,2.6795588,5.1107416,7.5401115,9.969481,12.400664,10.192475,7.9842873,5.7779117,3.5697234,1.3633479,1.3415923,1.3216497,1.3017071,1.2817645,1.261822,1.4141108,1.5682126,1.7205015,1.8727903,2.0250793,2.5544643,3.0856624,3.6150475,4.1444325,4.6756306,5.7072062,6.740595,7.7721705,8.805559,9.837135,8.582565,7.327995,6.071612,4.8170414,3.5624714,5.5893636,7.6180687,9.644961,11.671853,13.700559,11.990934,10.279498,8.569874,6.8602505,5.1506267,8.950596,12.750566,16.550535,20.350506,24.150475,21.117388,18.084301,15.053028,12.019942,8.9868555,8.109382,7.231908,6.354434,5.47696,4.599486,3.9450066,3.290527,2.6342347,1.9797552,1.3252757,1.0895905,0.8557183,0.6200332,0.38434806,0.15047589,0.13053331,0.11059072,0.09064813,0.07070554,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.052575916,0.054388877,0.058014803,0.059827764,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.10515183,0.21030366,0.3154555,0.42060733,0.52575916,0.44780177,0.36984438,0.291887,0.21574254,0.13778515,0.11240368,0.0870222,0.06164073,0.038072214,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.052575916,0.10515183,0.15772775,0.21030366,0.26287958,0.79226464,1.3216497,1.8528478,2.382233,2.911618,3.5751622,4.2368937,4.900438,5.562169,6.2257137,6.4777155,6.7297173,6.981719,7.2355337,7.4875355,15.007704,22.527874,30.048042,37.56821,45.08838,38.704937,32.32331,25.939869,19.55824,13.174799,10.656594,8.140202,5.621997,3.105605,0.5873999,0.581961,0.57833505,0.5728962,0.56745726,0.5620184,0.45686656,0.35171473,0.24837588,0.14322405,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.5058166,0.96087015,1.4159238,1.8691645,2.324218,2.5780327,2.8300345,3.0820365,3.3358512,3.587853,3.8851788,4.1825047,4.4798307,4.7771564,5.0744824,4.8079767,4.539658,4.273153,4.004834,3.738329,4.597673,5.4570174,6.3181744,7.177519,8.036863,9.458226,10.877775,12.297325,13.716875,15.138238,16.434505,17.732588,19.030668,20.326937,21.625017,22.872335,24.119654,25.366972,26.61429,27.861609,27.390238,26.917055,26.445684,25.972502,25.49932,24.163166,22.8252,21.487232,20.149265,18.813112,18.6155,18.417887,18.220274,18.022661,17.825048,16.748148,15.6694355,14.592536,13.515636,12.436923,12.714307,12.99169,13.270886,13.548269,13.825653,14.039582,14.255324,14.4692545,14.684997,14.90074,14.079468,13.260008,12.440549,11.619277,10.799818,8.841819,6.885632,4.9276323,2.9696326,1.0116332,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.0870222,0.11240368,0.13778515,0.16316663,0.18673515,0.2374981,0.28826106,0.33721104,0.387974,0.43692398,1.1874905,1.938057,2.6868105,3.437377,4.1879435,3.53709,2.8880494,2.2371957,1.5881553,0.93730164,0.7505665,0.5620184,0.37528324,0.18673515,0.0,0.0,0.0,0.0,0.0,0.0,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,0.22480737,0.19942589,0.17585737,0.15047589,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.12509441,0.25018883,0.37528324,0.50037766,0.62547207,2.8753586,5.125245,7.3751316,9.625018,11.874905,15.537089,19.199274,22.863272,26.525455,30.18764,27.26333,24.33721,21.4129,18.48678,15.56247,13.136727,10.712796,8.287052,5.863121,3.437377,2.7756457,2.1121013,1.4503701,0.7868258,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.8256533,3.6494937,5.475147,7.3008003,9.12464,7.362441,5.600241,3.8380418,2.0758421,0.31182957,3.1618068,6.011784,8.861761,11.711739,14.561715,11.862214,9.162713,6.4632115,3.7618973,1.062396,0.9880646,0.9119202,0.8375887,0.76325727,0.6871128,0.5747091,0.46230546,0.34990177,0.2374981,0.12509441,1.162109,2.1991236,3.2379513,4.274966,5.3119802,6.637256,7.9625316,9.287807,10.613083,11.938358,10.3502035,8.762048,7.175706,5.5875506,3.9993954,6.3616858,8.725789,11.088079,13.45037,15.812659,13.524701,11.236742,8.950596,6.6626377,4.3746786,8.675026,12.975373,17.27572,21.574255,25.874601,22.350203,18.825804,15.299591,11.775192,8.2507925,6.599184,4.949388,3.299592,1.649796,0.0,0.0,0.0,0.0,0.0,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.16316663,0.13778515,0.11240368,0.0870222,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06164073,0.12509441,0.18673515,0.25018883,0.31182957,0.5493277,0.7868258,1.0243238,1.261822,1.49932,2.712192,3.925064,5.137936,6.350808,7.5618668,15.937754,24.311829,32.687714,41.06179,49.437675,41.237648,33.037617,24.837587,16.637558,8.437528,6.7623506,5.087173,3.4119956,1.7368182,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.6000906,1.1367276,1.6751775,2.2118144,2.7502642,2.8626678,2.9750717,3.0874753,3.199879,3.3122826,3.7129474,4.1117992,4.512464,4.9131284,5.3119802,4.936697,4.5632267,4.1879435,3.8126602,3.437377,3.825351,4.213325,4.599486,4.98746,5.375434,6.200332,7.02523,7.850128,8.675026,9.499924,11.274815,13.049705,14.824595,16.599485,18.374376,20.149265,21.92597,23.70086,25.47575,27.25064,27.062092,26.875357,26.68681,26.500074,26.31334,25.20018,24.08702,22.975676,21.862516,20.749357,20.725788,20.700407,20.675026,20.649643,20.624262,19.275417,17.92476,16.574104,15.22526,13.874602,14.324218,14.775645,15.22526,15.674874,16.124489,16.537846,16.949387,17.362743,17.774284,18.187641,16.962078,15.736515,14.512766,13.287203,12.06164,9.737422,7.4113913,5.087173,2.762955,0.43692398,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.018129626,0.034446288,0.052575916,0.07070554,0.0870222,0.10333887,0.11784257,0.13234627,0.14684997,0.16316663,0.2030518,0.24293698,0.28282216,0.32270733,0.36259252,1.2455053,2.126605,3.009518,3.8924308,4.7753434,4.071914,3.3702974,2.666868,1.9652514,1.261822,1.0098201,0.75781834,0.5058166,0.2520018,0.0,0.0,0.0,0.0,0.0,0.0,0.04169814,0.08520924,0.12690738,0.17041849,0.21211663,0.19217403,0.17223145,0.15228885,0.13234627,0.11240368,0.092461094,0.072518505,0.052575916,0.032633327,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.099712946,0.19942589,0.2991388,0.40066472,0.50037766,2.3006494,4.099108,5.89938,7.699652,9.499924,12.429671,15.359419,18.289167,21.220728,24.150475,22.06738,19.984287,17.903006,15.819912,13.736817,11.651911,9.567003,7.4820967,5.3971896,3.3122826,2.6849976,2.0577126,1.4304274,0.8031424,0.17585737,0.16316663,0.15047589,0.13778515,0.12509441,0.11240368,0.10696479,0.10333887,0.09789998,0.092461094,0.0870222,0.15410182,0.2229944,0.29007402,0.35715362,0.42423326,0.34264994,0.25925365,0.17767033,0.09427405,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.2374981,0.4749962,0.7124943,0.9499924,1.1874905,2.4094272,3.633177,4.855114,6.0770507,7.3008003,5.8921285,4.4852695,3.0765975,1.6697385,0.26287958,2.5526514,4.842423,7.132195,9.421967,11.711739,9.539809,7.36788,5.1941376,3.0222087,0.85027945,0.79770356,0.7451276,0.69255173,0.6399758,0.5873999,0.968122,1.3470312,1.7277533,2.1066625,2.4873846,2.956942,3.4283123,3.8978696,4.367427,4.836984,5.9700856,7.1031876,8.234476,9.367578,10.500679,9.420154,8.339628,7.2591023,6.1803894,5.0998635,6.6100616,8.120259,9.630457,11.1406555,12.64904,10.859646,9.070251,7.2790446,5.4896507,3.7002566,7.0995617,10.500679,13.899984,17.29929,20.700407,17.879436,15.06028,12.23931,9.420154,6.599184,5.279347,3.9595103,2.6396735,1.3198367,0.0,0.0,0.0,0.0,0.0,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.13053331,0.11059072,0.09064813,0.07070554,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.018129626,0.034446288,0.052575916,0.07070554,0.0870222,0.2520018,0.4169814,0.581961,0.7469406,0.9119202,1.1331016,1.35247,1.5718386,1.79302,2.0123885,3.2578938,4.501586,5.7470913,6.9925966,8.238102,14.612478,20.986855,27.363045,33.73742,40.111797,33.44372,26.777458,20.10938,13.443117,6.775041,5.429823,4.0846047,2.7393866,1.3941683,0.05076295,0.04169814,0.034446288,0.027194439,0.01994259,0.012690738,0.09789998,0.18310922,0.26831847,0.35171473,0.43692398,0.39703882,0.35715362,0.31726846,0.27738327,0.2374981,0.19036107,0.14322405,0.09427405,0.047137026,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.072518505,0.14503701,0.21755551,0.29007402,0.36259252,0.8974165,1.4322405,1.9670644,2.5018883,3.0367124,3.1781235,3.3177216,3.4573197,3.5969179,3.738329,3.8543584,3.972201,4.0900435,4.207886,4.325729,4.07554,3.825351,3.5751622,3.3249733,3.0747845,3.4319382,3.7909048,4.1480584,4.505212,4.8623657,5.431636,6.002719,6.5719895,7.1430726,7.7123427,9.334945,10.957546,12.580148,14.202749,15.825351,17.364555,18.905573,20.444778,21.983984,23.525002,23.472427,23.419851,23.367275,23.3147,23.262123,22.31757,21.373016,20.42665,19.482096,18.537542,18.709774,18.882006,19.054237,19.228281,19.400513,18.457771,17.515032,16.57229,15.62955,14.68681,14.955129,15.223447,15.489952,15.758271,16.024776,16.708263,17.389936,18.073423,18.755098,19.436771,17.870373,16.30216,14.73576,13.167547,11.599335,10.274059,8.950596,7.6253204,6.300045,4.974769,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.11784257,0.12328146,0.12690738,0.13234627,0.13778515,0.16679256,0.19761293,0.22662032,0.2574407,0.28826106,1.3017071,2.3169663,3.3322253,4.347484,5.3627434,4.606738,3.8525455,3.0983531,2.3423476,1.5881553,1.2708868,0.95180535,0.6345369,0.31726846,0.0,0.0,0.0,0.0,0.0,0.0,0.034446288,0.07070554,0.10515183,0.13959812,0.17585737,0.15954071,0.14503701,0.13053331,0.11421664,0.099712946,0.08520924,0.07070554,0.054388877,0.03988518,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07433146,0.15047589,0.22480737,0.2991388,0.37528324,1.7241274,3.0747845,4.4254417,5.774286,7.124943,9.322253,11.519565,13.716875,15.914186,18.11331,16.873243,15.633177,14.39311,13.153044,11.912977,10.167094,8.423024,6.677141,4.933071,3.1871881,2.5943494,2.0033236,1.4104849,0.81764615,0.22480737,0.22480737,0.22480737,0.22480737,0.22480737,0.22480737,0.21574254,0.20486477,0.19579996,0.18492219,0.17585737,0.3100166,0.44417584,0.58014804,0.71430725,0.85027945,0.6852999,0.52032024,0.35534066,0.19036107,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.4749962,0.9499924,1.4249886,1.8999848,2.374981,2.9950142,3.6150475,4.2350807,4.855114,5.475147,4.421816,3.3702974,2.3169663,1.2654479,0.21211663,1.9416829,3.673062,5.4026284,7.132195,8.861761,7.217404,5.573047,3.926877,2.2825198,0.63816285,0.6073425,0.57833505,0.5475147,0.5166943,0.48768693,1.3597219,2.231757,3.105605,3.97764,4.8496747,4.751775,4.655688,4.557788,4.459888,4.361988,5.3029156,6.24203,7.1829576,8.122072,9.063,8.490104,7.9172077,7.344311,6.773228,6.200332,6.8566246,7.51473,8.172835,8.829127,9.487233,8.194591,6.9019485,5.6093063,4.3166637,3.0258346,5.524097,8.024173,10.524248,13.024323,15.524399,13.410484,11.294757,9.179029,7.065115,4.949388,3.9595103,2.9696326,1.9797552,0.9898776,0.0,0.0,0.0,0.0,0.0,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.09789998,0.08339628,0.06707962,0.052575916,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.034446288,0.07070554,0.10515183,0.13959812,0.17585737,0.44236287,0.7106813,0.97718686,1.2455053,1.5120108,1.7150626,1.9181144,2.1193533,2.322405,2.525457,3.8017826,5.0799212,6.35806,7.6343856,8.912524,13.287203,17.661882,22.038374,26.413052,30.787731,25.651608,20.517298,15.382988,10.246864,5.1125546,4.0972953,3.0820365,2.0667772,1.0533313,0.038072214,0.034446288,0.032633327,0.030820364,0.027194439,0.025381476,0.19579996,0.36440548,0.53482395,0.70524246,0.87566096,0.79589057,0.71430725,0.6345369,0.55476654,0.4749962,0.38072214,0.28463513,0.19036107,0.09427405,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13234627,0.26469254,0.39703882,0.5293851,0.66173136,1.1947423,1.7277533,2.2607644,2.7919624,3.3249733,3.491766,3.6603715,3.827164,3.9957695,4.162562,3.9975824,3.832603,3.6676233,3.5026438,3.3376641,3.2125697,3.0874753,2.962381,2.8372865,2.712192,3.0403383,3.3666716,3.6948178,4.022964,4.349297,4.664753,4.9802084,5.295664,5.6093063,5.924762,7.3950744,8.865387,10.3357,11.804199,13.274512,14.579845,15.885179,17.190512,18.494032,19.799364,19.882761,19.964344,20.04774,20.129324,20.212719,19.43496,18.657198,17.879436,17.101677,16.325727,16.695572,17.065416,17.43526,17.805105,18.17495,17.640125,17.105303,16.570478,16.035654,15.50083,15.584227,15.6694355,15.754644,15.839854,15.925063,16.87687,17.830486,18.782291,19.734098,20.687716,18.776854,16.867804,14.956942,13.047892,11.137029,10.812509,10.487988,10.161655,9.837135,9.512614,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.027194439,0.054388877,0.08339628,0.11059072,0.13778515,0.13234627,0.12690738,0.12328146,0.11784257,0.11240368,0.13234627,0.15228885,0.17223145,0.19217403,0.21211663,1.3597219,2.5073273,3.6549325,4.802538,5.9501433,5.143375,4.3347936,3.5280252,2.7194438,1.9126755,1.5301404,1.1476053,0.7650702,0.3825351,0.0,0.0,0.0,0.0,0.0,0.0,0.027194439,0.054388877,0.08339628,0.11059072,0.13778515,0.12690738,0.11784257,0.10696479,0.09789998,0.0870222,0.07795739,0.06707962,0.058014803,0.047137026,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,1.1494182,2.0504606,2.94969,3.8507326,4.749962,6.2148356,7.6797094,9.144584,10.609457,12.07433,11.677292,11.280253,10.883214,10.484363,10.087324,8.682278,7.2772317,5.8721857,4.4671397,3.0620937,2.5055144,1.9471219,1.3905423,0.8321498,0.2755703,0.28826106,0.2991388,0.31182957,0.3245203,0.33721104,0.32270733,0.30820364,0.291887,0.27738327,0.26287958,0.46411842,0.6671702,0.87022203,1.0732739,1.2745126,1.0279498,0.7795739,0.533011,0.28463513,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.7124943,1.4249886,2.137483,2.8499773,3.5624714,3.5806012,3.5969179,3.6150475,3.633177,3.6494937,2.953316,2.2553256,1.5573349,0.85934424,0.16316663,1.3325275,2.5018883,3.673062,4.842423,6.011784,4.894999,3.778214,2.659616,1.5428312,0.42423326,0.4169814,0.40972954,0.40247768,0.39522585,0.387974,1.7531348,3.1182957,4.4816437,5.846804,7.211965,6.546608,5.883064,5.217706,4.552349,3.8869917,4.6357455,5.382686,6.1296263,6.87838,7.6253204,7.560054,7.494787,7.4295206,7.364254,7.3008003,7.1050005,6.9092,6.7152133,6.5194135,6.3254266,5.529536,4.7354584,3.9395678,3.1454902,2.3495996,3.9504454,5.5494785,7.1503243,8.749357,10.3502035,8.939718,7.5292335,6.1205616,4.710077,3.299592,2.6396735,1.9797552,1.3198367,0.65991837,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.065266654,0.054388877,0.045324065,0.034446288,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.052575916,0.10515183,0.15772775,0.21030366,0.26287958,0.6327239,1.0025684,1.3724127,1.742257,2.1121013,2.2970235,2.4819458,2.666868,2.8517902,3.0367124,4.347484,5.658256,6.967215,8.2779875,9.5869465,11.961927,14.336908,16.71189,19.08687,21.461851,17.859495,14.257137,10.654781,7.0524244,3.4500678,2.764768,2.079468,1.3941683,0.7106813,0.025381476,0.027194439,0.030820364,0.032633327,0.034446288,0.038072214,0.291887,0.5475147,0.8031424,1.0569572,1.3125849,1.1929294,1.0732739,0.95180535,0.8321498,0.7124943,0.56927025,0.42785916,0.28463513,0.14322405,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.19217403,0.38434806,0.57833505,0.7705091,0.96268314,1.4920682,2.0232663,2.5526514,3.0820365,3.6132345,3.8072214,4.0030212,4.1970086,4.3928084,4.5867953,4.1408067,3.6930048,3.245203,2.7974012,2.3495996,2.3495996,2.3495996,2.3495996,2.3495996,2.3495996,2.6469254,2.9442513,3.24339,3.540716,3.8380418,3.8978696,3.9576974,4.017525,4.077353,4.137181,5.4552045,6.773228,8.089439,9.407463,10.725487,11.795135,12.864782,13.93443,15.004078,16.075539,16.293095,16.51065,16.728207,16.94576,17.163317,16.55235,15.9431925,15.332225,14.723069,14.112101,14.679558,15.247015,15.814472,16.38193,16.949387,16.82248,16.695572,16.566853,16.439945,16.313038,16.215137,16.117237,16.019337,15.92325,15.825351,17.047287,18.271036,19.492973,20.71491,21.936848,19.685148,17.431635,15.179935,12.928236,10.674724,11.349146,12.025381,12.699803,13.374225,14.05046,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.032633327,0.065266654,0.09789998,0.13053331,0.16316663,0.14684997,0.13234627,0.11784257,0.10333887,0.0870222,0.09789998,0.10696479,0.11784257,0.12690738,0.13778515,1.4177368,2.6976883,3.97764,5.2575917,6.5375433,5.678199,4.8170414,3.9576974,3.0983531,2.2371957,1.789394,1.3434052,0.89560354,0.44780177,0.0,0.0,0.0,0.0,0.0,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.09427405,0.09064813,0.08520924,0.07977036,0.07433146,0.07070554,0.065266654,0.059827764,0.054388877,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.5747091,1.0243238,1.4757515,1.9253663,2.374981,3.1074178,3.8398547,4.572292,5.3047285,6.037165,6.4831543,6.92733,7.3733187,7.817495,8.26167,7.1974616,6.1332526,5.06723,4.0030212,2.9369993,2.4148662,1.892733,1.3705997,0.8466535,0.3245203,0.34990177,0.37528324,0.40066472,0.42423326,0.44961473,0.42967212,0.40972954,0.38978696,0.36984438,0.34990177,0.6200332,0.8901646,1.1602961,1.4304274,1.7005589,1.3705997,1.0406405,0.7106813,0.38072214,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.9499924,1.8999848,2.8499773,3.7999697,4.749962,4.164375,3.5806012,2.9950142,2.4094272,1.8256533,1.4830034,1.1403534,0.79770356,0.4550536,0.11240368,0.72337204,1.3325275,1.9416829,2.5526514,3.1618068,2.572594,1.983381,1.3923552,0.8031424,0.21211663,0.22662032,0.24293698,0.2574407,0.27194437,0.28826106,2.1447346,4.0030212,5.859495,7.7177815,9.574255,8.343254,7.1104393,5.8776245,4.64481,3.4119956,3.966762,4.5233417,5.0781083,5.632875,6.187641,6.630004,7.072367,7.51473,7.957093,8.399456,7.3533764,6.305484,5.2575917,4.209699,3.1618068,2.864481,2.5671551,2.269829,1.9725033,1.6751775,2.374981,3.0747845,3.774588,4.4743915,5.1741953,4.4707656,3.7655232,3.0602808,2.3550384,1.649796,1.3198367,0.9898776,0.65991837,0.32995918,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.032633327,0.027194439,0.02175555,0.018129626,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07070554,0.13959812,0.21030366,0.27919623,0.34990177,0.823085,1.2944553,1.7676386,2.2408218,2.712192,2.8807976,3.04759,3.2143826,3.3829882,3.5497808,4.893186,6.2347784,7.5781837,8.919776,10.263181,10.636651,11.011934,11.3872175,11.762501,12.137785,10.067381,7.996978,5.9265747,3.8579843,1.7875811,1.4322405,1.0768998,0.72337204,0.3680314,0.012690738,0.01994259,0.027194439,0.034446288,0.04169814,0.05076295,0.38978696,0.7306239,1.0696479,1.4104849,1.7495089,1.5899682,1.4304274,1.2708868,1.1095331,0.9499924,0.75963134,0.56927025,0.38072214,0.19036107,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.2520018,0.5058166,0.75781834,1.0098201,1.261822,1.789394,2.3169663,2.8445382,3.3721104,3.8996825,4.122677,4.345671,4.5668526,4.7898474,5.0128417,4.2822175,3.5534067,2.8227828,2.0921588,1.3633479,1.4866294,1.6117238,1.7368182,1.8619126,1.987007,2.2553256,2.521831,2.7901495,3.056655,3.3249733,3.1291735,2.9351864,2.7393866,2.5453994,2.3495996,3.5153344,4.6792564,5.844991,7.0107265,8.174648,9.010424,9.844387,10.680162,11.514126,12.349901,12.701616,13.055143,13.406858,13.760386,14.112101,13.669738,13.227375,12.785012,12.342649,11.900287,12.665357,13.430427,14.195497,14.960567,15.725637,16.004833,16.285843,16.565039,16.844234,17.125244,16.844234,16.565039,16.285843,16.004833,15.725637,17.217705,18.709774,20.201841,21.695723,23.187792,20.591629,17.99728,15.40293,12.806767,10.212419,11.887595,13.562773,15.23795,16.913128,18.588305,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.16316663,0.13778515,0.11240368,0.0870222,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,1.4757515,2.8880494,4.3003473,5.712645,7.124943,6.2130227,5.2992897,4.3873696,3.4754493,2.561716,2.0504606,1.5373923,1.0243238,0.51306844,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.2872034,2.5744069,3.8634233,5.1506267,6.43783,5.712645,4.98746,4.262275,3.53709,2.811905,2.324218,1.8383441,1.3506571,0.8629702,0.37528324,0.41335547,0.44961473,0.48768693,0.52575916,0.5620184,0.53663695,0.51306844,0.48768693,0.46230546,0.43692398,0.774135,1.1131591,1.4503701,1.7875811,2.124792,1.7132497,1.2998942,0.8883517,0.4749962,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.1874905,2.374981,3.5624714,4.749962,5.9374523,4.749962,3.5624714,2.374981,1.1874905,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.11240368,0.16316663,0.21211663,0.26287958,0.31182957,0.25018883,0.18673515,0.12509441,0.06164073,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,2.5381477,4.8877473,7.2373466,9.5869465,11.938358,10.138086,8.337815,6.5375433,4.7372713,2.9369993,3.299592,3.6621845,4.024777,4.3873696,4.749962,5.6999545,6.6499467,7.5999393,8.549932,9.499924,7.5999393,5.6999545,3.7999697,1.8999848,0.0,0.19942589,0.40066472,0.6000906,0.7995165,1.0007553,0.7995165,0.6000906,0.40066472,0.19942589,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0870222,0.17585737,0.26287958,0.34990177,0.43692398,1.0116332,1.5881553,2.1628644,2.7375734,3.3122826,3.4627585,3.6132345,3.7618973,3.9123733,4.062849,5.4370747,6.813113,8.187339,9.563377,10.937603,9.313189,7.686961,6.0625467,4.4381323,2.811905,2.275268,1.7368182,1.2001812,0.66173136,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.48768693,0.9119202,1.3379664,1.7621996,2.1882458,1.987007,1.7875811,1.5881553,1.3869164,1.1874905,0.9499924,0.7124943,0.4749962,0.2374981,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.31182957,0.62547207,0.93730164,1.2491312,1.5627737,2.08672,2.612479,3.1382382,3.6621845,4.1879435,4.4381323,4.688321,4.936697,5.186886,5.4370747,4.4254417,3.4119956,2.4003625,1.3869164,0.37528324,0.62547207,0.87566096,1.1258497,1.3742256,1.6244144,1.8619126,2.0994108,2.3369088,2.5744069,2.811905,2.3622901,1.9126755,1.4630609,1.0116332,0.5620184,1.5754645,2.5870976,3.6005437,4.612177,5.6256227,6.2257137,6.825804,7.4258947,8.024173,8.624263,9.11195,9.599637,10.087324,10.57501,11.062697,10.7871275,10.51337,10.2378,9.96223,9.686659,10.649343,11.612025,12.574709,13.537392,14.500074,15.187187,15.8743,16.563227,17.25034,17.937452,17.475147,17.01284,16.550535,16.08823,15.624111,17.388124,19.150324,20.912523,22.674723,24.436922,21.499924,18.562923,15.624111,12.687112,9.750113,12.426045,15.100165,17.774284,20.450218,23.124338,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.045324065,0.09064813,0.13415924,0.1794833,0.22480737,0.21030366,0.19579996,0.1794833,0.16497959,0.15047589,0.4405499,0.7306239,1.020698,1.310772,1.6008459,2.420305,3.2397642,4.059223,4.880495,5.6999545,4.9693303,4.2405195,3.5098956,2.7792716,2.0504606,1.6407311,1.2291887,0.8194591,0.40972954,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.059827764,0.058014803,0.054388877,0.052575916,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.0297627,2.0595255,3.0892882,4.120864,5.1506267,4.5704784,3.9903307,3.4101827,2.8300345,2.2498865,1.8600996,1.4703126,1.0805258,0.69073874,0.2991388,0.32995918,0.36077955,0.38978696,0.42060733,0.44961473,0.43692398,0.42423326,0.41335547,0.40066472,0.387974,0.6526665,0.91735905,1.1820517,1.4467441,1.7132497,1.3905423,1.067835,0.7451276,0.4224203,0.099712946,0.08339628,0.065266654,0.047137026,0.030820364,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.9499924,1.8999848,2.8499773,3.7999697,4.749962,3.8906176,3.0294604,2.1701162,1.310772,0.44961473,0.36984438,0.29007402,0.21030366,0.13053331,0.05076295,0.09789998,0.14503701,0.19217403,0.23931105,0.28826106,0.23024625,0.17223145,0.11421664,0.058014803,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,2.030518,3.9105604,5.7906027,7.6706448,9.550687,8.265296,6.979906,5.6945157,4.409125,3.1255474,3.9450066,4.764466,5.5857377,6.4051967,7.224656,7.317117,7.409578,7.502039,7.5945,7.686961,6.149569,4.612177,3.0747845,1.5373923,0.0,0.15954071,0.3208944,0.48043507,0.6399758,0.7995165,0.64541465,0.4894999,0.33539808,0.1794833,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07070554,0.13959812,0.21030366,0.27919623,0.34990177,0.90466833,1.4594349,2.0142014,2.570781,3.1255474,3.290527,3.4555066,3.6204863,3.785466,3.9504454,4.9203806,5.8903155,6.8602505,7.8301854,8.80012,7.520169,6.240217,4.9602656,3.680314,2.4003625,1.9525607,1.504759,1.0569572,0.6091554,0.16316663,0.13053331,0.09789998,0.065266654,0.032633327,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.44236287,0.83577573,1.2273756,1.6207886,2.0123885,1.8220274,1.6316663,1.4431182,1.2527572,1.062396,0.85027945,0.63816285,0.42423326,0.21211663,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.25562772,0.5094425,0.7650702,1.020698,1.2745126,1.7150626,2.1556125,2.5943494,3.0348995,3.4754493,3.7909048,4.1045475,4.420003,4.7354584,5.049101,4.115425,3.1799364,2.2444477,1.310772,0.37528324,0.6091554,0.8448406,1.0805258,1.3143979,1.550083,1.7205015,1.8909199,2.0595255,2.229944,2.4003625,2.034144,1.6697385,1.305333,0.93911463,0.5747091,1.4630609,2.3495996,3.2379513,4.12449,5.0128417,5.522284,6.0317264,6.542982,7.0524244,7.5618668,7.9172077,8.272549,8.627889,8.98323,9.336758,9.180842,9.023115,8.865387,8.70766,8.549932,9.327692,10.1054535,10.883214,11.6591625,12.436923,13.180238,13.92174,14.665054,15.406556,16.14987,16.420002,16.690134,16.960264,17.230396,17.500528,19.112251,20.725788,22.337511,23.949236,25.562773,22.903156,20.241728,17.582111,14.922495,12.262879,13.987006,15.712947,17.437075,19.163015,20.887142,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.052575916,0.10515183,0.15772775,0.21030366,0.26287958,0.2574407,0.2520018,0.24837588,0.24293698,0.2374981,0.81764615,1.3977941,1.9779422,2.5580902,3.1382382,3.3648586,3.5932918,3.8199122,4.0483456,4.274966,3.727451,3.1799364,2.6324217,2.084907,1.5373923,1.2291887,0.922798,0.61459434,0.30820364,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.058014803,0.052575916,0.047137026,0.04169814,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.77232206,1.5446441,2.3169663,3.0892882,3.8616104,3.4283123,2.9932013,2.5580902,2.1229792,1.6878681,1.3941683,1.1022812,0.8103943,0.5166943,0.22480737,0.24837588,0.27013144,0.291887,0.3154555,0.33721104,0.33721104,0.33721104,0.33721104,0.33721104,0.33721104,0.5293851,0.72337204,0.9155461,1.1077201,1.2998942,1.067835,0.83577573,0.60190356,0.36984438,0.13778515,0.11421664,0.092461094,0.07070554,0.047137026,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.7124943,1.4249886,2.137483,2.8499773,3.5624714,3.0294604,2.4982624,1.9652514,1.4322405,0.89922947,0.726998,0.55476654,0.3825351,0.21030366,0.038072214,0.08339628,0.12690738,0.17223145,0.21755551,0.26287958,0.21030366,0.15772775,0.10515183,0.052575916,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,1.5228885,2.9315605,4.3420453,5.75253,7.1630154,6.392506,5.621997,4.853301,4.082792,3.3122826,4.590421,5.866747,7.1448855,8.423024,9.699349,8.934279,8.1692095,7.404139,6.640882,5.8758116,4.699199,3.5243993,2.3495996,1.1747998,0.0,0.11965553,0.23931105,0.36077955,0.48043507,0.6000906,0.4894999,0.38072214,0.27013144,0.15954071,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.052575916,0.10515183,0.15772775,0.21030366,0.26287958,0.79770356,1.3325275,1.8673514,2.4021754,2.9369993,3.1182957,3.2977788,3.4772623,3.6567454,3.8380418,4.401873,4.9675174,5.5331616,6.096993,6.6626377,5.727149,4.7916603,3.8579843,2.9224956,1.987007,1.6298534,1.2726997,0.9155461,0.55839247,0.19942589,0.15954071,0.11965553,0.07977036,0.03988518,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.39703882,0.75781834,1.1167849,1.4775645,1.8383441,1.6570477,1.4775645,1.2980812,1.1167849,0.93730164,0.7505665,0.5620184,0.37528324,0.18673515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.19761293,0.39522585,0.59283876,0.7904517,0.9880646,1.3434052,1.696933,2.0522738,2.4076142,2.762955,3.141864,3.5225863,3.9033084,4.2822175,4.6629395,3.8054085,2.9478772,2.0903459,1.2328146,0.37528324,0.5946517,0.81583315,1.0352017,1.2545701,1.4757515,1.5772774,1.6806163,1.7821422,1.8854811,1.987007,1.7078108,1.4268016,1.1476053,0.8684091,0.5873999,1.3506571,2.1121013,2.8753586,3.636803,4.40006,4.8206677,5.239462,5.660069,6.0806766,6.4994707,6.722465,6.94546,7.166641,7.3896356,7.61263,7.572745,7.5328593,7.4929743,7.453089,7.413204,8.00423,8.597069,9.189907,9.782746,10.375585,11.173288,11.969179,12.766883,13.564586,14.362289,15.364858,16.367426,17.369995,18.372562,19.375132,20.838192,22.29944,23.7625,25.225561,26.68681,24.304577,21.922344,19.540112,17.157877,14.775645,15.54978,16.325727,17.099863,17.87581,18.649946,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.059827764,0.11965553,0.1794833,0.23931105,0.2991388,0.3045777,0.3100166,0.3154555,0.3208944,0.3245203,1.1947423,2.0649643,2.9351864,3.8054085,4.6756306,4.309412,3.9450066,3.5806012,3.2143826,2.8499773,2.4855716,2.1193533,1.7549478,1.3905423,1.0243238,0.8194591,0.61459434,0.40972954,0.20486477,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.054388877,0.047137026,0.03988518,0.032633327,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.5148814,1.0297627,1.5446441,2.0595255,2.5744069,2.2843328,1.9942589,1.7041848,1.4141108,1.1258497,0.9300498,0.73424983,0.5402629,0.3444629,0.15047589,0.16497959,0.1794833,0.19579996,0.21030366,0.22480737,0.2374981,0.25018883,0.26287958,0.2755703,0.28826106,0.40791658,0.5275721,0.64722764,0.7668832,0.8883517,0.7451276,0.60190356,0.4604925,0.31726846,0.17585737,0.14684997,0.11965553,0.092461094,0.065266654,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.4749962,0.9499924,1.4249886,1.8999848,2.374981,2.1701162,1.9652514,1.7603867,1.5555218,1.3506571,1.0841516,0.8194591,0.55476654,0.29007402,0.025381476,0.06707962,0.11059072,0.15228885,0.19579996,0.2374981,0.19036107,0.14322405,0.09427405,0.047137026,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,1.015259,1.9543737,2.8953013,3.834416,4.7753434,4.519716,4.265901,4.0102735,3.7546456,3.5008307,5.235836,6.970841,8.705847,10.440851,12.175857,10.553255,8.930654,7.308052,5.6854506,4.062849,3.2506418,2.4384346,1.6244144,0.8122072,0.0,0.07977036,0.15954071,0.23931105,0.3208944,0.40066472,0.33539808,0.27013144,0.20486477,0.13959812,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.034446288,0.07070554,0.10515183,0.13959812,0.17585737,0.69073874,1.2056202,1.7205015,2.2353828,2.7502642,2.9442513,3.1400511,3.3358512,3.529838,3.7256382,3.8851788,4.0447197,4.2042603,4.365614,4.5251546,3.9341288,3.3449159,2.7557032,2.1646774,1.5754645,1.3071461,1.0406405,0.77232206,0.5058166,0.2374981,0.19036107,0.14322405,0.09427405,0.047137026,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.35171473,0.67986095,1.0080072,1.3343405,1.6624867,1.4920682,1.3216497,1.1530442,0.9826257,0.8122072,0.6508536,0.48768693,0.3245203,0.16316663,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13959812,0.27919623,0.42060733,0.56020546,0.69980353,0.969935,1.2400664,1.5101979,1.7803292,2.0504606,2.4946365,2.9406252,3.3848011,3.83079,4.274966,3.4953918,2.715818,1.9344311,1.1548572,0.37528324,0.58014804,0.7850128,0.9898776,1.1947423,1.3996071,1.4358664,1.4703126,1.504759,1.5392052,1.5754645,1.3796645,1.1856775,0.9898776,0.79589057,0.6000906,1.2382535,1.8746033,2.5127661,3.149116,3.787279,4.117238,4.4471974,4.7771564,5.1071157,5.4370747,5.527723,5.618371,5.7072062,5.7978544,5.8866897,5.964647,6.0426044,6.1205616,6.1967063,6.2746634,6.68258,7.0904965,7.498413,7.9045167,8.312433,9.164526,10.018432,10.870523,11.722616,12.574709,14.309713,16.04472,17.779724,19.514729,21.249735,22.562319,23.874905,25.187489,26.500074,27.812658,25.70781,23.60296,21.49811,19.393261,17.286598,17.112555,16.936697,16.762651,16.586794,16.41275,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06707962,0.13415924,0.2030518,0.27013144,0.33721104,0.35171473,0.3680314,0.3825351,0.39703882,0.41335547,1.5718386,2.7321346,3.8924308,5.0527267,6.2130227,5.2557783,4.2967215,3.339477,2.382233,1.4249886,1.2418793,1.0605831,0.8774739,0.69436467,0.51306844,0.40972954,0.30820364,0.20486477,0.10333887,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.052575916,0.04169814,0.032633327,0.02175555,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.2574407,0.5148814,0.77232206,1.0297627,1.2872034,1.1421664,0.99712944,0.8520924,0.7070554,0.5620184,0.46411842,0.3680314,0.27013144,0.17223145,0.07433146,0.08339628,0.09064813,0.09789998,0.10515183,0.11240368,0.13778515,0.16316663,0.18673515,0.21211663,0.2374981,0.28463513,0.33177215,0.38072214,0.42785916,0.4749962,0.4224203,0.36984438,0.31726846,0.26469254,0.21211663,0.1794833,0.14684997,0.11421664,0.08339628,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.2374981,0.4749962,0.7124943,0.9499924,1.1874905,1.310772,1.4322405,1.5555218,1.6769904,1.8002719,1.4431182,1.0841516,0.726998,0.36984438,0.012690738,0.052575916,0.092461094,0.13234627,0.17223145,0.21211663,0.17041849,0.12690738,0.08520924,0.04169814,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.5076295,0.97718686,1.4467441,1.9181144,2.3876717,2.6469254,2.907992,3.1672456,3.4283123,3.6875658,5.8794374,8.073122,10.264994,12.456866,14.650551,12.170418,9.690285,7.210152,4.7300196,2.2498865,1.8002719,1.3506571,0.89922947,0.44961473,0.0,0.03988518,0.07977036,0.11965553,0.15954071,0.19942589,0.1794833,0.15954071,0.13959812,0.11965553,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.018129626,0.034446288,0.052575916,0.07070554,0.0870222,0.581961,1.0768998,1.5718386,2.0667772,2.561716,2.7720199,2.9823234,3.1926272,3.4029307,3.6132345,3.3666716,3.1219215,2.8771715,2.6324217,2.3876717,2.1429217,1.8981718,1.651609,1.4068589,1.162109,0.98443866,0.80676836,0.629098,0.45324063,0.2755703,0.21936847,0.16497959,0.11059072,0.054388877,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.30820364,0.60190356,0.8974165,1.1929294,1.4866294,1.3270886,1.167548,1.0080072,0.8466535,0.6871128,0.5493277,0.41335547,0.2755703,0.13778515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08339628,0.16497959,0.24837588,0.32995918,0.41335547,0.5982776,0.78319985,0.968122,1.1530442,1.3379664,1.8474089,2.3568513,2.8681068,3.3775494,3.8869917,3.1853752,2.4819458,1.7803292,1.0768998,0.37528324,0.5656443,0.7541924,0.9445535,1.1349145,1.3252757,1.2926424,1.260009,1.2273756,1.1947423,1.162109,1.0533313,0.94274056,0.8321498,0.72337204,0.61278135,1.1258497,1.6371052,2.1501737,2.663242,3.1744974,3.4156215,3.6549325,3.8942437,4.135368,4.3746786,4.3329806,4.2894692,4.2477713,4.2042603,4.162562,4.358362,4.552349,4.748149,4.942136,5.137936,5.3591175,5.582112,5.805106,6.0281005,6.249282,7.157576,8.06587,8.972352,9.880646,10.7871275,13.254569,15.722012,18.189453,20.656897,23.124338,24.28826,25.450369,26.612478,27.774588,28.936695,27.10923,25.281763,23.454296,21.626831,19.799364,18.675327,17.549479,16.425442,15.299591,14.175554,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07433146,0.15047589,0.22480737,0.2991388,0.37528324,0.40066472,0.42423326,0.44961473,0.4749962,0.50037766,1.9507477,3.3993049,4.8496747,6.300045,7.750415,6.200332,4.650249,3.100166,1.550083,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.16316663,0.13778515,0.11240368,0.0870222,0.06164073,0.099712946,0.13778515,0.17585737,0.21211663,0.25018883,0.21211663,0.17585737,0.13778515,0.099712946,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.44961473,0.89922947,1.3506571,1.8002719,2.2498865,1.8002719,1.3506571,0.89922947,0.44961473,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.774135,1.550083,2.324218,3.100166,3.874301,6.5248523,9.175404,11.825955,14.474693,17.125244,13.7875805,10.449916,7.112252,3.774588,0.43692398,0.34990177,0.26287958,0.17585737,0.0870222,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.4749962,0.9499924,1.4249886,1.8999848,2.374981,2.5997884,2.8245957,3.049403,3.2742105,3.5008307,2.8499773,2.1991236,1.550083,0.89922947,0.25018883,0.34990177,0.44961473,0.5493277,0.6508536,0.7505665,0.66173136,0.5747091,0.48768693,0.40066472,0.31182957,0.25018883,0.18673515,0.12509441,0.06164073,0.0,0.0,0.0,0.0,0.0,0.0,0.26287958,0.52575916,0.7868258,1.0497054,1.3125849,1.162109,1.0116332,0.8629702,0.7124943,0.5620184,0.44961473,0.33721104,0.22480737,0.11240368,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.22480737,0.3245203,0.42423326,0.52575916,0.62547207,1.2001812,1.7748904,2.3495996,2.9243085,3.5008307,2.8753586,2.2498865,1.6244144,1.0007553,0.37528324,0.5493277,0.72518504,0.89922947,1.0750868,1.2491312,1.1494182,1.0497054,0.9499924,0.85027945,0.7505665,0.72518504,0.69980353,0.6744221,0.6508536,0.62547207,1.0116332,1.3996071,1.7875811,2.175555,2.561716,2.712192,2.8626678,3.0131438,3.1618068,3.3122826,3.1382382,2.962381,2.7883365,2.612479,2.4366217,2.7502642,3.0620937,3.3757362,3.6875658,3.9993954,4.0374675,4.07554,4.1117992,4.1498713,4.1879435,5.1506267,6.11331,7.07418,8.036863,8.999546,12.199425,15.401117,18.600996,21.799063,25.000753,26.012386,27.025833,28.037466,29.049099,30.062546,28.512463,26.96238,25.412296,23.862213,22.31213,20.238102,18.16226,16.08823,14.012388,11.938358,0.3245203,0.26287958,0.19942589,0.13778515,0.07433146,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.059827764,0.11965553,0.1794833,0.23931105,0.2991388,0.35715362,0.41516843,0.47318324,0.5293851,0.5873999,1.7096237,2.8318477,3.9558845,5.0781083,6.200332,4.9602656,3.720199,2.4801328,1.2400664,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.018129626,0.034446288,0.052575916,0.07070554,0.0870222,0.07070554,0.052575916,0.034446288,0.018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.13053331,0.11059072,0.09064813,0.07070554,0.05076295,0.07977036,0.11059072,0.13959812,0.17041849,0.19942589,0.17041849,0.13959812,0.11059072,0.07977036,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.36077955,0.7197462,1.0805258,1.4394923,1.8002719,1.4394923,1.0805258,0.7197462,0.36077955,0.0,0.43692398,0.87566096,1.3125849,1.7495089,2.1882458,1.7495089,1.3125849,0.87566096,0.43692398,0.0,0.18492219,0.36984438,0.55476654,0.73968875,0.9246109,0.73968875,0.55476654,0.36984438,0.18492219,0.0,0.6200332,1.2400664,1.8600996,2.4801328,3.100166,5.219519,7.3406854,9.460039,11.579392,13.700559,11.030065,8.3595705,5.6890764,3.0203958,0.34990177,0.27919623,0.21030366,0.13959812,0.07070554,0.0,0.0,0.0,0.0,0.0,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.045324065,0.09064813,0.13415924,0.1794833,0.22480737,0.1794833,0.13415924,0.09064813,0.045324065,0.0,0.0,0.0,0.0,0.0,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.18492219,0.27013144,0.35534066,0.4405499,0.52575916,1.0098201,1.4956942,1.9797552,2.465629,2.94969,2.9768846,3.005892,3.0330863,3.0602808,3.0874753,2.5127661,1.938057,1.3633479,0.7868258,0.21211663,0.291887,0.37165734,0.45324063,0.533011,0.61278135,0.5402629,0.46774435,0.39522585,0.32270733,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.0,0.0,0.0,0.0,0.0,0.21030366,0.42060733,0.629098,0.83940166,1.0497054,0.9499924,0.85027945,0.7505665,0.6508536,0.5493277,0.5529536,0.55476654,0.55839247,0.56020546,0.5620184,0.44961473,0.33721104,0.22480737,0.11240368,0.0,0.0,0.0,0.0,0.0,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.23568514,0.36984438,0.5058166,0.6399758,0.774135,1.5573349,2.3405347,3.1219215,3.9051213,4.688321,3.9341288,3.1817493,2.42937,1.6769904,0.9246109,1.017072,1.1095331,1.2019942,1.2944553,1.3869164,1.2491312,1.1131591,0.97537386,0.8375887,0.69980353,0.6671702,0.6345369,0.60190356,0.56927025,0.53663695,0.8520924,1.167548,1.4830034,1.7966459,2.1121013,2.2516994,2.3931105,2.5327086,2.6723068,2.811905,2.6976883,2.5816586,2.467442,2.3532255,2.2371957,2.520018,2.8028402,3.0856624,3.3666716,3.6494937,3.7093215,3.7691493,3.83079,3.8906176,3.9504454,4.8678045,5.7851634,6.7025228,7.6198816,8.537241,11.222239,13.907236,16.592234,19.277231,21.962229,23.220425,24.476809,25.735004,26.9932,28.249582,27.564283,26.880796,26.195496,25.510197,24.824896,23.01556,21.20441,19.395073,17.585737,15.774588,0.6508536,0.52575916,0.40066472,0.2755703,0.15047589,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.045324065,0.09064813,0.13415924,0.1794833,0.22480737,0.3154555,0.40429065,0.4949388,0.5855869,0.6744221,1.4703126,2.2643902,3.0602808,3.8543584,4.650249,3.720199,2.7901495,1.8600996,0.9300498,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.09064813,0.06707962,0.045324065,0.02175555,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.09789998,0.08339628,0.06707962,0.052575916,0.038072214,0.059827764,0.08339628,0.10515183,0.12690738,0.15047589,0.12690738,0.10515183,0.08339628,0.059827764,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.27013144,0.5402629,0.8103943,1.0805258,1.3506571,1.0805258,0.8103943,0.5402629,0.27013144,0.0,0.8375887,1.6751775,2.5127661,3.350355,4.1879435,3.350355,2.5127661,1.6751775,0.8375887,0.0,0.36984438,0.73968875,1.1095331,1.4793775,1.8492218,1.4793775,1.1095331,0.73968875,0.36984438,0.0,0.46411842,0.9300498,1.3941683,1.8600996,2.324218,3.9141862,5.504154,7.0959353,8.685904,10.275872,8.272549,6.2692246,4.267714,2.2643902,0.26287958,0.21030366,0.15772775,0.10515183,0.052575916,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.09064813,0.1794833,0.27013144,0.36077955,0.44961473,0.36077955,0.27013144,0.1794833,0.09064813,0.0,0.0,0.0,0.0,0.0,0.0,0.03988518,0.07977036,0.11965553,0.15954071,0.19942589,0.36984438,0.5402629,0.7106813,0.8792868,1.0497054,1.5446441,2.039583,2.5345216,3.0294604,3.5243993,3.3557937,3.1853752,3.0149567,2.8445382,2.6741197,2.175555,1.6751775,1.1747998,0.6744221,0.17585737,0.23568514,0.2955129,0.35534066,0.41516843,0.4749962,0.4169814,0.36077955,0.30276474,0.24474995,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.0,0.0,0.0,0.0,0.0,0.15772775,0.3154555,0.47318324,0.629098,0.7868258,0.73787576,0.6871128,0.63816285,0.5873999,0.53663695,0.6544795,0.77232206,0.8901646,1.0080072,1.1258497,0.89922947,0.6744221,0.44961473,0.22480737,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.24474995,0.41516843,0.5855869,0.7541924,0.9246109,1.9144884,2.904366,3.8942437,4.8841214,5.8758116,4.994712,4.115425,3.2343252,2.3550384,1.4757515,1.4848163,1.4956942,1.504759,1.5156367,1.5247015,1.3506571,1.1747998,1.0007553,0.824898,0.6508536,0.6091554,0.56927025,0.5293851,0.4894999,0.44961473,0.69255173,0.9354887,1.1766127,1.4195497,1.6624867,1.79302,1.9217403,2.0522738,2.182807,2.3133402,2.2571385,2.2027495,2.1483607,2.0921588,2.03777,2.2897718,2.5417736,2.7955883,3.04759,3.299592,3.3829882,3.4645715,3.5479677,3.6295512,3.7129474,4.5849824,5.4570174,6.3308654,7.2029004,8.074935,10.245051,12.415168,14.585284,16.7554,18.925516,20.428463,21.929596,23.43254,24.935488,26.43662,26.617916,26.7974,26.976883,27.15818,27.337664,25.793018,24.246561,22.701918,21.157274,19.612629,0.97537386,0.7868258,0.6000906,0.41335547,0.22480737,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.27194437,0.39522585,0.5166943,0.6399758,0.76325727,1.2291887,1.696933,2.1646774,2.6324217,3.100166,2.4801328,1.8600996,1.2400664,0.6200332,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.027194439,0.054388877,0.08339628,0.11059072,0.13778515,0.11059072,0.08339628,0.054388877,0.027194439,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.065266654,0.054388877,0.045324065,0.034446288,0.025381476,0.03988518,0.054388877,0.07070554,0.08520924,0.099712946,0.08520924,0.07070554,0.054388877,0.03988518,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1794833,0.36077955,0.5402629,0.7197462,0.89922947,0.7197462,0.5402629,0.36077955,0.1794833,0.0,1.2382535,2.474694,3.7129474,4.949388,6.187641,4.949388,3.7129474,2.474694,1.2382535,0.0,0.55476654,1.1095331,1.6642996,2.220879,2.7756457,2.220879,1.6642996,1.1095331,0.55476654,0.0,0.3100166,0.6200332,0.9300498,1.2400664,1.550083,2.610666,3.6694362,4.7300196,5.7906027,6.849373,5.5150323,4.1806917,2.8445382,1.5101979,0.17585737,0.13959812,0.10515183,0.07070554,0.034446288,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13415924,0.27013144,0.40429065,0.5402629,0.6744221,0.5402629,0.40429065,0.27013144,0.13415924,0.0,0.0,0.0,0.0,0.0,0.0,0.059827764,0.11965553,0.1794833,0.23931105,0.2991388,0.55476654,0.8103943,1.064209,1.3198367,1.5754645,2.079468,2.5852847,3.0892882,3.5951047,4.099108,3.73289,3.3648586,2.9968271,2.6306088,2.2625773,1.8383441,1.4122978,0.9880646,0.5620184,0.13778515,0.17767033,0.21755551,0.2574407,0.29732585,0.33721104,0.2955129,0.2520018,0.21030366,0.16679256,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.10515183,0.21030366,0.3154555,0.42060733,0.52575916,0.52575916,0.52575916,0.52575916,0.52575916,0.52575916,0.75781834,0.9898776,1.2219368,1.455809,1.6878681,1.3506571,1.0116332,0.6744221,0.33721104,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.25562772,0.4604925,0.6653573,0.87022203,1.0750868,2.2734551,3.4700103,4.668379,5.864934,7.063302,6.055295,5.047288,4.0392804,3.0330863,2.0250793,1.9525607,1.8800422,1.8075237,1.7350051,1.6624867,1.4503701,1.2382535,1.0243238,0.8122072,0.6000906,0.5529536,0.5058166,0.45686656,0.40972954,0.36259252,0.533011,0.7016165,0.872035,1.0424535,1.2128719,1.3325275,1.452183,1.5718386,1.693307,1.8129625,1.8184015,1.8220274,1.8274662,1.8329052,1.8383441,2.0595255,2.2825198,2.5055144,2.7266958,2.94969,3.054842,3.159994,3.2651455,3.3702974,3.4754493,4.3021603,5.130684,5.957395,6.784106,7.61263,9.267865,10.9230995,12.578335,14.231756,15.8869915,17.634687,19.382383,21.13008,22.877775,24.625471,25.669737,26.715816,27.760082,28.80435,29.85043,28.570477,27.290525,26.010574,24.730623,23.45067,1.2998942,1.0497054,0.7995165,0.5493277,0.2991388,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.23024625,0.38434806,0.5402629,0.69436467,0.85027945,0.9898776,1.1294757,1.2708868,1.4104849,1.550083,1.2400664,0.9300498,0.6200332,0.3100166,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.032633327,0.065266654,0.09789998,0.13053331,0.16316663,0.13053331,0.09789998,0.065266654,0.032633327,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.032633327,0.027194439,0.02175555,0.018129626,0.012690738,0.01994259,0.027194439,0.034446288,0.04169814,0.05076295,0.04169814,0.034446288,0.027194439,0.01994259,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.09064813,0.1794833,0.27013144,0.36077955,0.44961473,0.36077955,0.27013144,0.1794833,0.09064813,0.0,1.6371052,3.2742105,4.9131284,6.550234,8.187339,6.550234,4.9131284,3.2742105,1.6371052,0.0,0.73968875,1.4793775,2.220879,2.960568,3.7002566,2.960568,2.220879,1.4793775,0.73968875,0.0,0.15410182,0.3100166,0.46411842,0.6200332,0.774135,1.305333,1.8347181,2.3641033,2.8953013,3.4246864,2.7575161,2.0903459,1.4231756,0.7541924,0.0870222,0.07070554,0.052575916,0.034446288,0.018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1794833,0.36077955,0.5402629,0.7197462,0.89922947,0.7197462,0.5402629,0.36077955,0.1794833,0.0,0.0,0.0,0.0,0.0,0.0,0.07977036,0.15954071,0.23931105,0.3208944,0.40066472,0.73968875,1.0805258,1.4195497,1.7603867,2.0994108,2.6142921,3.1291735,3.6458678,4.160749,4.6756306,4.1099863,3.5443418,2.9805105,2.4148662,1.8492218,1.49932,1.1494182,0.7995165,0.44961473,0.099712946,0.11965553,0.13959812,0.15954071,0.1794833,0.19942589,0.17223145,0.14503701,0.11784257,0.09064813,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.052575916,0.10515183,0.15772775,0.21030366,0.26287958,0.31182957,0.36259252,0.41335547,0.46230546,0.51306844,0.85934424,1.2074331,1.5555218,1.9017978,2.2498865,1.8002719,1.3506571,0.89922947,0.44961473,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.26469254,0.5058166,0.7451276,0.98443866,1.2255627,2.6306088,4.0356545,5.4407005,6.8457465,8.2507925,7.114065,5.979151,4.844236,3.7093215,2.5744069,2.420305,2.2643902,2.1102884,1.9543737,1.8002719,1.550083,1.2998942,1.0497054,0.7995165,0.5493277,0.4949388,0.4405499,0.38434806,0.32995918,0.2755703,0.37165734,0.46955732,0.56745726,0.6653573,0.76325727,0.872035,0.9826257,1.0932164,1.2019942,1.3125849,1.3778516,1.4431182,1.5083848,1.5718386,1.6371052,1.8292793,2.0232663,2.2154403,2.4076142,2.5997884,2.7266958,2.855416,2.9823234,3.1092308,3.2379513,4.019338,4.802538,5.5857377,6.3671246,7.1503243,8.290678,9.429218,10.5695715,11.709926,12.850279,14.842725,16.83517,18.827616,20.820063,22.812508,24.723372,26.63242,28.543283,30.452332,32.363194,31.347937,30.332678,29.317417,28.302158,27.2869,1.6244144,1.3125849,1.0007553,0.6871128,0.37528324,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.18673515,0.37528324,0.5620184,0.7505665,0.93730164,0.7505665,0.5620184,0.37528324,0.18673515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.03777,4.07554,6.11331,8.149267,10.1870365,8.149267,6.11331,4.07554,2.03777,0.0,0.9246109,1.8492218,2.7756457,3.7002566,4.6248674,3.7002566,2.7756457,1.8492218,0.9246109,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.22480737,0.44961473,0.6744221,0.89922947,1.1258497,0.89922947,0.6744221,0.44961473,0.22480737,0.0,0.0,0.0,0.0,0.0,0.0,0.099712946,0.19942589,0.2991388,0.40066472,0.50037766,0.9246109,1.3506571,1.7748904,2.1991236,2.6251698,3.150929,3.6748753,4.2006345,4.7245803,5.2503395,4.4870825,3.7256382,2.962381,2.1991236,1.4376793,1.162109,0.8883517,0.61278135,0.33721104,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.099712946,0.19942589,0.2991388,0.40066472,0.50037766,0.96268314,1.4249886,1.887294,2.3495996,2.811905,2.2498865,1.6878681,1.1258497,0.5620184,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.2755703,0.5493277,0.824898,1.1004683,1.3742256,2.9877625,4.599486,6.2130227,7.8247466,9.438283,8.174648,6.9128265,5.6491914,4.3873696,3.1255474,2.8880494,2.6505513,2.4130533,2.175555,1.938057,1.649796,1.3633479,1.0750868,0.7868258,0.50037766,0.43692398,0.37528324,0.31182957,0.25018883,0.18673515,0.21211663,0.2374981,0.26287958,0.28826106,0.31182957,0.41335547,0.51306844,0.61278135,0.7124943,0.8122072,0.93730164,1.062396,1.1874905,1.3125849,1.4376793,1.6008459,1.7621996,1.9253663,2.08672,2.2498865,2.4003625,2.5508385,2.6995013,2.8499773,3.000453,3.738329,4.4743915,5.2122674,5.9501433,6.688019,7.311678,7.93715,8.562622,9.188094,9.811753,12.050762,14.287958,16.525154,18.76235,20.999546,23.77519,26.550837,29.324669,32.100315,34.87415,34.125393,33.37483,32.62426,31.875507,31.12494,1.4757515,1.1893034,0.90466833,0.6200332,0.33539808,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.065266654,0.13053331,0.19579996,0.25925365,0.3245203,0.26831847,0.21030366,0.15228885,0.09427405,0.038072214,0.83940166,1.6425442,2.4456866,3.247016,4.0501585,3.4083695,2.764768,2.1229792,1.4793775,0.8375887,0.7016165,0.56745726,0.43329805,0.29732585,0.16316663,0.17767033,0.19217403,0.20667773,0.2229944,0.2374981,0.34083697,0.44236287,0.54570174,0.64722764,0.7505665,0.60190356,0.4550536,0.30820364,0.15954071,0.012690738,0.35534066,0.6979906,1.0406405,1.3832904,1.7259403,1.3905423,1.0551442,0.7197462,0.38434806,0.05076295,0.09064813,0.13053331,0.17041849,0.21030366,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.07433146,0.15047589,0.22480737,0.2991388,0.37528324,0.3245203,0.2755703,0.22480737,0.17585737,0.12509441,0.10333887,0.07977036,0.058014803,0.034446288,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.6298534,3.2597067,4.88956,6.5194135,8.149267,6.5194135,4.88956,3.2597067,1.6298534,0.0,0.73968875,1.4793775,2.220879,2.960568,3.7002566,2.960568,2.220879,1.4793775,0.73968875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.28463513,0.56927025,0.8557183,1.1403534,1.4249886,1.4830034,1.5392052,1.5972201,1.6552348,1.7132497,1.3778516,1.0424535,0.7070554,0.37165734,0.038072214,1.0805258,2.1229792,3.1654327,4.207886,5.2503395,4.9657044,4.6792564,4.3946214,4.1099863,3.825351,4.267714,4.710077,5.1524396,5.5948024,6.037165,5.576673,5.1179934,4.6575007,4.1970086,3.738329,3.000453,2.2625773,1.5247015,0.7868258,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07977036,0.15954071,0.23931105,0.3208944,0.40066472,0.7705091,1.1403534,1.5101979,1.8800422,2.2498865,1.8002719,1.3506571,0.89922947,0.44961473,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.22480737,0.44961473,0.6744221,0.89922947,1.1258497,2.5834718,4.0392804,5.4969025,6.9545245,8.412147,7.2826705,6.153195,5.0219064,3.8924308,2.762955,2.5272698,2.2933977,2.0577126,1.8220274,1.5881553,1.3542831,1.1222239,0.8901646,0.65810543,0.42423326,0.37528324,0.3245203,0.2755703,0.22480737,0.17585737,0.19761293,0.21936847,0.24293698,0.26469254,0.28826106,0.36984438,0.45324063,0.53482395,0.61822027,0.69980353,0.80676836,0.9155461,1.0225109,1.1294757,1.2382535,1.3651608,1.4920682,1.6207886,1.7476959,1.8746033,2.0268922,2.179181,2.333283,2.4855716,2.6378605,3.2506418,3.8634233,4.4743915,5.087173,5.6999545,6.510349,7.320743,8.129324,8.939718,9.750113,11.479679,13.211059,14.940624,16.67019,18.399757,21.050308,23.70086,26.349598,29.000149,31.650702,31.554613,31.46034,31.364252,31.26998,31.175705,1.3252757,1.067835,0.8103943,0.5529536,0.2955129,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.13053331,0.25925365,0.38978696,0.52032024,0.6508536,0.53482395,0.42060733,0.3045777,0.19036107,0.07433146,1.6806163,3.2850883,4.88956,6.495845,8.100317,6.814926,5.529536,4.2441454,2.960568,1.6751775,1.405046,1.1349145,0.86478317,0.5946517,0.3245203,0.35534066,0.38434806,0.41516843,0.44417584,0.4749962,0.49312583,0.5094425,0.5275721,0.54570174,0.5620184,0.4550536,0.3480888,0.23931105,0.13234627,0.025381476,0.7106813,1.3941683,2.079468,2.764768,3.4500678,2.7792716,2.1102884,1.4394923,0.7705091,0.099712946,0.1794833,0.25925365,0.34083697,0.42060733,0.50037766,0.40066472,0.2991388,0.19942589,0.099712946,0.0,0.11240368,0.22480737,0.33721104,0.44961473,0.5620184,0.50037766,0.43692398,0.37528324,0.31182957,0.25018883,0.20486477,0.15954071,0.11421664,0.07070554,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.2219368,2.4456866,3.6676233,4.88956,6.11331,4.88956,3.6676233,2.4456866,1.2219368,0.0,0.55476654,1.1095331,1.6642996,2.220879,2.7756457,2.220879,1.6642996,1.1095331,0.55476654,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.3444629,0.69073874,1.0352017,1.3796645,1.7241274,2.0649643,2.4058013,2.7448254,3.0856624,3.4246864,2.7557032,2.084907,1.4141108,0.7451276,0.07433146,2.0595255,4.0447197,6.0299134,8.015107,10.000301,9.004985,8.009668,7.0143523,6.0208488,5.0255322,5.384499,5.7452784,6.104245,6.4650245,6.825804,6.6680765,6.510349,6.352621,6.1948934,6.037165,4.836984,3.636803,2.4366217,1.2382535,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.059827764,0.11965553,0.1794833,0.23931105,0.2991388,0.57833505,0.8557183,1.1331016,1.4104849,1.6878681,1.3506571,1.0116332,0.6744221,0.33721104,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.17585737,0.34990177,0.52575916,0.69980353,0.87566096,2.1773682,3.4790752,4.782595,6.0843024,7.3878226,6.390693,5.391751,4.3946214,3.397492,2.4003625,2.1683033,1.9344311,1.7023718,1.4703126,1.2382535,1.0605831,0.88291276,0.70524246,0.5275721,0.34990177,0.31182957,0.2755703,0.2374981,0.19942589,0.16316663,0.18310922,0.2030518,0.2229944,0.24293698,0.26287958,0.32814622,0.3934129,0.45686656,0.52213323,0.5873999,0.678048,0.7668832,0.8575313,0.9481794,1.0370146,1.1294757,1.2219368,1.3143979,1.4068589,1.49932,1.6552348,1.8093367,1.9652514,2.1193533,2.275268,2.762955,3.2506418,3.738329,4.2242026,4.7118897,5.7072062,6.7025228,7.6978393,8.693155,9.686659,10.910409,12.132345,13.354282,14.5780325,15.799969,18.325426,20.850883,23.374527,25.899984,28.42544,28.985645,29.54585,30.104244,30.66445,31.224655,1.1747998,0.9445535,0.71430725,0.48587397,0.25562772,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.19579996,0.38978696,0.5855869,0.7795739,0.97537386,0.8031424,0.629098,0.45686656,0.28463513,0.11240368,2.520018,4.9276323,7.3352466,9.742861,12.1504755,10.223296,8.294304,6.3671246,4.439945,2.5127661,2.1066625,1.7023718,1.2980812,0.8919776,0.48768693,0.533011,0.57833505,0.62184614,0.6671702,0.7124943,0.64541465,0.57833505,0.5094425,0.44236287,0.37528324,0.30820364,0.23931105,0.17223145,0.10515183,0.038072214,1.064209,2.0921588,3.1201086,4.1480584,5.1741953,4.169814,3.1654327,2.1592383,1.1548572,0.15047589,0.27013144,0.38978696,0.5094425,0.629098,0.7505665,0.6000906,0.44961473,0.2991388,0.15047589,0.0,0.15047589,0.2991388,0.44961473,0.6000906,0.7505665,0.6744221,0.6000906,0.52575916,0.44961473,0.37528324,0.30820364,0.23931105,0.17223145,0.10515183,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.81583315,1.6298534,2.4456866,3.2597067,4.07554,3.2597067,2.4456866,1.6298534,0.81583315,0.0,0.36984438,0.73968875,1.1095331,1.4793775,1.8492218,1.4793775,1.1095331,0.73968875,0.36984438,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.40429065,0.8103943,1.214685,1.6207886,2.0250793,2.6469254,3.2705846,3.8924308,4.514277,5.137936,4.1317415,3.1273603,2.1229792,1.1167849,0.11240368,3.0403383,5.9682727,8.894395,11.822329,14.750263,13.044266,11.340081,9.634083,7.9298983,6.2257137,6.5030966,6.78048,7.057863,7.3352466,7.61263,7.757667,7.902704,8.047741,8.192778,8.337815,6.6753283,5.0128417,3.350355,1.6878681,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03988518,0.07977036,0.11965553,0.15954071,0.19942589,0.38434806,0.56927025,0.7541924,0.93911463,1.1258497,0.89922947,0.6744221,0.44961473,0.22480737,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.12509441,0.25018883,0.37528324,0.50037766,0.62547207,1.7730774,2.9206827,4.068288,5.2140803,6.3616858,5.4969025,4.632119,3.7673361,2.902553,2.03777,1.8075237,1.5772774,1.3470312,1.1167849,0.8883517,0.7650702,0.6417888,0.52032024,0.39703882,0.2755703,0.25018883,0.22480737,0.19942589,0.17585737,0.15047589,0.16679256,0.18492219,0.2030518,0.21936847,0.2374981,0.28463513,0.33177215,0.38072214,0.42785916,0.4749962,0.5475147,0.6200332,0.69255173,0.7650702,0.8375887,0.89560354,0.95180535,1.0098201,1.067835,1.1258497,1.2817645,1.4394923,1.5972201,1.7549478,1.9126755,2.275268,2.6378605,3.000453,3.3630457,3.7256382,4.9058766,6.0843024,7.264541,8.444779,9.625018,10.339326,11.055446,11.769753,12.485873,13.200181,15.600543,18.000906,20.399454,22.799818,25.20018,26.414865,27.629549,28.844234,30.060732,31.275417,1.0243238,0.823085,0.6200332,0.4169814,0.21574254,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.25925365,0.52032024,0.7795739,1.0406405,1.2998942,1.0696479,0.83940166,0.6091554,0.38072214,0.15047589,3.3594196,6.5701766,9.780933,12.989877,16.200634,13.629852,11.060884,8.490104,5.919323,3.350355,2.810092,2.269829,1.7295663,1.1893034,0.6508536,0.7106813,0.7705091,0.83033687,0.8901646,0.9499924,0.79770356,0.64541465,0.49312583,0.34083697,0.18673515,0.15954071,0.13234627,0.10515183,0.07795739,0.05076295,1.4195497,2.7901495,4.160749,5.529536,6.9001355,5.560356,4.220577,2.8807976,1.5392052,0.19942589,0.36077955,0.52032024,0.67986095,0.83940166,1.0007553,0.7995165,0.6000906,0.40066472,0.19942589,0.0,0.18673515,0.37528324,0.5620184,0.7505665,0.93730164,0.85027945,0.76325727,0.6744221,0.5873999,0.50037766,0.40972954,0.3208944,0.23024625,0.13959812,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.40791658,0.81583315,1.2219368,1.6298534,2.03777,1.6298534,1.2219368,0.81583315,0.40791658,0.0,0.18492219,0.36984438,0.55476654,0.73968875,0.9246109,0.73968875,0.55476654,0.36984438,0.18492219,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.4659314,0.9300498,1.3941683,1.8600996,2.324218,3.2306993,4.135368,5.040036,5.9447045,6.849373,5.5095935,4.169814,2.8300345,1.4902552,0.15047589,4.021151,7.890013,11.760688,15.62955,19.500225,17.08536,14.670493,12.255627,9.840761,7.4258947,7.6198816,7.8156815,8.009668,8.205468,8.399456,8.847258,9.295059,9.742861,10.190662,10.636651,8.511859,6.3870673,4.262275,2.137483,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.19217403,0.28463513,0.3770962,0.46955732,0.5620184,0.44961473,0.33721104,0.22480737,0.11240368,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07433146,0.15047589,0.22480737,0.2991388,0.37528324,1.3669738,2.3604772,3.3521678,4.345671,5.337362,4.604925,3.872488,3.1400511,2.4076142,1.6751775,1.4467441,1.2201238,0.9916905,0.7650702,0.53663695,0.46955732,0.40247768,0.33539808,0.26831847,0.19942589,0.18673515,0.17585737,0.16316663,0.15047589,0.13778515,0.15228885,0.16679256,0.18310922,0.19761293,0.21211663,0.24293698,0.27194437,0.30276474,0.33177215,0.36259252,0.4169814,0.47318324,0.5275721,0.581961,0.63816285,0.65991837,0.68167394,0.70524246,0.726998,0.7505665,0.9101072,1.0696479,1.2291887,1.3905423,1.550083,1.7875811,2.0250793,2.2625773,2.5000753,2.7375734,4.102734,5.467895,6.833056,8.198216,9.563377,9.770056,9.976733,10.185224,10.391902,10.600392,12.87566,15.1509285,17.424383,19.699652,21.97492,23.845898,25.715061,27.584227,29.455204,31.324368,0.87566096,0.69980353,0.52575916,0.34990177,0.17585737,0.0,0.0,0.0,0.0,0.0,0.0,0.3245203,0.6508536,0.97537386,1.2998942,1.6244144,1.3379664,1.0497054,0.76325727,0.4749962,0.18673515,4.2006345,8.212721,12.224807,16.236893,20.250792,17.038223,13.825653,10.613083,7.400513,4.1879435,3.5117085,2.8372865,2.1628644,1.4866294,0.8122072,0.8883517,0.96268314,1.0370146,1.1131591,1.1874905,0.9499924,0.7124943,0.4749962,0.2374981,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,1.7748904,3.48814,5.199577,6.9128265,8.624263,6.9508986,5.275721,3.6005437,1.9253663,0.25018883,0.44961473,0.6508536,0.85027945,1.0497054,1.2491312,1.0007553,0.7505665,0.50037766,0.25018883,0.0,0.22480737,0.44961473,0.6744221,0.89922947,1.1258497,1.0243238,0.9246109,0.824898,0.72518504,0.62547207,0.51306844,0.40066472,0.28826106,0.17585737,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.52575916,1.0497054,1.5754645,2.0994108,2.6251698,3.8126602,5.0001507,6.187641,7.3751316,8.562622,6.887445,5.2122674,3.53709,1.8619126,0.18673515,5.0001507,9.811753,14.625169,19.436771,24.250187,21.12464,18.000906,14.875358,11.74981,8.624263,8.736667,8.8508835,8.963287,9.07569,9.188094,9.936848,10.687414,11.437981,12.186734,12.937301,10.3502035,7.763106,5.1741953,2.5870976,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.96268314,1.8002719,2.6378605,3.4754493,4.313038,3.7129474,3.1128569,2.5127661,1.9126755,1.3125849,1.0877775,0.8629702,0.63816285,0.41335547,0.18673515,0.17585737,0.16316663,0.15047589,0.13778515,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.13778515,0.15047589,0.16316663,0.17585737,0.18673515,0.19942589,0.21211663,0.22480737,0.2374981,0.25018883,0.28826106,0.3245203,0.36259252,0.40066472,0.43692398,0.42423326,0.41335547,0.40066472,0.387974,0.37528324,0.53663695,0.69980353,0.8629702,1.0243238,1.1874905,1.2998942,1.4122978,1.5247015,1.6371052,1.7495089,3.299592,4.8496747,6.399758,7.949841,9.499924,9.200785,8.899834,8.600695,8.299743,8.000604,10.150778,12.300951,14.449312,16.599485,18.749659,21.275116,23.800573,26.324217,28.849674,31.37513,0.8375887,0.67079616,0.50219065,0.33539808,0.16679256,0.0,0.04169814,0.08520924,0.12690738,0.17041849,0.21211663,0.4550536,0.6979906,0.93911463,1.1820517,1.4249886,1.1693609,0.9155461,0.65991837,0.40429065,0.15047589,3.3594196,6.5701766,9.780933,12.989877,16.200634,13.629852,11.060884,8.490104,5.919323,3.350355,2.810092,2.269829,1.7295663,1.1893034,0.6508536,0.7106813,0.7705091,0.83033687,0.8901646,0.9499924,0.7795739,0.6091554,0.4405499,0.27013144,0.099712946,0.39159992,0.6852999,0.97718686,1.2708868,1.5627737,2.762955,3.9631362,5.163317,6.3616858,7.5618668,6.2347784,4.9076896,3.5806012,2.2516994,0.9246109,1.4231756,1.9199274,2.4166791,2.9152439,3.4119956,2.9279346,2.4420607,1.9579996,1.4721256,0.9880646,0.9808127,0.97174793,0.9644961,0.9572442,0.9499924,0.91917205,0.8901646,0.85934424,0.83033687,0.7995165,0.678048,0.55476654,0.43329805,0.3100166,0.18673515,0.15228885,0.11784257,0.08339628,0.047137026,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.034446288,0.07070554,0.10515183,0.13959812,0.17585737,0.13959812,0.10515183,0.07070554,0.034446288,0.0,0.027194439,0.054388877,0.08339628,0.11059072,0.13778515,0.11059072,0.08339628,0.054388877,0.027194439,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.53482395,0.9572442,1.3796645,1.8020848,2.2245052,3.9123733,5.600241,7.28811,8.974165,10.662033,9.066626,7.473032,5.8776245,4.2822175,2.6868105,6.1731377,9.657652,13.142166,16.62668,20.113007,18.042604,15.9722,13.901797,11.833207,9.762803,10.190662,10.616709,11.044568,11.472427,11.900287,11.833207,11.764315,11.697234,11.630155,11.563075,9.3150015,7.066928,4.8206677,2.572594,0.3245203,0.5293851,0.73424983,0.94092757,1.1457924,1.3506571,2.035957,2.7194438,3.4047437,4.0900435,4.7753434,4.844236,4.914942,4.985647,5.0545397,5.125245,4.209699,3.295966,2.38042,1.4648738,0.5493277,0.44961473,0.34990177,0.25018883,0.15047589,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.8448406,1.5899682,2.335096,3.0802233,3.825351,3.2796493,2.7357605,2.1900587,1.6443571,1.1004683,0.91735905,0.73424983,0.5529536,0.36984438,0.18673515,0.17223145,0.15772775,0.14322405,0.12690738,0.11240368,0.11421664,0.11784257,0.11965553,0.12328146,0.12509441,0.13234627,0.13959812,0.14684997,0.15410182,0.16316663,0.17585737,0.18673515,0.19942589,0.21211663,0.22480737,0.2574407,0.29007402,0.32270733,0.35534066,0.387974,0.37528324,0.36259252,0.34990177,0.33721104,0.3245203,0.45686656,0.58921283,0.72337204,0.8557183,0.9880646,1.2074331,1.4268016,1.647983,1.8673514,2.08672,3.3050308,4.5233417,5.7398396,6.9581504,8.174648,7.895452,7.614443,7.3352466,7.0542374,6.775041,8.798307,10.81976,12.843027,14.86448,16.887747,19.237347,21.586945,23.938358,26.287958,28.637556,0.7995165,0.6399758,0.48043507,0.3208944,0.15954071,0.0,0.08520924,0.17041849,0.25562772,0.34083697,0.42423326,0.5855869,0.7451276,0.90466833,1.064209,1.2255627,1.0025684,0.7795739,0.55839247,0.33539808,0.11240368,2.520018,4.9276323,7.3352466,9.742861,12.1504755,10.223296,8.294304,6.3671246,4.439945,2.5127661,2.1066625,1.7023718,1.2980812,0.8919776,0.48768693,0.533011,0.57833505,0.62184614,0.6671702,0.7124943,0.6091554,0.5076295,0.40429065,0.30276474,0.19942589,0.77232206,1.3452182,1.9181144,2.4891977,3.0620937,3.7492065,4.4381323,5.125245,5.812358,6.4994707,5.520471,4.539658,3.5606585,2.5798457,1.6008459,2.3949237,3.1908143,3.9848917,4.780782,5.57486,4.855114,4.135368,3.4156215,2.6958754,1.9743162,1.7350051,1.4956942,1.2545701,1.015259,0.774135,0.81583315,0.8557183,0.89560354,0.9354887,0.97537386,0.8430276,0.7106813,0.57833505,0.44417584,0.31182957,0.25562772,0.19761293,0.13959812,0.08339628,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07070554,0.13959812,0.21030366,0.27919623,0.34990177,0.27919623,0.21030366,0.13959812,0.07070554,0.0,0.054388877,0.11059072,0.16497959,0.21936847,0.2755703,0.21936847,0.16497959,0.11059072,0.054388877,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.045324065,0.09064813,0.13415924,0.1794833,0.22480737,0.54570174,0.86478317,1.1856775,1.504759,1.8256533,4.0120864,6.200332,8.386765,10.57501,12.763257,11.24762,9.731983,8.21816,6.7025228,5.186886,7.344311,9.501737,11.6591625,13.8184,15.975826,14.960567,13.945308,12.930049,11.91479,10.899531,11.642846,12.384347,13.127662,13.8691635,14.612478,13.727753,12.843027,11.958302,11.071762,10.1870365,8.2798,6.3725634,4.465327,2.5580902,0.6508536,1.0605831,1.4703126,1.8800422,2.2897718,2.6995013,4.070101,5.4407005,6.8094873,8.180087,9.550687,9.690285,9.829884,9.969481,10.110892,10.25049,8.419398,6.590119,4.76084,2.9297476,1.1004683,0.89922947,0.69980353,0.50037766,0.2991388,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.726998,1.3796645,2.032331,2.6849976,3.3376641,2.8481643,2.3568513,1.8673514,1.3778516,0.8883517,0.7469406,0.6073425,0.46774435,0.32814622,0.18673515,0.17041849,0.15228885,0.13415924,0.11784257,0.099712946,0.10515183,0.11059072,0.11421664,0.11965553,0.12509441,0.12690738,0.13053331,0.13234627,0.13415924,0.13778515,0.15047589,0.16316663,0.17585737,0.18673515,0.19942589,0.22662032,0.25562772,0.28282216,0.3100166,0.33721104,0.3245203,0.31182957,0.2991388,0.28826106,0.2755703,0.3770962,0.48043507,0.581961,0.6852999,0.7868258,1.114972,1.4431182,1.7694515,2.0975976,2.4257438,3.3104696,4.195195,5.0799212,5.964647,6.849373,6.590119,6.3290524,6.069799,5.810545,5.5494785,7.4458375,9.340384,11.234929,13.129475,15.025834,17.199575,19.375132,21.550686,23.724428,25.899984,0.76325727,0.6091554,0.45686656,0.3045777,0.15228885,0.0,0.12690738,0.25562772,0.3825351,0.5094425,0.63816285,0.71430725,0.79226464,0.87022203,0.9481794,1.0243238,0.83577573,0.64541465,0.4550536,0.26469254,0.07433146,1.6806163,3.2850883,4.88956,6.495845,8.100317,6.814926,5.529536,4.2441454,2.960568,1.6751775,1.405046,1.1349145,0.86478317,0.5946517,0.3245203,0.35534066,0.38434806,0.41516843,0.44417584,0.4749962,0.4405499,0.40429065,0.36984438,0.33539808,0.2991388,1.1530442,2.0051367,2.857229,3.7093215,4.5632267,4.7372713,4.9131284,5.087173,5.2630305,5.4370747,4.804351,4.171627,3.540716,2.907992,2.275268,3.3666716,4.459888,5.5531044,6.644508,7.7377243,6.782293,5.826862,4.8732433,3.917812,2.962381,2.4891977,2.0178273,1.5446441,1.0732739,0.6000906,0.7106813,0.8194591,0.9300498,1.0406405,1.1494182,1.0080072,0.86478317,0.72337204,0.58014804,0.43692398,0.35715362,0.27738327,0.19761293,0.11784257,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.09064813,0.06707962,0.045324065,0.02175555,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.10515183,0.21030366,0.3154555,0.42060733,0.52575916,0.42060733,0.3154555,0.21030366,0.10515183,0.0,0.08339628,0.16497959,0.24837588,0.32995918,0.41335547,0.32995918,0.24837588,0.16497959,0.08339628,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06707962,0.13415924,0.2030518,0.27013144,0.33721104,0.55476654,0.77232206,0.9898776,1.2074331,1.4249886,4.1117992,6.8004227,9.487233,12.175857,14.862667,13.426801,11.992747,10.556881,9.122828,7.686961,8.517298,9.347635,10.177972,11.008308,11.836833,11.876718,11.918416,11.958302,11.998186,12.038072,13.095029,14.151986,15.210756,16.267714,17.32467,15.622298,13.919927,12.217555,10.515183,8.812811,7.2445984,5.678199,4.1099863,2.5417736,0.97537386,1.5899682,2.2045624,2.819157,3.435564,4.0501585,6.104245,8.160145,10.2142315,12.270131,14.324218,14.534521,14.744824,14.955129,15.165432,15.375735,12.629097,9.884272,7.1394467,4.3946214,1.649796,1.3506571,1.0497054,0.7505665,0.44961473,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.6091554,1.1693609,1.7295663,2.2897718,2.8499773,2.4148662,1.9797552,1.5446441,1.1095331,0.6744221,0.57833505,0.48043507,0.3825351,0.28463513,0.18673515,0.16679256,0.14684997,0.12690738,0.10696479,0.0870222,0.09427405,0.10333887,0.11059072,0.11784257,0.12509441,0.12328146,0.11965553,0.11784257,0.11421664,0.11240368,0.12509441,0.13778515,0.15047589,0.16316663,0.17585737,0.19761293,0.21936847,0.24293698,0.26469254,0.28826106,0.2755703,0.26287958,0.25018883,0.2374981,0.22480737,0.29732585,0.36984438,0.44236287,0.5148814,0.5873999,1.0225109,1.4576219,1.892733,2.327844,2.762955,3.3159087,3.8670492,4.420003,4.972956,5.52591,5.2847857,5.045475,4.804351,4.5650396,4.325729,6.093367,7.861006,9.626831,11.39447,13.162108,15.161806,17.163317,19.163015,21.162712,23.16241,0.72518504,0.58014804,0.43511102,0.29007402,0.14503701,0.0,0.17041849,0.34083697,0.5094425,0.67986095,0.85027945,0.8448406,0.83940166,0.83577573,0.83033687,0.824898,0.6671702,0.5094425,0.35171473,0.19579996,0.038072214,0.83940166,1.6425442,2.4456866,3.247016,4.0501585,3.4065566,2.764768,2.1229792,1.4793775,0.8375887,0.7016165,0.56745726,0.43329805,0.29732585,0.16316663,0.17767033,0.19217403,0.20667773,0.2229944,0.2374981,0.27013144,0.30276474,0.33539808,0.3680314,0.40066472,1.5319533,2.665055,3.7981565,4.9294453,6.0625467,5.7253356,5.388125,5.049101,4.7118897,4.3746786,4.0900435,3.8054085,3.5207734,3.2343252,2.94969,4.3402324,5.730775,7.119504,8.510046,9.900589,8.709473,7.520169,6.3308654,5.139749,3.9504454,3.245203,2.5399606,1.8347181,1.1294757,0.42423326,0.6055295,0.7850128,0.9644961,1.1457924,1.3252757,1.1729867,1.020698,0.8665961,0.71430725,0.5620184,0.4604925,0.35715362,0.25562772,0.15228885,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13959812,0.27919623,0.42060733,0.56020546,0.69980353,0.56020546,0.42060733,0.27919623,0.13959812,0.0,0.11059072,0.21936847,0.32995918,0.4405499,0.5493277,0.4405499,0.32995918,0.21936847,0.11059072,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.09064813,0.1794833,0.27013144,0.36077955,0.44961473,0.5656443,0.67986095,0.79589057,0.9101072,1.0243238,4.213325,7.400513,10.587702,13.77489,16.962078,15.607795,14.2516985,12.897416,11.543133,10.1870365,9.690285,9.19172,8.694968,8.198216,7.699652,8.794682,9.88971,10.98474,12.07977,13.174799,14.547212,15.919624,17.292038,18.66445,20.036863,17.516844,14.996826,12.476809,9.956791,7.4367723,6.209397,4.9820213,3.7546456,2.5272698,1.2998942,2.1193533,2.9406252,3.7600844,4.5795436,5.4008155,8.140202,10.879588,13.620788,16.360174,19.099562,19.38057,19.659767,19.940775,20.219973,20.50098,16.840609,13.180238,9.519867,5.859495,2.1991236,1.8002719,1.3996071,1.0007553,0.6000906,0.19942589,0.15954071,0.11965553,0.07977036,0.03988518,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.49312583,0.96087015,1.4268016,1.8945459,2.3622901,1.9815681,1.6026589,1.2219368,0.8430276,0.46230546,0.40791658,0.35171473,0.29732585,0.24293698,0.18673515,0.16497959,0.14322405,0.11965553,0.09789998,0.07433146,0.08520924,0.09427405,0.10515183,0.11421664,0.12509441,0.11784257,0.11059072,0.10333887,0.09427405,0.0870222,0.099712946,0.11240368,0.12509441,0.13778515,0.15047589,0.16679256,0.18492219,0.2030518,0.21936847,0.2374981,0.22480737,0.21211663,0.19942589,0.18673515,0.17585737,0.21755551,0.25925365,0.30276474,0.3444629,0.387974,0.9300498,1.4721256,2.0142014,2.5580902,3.100166,3.3195345,3.540716,3.7600844,3.9794528,4.2006345,3.9794528,3.7600844,3.540716,3.3195345,3.100166,4.740897,6.379815,8.020547,9.659465,11.300196,13.125849,14.94969,16.775343,18.599184,20.424837,0.6871128,0.5493277,0.41335547,0.2755703,0.13778515,0.0,0.21211663,0.42423326,0.63816285,0.85027945,1.062396,0.97537386,0.8883517,0.7995165,0.7124943,0.62547207,0.50037766,0.37528324,0.25018883,0.12509441,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.099712946,0.19942589,0.2991388,0.40066472,0.50037766,1.9126755,3.3249733,4.7372713,6.149569,7.5618668,6.7134004,5.863121,5.0128417,4.162562,3.3122826,3.3757362,3.437377,3.5008307,3.5624714,3.6241121,5.3119802,6.9998484,8.6877165,10.375585,12.06164,10.636651,9.211663,7.7866745,6.3616858,4.936697,3.9993954,3.0620937,2.124792,1.1874905,0.25018883,0.50037766,0.7505665,1.0007553,1.2491312,1.49932,1.3379664,1.1747998,1.0116332,0.85027945,0.6871128,0.5620184,0.43692398,0.31182957,0.18673515,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.17585737,0.34990177,0.52575916,0.69980353,0.87566096,0.69980353,0.52575916,0.34990177,0.17585737,0.0,0.13778515,0.2755703,0.41335547,0.5493277,0.6871128,0.5493277,0.41335547,0.2755703,0.13778515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.11240368,0.22480737,0.33721104,0.44961473,0.5620184,0.5747091,0.5873999,0.6000906,0.61278135,0.62547207,4.313038,8.000604,11.6881695,15.375735,19.063301,17.786976,16.512463,15.23795,13.961625,12.687112,10.863272,9.037619,7.211965,5.388125,3.5624714,5.712645,7.8628187,10.012992,12.163166,14.313339,15.999394,17.687263,19.375132,21.063,22.750868,19.413204,16.075539,12.737875,9.400211,6.0625467,5.1741953,4.2876563,3.3993049,2.5127661,1.6244144,2.6505513,3.6748753,4.699199,5.7253356,6.7496595,10.174346,13.599032,17.025532,20.450218,23.874905,24.224806,24.574707,24.92461,25.274511,25.624413,21.050308,16.474392,11.900287,7.326182,2.7502642,2.2498865,1.7495089,1.2491312,0.7505665,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.37528324,0.7505665,1.1258497,1.49932,1.8746033,1.550083,1.2255627,0.89922947,0.5747091,0.25018883,0.2374981,0.22480737,0.21211663,0.19942589,0.18673515,0.16316663,0.13778515,0.11240368,0.0870222,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.13778515,0.15047589,0.16316663,0.17585737,0.18673515,0.17585737,0.16316663,0.15047589,0.13778515,0.12509441,0.13778515,0.15047589,0.16316663,0.17585737,0.18673515,0.8375887,1.4884423,2.137483,2.7883365,3.437377,3.3249733,3.2125697,3.100166,2.9877625,2.8753586,2.6741197,2.474694,2.275268,2.0758421,1.8746033,3.388427,4.900438,6.412449,7.9244595,9.438283,11.088079,12.737875,14.387671,16.037468,17.687263,0.5493277,0.44780177,0.3444629,0.24293698,0.13959812,0.038072214,0.19942589,0.36259252,0.52575916,0.6871128,0.85027945,0.7795739,0.7106813,0.6399758,0.56927025,0.50037766,0.40066472,0.2991388,0.19942589,0.099712946,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08339628,0.16497959,0.24837588,0.32995918,0.41335547,1.5899682,2.7665808,3.9450066,5.121619,6.300045,5.5857377,4.8696175,4.15531,3.43919,2.7248828,3.0421512,3.3594196,3.6766882,3.9957695,4.313038,5.389938,6.4668374,7.5455503,8.62245,9.699349,8.584378,7.4694057,6.354434,5.239462,4.12449,3.5044568,2.8844235,2.2643902,1.6443571,1.0243238,1.3071461,1.5899682,1.8727903,2.1556125,2.4366217,2.1030366,1.7676386,1.4322405,1.0968424,0.76325727,0.9880646,1.2128719,1.4376793,1.6624867,1.887294,1.7621996,1.6371052,1.5120108,1.3869164,1.261822,1.017072,0.77232206,0.5275721,0.28282216,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.12328146,0.09427405,0.06707962,0.03988518,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13959812,0.27919623,0.42060733,0.56020546,0.69980353,0.56020546,0.42060733,0.27919623,0.13959812,0.0,0.11059072,0.21936847,0.32995918,0.4405499,0.5493277,0.4405499,0.32995918,0.21936847,0.11059072,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.045324065,0.09064813,0.13415924,0.1794833,0.22480737,0.38072214,0.53482395,0.69073874,0.8448406,1.0007553,1.5446441,2.0903459,2.6342347,3.1799364,3.7256382,6.7986097,9.869768,12.9427395,16.01571,19.08687,17.705393,16.322102,14.940624,13.557334,12.175857,11.037316,9.900589,8.762048,7.6253204,6.48678,7.8247466,9.162713,10.500679,11.836833,13.174799,14.257137,15.339477,16.421816,17.504154,18.588305,15.859797,13.1331005,10.4045925,7.6778965,4.949388,4.6357455,4.3202896,4.004834,3.6893787,3.3757362,3.8126602,4.249584,4.688321,5.125245,5.562169,8.830941,12.097899,15.364858,18.631817,21.900587,22.042,22.185223,22.326633,22.469858,22.613083,19.101374,15.593291,12.081583,8.5735,5.0617914,4.265901,3.4681973,2.6704938,1.8727903,1.0750868,0.85934424,0.64541465,0.42967212,0.21574254,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.01994259,0.027194439,0.034446288,0.04169814,0.05076295,0.34083697,0.629098,0.91917205,1.209246,1.49932,1.2400664,0.9808127,0.7197462,0.4604925,0.19942589,0.27013144,0.34083697,0.40972954,0.48043507,0.5493277,0.45324063,0.35534066,0.2574407,0.15954071,0.06164073,0.07070554,0.07795739,0.08520924,0.092461094,0.099712946,0.09064813,0.07977036,0.07070554,0.059827764,0.05076295,0.065266654,0.07977036,0.09427405,0.11059072,0.12509441,0.16497959,0.20486477,0.24474995,0.28463513,0.3245203,0.3444629,0.36440548,0.38434806,0.40429065,0.42423326,0.43329805,0.4405499,0.44780177,0.4550536,0.46230546,0.98443866,1.5083848,2.030518,2.5526514,3.0747845,3.0203958,2.9641938,2.909805,2.855416,2.7992141,2.570781,2.3405347,2.1102884,1.8800422,1.649796,3.2869012,4.9258194,6.5629244,8.200029,9.837135,11.664601,13.492067,15.319533,17.147,18.974466,0.41335547,0.3444629,0.27738327,0.21030366,0.14322405,0.07433146,0.18673515,0.2991388,0.41335547,0.52575916,0.63816285,0.5855869,0.533011,0.48043507,0.42785916,0.37528324,0.2991388,0.22480737,0.15047589,0.07433146,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.065266654,0.13053331,0.19579996,0.25925365,0.3245203,1.2672608,2.2100015,3.152742,4.0954823,5.038223,4.458075,3.877927,3.2977788,2.7176309,2.137483,2.7103791,3.2832751,3.8543584,4.4272547,5.0001507,5.467895,5.9356394,6.4033837,6.869315,7.3370595,6.532104,5.727149,4.9221935,4.117238,3.3122826,3.009518,2.7067533,2.4058013,2.1030366,1.8002719,2.1157274,2.42937,2.7448254,3.0602808,3.3757362,2.8681068,2.3604772,1.8528478,1.3452182,0.8375887,1.4122978,1.987007,2.561716,3.1382382,3.7129474,3.4754493,3.2379513,3.000453,2.762955,2.525457,2.034144,1.5446441,1.0551442,0.5656443,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.09427405,0.07795739,0.059827764,0.04169814,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.10515183,0.21030366,0.3154555,0.42060733,0.52575916,0.42060733,0.3154555,0.21030366,0.10515183,0.0,0.08339628,0.16497959,0.24837588,0.32995918,0.41335547,0.32995918,0.24837588,0.16497959,0.08339628,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.09064813,0.1794833,0.27013144,0.36077955,0.44961473,0.64722764,0.8448406,1.0424535,1.2400664,1.4376793,2.514579,3.5932918,4.670192,5.7470913,6.825804,9.282369,11.740746,14.19731,16.655687,19.112251,17.621996,16.13174,14.643299,13.153044,11.662788,11.213174,10.761745,10.312131,9.862516,9.412902,9.936848,10.462607,10.988366,11.512312,12.038072,12.514881,12.99169,13.470312,13.947122,14.425743,12.308203,10.190662,8.073122,5.955582,3.8380418,4.0954823,4.3529234,4.610364,4.8678045,5.125245,4.974769,4.8242936,4.6756306,4.5251546,4.3746786,7.4857225,10.594954,13.704185,16.815228,19.92446,19.859192,19.795738,19.730473,19.665205,19.59994,17.154251,14.710379,12.264692,9.820818,7.3751316,6.2801023,5.185073,4.0900435,2.9950142,1.8999848,1.5192627,1.1403534,0.75963134,0.38072214,0.0,0.0,0.0,0.0,0.0,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.03988518,0.054388877,0.07070554,0.08520924,0.099712946,0.3045777,0.5094425,0.71430725,0.91917205,1.1258497,0.9300498,0.73424983,0.5402629,0.3444629,0.15047589,0.30276474,0.4550536,0.6073425,0.75963134,0.9119202,0.7433147,0.5728962,0.40247768,0.23205921,0.06164073,0.065266654,0.06707962,0.07070554,0.072518505,0.07433146,0.06707962,0.059827764,0.052575916,0.045324065,0.038072214,0.054388877,0.072518505,0.09064813,0.10696479,0.12509441,0.19217403,0.25925365,0.32814622,0.39522585,0.46230546,0.5148814,0.56745726,0.6200332,0.6726091,0.72518504,0.726998,0.7306239,0.7324369,0.73424983,0.73787576,1.1331016,1.5283275,1.9217403,2.3169663,2.712192,2.715818,2.7176309,2.7194438,2.72307,2.7248828,2.465629,2.2045624,1.9453088,1.6842422,1.4249886,3.1871881,4.949388,6.7134004,8.4756,10.2378,12.242936,14.248073,16.25321,18.256533,20.26167,0.2755703,0.24293698,0.21030366,0.17767033,0.14503701,0.11240368,0.17585737,0.2374981,0.2991388,0.36259252,0.42423326,0.38978696,0.35534066,0.3208944,0.28463513,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.047137026,0.09427405,0.14322405,0.19036107,0.2374981,0.9445535,1.651609,2.3604772,3.0675328,3.774588,3.3304121,2.8844235,2.4402475,1.9942589,1.550083,2.3767939,3.2053177,4.0320287,4.860553,5.6872635,5.5458527,5.4026284,5.2594047,5.1179934,4.974769,4.4798307,3.9848917,3.489953,2.9950142,2.5000753,2.514579,2.5308957,2.5453994,2.5599031,2.5744069,2.9224956,3.2705846,3.6168604,3.9649491,4.313038,3.633177,2.953316,2.2716422,1.5917811,0.9119202,1.8383441,2.762955,3.6875658,4.612177,5.5367875,5.186886,4.836984,4.4870825,4.137181,3.787279,3.053029,2.3169663,1.5827163,0.8466535,0.11240368,0.09064813,0.06707962,0.045324065,0.02175555,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.06707962,0.059827764,0.052575916,0.045324065,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07070554,0.13959812,0.21030366,0.27919623,0.34990177,0.27919623,0.21030366,0.13959812,0.07070554,0.0,0.054388877,0.11059072,0.16497959,0.21936847,0.2755703,0.21936847,0.16497959,0.11059072,0.054388877,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13415924,0.27013144,0.40429065,0.5402629,0.6744221,0.9155461,1.1548572,1.3941683,1.6352923,1.8746033,3.484514,5.0944247,6.7043357,8.314246,9.924157,11.7679405,13.60991,15.45188,17.295664,19.137632,17.540413,15.9431925,14.34416,12.74694,11.14972,11.3872175,11.624716,11.862214,12.099712,12.337211,12.050762,11.762501,11.47424,11.187792,10.899531,10.772624,10.645717,10.516996,10.390089,10.263181,8.754796,7.2482243,5.7398396,4.233268,2.7248828,3.5552197,4.3855567,5.2158933,6.0444174,6.874754,6.1368785,5.4008155,4.6629395,3.925064,3.1871881,6.1405044,9.092008,12.045323,14.996826,17.950142,17.678198,17.40444,17.132496,16.860552,16.586794,15.20713,13.827466,12.447801,11.068136,9.686659,8.294304,6.9019485,5.5095935,4.117238,2.7248828,2.179181,1.6352923,1.0895905,0.54570174,0.0,0.0,0.0,0.0,0.0,0.0,0.045324065,0.09064813,0.13415924,0.1794833,0.22480737,0.1794833,0.13415924,0.09064813,0.045324065,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.059827764,0.08339628,0.10515183,0.12690738,0.15047589,0.27013144,0.38978696,0.5094425,0.629098,0.7505665,0.6200332,0.4894999,0.36077955,0.23024625,0.099712946,0.33539808,0.56927025,0.80495536,1.0406405,1.2745126,1.0333886,0.7904517,0.5475147,0.3045777,0.06164073,0.059827764,0.058014803,0.054388877,0.052575916,0.05076295,0.045324065,0.03988518,0.034446288,0.030820364,0.025381476,0.045324065,0.065266654,0.08520924,0.10515183,0.12509441,0.21936847,0.3154555,0.40972954,0.5058166,0.6000906,0.6852999,0.7705091,0.8557183,0.93911463,1.0243238,1.0225109,1.020698,1.017072,1.015259,1.0116332,1.2799516,1.54827,1.8147756,2.0830941,2.3495996,2.4094272,2.469255,2.5308957,2.5907235,2.6505513,2.3604772,2.0704033,1.7803292,1.4902552,1.2001812,3.0874753,4.974769,6.8620634,8.749357,10.636651,12.819458,15.002265,17.185072,19.36788,21.550686,0.13778515,0.13959812,0.14322405,0.14503701,0.14684997,0.15047589,0.16316663,0.17585737,0.18673515,0.19942589,0.21211663,0.19579996,0.17767033,0.15954071,0.14322405,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.62184614,1.0950294,1.5682126,2.039583,2.5127661,2.2027495,1.892733,1.5827163,1.2726997,0.96268314,2.0450218,3.1273603,4.209699,5.292038,6.3743763,5.621997,4.8696175,4.117238,3.3648586,2.612479,2.427557,2.2426348,2.0577126,1.8727903,1.6878681,2.0196402,2.3532255,2.6849976,3.0167696,3.350355,3.729264,4.1099863,4.4907084,4.8696175,5.2503395,4.3982472,3.5443418,2.6922495,1.840157,0.9880646,2.2625773,3.53709,4.8134155,6.0879283,7.362441,6.9001355,6.43783,5.975525,5.5132194,5.050914,4.070101,3.0892882,2.1102884,1.1294757,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.03988518,0.04169814,0.045324065,0.047137026,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.034446288,0.07070554,0.10515183,0.13959812,0.17585737,0.13959812,0.10515183,0.07070554,0.034446288,0.0,0.027194439,0.054388877,0.08339628,0.11059072,0.13778515,0.11059072,0.08339628,0.054388877,0.027194439,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1794833,0.36077955,0.5402629,0.7197462,0.89922947,1.1820517,1.4648738,1.7476959,2.030518,2.3133402,4.454449,6.5973706,8.740293,10.883214,13.024323,14.253511,15.480887,16.708263,17.935638,19.163015,17.457016,15.752831,14.046834,12.342649,10.636651,11.563075,12.487686,13.412297,14.336908,15.263332,14.162864,13.062395,11.961927,10.863272,9.762803,9.030367,8.29793,7.5654926,6.833056,6.1006193,5.2032027,4.305786,3.4065566,2.5091403,1.6117238,3.0149567,4.41819,5.81961,7.2228427,8.624263,7.3008003,5.975525,4.650249,3.3249733,1.9996977,4.795286,7.5890613,10.384649,13.180238,15.975826,15.495391,15.014956,14.534521,14.054086,13.575464,13.260008,12.944552,12.629097,12.3154545,11.999999,10.310318,8.620637,6.929143,5.239462,3.5497808,2.8390994,2.1302311,1.4195497,0.7106813,0.0,0.0,0.0,0.0,0.0,0.0,0.059827764,0.11965553,0.1794833,0.23931105,0.2991388,0.23931105,0.1794833,0.11965553,0.059827764,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.07977036,0.11059072,0.13959812,0.17041849,0.19942589,0.23568514,0.27013144,0.3045777,0.34083697,0.37528324,0.3100166,0.24474995,0.1794833,0.11421664,0.05076295,0.3680314,0.6852999,1.0025684,1.3198367,1.6371052,1.3216497,1.0080072,0.69255173,0.3770962,0.06164073,0.054388877,0.047137026,0.03988518,0.032633327,0.025381476,0.02175555,0.01994259,0.018129626,0.014503701,0.012690738,0.034446288,0.058014803,0.07977036,0.10333887,0.12509441,0.24837588,0.36984438,0.49312583,0.61459434,0.73787576,0.8557183,0.97174793,1.0895905,1.2074331,1.3252757,1.3180238,1.310772,1.3017071,1.2944553,1.2872034,1.4268016,1.5682126,1.7078108,1.8474089,1.987007,2.1048496,2.222692,2.3405347,2.4583774,2.5744069,2.2553256,1.9344311,1.6153497,1.2944553,0.97537386,2.9877625,5.0001507,7.0125394,9.024928,11.037316,13.397794,15.758271,18.116936,20.477413,22.837889,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.2991388,0.53663695,0.774135,1.0116332,1.2491312,1.0750868,0.89922947,0.72518504,0.5493277,0.37528324,1.7132497,3.049403,4.3873696,5.7253356,7.063302,5.6999545,4.3384194,2.9750717,1.6117238,0.25018883,0.37528324,0.50037766,0.62547207,0.7505665,0.87566096,1.5247015,2.175555,2.8245957,3.4754493,4.12449,4.537845,4.949388,5.3627434,5.774286,6.187641,5.163317,4.137181,3.1128569,2.08672,1.062396,2.6868105,4.313038,5.9374523,7.5618668,9.188094,8.613385,8.036863,7.462154,6.887445,6.3127356,5.087173,3.8634233,2.6378605,1.4122978,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.22480737,0.44961473,0.6744221,0.89922947,1.1258497,1.4503701,1.7748904,2.0994108,2.4257438,2.7502642,5.424384,8.100317,10.774437,13.45037,16.124489,16.73727,17.350052,17.962833,18.575615,19.188396,17.375433,15.56247,13.749508,11.938358,10.125396,11.73712,13.3506565,14.96238,16.575916,18.187641,16.274965,14.362289,12.449615,10.536939,8.624263,7.28811,5.9501433,4.612177,3.2742105,1.938057,1.649796,1.3633479,1.0750868,0.7868258,0.50037766,2.474694,4.4508233,6.4251394,8.399456,10.375585,8.46291,6.550234,4.6375585,2.7248828,0.8122072,3.4500678,6.0879283,8.725789,11.361836,13.999697,13.312584,12.625471,11.938358,11.249433,10.56232,11.312886,12.06164,12.812206,13.562773,14.313339,12.32452,10.337513,8.350506,6.3634987,4.3746786,3.5008307,2.6251698,1.7495089,0.87566096,0.0,0.0,0.0,0.0,0.0,0.0,0.07433146,0.15047589,0.22480737,0.2991388,0.37528324,0.2991388,0.22480737,0.15047589,0.07433146,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.099712946,0.13778515,0.17585737,0.21211663,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.0,0.0,0.0,0.0,0.0,0.40066472,0.7995165,1.2001812,1.6008459,1.9996977,1.6117238,1.2255627,0.8375887,0.44961473,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.2755703,0.42423326,0.5747091,0.72518504,0.87566096,1.0243238,1.1747998,1.3252757,1.4757515,1.6244144,1.6117238,1.6008459,1.5881553,1.5754645,1.5627737,1.5754645,1.5881553,1.6008459,1.6117238,1.6244144,1.8002719,1.9743162,2.1501737,2.324218,2.5000753,2.1501737,1.8002719,1.4503701,1.1004683,0.7505665,2.8880494,5.0255322,7.1630154,9.300498,11.437981,13.974316,16.512463,19.050611,21.586945,24.125093,0.038072214,0.072518505,0.10696479,0.14322405,0.17767033,0.21211663,0.34264994,0.47318324,0.60190356,0.7324369,0.8629702,0.7197462,0.57833505,0.43511102,0.291887,0.15047589,0.291887,0.43511102,0.57833505,0.7197462,0.8629702,0.7850128,0.7070554,0.630911,0.5529536,0.4749962,1.8854811,3.294153,4.704638,6.115123,7.5256076,6.207584,4.88956,3.5733492,2.2553256,0.93730164,0.7505665,0.5620184,0.37528324,0.18673515,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.23931105,0.42967212,0.6200332,0.8103943,1.0007553,0.85934424,0.7197462,0.58014804,0.4405499,0.2991388,1.3705997,2.4402475,3.5098956,4.5795436,5.6491914,4.5632267,3.4754493,2.3876717,1.2998942,0.21211663,0.35171473,0.49312583,0.6327239,0.77232206,0.9119202,1.403233,1.892733,2.382233,2.8717327,3.3630457,3.6966307,4.0320287,4.367427,4.702825,5.038223,4.25321,3.4681973,2.6831846,1.8981718,1.1131591,2.4366217,3.7618973,5.087173,6.412449,7.7377243,7.2029004,6.6680765,6.1332526,5.5966153,5.0617914,4.0846047,3.1074178,2.1302311,1.1530442,0.17585737,0.14684997,0.11965553,0.092461094,0.065266654,0.038072214,0.032633327,0.027194439,0.02175555,0.018129626,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.06707962,0.059827764,0.052575916,0.045324065,0.038072214,0.034446288,0.032633327,0.030820364,0.027194439,0.025381476,0.054388877,0.08520924,0.11421664,0.14503701,0.17585737,0.17767033,0.1794833,0.18310922,0.18492219,0.18673515,0.15954071,0.13234627,0.10515183,0.07795739,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.12328146,0.24474995,0.3680314,0.4894999,0.61278135,0.4894999,0.3680314,0.24474995,0.12328146,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.2374981,0.46230546,0.6871128,0.9119202,1.1367276,1.5827163,2.0268922,2.472881,2.9170568,3.3630457,5.674573,7.987913,10.29944,12.612781,14.924308,15.798156,16.67019,17.542227,18.41426,19.288109,17.397188,15.508082,13.617162,11.728055,9.837135,11.088079,12.337211,13.588155,14.837286,16.08823,14.498261,12.908294,11.318325,9.728357,8.138389,7.1630154,6.187641,5.2122674,4.2368937,3.2633326,2.9351864,2.6070402,2.280707,1.9525607,1.6244144,3.5080826,5.389938,7.271793,9.155461,11.037316,9.157274,7.2772317,5.3971896,3.5171473,1.6371052,3.825351,6.011784,8.200029,10.388275,12.574709,11.920229,11.26575,10.609457,9.954978,9.300498,10.31757,11.334642,12.351714,13.370599,14.387671,12.7777605,11.16785,9.557939,7.948028,6.338117,5.2140803,4.0918565,2.9696326,1.8474089,0.72518504,0.63816285,0.5493277,0.46230546,0.37528324,0.28826106,0.29007402,0.291887,0.2955129,0.29732585,0.2991388,0.4550536,0.6091554,0.7650702,0.91917205,1.0750868,1.1059072,1.1349145,1.1657349,1.1947423,1.2255627,1.2872034,1.3506571,1.4122978,1.4757515,1.5373923,1.4322405,1.3270886,1.2219368,1.1167849,1.0116332,0.90466833,0.79770356,0.69073874,0.581961,0.4749962,0.7850128,1.0950294,1.405046,1.7150626,2.0250793,1.6624867,1.2998942,0.93730164,0.5747091,0.21211663,0.17223145,0.13234627,0.092461094,0.052575916,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.03988518,0.06707962,0.09427405,0.12328146,0.15047589,0.30820364,0.46411842,0.62184614,0.7795739,0.93730164,1.0279498,1.1167849,1.2074331,1.2980812,1.3869164,1.3778516,1.3669738,1.357909,1.3470312,1.3379664,1.4304274,1.5228885,1.6153497,1.7078108,1.8002719,2.0667772,2.335096,2.6034143,2.8699198,3.1382382,2.8880494,2.6378605,2.3876717,2.137483,1.887294,3.9069343,5.9283876,7.948028,9.967669,11.9873085,14.329657,16.672005,19.01435,21.356699,23.70086,0.07433146,0.10696479,0.13959812,0.17223145,0.20486477,0.2374981,0.53482395,0.8321498,1.1294757,1.4268016,1.7241274,1.4394923,1.1548572,0.87022203,0.5855869,0.2991388,0.5855869,0.87022203,1.1548572,1.4394923,1.7241274,1.5700256,1.4141108,1.260009,1.1059072,0.9499924,3.7691493,6.590119,9.409276,12.230246,15.049402,12.415168,9.780933,7.1448855,4.510651,1.8746033,1.49932,1.1258497,0.7505665,0.37528324,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.1794833,0.32270733,0.46411842,0.6073425,0.7505665,0.64541465,0.5402629,0.43511102,0.32995918,0.22480737,1.0279498,1.8292793,2.6324217,3.435564,4.2368937,3.4246864,2.612479,1.8002719,0.9880646,0.17585737,0.32995918,0.48587397,0.6399758,0.79589057,0.9499924,1.2799516,1.6099107,1.93987,2.269829,2.5997884,2.857229,3.1146698,3.3721104,3.6295512,3.8869917,3.343103,2.7974012,2.2516994,1.7078108,1.162109,2.1882458,3.2125697,4.2368937,5.2630305,6.2873545,5.7924156,5.297477,4.802538,4.307599,3.8126602,3.0820365,2.3532255,1.6226015,0.8919776,0.16316663,0.14503701,0.12690738,0.11059072,0.092461094,0.07433146,0.065266654,0.054388877,0.045324065,0.034446288,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.13415924,0.11965553,0.10515183,0.09064813,0.07433146,0.07070554,0.065266654,0.059827764,0.054388877,0.05076295,0.09789998,0.14503701,0.19217403,0.23931105,0.28826106,0.3045777,0.32270733,0.34083697,0.35715362,0.37528324,0.3208944,0.26469254,0.21030366,0.15410182,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.24474995,0.4894999,0.73424983,0.9808127,1.2255627,0.9808127,0.73424983,0.4894999,0.24474995,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.25018883,0.4749962,0.69980353,0.9246109,1.1494182,1.7150626,2.280707,2.8445382,3.4101827,3.975827,5.924762,7.8755093,9.824444,11.775192,13.724127,14.857228,15.99033,17.123432,18.25472,19.387821,17.420757,15.45188,13.484816,11.517752,9.550687,10.437225,11.325577,12.212116,13.100468,13.987006,12.719746,11.452485,10.185224,8.917963,7.650702,7.037921,6.4251394,5.812358,5.199577,4.5867953,4.220577,3.8525455,3.484514,3.1182957,2.7502642,4.539658,6.3290524,8.120259,9.909654,11.700861,9.851639,8.00423,6.156821,4.309412,2.4620032,4.2006345,5.9374523,7.6742706,9.412902,11.14972,10.527874,9.904215,9.282369,8.660522,8.036863,9.322253,10.607644,11.893035,13.176612,14.462003,13.229188,11.998186,10.765372,9.5325575,8.299743,6.929143,5.560356,4.1897564,2.8209698,1.4503701,1.2745126,1.1004683,0.9246109,0.7505665,0.5747091,0.5058166,0.43511102,0.36440548,0.2955129,0.22480737,0.6091554,0.99531645,1.3796645,1.7658255,2.1501737,2.1973107,2.2444477,2.2933977,2.3405347,2.3876717,2.474694,2.561716,2.6505513,2.7375734,2.8245957,2.665055,2.5055144,2.3441606,2.18462,2.0250793,1.8093367,1.5954071,1.3796645,1.1657349,0.9499924,1.1693609,1.3905423,1.6099107,1.8292793,2.0504606,1.7132497,1.3742256,1.0370146,0.69980353,0.36259252,0.2955129,0.22662032,0.15954071,0.092461094,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.054388877,0.08520924,0.11421664,0.14503701,0.17585737,0.34083697,0.5058166,0.67079616,0.83577573,1.0007553,1.0297627,1.0605831,1.0895905,1.1204109,1.1494182,1.1421664,1.1349145,1.1276628,1.1204109,1.1131591,1.2853905,1.4576219,1.6298534,1.8020848,1.9743162,2.335096,2.6958754,3.054842,3.4156215,3.774588,3.6241121,3.4754493,3.3249733,3.1744974,3.0258346,4.9276323,6.82943,8.733041,10.634838,12.536636,14.684997,16.833357,18.979906,21.128265,23.274813,0.11240368,0.14322405,0.17223145,0.2030518,0.23205921,0.26287958,0.726998,1.1929294,1.6570477,2.1229792,2.5870976,2.1592383,1.7331922,1.305333,0.8774739,0.44961473,0.8774739,1.305333,1.7331922,2.1592383,2.5870976,2.3550384,2.1229792,1.889107,1.6570477,1.4249886,5.65463,9.884272,14.115726,18.345367,22.57501,18.622751,14.670493,10.718235,6.7641635,2.811905,2.2498865,1.6878681,1.1258497,0.5620184,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.11965553,0.21574254,0.3100166,0.40429065,0.50037766,0.42967212,0.36077955,0.29007402,0.21936847,0.15047589,0.6852999,1.2201238,1.7549478,2.2897718,2.8245957,2.2879589,1.7495089,1.2128719,0.6744221,0.13778515,0.30820364,0.47680917,0.64722764,0.81764615,0.9880646,1.1566701,1.3270886,1.4975071,1.6679256,1.8383441,2.0178273,2.1973107,2.3767939,2.5580902,2.7375734,2.4329958,2.128418,1.8220274,1.5174497,1.2128719,1.938057,2.663242,3.388427,4.1117992,4.836984,4.3819304,3.926877,3.4718235,3.0167696,2.561716,2.079468,1.5972201,1.114972,0.6327239,0.15047589,0.14322405,0.13415924,0.12690738,0.11965553,0.11240368,0.09789998,0.08339628,0.06707962,0.052575916,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.045324065,0.09064813,0.13415924,0.1794833,0.22480737,0.2030518,0.1794833,0.15772775,0.13415924,0.11240368,0.10515183,0.09789998,0.09064813,0.08339628,0.07433146,0.13959812,0.20486477,0.27013144,0.33539808,0.40066472,0.43329805,0.46411842,0.49675176,0.5293851,0.5620184,0.48043507,0.39703882,0.3154555,0.23205921,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.3680314,0.73424983,1.1022812,1.4703126,1.8383441,1.4703126,1.1022812,0.73424983,0.3680314,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.26287958,0.48768693,0.7124943,0.93730164,1.162109,1.8474089,2.5327086,3.2180085,3.9033084,4.5867953,6.1749506,7.763106,9.349448,10.937603,12.525759,13.918114,15.310469,16.702824,18.095179,19.487535,17.442513,15.397491,13.352469,11.307447,9.262425,9.788185,10.312131,10.837891,11.361836,11.887595,10.943042,9.9966755,9.052122,8.107569,7.1630154,6.9128265,6.6626377,6.412449,6.16226,5.9120708,5.504154,5.0980506,4.690134,4.2822175,3.874301,5.573047,7.26998,8.966913,10.665659,12.362592,10.547816,8.733041,6.9182653,5.101677,3.2869012,4.5759177,5.863121,7.1503243,8.437528,9.724731,9.135518,8.544493,7.95528,7.364254,6.775041,8.326937,9.880646,11.432542,12.984438,14.538147,13.682428,12.826711,11.972805,11.117086,10.263181,8.644206,7.027043,5.40988,3.7927177,2.175555,1.9126755,1.649796,1.3869164,1.1258497,0.8629702,0.7197462,0.57833505,0.43511102,0.291887,0.15047589,0.7650702,1.3796645,1.9942589,2.610666,3.2252605,3.290527,3.3557937,3.4192474,3.484514,3.5497808,3.6621845,3.774588,3.8869917,3.9993954,4.1117992,3.8978696,3.682127,3.4681973,3.2524548,3.0367124,2.715818,2.3931105,2.0704033,1.7476959,1.4249886,1.5555218,1.6842422,1.8147756,1.9453088,2.0758421,1.7621996,1.4503701,1.1367276,0.824898,0.51306844,0.4169814,0.32270733,0.22662032,0.13234627,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.07070554,0.10333887,0.13415924,0.16679256,0.19942589,0.37165734,0.54570174,0.7179332,0.8901646,1.062396,1.0333886,1.0025684,0.97174793,0.94274056,0.9119202,0.90829426,0.90285534,0.8974165,0.8919776,0.8883517,1.1403534,1.3923552,1.6443571,1.8981718,2.1501737,2.6034143,3.054842,3.5080826,3.9595103,4.4127507,4.361988,4.313038,4.262275,4.213325,4.162562,5.9483304,7.7322855,9.518054,11.302009,13.087777,15.040338,16.992899,18.94546,20.89802,22.85058,0.15047589,0.17767033,0.20486477,0.23205921,0.25925365,0.28826106,0.91917205,1.551896,2.18462,2.817344,3.4500678,2.8807976,2.3097143,1.7404441,1.1693609,0.6000906,1.1693609,1.7404441,2.3097143,2.8807976,3.4500678,3.1400511,2.8300345,2.520018,2.2100015,1.8999848,7.5401115,13.180238,18.820364,24.460491,30.100618,24.830336,19.560053,14.289771,9.019489,3.7492065,3.000453,2.2498865,1.49932,0.7505665,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.059827764,0.10696479,0.15410182,0.2030518,0.25018883,0.21574254,0.1794833,0.14503701,0.11059072,0.07433146,0.34264994,0.6091554,0.8774739,1.1457924,1.4122978,1.1494182,0.8883517,0.62547207,0.36259252,0.099712946,0.28463513,0.46955732,0.6544795,0.83940166,1.0243238,1.0352017,1.0442665,1.0551442,1.064209,1.0750868,1.1766127,1.2799516,1.3832904,1.4848163,1.5881553,1.5228885,1.4576219,1.3923552,1.3270886,1.261822,1.6878681,2.1121013,2.5381477,2.962381,3.386614,2.9732587,2.5580902,2.1429217,1.7277533,1.3125849,1.0768998,0.8430276,0.6073425,0.37165734,0.13778515,0.13959812,0.14322405,0.14503701,0.14684997,0.15047589,0.13053331,0.11059072,0.09064813,0.07070554,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.059827764,0.11965553,0.1794833,0.23931105,0.2991388,0.27013144,0.23931105,0.21030366,0.1794833,0.15047589,0.13959812,0.13053331,0.11965553,0.11059072,0.099712946,0.18310922,0.26469254,0.3480888,0.42967212,0.51306844,0.56020546,0.6073425,0.6544795,0.7016165,0.7505665,0.6399758,0.5293851,0.42060733,0.3100166,0.19942589,0.15954071,0.11965553,0.07977036,0.03988518,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.4894999,0.9808127,1.4703126,1.9598125,2.4493124,1.9598125,1.4703126,0.9808127,0.4894999,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.2755703,0.50037766,0.72518504,0.9499924,1.1747998,1.9797552,2.7847104,3.589666,4.3946214,5.199577,6.4251394,7.650702,8.874452,10.100015,11.325577,12.977186,14.630608,16.282217,17.935638,19.587248,17.464268,15.343102,13.220123,11.097144,8.974165,9.137331,9.300498,9.461852,9.625018,9.788185,9.164526,8.54268,7.9208336,7.2971745,6.6753283,6.787732,6.9001355,7.0125394,7.124943,7.2373466,6.789545,6.341743,5.8957543,5.4479527,5.0001507,6.604623,8.209095,9.815379,11.419851,13.024323,11.242181,9.460039,7.6778965,5.8957543,4.1117992,4.949388,5.7869763,6.624565,7.462154,8.299743,7.743163,7.1847706,6.628191,6.069799,5.5132194,7.3334336,9.151835,10.97205,12.792264,14.612478,14.13567,13.657047,13.180238,12.703429,12.224807,10.359268,8.495543,6.630004,4.764466,2.9007401,2.5508385,2.1991236,1.8492218,1.49932,1.1494182,0.9354887,0.7197462,0.5058166,0.29007402,0.07433146,0.91917205,1.7658255,2.610666,3.4555066,4.3003473,4.3819304,4.465327,4.5469103,4.6303062,4.7118897,4.8496747,4.98746,5.125245,5.2630305,5.4008155,5.130684,4.860553,4.590421,4.3202896,4.0501585,3.6204863,3.1908143,2.759329,2.3296568,1.8999848,1.93987,1.9797552,2.0196402,2.0595255,2.0994108,1.8129625,1.5247015,1.2382535,0.9499924,0.66173136,0.5402629,0.4169814,0.2955129,0.17223145,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.08520924,0.11965553,0.15410182,0.19036107,0.22480737,0.40429065,0.5855869,0.7650702,0.9445535,1.1258497,1.0352017,0.9445535,0.8557183,0.7650702,0.6744221,0.6726091,0.67079616,0.6671702,0.6653573,0.66173136,0.99531645,1.3270886,1.6606737,1.9924458,2.324218,2.8699198,3.4156215,3.9595103,4.505212,5.050914,5.0998635,5.1506267,5.199577,5.2503395,5.2992897,6.967215,8.63514,10.303066,11.969179,13.637105,15.3956785,17.15244,18.9092,20.667774,22.424534,0.18673515,0.21211663,0.2374981,0.26287958,0.28826106,0.31182957,1.1131591,1.9126755,2.712192,3.5117085,4.313038,3.6005437,2.8880494,2.175555,1.4630609,0.7505665,1.4630609,2.175555,2.8880494,3.6005437,4.313038,3.925064,3.53709,3.149116,2.762955,2.374981,9.425592,16.474392,23.525002,30.575613,37.624413,31.03792,24.449614,17.863121,11.274815,4.688321,3.7492065,2.811905,1.8746033,0.93730164,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.26287958,0.46230546,0.66173136,0.8629702,1.062396,0.9119202,0.76325727,0.61278135,0.46230546,0.31182957,0.33721104,0.36259252,0.387974,0.41335547,0.43692398,0.61278135,0.7868258,0.96268314,1.1367276,1.3125849,1.4376793,1.5627737,1.6878681,1.8129625,1.938057,1.5627737,1.1874905,0.8122072,0.43692398,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.13778515,0.15047589,0.16316663,0.17585737,0.18673515,0.16316663,0.13778515,0.11240368,0.0870222,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07433146,0.15047589,0.22480737,0.2991388,0.37528324,0.33721104,0.2991388,0.26287958,0.22480737,0.18673515,0.17585737,0.16316663,0.15047589,0.13778515,0.12509441,0.22480737,0.3245203,0.42423326,0.52575916,0.62547207,0.6871128,0.7505665,0.8122072,0.87566096,0.93730164,0.7995165,0.66173136,0.52575916,0.387974,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.61278135,1.2255627,1.8383441,2.4493124,3.0620937,2.4493124,1.8383441,1.2255627,0.61278135,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.28826106,0.51306844,0.73787576,0.96268314,1.1874905,2.1121013,3.0367124,3.9631362,4.8877473,5.812358,6.6753283,7.5382986,8.399456,9.262425,10.125396,12.038072,13.9507475,15.863422,17.774284,19.68696,17.487837,15.2869005,13.087777,10.88684,8.6877165,8.488291,8.287052,8.087626,7.8882003,7.686961,7.3878226,7.0868707,6.787732,6.48678,6.187641,6.6626377,7.137634,7.61263,8.087626,8.562622,8.074935,7.5872483,7.0995617,6.6118746,6.1241875,7.6380115,9.1500225,10.662033,12.175857,13.687867,11.936545,10.1870365,8.437528,6.688019,4.936697,5.3246713,5.712645,6.1006193,6.48678,6.874754,6.350808,5.825049,5.2992897,4.7753434,4.249584,6.338117,8.424837,10.51337,12.60009,14.68681,14.587097,14.487384,14.387671,14.287958,14.188245,12.07433,9.96223,7.850128,5.7380266,3.6241121,3.1871881,2.7502642,2.3133402,1.8746033,1.4376793,1.1494182,0.8629702,0.5747091,0.28826106,0.0,1.0750868,2.1501737,3.2252605,4.3003473,5.375434,5.475147,5.57486,5.674573,5.774286,5.8758116,6.037165,6.200332,6.3616858,6.5248523,6.688019,6.3616858,6.037165,5.712645,5.388125,5.0617914,4.5251546,3.9867048,3.4500678,2.913431,2.374981,2.324218,2.275268,2.2245052,2.175555,2.124792,1.8619126,1.6008459,1.3379664,1.0750868,0.8122072,0.66173136,0.51306844,0.36259252,0.21211663,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.099712946,0.13778515,0.17585737,0.21211663,0.25018883,0.43692398,0.62547207,0.8122072,1.0007553,1.1874905,1.0370146,0.8883517,0.73787576,0.5873999,0.43692398,0.43692398,0.43692398,0.43692398,0.43692398,0.43692398,0.85027945,1.261822,1.6751775,2.08672,2.5000753,3.1382382,3.774588,4.4127507,5.049101,5.6872635,5.8377395,5.9882154,6.1368785,6.2873545,6.43783,7.987913,9.537996,11.088079,12.638163,14.188245,15.749206,17.31198,18.874754,20.437527,22.000301,0.69980353,0.61459434,0.5293851,0.44417584,0.36077955,0.2755703,0.9101072,1.5446441,2.179181,2.8155308,3.4500678,2.8807976,2.3097143,1.7404441,1.1693609,0.6000906,1.3851035,2.1701162,2.955129,3.7401419,4.5251546,4.0574102,3.589666,3.1219215,2.6541772,2.1882458,7.783048,13.377851,18.972654,24.567455,30.162258,24.879286,19.598125,14.315152,9.03218,3.7492065,3.0602808,2.3695421,1.6806163,0.9898776,0.2991388,0.23931105,0.1794833,0.11965553,0.059827764,0.0,0.0,0.0,0.0,0.0,0.0,0.018129626,0.034446288,0.052575916,0.07070554,0.0870222,0.16679256,0.24837588,0.32814622,0.40791658,0.48768693,1.3724127,2.2571385,3.141864,4.028403,4.9131284,4.1117992,3.3122826,2.5127661,1.7132497,0.9119202,1.0333886,1.1530442,1.2726997,1.3923552,1.5120108,1.5156367,1.5174497,1.5192627,1.5228885,1.5247015,1.4666867,1.4104849,1.35247,1.2944553,1.2382535,1.3252757,1.4122978,1.49932,1.5881553,1.6751775,1.4576219,1.2400664,1.0225109,0.80495536,0.5873999,1.0877775,1.5881553,2.08672,2.5870976,3.0874753,3.1128569,3.1382382,3.1618068,3.1871881,3.2125697,2.8699198,2.5272698,2.18462,1.84197,1.49932,1.2273756,0.9554313,0.68167394,0.40972954,0.13778515,0.11059072,0.08339628,0.054388877,0.027194439,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06707962,0.13415924,0.2030518,0.27013144,0.33721104,0.6526665,0.968122,1.2817645,1.5972201,1.9126755,1.6099107,1.3071461,1.0043813,0.7016165,0.40066472,0.4550536,0.5094425,0.5656443,0.6200332,0.6744221,0.7179332,0.75963134,0.8031424,0.8448406,0.8883517,0.7668832,0.64722764,0.5275721,0.40791658,0.28826106,0.23024625,0.17223145,0.11421664,0.058014803,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.5275721,1.0297627,1.5319533,2.034144,2.5381477,2.13567,1.7331922,1.3307146,0.92823684,0.52575916,0.52575916,0.52575916,0.52575916,0.52575916,0.52575916,0.42060733,0.3154555,0.21030366,0.10515183,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.23024625,0.40972954,0.58921283,0.7705091,0.9499924,1.7821422,2.6142921,3.4482548,4.2804046,5.1125546,6.16226,7.211965,8.26167,9.313189,10.362894,11.91479,13.466686,15.020395,16.57229,18.124187,16.095482,14.064963,12.034446,10.00574,7.9752226,7.723221,7.4694057,7.217404,6.965402,6.7115874,6.814926,6.9182653,7.019791,7.12313,7.224656,7.6198816,8.015107,8.410334,8.805559,9.200785,8.432089,7.665206,6.8983226,6.1296263,5.3627434,7.382384,9.402024,11.423477,13.443117,15.462758,13.383289,11.302009,9.222541,7.1430726,5.0617914,6.0879283,7.112252,8.138389,9.162713,10.1870365,9.690285,9.19172,8.694968,8.198216,7.699652,8.716724,9.735609,10.752681,11.769753,12.786825,13.722314,14.657803,15.593291,16.526966,17.462456,14.549025,11.637406,8.725789,5.812358,2.9007401,2.5508385,2.1991236,1.8492218,1.49932,1.1494182,0.91917205,0.69073874,0.4604925,0.23024625,0.0,0.85934424,1.7205015,2.5798457,3.43919,4.3003473,4.3801174,4.459888,4.539658,4.6194286,4.699199,4.860553,5.0200934,5.179634,5.3391747,5.5005283,5.2140803,4.9294453,4.64481,4.360175,4.07554,3.6422417,3.2107568,2.7774587,2.3441606,1.9126755,1.8782293,1.84197,1.8075237,1.7730774,1.7368182,1.5754645,1.4122978,1.2491312,1.0877775,0.9246109,0.75781834,0.58921283,0.4224203,0.25562772,0.0870222,0.092461094,0.09789998,0.10333887,0.10696479,0.11240368,0.15047589,0.18673515,0.22480737,0.26287958,0.2991388,0.46955732,0.6399758,0.8103943,0.9808127,1.1494182,1.0225109,0.89560354,0.7668832,0.6399758,0.51306844,0.5620184,0.61278135,0.66173136,0.7124943,0.76325727,1.1476053,1.5319533,1.9181144,2.3024626,2.6868105,3.2016919,3.7183862,4.233268,4.748149,5.2630305,5.504154,5.7470913,5.9900284,6.2329655,6.4759026,8.029612,9.585134,11.1406555,12.694364,14.249886,14.9877615,15.725637,16.4617,17.199575,17.937452,1.2128719,1.017072,0.823085,0.62728506,0.43329805,0.2374981,0.7070554,1.1766127,1.647983,2.1175404,2.5870976,2.1592383,1.7331922,1.305333,0.8774739,0.44961473,1.3071461,2.1646774,3.0222087,3.87974,4.7372713,4.1897564,3.6422417,3.094727,2.5472124,1.9996977,6.1405044,10.279498,14.420304,18.559298,22.700104,18.722466,14.744824,10.767185,6.789545,2.811905,2.3695421,1.9271792,1.4848163,1.0424535,0.6000906,0.48043507,0.36077955,0.23931105,0.11965553,0.0,0.0,0.0,0.0,0.0,0.0,0.034446288,0.07070554,0.10515183,0.13959812,0.17585737,0.33539808,0.4949388,0.6544795,0.81583315,0.97537386,2.7321346,4.4907084,6.247469,8.00423,9.762803,7.9625316,6.16226,4.361988,2.561716,0.76325727,1.1530442,1.5428312,1.9326181,2.322405,2.712192,2.6922495,2.6723068,2.6523643,2.6324217,2.612479,2.322405,2.032331,1.742257,1.452183,1.162109,1.2128719,1.261822,1.3125849,1.3633479,1.4122978,1.35247,1.2926424,1.2328146,1.1729867,1.1131591,2.0994108,3.0874753,4.07554,5.0617914,6.049856,6.0879283,6.1241875,6.16226,6.200332,6.2384043,5.576673,4.9167547,4.256836,3.5969179,2.9369993,2.4058013,1.8727903,1.3397794,0.80676836,0.2755703,0.21936847,0.16497959,0.11059072,0.054388877,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.059827764,0.11965553,0.1794833,0.23931105,0.2991388,0.968122,1.6352923,2.3024626,2.9696326,3.636803,3.045777,2.4529383,1.8600996,1.2672608,0.6744221,0.6852999,0.69436467,0.70524246,0.71430725,0.72518504,0.7469406,0.7705091,0.79226464,0.81583315,0.8375887,0.73424983,0.6327239,0.5293851,0.42785916,0.3245203,0.25925365,0.19579996,0.13053331,0.065266654,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.44236287,0.83577573,1.2273756,1.6207886,2.0123885,1.8202144,1.6280404,1.4358664,1.2418793,1.0497054,1.0497054,1.0497054,1.0497054,1.0497054,1.0497054,0.83940166,0.630911,0.42060733,0.21030366,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.17223145,0.30820364,0.44236287,0.57833505,0.7124943,1.452183,2.1918716,2.9333735,3.673062,4.4127507,5.6491914,6.887445,8.125698,9.362139,10.600392,11.793322,12.984438,14.177367,15.3702965,16.563227,14.703127,12.843027,10.982927,9.122828,7.262728,6.9581504,6.6517596,6.347182,6.0426044,5.7380266,6.24203,6.7478466,7.25185,7.757667,8.26167,8.577126,8.892582,9.208037,9.52168,9.837135,8.789243,7.743163,6.695271,5.6473784,4.599486,7.1267557,9.654026,12.183108,14.710379,17.237648,14.828221,12.416981,10.007553,7.5981264,5.186886,6.849373,8.511859,10.174346,11.836833,13.499319,13.029762,12.5602045,12.090648,11.619277,11.14972,11.097144,11.044568,10.991992,10.939416,10.88684,12.857531,14.828221,16.797098,18.767788,20.736666,17.025532,13.312584,9.599637,5.8885026,2.175555,1.9126755,1.649796,1.3869164,1.1258497,0.8629702,0.69073874,0.5166943,0.3444629,0.17223145,0.0,0.64541465,1.2908293,1.9344311,2.5798457,3.2252605,3.2850883,3.3449159,3.4047437,3.4645715,3.5243993,3.682127,3.8398547,3.9975824,4.15531,4.313038,4.068288,3.8217251,3.576975,3.3322253,3.0874753,2.759329,2.4329958,2.1048496,1.7767034,1.4503701,1.4304274,1.4104849,1.3905423,1.3705997,1.3506571,1.2872034,1.2255627,1.162109,1.1004683,1.0370146,0.8520924,0.6671702,0.48224804,0.29732585,0.11240368,0.12328146,0.13234627,0.14322405,0.15228885,0.16316663,0.19942589,0.2374981,0.2755703,0.31182957,0.34990177,0.50219065,0.6544795,0.80676836,0.96087015,1.1131591,1.0080072,0.90285534,0.79770356,0.69255173,0.5873999,0.6871128,0.7868258,0.8883517,0.9880646,1.0877775,1.4449311,1.8020848,2.1592383,2.518205,2.8753586,3.2669585,3.6603715,4.0519714,4.445384,4.836984,5.1723824,5.5077806,5.8431783,6.1767635,6.5121617,8.073122,9.63227,11.193231,12.752378,14.313339,14.224504,14.137483,14.05046,13.961625,13.874602,1.7241274,1.4195497,1.114972,0.8103943,0.5058166,0.19942589,0.5058166,0.8103943,1.114972,1.4195497,1.7241274,1.4394923,1.1548572,0.87022203,0.5855869,0.2991388,1.2291887,2.1592383,3.0892882,4.019338,4.949388,4.322103,3.6948178,3.0675328,2.4402475,1.8129625,4.49796,7.1829576,9.867955,12.552953,15.23795,12.565643,9.893337,7.219217,4.5469103,1.8746033,1.6806163,1.4848163,1.2908293,1.0950294,0.89922947,0.7197462,0.5402629,0.36077955,0.1794833,0.0,0.0,0.0,0.0,0.0,0.0,0.052575916,0.10515183,0.15772775,0.21030366,0.26287958,0.50219065,0.7433147,0.9826257,1.2219368,1.4630609,4.0918565,6.722465,9.353074,11.98187,14.612478,11.813264,9.012237,6.2130227,3.4119956,0.61278135,1.2726997,1.9326181,2.5925364,3.2524548,3.9123733,3.870675,3.827164,3.785466,3.7419548,3.7002566,3.1781235,2.6541772,2.132044,1.6099107,1.0877775,1.1004683,1.1131591,1.1258497,1.1367276,1.1494182,1.2473183,1.3452182,1.4431182,1.5392052,1.6371052,3.1128569,4.5867953,6.0625467,7.5382986,9.012237,9.063,9.11195,9.162713,9.211663,9.262425,8.285239,7.308052,6.3290524,5.351866,4.3746786,3.5824142,2.7901495,1.9978848,1.2056202,0.41335547,0.32995918,0.24837588,0.16497959,0.08339628,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.052575916,0.10515183,0.15772775,0.21030366,0.26287958,1.2817645,2.3024626,3.3231604,4.3420453,5.3627434,4.4798307,3.5969179,2.715818,1.8329052,0.9499924,0.9155461,0.8792868,0.8448406,0.8103943,0.774135,0.7777609,0.7795739,0.78319985,0.7850128,0.7868258,0.7016165,0.61822027,0.533011,0.44780177,0.36259252,0.29007402,0.21755551,0.14503701,0.072518505,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.35715362,0.6399758,0.922798,1.2056202,1.4866294,1.504759,1.5228885,1.5392052,1.5573349,1.5754645,1.5754645,1.5754645,1.5754645,1.5754645,1.5754645,1.260009,0.9445535,0.629098,0.3154555,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.11421664,0.20486477,0.2955129,0.38434806,0.4749962,1.1222239,1.7694515,2.4166791,3.0657198,3.7129474,5.137936,6.5629244,7.987913,9.412902,10.837891,11.67004,12.50219,13.33434,14.168303,15.000452,13.310771,11.619277,9.929596,8.239915,6.550234,6.19308,5.8341136,5.47696,5.1198063,4.762653,5.670947,6.5774283,7.4857225,8.392203,9.300498,9.53437,9.770056,10.00574,10.239613,10.475298,9.14821,7.819308,6.492219,5.1651306,3.8380418,6.872941,9.907841,12.9427395,15.977639,19.012539,16.273151,13.531953,10.792566,8.05318,5.3119802,7.61263,9.91328,12.212116,14.512766,16.811602,16.36924,15.926876,15.484513,15.0421505,14.599788,13.477564,12.35534,11.233116,10.110892,8.9868555,11.992747,14.996826,18.002718,21.006798,24.01269,19.500225,14.9877615,10.475298,5.962834,1.4503701,1.2745126,1.1004683,0.9246109,0.7505665,0.5747091,0.4604925,0.3444629,0.23024625,0.11421664,0.0,0.42967212,0.85934424,1.2908293,1.7205015,2.1501737,2.1900587,2.229944,2.269829,2.3097143,2.3495996,2.5055144,2.659616,2.8155308,2.9696326,3.1255474,2.9206827,2.715818,2.5091403,2.3042755,2.0994108,1.8782293,1.6552348,1.4322405,1.209246,0.9880646,0.9826257,0.97718686,0.97174793,0.968122,0.96268314,1.0007553,1.0370146,1.0750868,1.1131591,1.1494182,0.9481794,0.7451276,0.5420758,0.34083697,0.13778515,0.15228885,0.16679256,0.18310922,0.19761293,0.21211663,0.25018883,0.28826106,0.3245203,0.36259252,0.40066472,0.53482395,0.67079616,0.80495536,0.93911463,1.0750868,0.9916905,0.9101072,0.82671094,0.7451276,0.66173136,0.8122072,0.96268314,1.1131591,1.261822,1.4122978,1.742257,2.0722163,2.4021754,2.7321346,3.0620937,3.3322253,3.6023567,3.872488,4.1426196,4.4127507,4.84061,5.2666564,5.6945157,6.1223745,6.550234,8.1148205,9.679407,11.245807,12.810393,14.37498,13.46306,12.549327,11.637406,10.725487,9.811753,2.2371957,1.8220274,1.4068589,0.9916905,0.57833505,0.16316663,0.30276474,0.44236287,0.581961,0.72337204,0.8629702,0.7197462,0.57833505,0.43511102,0.291887,0.15047589,1.1530442,2.1556125,3.1581807,4.160749,5.163317,4.454449,3.7473936,3.0403383,2.333283,1.6244144,2.855416,4.0846047,5.315606,6.544795,7.7739835,6.4070096,5.040036,3.673062,2.3042755,0.93730164,0.9898776,1.0424535,1.0950294,1.1476053,1.2001812,0.96087015,0.7197462,0.48043507,0.23931105,0.0,0.0,0.0,0.0,0.0,0.0,0.07070554,0.13959812,0.21030366,0.27919623,0.34990177,0.67079616,0.9898776,1.310772,1.6298534,1.9507477,5.4515786,8.954222,12.456866,15.95951,19.462152,15.662184,11.862214,8.062244,4.262275,0.46230546,1.3923552,2.322405,3.2524548,4.1825047,5.1125546,5.047288,4.9820213,4.9167547,4.853301,4.788034,4.0320287,3.2778363,2.521831,1.7676386,1.0116332,0.9880646,0.96268314,0.93730164,0.9119202,0.8883517,1.1421664,1.3977941,1.651609,1.9072367,2.1628644,4.12449,6.0879283,8.049554,10.012992,11.974618,12.038072,12.099712,12.163166,12.224807,12.28826,10.991992,9.697536,8.403082,7.1068134,5.812358,4.76084,3.7075086,2.6541772,1.6026589,0.5493277,0.4405499,0.32995918,0.21936847,0.11059072,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.045324065,0.09064813,0.13415924,0.1794833,0.22480737,1.5972201,2.9696326,4.3420453,5.714458,7.0868707,5.915697,4.74271,3.5697234,2.3967366,1.2255627,1.1457924,1.064209,0.98443866,0.90466833,0.824898,0.80676836,0.7904517,0.77232206,0.7541924,0.73787576,0.67079616,0.60190356,0.53482395,0.46774435,0.40066472,0.3208944,0.23931105,0.15954071,0.07977036,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.27194437,0.44417584,0.61822027,0.7904517,0.96268314,1.1893034,1.4177368,1.6443571,1.8727903,2.0994108,2.0994108,2.0994108,2.0994108,2.0994108,2.0994108,1.6806163,1.260009,0.83940166,0.42060733,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.058014803,0.10333887,0.14684997,0.19217403,0.2374981,0.79226464,1.3470312,1.9017978,2.4583774,3.0131438,4.6248674,6.2365913,7.850128,9.461852,11.075388,11.546759,12.019942,12.493125,12.964496,13.437678,11.916603,10.397341,8.8780775,7.3570023,5.8377395,5.42801,5.0182805,4.606738,4.1970086,3.787279,5.0980506,6.4070096,7.7177815,9.026741,10.337513,10.493427,10.64753,10.801631,10.957546,11.111648,9.5053625,7.897265,6.2891674,4.6828823,3.0747845,6.6173134,10.1598425,13.702372,17.2449,20.78743,17.718082,14.646925,11.5775795,8.508233,5.4370747,8.375887,11.312886,14.249886,17.186886,20.125698,19.71053,19.29536,18.880192,18.465023,18.049856,15.857984,13.664299,11.472427,9.280556,7.0868707,11.127964,15.167245,19.208338,23.24762,27.2869,21.97492,16.66294,11.349146,6.037165,0.72518504,0.63816285,0.5493277,0.46230546,0.37528324,0.28826106,0.23024625,0.17223145,0.11421664,0.058014803,0.0,0.21574254,0.42967212,0.64541465,0.85934424,1.0750868,1.0950294,1.114972,1.1349145,1.1548572,1.1747998,1.3270886,1.4793775,1.6316663,1.7857682,1.938057,1.7730774,1.6080978,1.4431182,1.2781386,1.1131591,0.99531645,0.8774739,0.75963134,0.6417888,0.52575916,0.53482395,0.54570174,0.55476654,0.5656443,0.5747091,0.7124943,0.85027945,0.9880646,1.1258497,1.261822,1.0424535,0.823085,0.60190356,0.3825351,0.16316663,0.18310922,0.2030518,0.2229944,0.24293698,0.26287958,0.2991388,0.33721104,0.37528324,0.41335547,0.44961473,0.56745726,0.6852999,0.8031424,0.91917205,1.0370146,0.97718686,0.91735905,0.8575313,0.79770356,0.73787576,0.93730164,1.1367276,1.3379664,1.5373923,1.7368182,2.039583,2.3423476,2.6451125,2.9478772,3.2506418,3.397492,3.5443418,3.6930048,3.8398547,3.9867048,4.507025,5.027345,5.5476656,6.0679855,6.588306,8.158332,9.728357,11.298383,12.866595,14.436621,12.699803,10.962985,9.224354,7.4875355,5.750717,2.7502642,2.2245052,1.7005589,1.1747998,0.6508536,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,1.0750868,2.1501737,3.2252605,4.3003473,5.375434,4.5867953,3.7999697,3.0131438,2.2245052,1.4376793,1.2128719,0.9880646,0.76325727,0.53663695,0.31182957,0.25018883,0.18673515,0.12509441,0.06164073,0.0,0.2991388,0.6000906,0.89922947,1.2001812,1.49932,1.2001812,0.89922947,0.6000906,0.2991388,0.0,0.0,0.0,0.0,0.0,0.0,0.0870222,0.17585737,0.26287958,0.34990177,0.43692398,0.8375887,1.2382535,1.6371052,2.03777,2.4366217,6.813113,11.187792,15.56247,19.93715,24.311829,19.512917,14.712192,9.911467,5.1125546,0.31182957,1.5120108,2.712192,3.9123733,5.1125546,6.3127356,6.2257137,6.1368785,6.049856,5.962834,5.8758116,4.8877473,3.8996825,2.911618,1.9253663,0.93730164,0.87566096,0.8122072,0.7505665,0.6871128,0.62547207,1.0370146,1.4503701,1.8619126,2.275268,2.6868105,5.137936,7.5872483,10.038374,12.487686,14.936998,15.013144,15.087475,15.161806,15.23795,15.312282,13.700559,12.087022,10.475298,8.861761,7.250037,5.9374523,4.6248674,3.3122826,1.9996977,0.6871128,0.5493277,0.41335547,0.2755703,0.13778515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,1.9126755,3.636803,5.3627434,7.0868707,8.812811,7.3497505,5.8866897,4.4254417,2.962381,1.49932,1.3742256,1.2491312,1.1258497,1.0007553,0.87566096,0.8375887,0.7995165,0.76325727,0.72518504,0.6871128,0.63816285,0.5873999,0.53663695,0.48768693,0.43692398,0.34990177,0.26287958,0.17585737,0.0870222,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.18673515,0.25018883,0.31182957,0.37528324,0.43692398,0.87566096,1.3125849,1.7495089,2.1882458,2.6251698,2.6251698,2.6251698,2.6251698,2.6251698,2.6251698,2.0994108,1.5754645,1.0497054,0.52575916,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.46230546,0.9246109,1.3869164,1.8492218,2.3133402,4.1117992,5.9120708,7.7123427,9.512614,11.312886,11.42529,11.537694,11.650098,11.762501,11.874905,10.524248,9.175404,7.8247466,6.474089,5.125245,4.6629395,4.2006345,3.738329,3.2742105,2.811905,4.5251546,6.2365913,7.949841,9.663091,11.374527,11.450671,11.525003,11.599335,11.675479,11.74981,9.862516,7.9752226,6.0879283,4.2006345,2.3133402,6.3634987,10.411844,14.462003,18.512161,22.562319,19.163015,15.761897,12.362592,8.963287,5.562169,9.137331,12.712494,16.287657,19.862818,23.43798,23.050007,22.662033,22.275871,21.887897,21.499924,18.236591,14.975071,11.711739,8.450218,5.186886,10.263181,15.337664,20.412146,25.486628,30.562923,24.449614,18.338116,12.224807,6.11331,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.15047589,0.2991388,0.44961473,0.6000906,0.7505665,0.62547207,0.50037766,0.37528324,0.25018883,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.0870222,0.11240368,0.13778515,0.16316663,0.18673515,0.42423326,0.66173136,0.89922947,1.1367276,1.3742256,1.1367276,0.89922947,0.66173136,0.42423326,0.18673515,0.21211663,0.2374981,0.26287958,0.28826106,0.31182957,0.34990177,0.387974,0.42423326,0.46230546,0.50037766,0.6000906,0.69980353,0.7995165,0.89922947,1.0007553,0.96268314,0.9246109,0.8883517,0.85027945,0.8122072,1.062396,1.3125849,1.5627737,1.8129625,2.0631514,2.3369088,2.612479,2.8880494,3.1618068,3.437377,3.4627585,3.48814,3.5117085,3.53709,3.5624714,4.175253,4.788034,5.4008155,6.011784,6.624565,8.200029,9.775495,11.349146,12.92461,14.500074,11.936545,9.374829,6.813113,4.249584,1.6878681,2.2118144,1.789394,1.3669738,0.9445535,0.52213323,0.099712946,0.0870222,0.07433146,0.06164073,0.05076295,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.85934424,1.7205015,2.5798457,3.43919,4.3003473,3.6694362,3.0403383,2.4094272,1.7803292,1.1494182,1.0569572,0.9644961,0.872035,0.7795739,0.6871128,2.5018883,4.3166637,6.1332526,7.948028,9.762803,8.520925,7.2772317,6.035352,4.7916603,3.5497808,3.3267863,3.105605,2.8826106,2.659616,2.4384346,2.08672,1.7368182,1.3869164,1.0370146,0.6871128,0.6417888,0.5982776,0.5529536,0.5076295,0.46230546,0.824898,1.1874905,1.550083,1.9126755,2.275268,5.709019,9.144584,12.580148,16.01571,19.449463,15.609608,11.769753,7.9298983,4.0900435,0.25018883,1.209246,2.1701162,3.1291735,4.0900435,5.049101,4.9802084,4.9095025,4.84061,4.7699046,4.699199,3.9105604,3.1201086,2.3296568,1.5392052,0.7505665,0.7324369,0.71430725,0.6979906,0.67986095,0.66173136,1.2019942,1.742257,2.2825198,2.8227828,3.3630457,5.23221,7.1031876,8.972352,10.843329,12.712494,13.062395,13.412297,13.762199,14.112101,14.462003,13.020698,11.5775795,10.13446,8.693155,7.250037,6.2257137,5.199577,4.175253,3.149116,2.124792,2.1501737,2.175555,2.2009366,2.2245052,2.2498865,2.0595255,1.8691645,1.6806163,1.4902552,1.2998942,1.1548572,1.0098201,0.86478317,0.7197462,0.5747091,0.54570174,0.5148814,0.48587397,0.4550536,0.42423326,0.47318324,0.52032024,0.56745726,0.61459434,0.66173136,0.63816285,0.61278135,0.5873999,0.5620184,0.53663695,0.50037766,0.46230546,0.42423326,0.387974,0.34990177,0.52032024,0.69073874,0.85934424,1.0297627,1.2001812,2.4076142,3.6150475,4.8224807,6.0299134,7.2373466,6.0770507,4.9167547,3.7582715,2.5979755,1.4376793,1.4195497,1.403233,1.3851035,1.3669738,1.3506571,1.3270886,1.305333,1.2817645,1.260009,1.2382535,1.1421664,1.0478923,0.95180535,0.8575313,0.76325727,0.65991837,0.55839247,0.4550536,0.35171473,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.15954071,0.21936847,0.27919623,0.34083697,0.40066472,0.78319985,1.1657349,1.54827,1.9308052,2.3133402,2.4148662,2.518205,2.619731,2.72307,2.8245957,2.427557,2.030518,1.6316663,1.2346275,0.8375887,0.678048,0.5166943,0.35715362,0.19761293,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.21574254,0.42967212,0.64541465,0.85934424,1.0750868,0.85934424,0.64541465,0.42967212,0.21574254,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.40066472,0.7995165,1.2001812,1.6008459,1.9996977,3.6549325,5.3101673,6.965402,8.620637,10.275872,10.303066,10.330261,10.357455,10.384649,10.411844,9.460039,8.508233,7.554615,6.60281,5.6491914,5.335549,5.0200934,4.704638,4.3891826,4.07554,5.317419,6.5592985,7.802991,9.04487,10.28675,10.319383,10.352016,10.384649,10.417283,10.449916,8.939718,7.4295206,5.919323,4.409125,2.9007401,6.202145,9.5053625,12.806767,16.109985,19.413204,16.92038,14.427556,11.934732,9.441909,6.9508986,9.452786,11.954676,14.458377,16.960264,19.462152,19.124943,18.787731,18.45052,18.11331,17.774284,15.332225,12.890164,10.448103,8.0060425,5.562169,9.724731,13.887294,18.049856,22.212418,26.374979,21.539808,16.704638,11.869466,7.036108,2.2009366,2.0595255,1.9199274,1.7803292,1.6407311,1.49932,1.2183108,0.9354887,0.6526665,0.36984438,0.0870222,0.07433146,0.06164073,0.05076295,0.038072214,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.2030518,0.38072214,0.55839247,0.73424983,0.9119202,0.823085,0.7324369,0.6417888,0.5529536,0.46230546,0.40972954,0.35715362,0.3045777,0.2520018,0.19942589,0.23205921,0.26469254,0.29732585,0.32995918,0.36259252,0.5873999,0.8122072,1.0370146,1.261822,1.4866294,1.35247,1.2183108,1.0823387,0.9481794,0.8122072,0.8430276,0.872035,0.90285534,0.9318628,0.96268314,0.8774739,0.79226464,0.7070554,0.62184614,0.53663695,0.6744221,0.8122072,0.9499924,1.0877775,1.2255627,1.2672608,1.310772,1.35247,1.3941683,1.4376793,1.6117238,1.7875811,1.9616255,2.137483,2.3133402,2.5979755,2.8826106,3.1672456,3.4518807,3.738329,3.7492065,3.7618973,3.774588,3.787279,3.7999697,4.2804046,4.76084,5.239462,5.719897,6.200332,7.5654926,8.930654,10.2958145,11.6591625,13.024323,10.798005,8.569874,6.341743,4.115425,1.887294,1.6751775,1.3542831,1.0352017,0.71430725,0.39522585,0.07433146,0.07433146,0.07433146,0.07433146,0.07433146,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.64541465,1.2908293,1.9344311,2.5798457,3.2252605,2.752077,2.280707,1.8075237,1.3343405,0.8629702,0.90285534,0.94274056,0.9826257,1.0225109,1.062396,4.7554007,8.446592,12.139598,15.8326025,19.525606,16.740896,13.954373,11.169662,8.384952,5.600241,5.4552045,5.3101673,5.1651306,5.0200934,4.8750563,4.175253,3.4754493,2.7756457,2.0758421,1.3742256,1.1983683,1.020698,0.8430276,0.6653573,0.48768693,0.8122072,1.1367276,1.4630609,1.7875811,2.1121013,4.606738,7.1031876,9.597824,12.092461,14.587097,11.708113,8.827314,5.9465175,3.0675328,0.18673515,0.90829426,1.6280404,2.3477864,3.0675328,3.787279,3.7347028,3.682127,3.6295512,3.576975,3.5243993,2.9333735,2.3405347,1.7476959,1.1548572,0.5620184,0.58921283,0.61822027,0.64541465,0.6726091,0.69980353,1.3669738,2.034144,2.7031271,3.3702974,4.0374675,5.328297,6.6173134,7.9081426,9.197159,10.487988,11.111648,11.73712,12.362592,12.988064,13.611723,12.340837,11.068136,9.795437,8.5227375,7.250037,6.5121617,5.774286,5.038223,4.3003473,3.5624714,3.7492065,3.9377546,4.12449,4.313038,4.499773,4.120864,3.7401419,3.3594196,2.9805105,2.5997884,2.3097143,2.0196402,1.7295663,1.4394923,1.1494182,1.0895905,1.0297627,0.969935,0.9101072,0.85027945,0.9445535,1.0406405,1.1349145,1.2291887,1.3252757,1.2745126,1.2255627,1.1747998,1.1258497,1.0750868,1.0007553,0.9246109,0.85027945,0.774135,0.69980353,1.0025684,1.305333,1.6080978,1.9108626,2.2118144,2.902553,3.5932918,4.2822175,4.972956,5.661882,4.804351,3.9468195,3.0892882,2.231757,1.3742256,1.4648738,1.5555218,1.6443571,1.7350051,1.8256533,1.8184015,1.8093367,1.8020848,1.794833,1.7875811,1.647983,1.5083848,1.3669738,1.2273756,1.0877775,0.969935,0.8520924,0.73424983,0.61822027,0.50037766,0.40066472,0.2991388,0.19942589,0.099712946,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.13234627,0.19036107,0.24837588,0.3045777,0.36259252,0.69073874,1.017072,1.3452182,1.6733645,1.9996977,2.2045624,2.4094272,2.6142921,2.819157,3.0258346,2.7557032,2.4855716,2.2154403,1.9453088,1.6751775,1.3542831,1.0352017,0.71430725,0.39522585,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.42967212,0.85934424,1.2908293,1.7205015,2.1501737,1.7205015,1.2908293,0.85934424,0.42967212,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.33721104,0.6744221,1.0116332,1.3506571,1.6878681,3.198066,4.708264,6.2166486,7.7268467,9.237044,9.180842,9.122828,9.064813,9.006798,8.950596,8.39583,7.83925,7.2844834,6.7297173,6.1749506,6.008158,5.8395524,5.67276,5.504154,5.337362,6.109684,6.882006,7.654328,8.42665,9.200785,9.189907,9.180842,9.169965,9.159087,9.1500225,8.01692,6.885632,5.75253,4.6194286,3.48814,6.0426044,8.597069,11.153346,13.70781,16.262274,14.677745,13.093216,11.506873,9.922344,8.337815,9.768243,11.1968565,12.627284,14.057712,15.488139,15.199879,14.911617,14.625169,14.336908,14.05046,12.427858,10.805257,9.182655,7.560054,5.9374523,9.188094,12.436923,15.687565,18.936394,22.187037,18.630003,15.072971,11.514126,7.957093,4.40006,4.120864,3.8398547,3.5606585,3.2796493,3.000453,2.4348087,1.8691645,1.305333,0.73968875,0.17585737,0.15047589,0.12509441,0.099712946,0.07433146,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.25562772,0.4604925,0.6653573,0.87022203,1.0750868,1.020698,0.9644961,0.9101072,0.8557183,0.7995165,0.7070554,0.61459434,0.52213323,0.42967212,0.33721104,0.3770962,0.4169814,0.45686656,0.49675176,0.53663695,0.7505665,0.96268314,1.1747998,1.3869164,1.6008459,1.5682126,1.5355793,1.502946,1.4703126,1.4376793,1.4721256,1.5083848,1.5428312,1.5772774,1.6117238,1.405046,1.1983683,0.9898776,0.78319985,0.5747091,0.7505665,0.9246109,1.1004683,1.2745126,1.4503701,1.5718386,1.69512,1.8184015,1.93987,2.0631514,2.1628644,2.2625773,2.3622901,2.4620032,2.561716,2.857229,3.152742,3.4482548,3.7419548,4.0374675,4.0374675,4.0374675,4.0374675,4.0374675,4.0374675,4.3855567,4.7318325,5.0799212,5.42801,5.774286,6.930956,8.0858135,9.24067,10.395528,11.5503845,9.657652,7.764919,5.8721857,3.9794528,2.08672,1.1367276,0.91917205,0.7016165,0.48587397,0.26831847,0.05076295,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.09064813,0.06707962,0.045324065,0.02175555,0.0,0.42967212,0.85934424,1.2908293,1.7205015,2.1501737,1.8347181,1.5192627,1.2056202,0.8901646,0.5747091,0.7469406,0.91917205,1.0932164,1.2654479,1.4376793,7.0071006,12.576522,18.147755,23.717176,29.286598,24.960869,20.633327,16.303972,11.978244,7.650702,7.5818095,7.51473,7.4476504,7.380571,7.311678,6.261973,5.2122674,4.162562,3.1128569,2.0631514,1.7531348,1.4431182,1.1331016,0.823085,0.51306844,0.7995165,1.0877775,1.3742256,1.6624867,1.9507477,3.5044568,5.0599785,6.6155005,8.1692095,9.724731,7.804804,5.8848767,3.9649491,2.0450218,0.12509441,0.6055295,1.0841516,1.5645868,2.0450218,2.525457,2.4891977,2.4547513,2.420305,2.3858588,2.3495996,1.9543737,1.5591478,1.1657349,0.7705091,0.37528324,0.44780177,0.52032024,0.59283876,0.6653573,0.73787576,1.5319533,2.327844,3.1219215,3.917812,4.7118897,5.422571,6.1332526,6.8421206,7.552802,8.26167,9.162713,10.061942,10.962985,11.862214,12.763257,11.6591625,10.556881,9.4546,8.352319,7.250037,6.8004227,6.350808,5.89938,5.4497657,5.0001507,5.3500524,5.6999545,6.049856,6.399758,6.7496595,6.1803894,5.6093063,5.040036,4.4707656,3.8996825,3.4645715,3.0294604,2.5943494,2.1592383,1.7241274,1.6352923,1.5446441,1.455809,1.3651608,1.2745126,1.4177368,1.5591478,1.7023718,1.845596,1.987007,1.9126755,1.8383441,1.7621996,1.6878681,1.6117238,1.49932,1.3869164,1.2745126,1.162109,1.0497054,1.4848163,1.9199274,2.3550384,2.7901495,3.2252605,3.397492,3.5697234,3.7419548,3.9141862,4.0882306,3.531651,2.9768846,2.422118,1.8673514,1.3125849,1.5101979,1.7078108,1.9054236,2.1030366,2.3006494,2.3079014,2.3151531,2.322405,2.3296568,2.3369088,2.1519866,1.9670644,1.7821422,1.5972201,1.4122978,1.2799516,1.1476053,1.015259,0.88291276,0.7505665,0.6000906,0.44961473,0.2991388,0.15047589,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.10515183,0.15954071,0.21574254,0.27013144,0.3245203,0.5982776,0.87022203,1.1421664,1.4141108,1.6878681,1.9942589,2.3024626,2.610666,2.9170568,3.2252605,3.0820365,2.9406252,2.7974012,2.6541772,2.5127661,2.032331,1.551896,1.0732739,0.59283876,0.11240368,0.09064813,0.06707962,0.045324065,0.02175555,0.0,0.64541465,1.2908293,1.9344311,2.5798457,3.2252605,2.5798457,1.9344311,1.2908293,0.64541465,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.2755703,0.5493277,0.824898,1.1004683,1.3742256,2.7393866,4.1045475,5.469708,6.834869,8.200029,8.056806,7.915395,7.7721705,7.6307597,7.4875355,7.3298078,7.17208,7.0143523,6.8566246,6.70071,6.680767,6.6608243,6.640882,6.6191263,6.599184,6.9019485,7.2047133,7.507478,7.8102427,8.113008,8.0604315,8.007855,7.95528,7.902704,7.850128,7.0941224,6.33993,5.5857377,4.8297324,4.07554,5.883064,7.690587,9.498111,11.3056345,13.113158,12.43511,11.757062,11.080828,10.40278,9.724731,10.081885,10.440851,10.798005,11.155159,11.512312,11.274815,11.037316,10.799818,10.56232,10.324821,9.52168,8.72035,7.9172077,7.115878,6.3127356,8.649645,10.986553,13.325275,15.662184,18.000906,15.720199,13.439491,11.160598,8.87989,6.599184,6.1803894,5.7597823,5.3391747,4.9203806,4.499773,3.6531196,2.8046532,1.9579996,1.1095331,0.26287958,0.22480737,0.18673515,0.15047589,0.11240368,0.07433146,0.07433146,0.07433146,0.07433146,0.07433146,0.07433146,0.30820364,0.5402629,0.77232206,1.0043813,1.2382535,1.2183108,1.1983683,1.1766127,1.1566701,1.1367276,1.0043813,0.872035,0.73968875,0.6073425,0.4749962,0.52213323,0.56927025,0.61822027,0.6653573,0.7124943,0.9119202,1.1131591,1.3125849,1.5120108,1.7132497,1.7821422,1.8528478,1.9217403,1.9924458,2.0631514,2.1030366,2.1429217,2.182807,2.222692,2.2625773,1.9326181,1.6026589,1.2726997,0.94274056,0.61278135,0.824898,1.0370146,1.2491312,1.4630609,1.6751775,1.8782293,2.079468,2.2825198,2.4855716,2.6868105,2.712192,2.7375734,2.762955,2.7883365,2.811905,3.1182957,3.4228733,3.727451,4.0320287,4.3366065,4.325729,4.313038,4.3003473,4.2876563,4.274966,4.4907084,4.704638,4.9203806,5.1343102,5.3500524,6.294606,7.2409725,8.185526,9.130079,10.074633,8.517298,6.9599633,5.4026284,3.8452935,2.2879589,0.6000906,0.48587397,0.36984438,0.25562772,0.13959812,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.21574254,0.42967212,0.64541465,0.85934424,1.0750868,0.91735905,0.75963134,0.60190356,0.44417584,0.28826106,0.59283876,0.8974165,1.2019942,1.5083848,1.8129625,9.2606125,16.70645,24.155914,31.603563,39.0494,33.18084,27.310469,21.440096,15.569723,9.699349,9.710228,9.719293,9.73017,9.739235,9.750113,8.350506,6.9508986,5.5494785,4.1498713,2.7502642,2.3079014,1.8655385,1.4231756,0.9808127,0.53663695,0.7868258,1.0370146,1.2872034,1.5373923,1.7875811,2.4021754,3.0167696,3.633177,4.2477713,4.8623657,3.9033084,2.9424384,1.9815681,1.0225109,0.06164073,0.30276474,0.5420758,0.78319985,1.0225109,1.261822,1.2455053,1.2273756,1.209246,1.1929294,1.1747998,0.97718686,0.7795739,0.581961,0.38434806,0.18673515,0.3045777,0.4224203,0.5402629,0.65810543,0.774135,1.696933,2.619731,3.5425289,4.465327,5.388125,5.516845,5.6473784,5.7779117,5.906632,6.037165,7.211965,8.386765,9.563377,10.738177,11.912977,10.979301,10.047439,9.115576,8.1819,7.250037,7.0868707,6.925517,6.7623506,6.599184,6.43783,6.9508986,7.462154,7.9752226,8.488291,8.999546,8.239915,7.4802837,6.720652,5.959208,5.199577,4.6194286,4.0392804,3.4591327,2.8807976,2.3006494,2.179181,2.0595255,1.93987,1.8202144,1.7005589,1.889107,2.079468,2.269829,2.4601903,2.6505513,2.5508385,2.4493124,2.3495996,2.2498865,2.1501737,1.9996977,1.8492218,1.7005589,1.550083,1.3996071,1.9670644,2.5345216,3.101979,3.6694362,4.2368937,3.8924308,3.5479677,3.2016919,2.857229,2.5127661,2.2607644,2.0069497,1.7549478,1.502946,1.2491312,1.5555218,1.8600996,2.1646774,2.469255,2.7756457,2.7974012,2.819157,2.8427253,2.864481,2.8880494,2.657803,2.427557,2.1973107,1.9670644,1.7368182,1.5899682,1.4431182,1.2944553,1.1476053,1.0007553,0.7995165,0.6000906,0.40066472,0.19942589,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.07795739,0.13053331,0.18310922,0.23568514,0.28826106,0.5058166,0.72337204,0.93911463,1.1566701,1.3742256,1.7857682,2.1954978,2.6052272,3.0149567,3.4246864,3.4101827,3.395679,3.3793623,3.3648586,3.350355,2.7103791,2.0704033,1.4304274,0.7904517,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.85934424,1.7205015,2.5798457,3.43919,4.3003473,3.43919,2.5798457,1.7205015,0.85934424,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.21211663,0.42423326,0.63816285,0.85027945,1.062396,2.2825198,3.5026438,4.7227674,5.942891,7.1630154,6.9345818,6.7079616,6.4795284,6.2529078,6.0244746,6.265599,6.5049095,6.7442207,6.985345,7.224656,7.3533764,7.4802837,7.607191,7.7359114,7.8628187,7.6942134,7.5274205,7.360628,7.192023,7.02523,6.929143,6.834869,6.740595,6.644508,6.550234,6.1731377,5.7942286,5.4171324,5.040036,4.6629395,5.7217097,6.782293,7.842876,8.901647,9.96223,10.192475,10.422722,10.652968,10.883214,11.111648,10.397341,9.683033,8.966913,8.252605,7.5382986,7.3497505,7.1630154,6.9744673,6.787732,6.599184,6.6173134,6.635443,6.6517596,6.6698895,6.688019,8.113008,9.537996,10.962985,12.387974,13.812962,12.810393,11.807825,10.805257,9.802689,8.80012,8.239915,7.6797094,7.119504,6.5592985,6.000906,4.8696175,3.7401419,2.610666,1.4793775,0.34990177,0.2991388,0.25018883,0.19942589,0.15047589,0.099712946,0.099712946,0.099712946,0.099712946,0.099712946,0.099712946,0.36077955,0.6200332,0.8792868,1.1403534,1.3996071,1.4141108,1.4304274,1.4449311,1.4594349,1.4757515,1.3017071,1.1294757,0.9572442,0.7850128,0.61278135,0.6671702,0.72337204,0.7777609,0.8321498,0.8883517,1.0750868,1.261822,1.4503701,1.6371052,1.8256533,1.9978848,2.1701162,2.3423476,2.514579,2.6868105,2.7321346,2.7774587,2.8227828,2.8681068,2.911618,2.4601903,2.0069497,1.5555218,1.1022812,0.6508536,0.89922947,1.1494182,1.3996071,1.649796,1.8999848,2.182807,2.465629,2.7466383,3.0294604,3.3122826,3.2633326,3.2125697,3.1618068,3.1128569,3.0620937,3.3775494,3.6930048,4.006647,4.322103,4.6375585,4.612177,4.5867953,4.5632267,4.537845,4.512464,4.59586,4.6774435,4.76084,4.842423,4.9258194,5.660069,6.394319,7.130382,7.8646317,8.600695,7.3769445,6.155008,4.933071,3.7093215,2.4873846,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.43692398,0.87566096,1.3125849,1.7495089,2.1882458,11.512312,20.836378,30.162258,39.488136,48.812206,41.400814,33.98761,26.574406,19.163015,11.74981,11.836833,11.925668,12.012691,12.099712,12.186734,10.437225,8.6877165,6.9382076,5.186886,3.437377,2.8626678,2.2879589,1.7132497,1.1367276,0.5620184,0.774135,0.9880646,1.2001812,1.4122978,1.6244144,1.2998942,0.97537386,0.6508536,0.3245203,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.16316663,0.3245203,0.48768693,0.6508536,0.8122072,1.8619126,2.911618,3.9631362,5.0128417,6.0625467,5.612932,5.163317,4.7118897,4.262275,3.8126602,5.2630305,6.7115874,8.161958,9.612328,11.062697,10.29944,9.537996,8.774739,8.013294,7.250037,7.3751316,7.500226,7.6253204,7.750415,7.8755093,8.549932,9.224354,9.900589,10.57501,11.249433,10.29944,9.349448,8.399456,7.4494634,6.4994707,5.774286,5.050914,4.325729,3.6005437,2.8753586,2.7248828,2.5744069,2.4257438,2.275268,2.124792,2.3622901,2.5997884,2.8372865,3.0747845,3.3122826,3.1871881,3.0620937,2.9369993,2.811905,2.6868105,2.5000753,2.3133402,2.124792,1.938057,1.7495089,2.4493124,3.149116,3.8507326,4.550536,5.2503395,4.3873696,3.5243993,2.663242,1.8002719,0.93730164,0.9880646,1.0370146,1.0877775,1.1367276,1.1874905,1.6008459,2.0123885,2.4257438,2.8372865,3.2506418,3.2869012,3.3249733,3.3630457,3.3993049,3.437377,3.1618068,2.8880494,2.612479,2.3369088,2.0631514,1.8999848,1.7368182,1.5754645,1.4122978,1.2491312,1.0007553,0.7505665,0.50037766,0.25018883,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,0.41335547,0.5747091,0.73787576,0.89922947,1.062396,1.5754645,2.08672,2.5997884,3.1128569,3.6241121,3.738329,3.8507326,3.9631362,4.07554,4.1879435,3.386614,2.5870976,1.7875811,0.9880646,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,1.0750868,2.1501737,3.2252605,4.3003473,5.375434,4.3003473,3.2252605,2.1501737,1.0750868,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.15047589,0.2991388,0.44961473,0.6000906,0.7505665,1.8256533,2.9007401,3.975827,5.050914,6.1241875,5.812358,5.5005283,5.186886,4.8750563,4.5632267,5.199577,5.8377395,6.4759026,7.112252,7.750415,8.024173,8.299743,8.575313,8.8508835,9.12464,8.488291,7.850128,7.211965,6.5756154,5.9374523,5.7996674,5.661882,5.524097,5.388125,5.2503395,5.2503395,5.2503395,5.2503395,5.2503395,5.2503395,5.562169,5.8758116,6.187641,6.4994707,6.813113,7.949841,9.086569,10.225109,11.361836,12.500377,10.712796,8.925215,7.137634,5.3500524,3.5624714,3.4246864,3.2869012,3.149116,3.0131438,2.8753586,3.7129474,4.550536,5.388125,6.2257137,7.063302,7.574558,8.087626,8.600695,9.11195,9.625018,9.900589,10.174346,10.449916,10.725487,10.999244,10.29944,9.599637,8.899834,8.200029,7.500226,6.0879283,4.6756306,3.2633326,1.8492218,0.43692398,0.37528324,0.31182957,0.25018883,0.18673515,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.41335547,0.69980353,0.9880646,1.2745126,1.5627737,1.6117238,1.6624867,1.7132497,1.7621996,1.8129625,1.6008459,1.3869164,1.1747998,0.96268314,0.7505665,0.8122072,0.87566096,0.93730164,1.0007553,1.062396,1.2382535,1.4122978,1.5881553,1.7621996,1.938057,2.2118144,2.4873846,2.762955,3.0367124,3.3122826,3.3630457,3.4119956,3.4627585,3.5117085,3.5624714,2.9877625,2.4130533,1.8383441,1.261822,0.6871128,0.97537386,1.261822,1.550083,1.8383441,2.124792,2.4873846,2.8499773,3.2125697,3.5751622,3.9377546,3.8126602,3.6875658,3.5624714,3.437377,3.3122826,3.636803,3.9631362,4.2876563,4.612177,4.936697,4.900438,4.8623657,4.8242936,4.788034,4.749962,4.699199,4.650249,4.599486,4.550536,4.499773,5.0255322,5.5494785,6.0752378,6.599184,7.124943,6.2365913,5.3500524,4.461701,3.5751622,2.6868105,0.42423326,0.4224203,0.42060733,0.4169814,0.41516843,0.41335547,0.43511102,0.45686656,0.48043507,0.50219065,0.52575916,0.45324063,0.38072214,0.30820364,0.23568514,0.16316663,0.13053331,0.09789998,0.065266654,0.032633327,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.40066472,0.73787576,1.0750868,1.4122978,1.7495089,9.229793,16.710075,24.19036,31.670643,39.149113,33.200783,27.25064,21.300497,15.350354,9.400211,9.469104,9.539809,9.610515,9.679407,9.750113,8.350506,6.9508986,5.5494785,4.1498713,2.7502642,2.5599031,2.3695421,2.179181,1.9906329,1.8002719,1.7603867,1.7205015,1.6806163,1.6407311,1.6008459,1.9543737,2.3097143,2.665055,3.0203958,3.3757362,3.0693457,2.764768,2.4601903,2.1556125,1.8492218,1.8619126,1.8746033,1.887294,1.8999848,1.9126755,1.6570477,1.403233,1.1476053,0.8919776,0.63816285,0.52032024,0.40247768,0.28463513,0.16679256,0.05076295,0.17041849,0.29007402,0.40972954,0.5293851,0.6508536,1.4902552,2.3296568,3.1708715,4.0102735,4.8496747,4.4907084,4.1299286,3.7691493,3.4101827,3.049403,4.209699,5.369995,6.530291,7.690587,8.849071,8.239915,7.6307597,7.019791,6.4106355,5.7996674,5.89938,5.999093,6.1006193,6.200332,6.300045,6.8421206,7.3841968,7.9280853,8.470161,9.012237,8.540867,8.067683,7.5945,7.12313,6.6499467,6.060734,5.469708,4.880495,4.2894692,3.7002566,3.531651,3.3648586,3.198066,3.0294604,2.8626678,2.8626678,2.8626678,2.8626678,2.8626678,2.8626678,2.7883365,2.712192,2.6378605,2.561716,2.4873846,2.2897718,2.0921588,1.8945459,1.696933,1.49932,2.0522738,2.6052272,3.1581807,3.7093215,4.262275,3.8543584,3.4482548,3.0403383,2.6324217,2.2245052,2.0504606,1.8746033,1.7005589,1.5247015,1.3506571,1.7404441,2.1302311,2.520018,2.909805,3.299592,3.199879,3.100166,3.000453,2.9007401,2.7992141,2.570781,2.3405347,2.1102884,1.8800422,1.649796,1.5228885,1.3941683,1.2672608,1.1403534,1.0116332,0.8122072,0.61278135,0.41335547,0.21211663,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.19942589,0.387974,0.5747091,0.76325727,0.9499924,0.76325727,0.5747091,0.387974,0.19942589,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.07977036,0.13415924,0.19036107,0.24474995,0.2991388,0.5058166,0.7106813,0.9155461,1.1204109,1.3252757,1.7023718,2.079468,2.4583774,2.8354735,3.2125697,3.339477,3.4681973,3.5951047,3.7220123,3.8507326,3.1219215,2.3949237,1.6679256,0.93911463,0.21211663,0.17223145,0.13234627,0.092461094,0.052575916,0.012690738,0.9354887,1.8582866,2.7792716,3.7020695,4.6248674,3.7727752,2.9206827,2.0667772,1.214685,0.36259252,0.30276474,0.24293698,0.18310922,0.12328146,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13053331,0.25925365,0.38978696,0.52032024,0.6508536,1.7041848,2.759329,3.8144734,4.8696175,5.924762,5.7470913,5.569421,5.391751,5.2158933,5.038223,5.6655083,6.2927933,6.9200783,7.5473633,8.174648,8.160145,8.145641,8.129324,8.1148205,8.100317,7.9244595,7.750415,7.574558,7.400513,7.224656,7.079619,6.9345818,6.789545,6.644508,6.4994707,6.4704633,6.439643,6.4106355,6.379815,6.350808,6.6082487,6.8656893,7.12313,7.380571,7.6380115,8.602508,9.567003,10.533313,11.497808,12.462305,10.939416,9.418341,7.895452,6.3725634,4.8496747,4.5432844,4.2350807,3.926877,3.6204863,3.3122826,3.9867048,4.6629395,5.337362,6.011784,6.688019,7.0850577,7.4820967,7.8791356,8.2779875,8.675026,8.709473,8.745731,8.780178,8.814624,8.849071,8.357758,7.8646317,7.3733187,6.880193,6.3870673,5.2865987,4.1879435,3.0874753,1.987007,0.8883517,0.7705091,0.6526665,0.53482395,0.4169814,0.2991388,0.26831847,0.23568514,0.2030518,0.17041849,0.13778515,0.37528324,0.61278135,0.85027945,1.0877775,1.3252757,1.357909,1.3905423,1.4231756,1.455809,1.4866294,1.3705997,1.2527572,1.1349145,1.017072,0.89922947,0.9572442,1.015259,1.0732739,1.1294757,1.1874905,1.2853905,1.3832904,1.4793775,1.5772774,1.6751775,1.9471219,2.220879,2.4928236,2.764768,3.0367124,3.147303,3.2578938,3.3666716,3.4772623,3.587853,3.0874753,2.5870976,2.08672,1.5881553,1.0877775,1.2672608,1.4467441,1.6280404,1.8075237,1.987007,2.277081,2.5671551,2.857229,3.147303,3.437377,3.3721104,3.3068438,3.24339,3.1781235,3.1128569,3.4591327,3.8072214,4.15531,4.501586,4.8496747,4.6828823,4.514277,4.347484,4.1806917,4.0120864,3.9903307,3.966762,3.9450066,3.923251,3.8996825,4.3547363,4.8097897,5.2648435,5.719897,6.1749506,5.529536,4.8841214,4.2405195,3.5951047,2.94969,0.7868258,0.79589057,0.8031424,0.8103943,0.81764615,0.824898,0.8321498,0.83940166,0.8466535,0.8557183,0.8629702,0.7541924,0.64722764,0.5402629,0.43329805,0.3245203,0.25925365,0.19579996,0.13053331,0.065266654,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.36259252,0.6000906,0.8375887,1.0750868,1.3125849,6.947273,12.581961,18.21846,23.85315,29.487837,25.000753,20.511858,16.024776,11.537694,7.0506115,7.1031876,7.155763,7.208339,7.2591023,7.311678,6.261973,5.2122674,4.162562,3.1128569,2.0631514,2.2571385,2.4529383,2.6469254,2.8427253,3.0367124,2.7448254,2.4529383,2.1592383,1.8673514,1.5754645,2.610666,3.6458678,4.6792564,5.714458,6.7496595,6.1405044,5.529536,4.9203806,4.309412,3.7002566,3.7256382,3.7492065,3.774588,3.7999697,3.825351,3.3159087,2.8046532,2.2952106,1.7857682,1.2745126,1.0406405,0.80495536,0.56927025,0.33539808,0.099712946,0.17767033,0.25562772,0.33177215,0.40972954,0.48768693,1.1167849,1.7476959,2.3767939,3.007705,3.636803,3.3666716,3.0983531,2.8282216,2.5580902,2.2879589,3.1581807,4.02659,4.896812,5.767034,6.637256,6.1803894,5.7217097,5.2648435,4.8079767,4.349297,4.4254417,4.499773,4.574105,4.650249,4.7245803,5.1343102,5.5458527,5.955582,6.3653116,6.775041,6.78048,6.784106,6.789545,6.794984,6.8004227,6.345369,5.8903155,5.4352617,4.9802084,4.5251546,4.3402324,4.15531,3.9703882,3.785466,3.6005437,3.3630457,3.1255474,2.8880494,2.6505513,2.4130533,2.3876717,2.3622901,2.3369088,2.3133402,2.2879589,2.079468,1.8727903,1.6642996,1.4576219,1.2491312,1.6552348,2.0595255,2.465629,2.8699198,3.2742105,3.3231604,3.3702974,3.4174345,3.4645715,3.5117085,3.1128569,2.712192,2.3133402,1.9126755,1.5120108,1.8800422,2.2480736,2.6142921,2.9823234,3.350355,3.1128569,2.8753586,2.6378605,2.4003625,2.1628644,1.9779422,1.79302,1.6080978,1.4231756,1.2382535,1.1457924,1.0533313,0.96087015,0.8665961,0.774135,0.62547207,0.4749962,0.3245203,0.17585737,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.40066472,0.774135,1.1494182,1.5247015,1.8999848,1.5247015,1.1494182,0.774135,0.40066472,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.11059072,0.17041849,0.23024625,0.29007402,0.34990177,0.5982776,0.8448406,1.0932164,1.3397794,1.5881553,1.8292793,2.0722163,2.3151531,2.5580902,2.7992141,2.9424384,3.0856624,3.2270734,3.3702974,3.5117085,2.857229,2.2027495,1.54827,0.8919776,0.2374981,0.19579996,0.15228885,0.11059072,0.06707962,0.025381476,0.79589057,1.5645868,2.335096,3.105605,3.874301,3.245203,2.6142921,1.9851941,1.3542831,0.72518504,0.6055295,0.48587397,0.36440548,0.24474995,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.11059072,0.21936847,0.32995918,0.4405499,0.5493277,1.5845293,2.619731,3.6549325,4.690134,5.7253356,5.6818247,5.6401267,5.5966153,5.5549173,5.5132194,6.1296263,6.7478466,7.364254,7.9824743,8.600695,8.294304,7.989726,7.6851482,7.380571,7.07418,7.362441,7.650702,7.93715,8.225411,8.511859,8.3595705,8.207282,8.054993,7.902704,7.750415,7.690587,7.6307597,7.569119,7.509291,7.4494634,7.652515,7.855567,8.056806,8.259857,8.46291,9.255174,10.047439,10.839704,11.631968,12.4242325,11.16785,9.909654,8.653271,7.3950744,6.1368785,5.660069,5.18326,4.704638,4.227829,3.7492065,4.262275,4.7753434,5.2884116,5.7996674,6.3127356,6.5955577,6.87838,7.159389,7.4422116,7.7250338,7.520169,7.315304,7.1104393,6.9055743,6.70071,6.414262,6.1296263,5.844991,5.560356,5.275721,4.4870825,3.7002566,2.911618,2.124792,1.3379664,1.1657349,0.9916905,0.8194591,0.64722764,0.4749962,0.40972954,0.3444629,0.27919623,0.21574254,0.15047589,0.33721104,0.52575916,0.7124943,0.89922947,1.0877775,1.1022812,1.1167849,1.1331016,1.1476053,1.162109,1.1403534,1.1167849,1.0950294,1.0732739,1.0497054,1.1022812,1.1548572,1.2074331,1.260009,1.3125849,1.3325275,1.35247,1.3724127,1.3923552,1.4122978,1.6824293,1.9525607,2.222692,2.4928236,2.762955,2.9333735,3.101979,3.2723975,3.442816,3.6132345,3.1871881,2.762955,2.3369088,1.9126755,1.4866294,1.5591478,1.6316663,1.7041848,1.7767034,1.8492218,2.0667772,2.2843328,2.5018883,2.7194438,2.9369993,2.9333735,2.9279346,2.9224956,2.9170568,2.911618,3.2832751,3.6531196,4.022964,4.3928084,4.762653,4.465327,4.168001,3.870675,3.5733492,3.2742105,3.2796493,3.2850883,3.290527,3.294153,3.299592,3.6857529,4.070101,4.454449,4.84061,5.224958,4.8224807,4.420003,4.017525,3.6150475,3.2125697,1.1494182,1.167548,1.1856775,1.2019942,1.2201238,1.2382535,1.2291887,1.2219368,1.214685,1.2074331,1.2001812,1.0569572,0.9155461,0.77232206,0.629098,0.48768693,0.38978696,0.291887,0.19579996,0.09789998,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.3245203,0.46230546,0.6000906,0.73787576,0.87566096,4.664753,8.455658,12.244749,16.035654,19.824745,16.800724,13.77489,10.749055,7.7250338,4.699199,4.7354584,4.7699046,4.804351,4.84061,4.8750563,4.175253,3.4754493,2.7756457,2.0758421,1.3742256,1.9543737,2.5345216,3.1146698,3.6948178,4.274966,3.729264,3.1853752,2.6396735,2.0957847,1.550083,3.2651455,4.9802084,6.695271,8.410334,10.125396,9.20985,8.294304,7.380571,6.4650245,5.5494785,5.5875506,5.6256227,5.661882,5.6999545,5.7380266,4.972956,4.207886,3.442816,2.6777458,1.9126755,1.5591478,1.2074331,0.8557183,0.50219065,0.15047589,0.18492219,0.21936847,0.25562772,0.29007402,0.3245203,0.7451276,1.1657349,1.5845293,2.0051367,2.4257438,2.2444477,2.0649643,1.8854811,1.7041848,1.5247015,2.1048496,2.6849976,3.2651455,3.8452935,4.4254417,4.120864,3.8144734,3.5098956,3.2053177,2.9007401,2.94969,3.000453,3.049403,3.100166,3.149116,3.4283123,3.7056956,3.9830787,4.2604623,4.537845,5.0200934,5.5023413,5.9845896,6.4668374,6.9508986,6.630004,6.3091097,5.9900284,5.669134,5.3500524,5.147001,4.945762,4.74271,4.539658,4.3366065,3.8616104,3.386614,2.911618,2.4366217,1.9616255,1.987007,2.0123885,2.03777,2.0631514,2.08672,1.8691645,1.651609,1.4358664,1.2183108,1.0007553,1.258196,1.5156367,1.7730774,2.030518,2.2879589,2.7901495,3.29234,3.7945306,4.2967215,4.800725,4.175253,3.5497808,2.9243085,2.3006494,1.6751775,2.0196402,2.3641033,2.7103791,3.054842,3.3993049,3.0258346,2.6505513,2.275268,1.8999848,1.5247015,1.3851035,1.2455053,1.1040943,0.9644961,0.824898,0.7668832,0.7106813,0.6526665,0.5946517,0.53663695,0.43692398,0.33721104,0.2374981,0.13778515,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.6000906,1.162109,1.7241274,2.2879589,2.8499773,2.2879589,1.7241274,1.162109,0.6000906,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.13959812,0.20486477,0.27013144,0.33539808,0.40066472,0.69073874,0.9808127,1.2708868,1.5591478,1.8492218,1.9579996,2.0649643,2.1719291,2.280707,2.3876717,2.5453994,2.7031271,2.8608549,3.0167696,3.1744974,2.5925364,2.0105755,1.4268016,0.8448406,0.26287958,0.21755551,0.17223145,0.12690738,0.08339628,0.038072214,0.6544795,1.2726997,1.8909199,2.5073273,3.1255474,2.7176309,2.3097143,1.9017978,1.4956942,1.0877775,0.90829426,0.726998,0.5475147,0.3680314,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.09064813,0.1794833,0.27013144,0.36077955,0.44961473,1.4648738,2.4801328,3.4953918,4.510651,5.524097,5.618371,5.710832,5.803293,5.8957543,5.9882154,6.5955577,7.2029004,7.8102427,8.417585,9.024928,8.430276,7.835624,7.2391596,6.644508,6.049856,6.8004227,7.549176,8.299743,9.050309,9.800876,9.639522,9.479981,9.32044,9.159087,8.999546,8.910711,8.820063,8.729415,8.640579,8.549932,8.696781,8.845445,8.992294,9.139144,9.287807,9.907841,10.527874,11.147907,11.7679405,12.387974,11.39447,10.40278,9.409276,8.417585,7.4258947,6.776854,6.1296263,5.482399,4.835171,4.1879435,4.537845,4.8877473,5.237649,5.5875506,5.9374523,6.104245,6.2728505,6.439643,6.6082487,6.775041,6.3308654,5.8848767,5.4407005,4.994712,4.550536,4.4725785,4.3946214,4.3166637,4.2405195,4.162562,3.6875658,3.2125697,2.7375734,2.2625773,1.7875811,1.5591478,1.3325275,1.1040943,0.8774739,0.6508536,0.5529536,0.4550536,0.35715362,0.25925365,0.16316663,0.2991388,0.43692398,0.5747091,0.7124943,0.85027945,0.8466535,0.8448406,0.8430276,0.83940166,0.8375887,0.9101072,0.9826257,1.0551442,1.1276628,1.2001812,1.2473183,1.2944553,1.3434052,1.3905423,1.4376793,1.3796645,1.3216497,1.2654479,1.2074331,1.1494182,1.4177368,1.6842422,1.9525607,2.220879,2.4873846,2.7176309,2.9478772,3.1781235,3.4083695,3.636803,3.2869012,2.9369993,2.5870976,2.2371957,1.887294,1.8528478,1.8165885,1.7821422,1.7476959,1.7132497,1.8582866,2.0033236,2.1483607,2.2933977,2.4366217,2.4928236,2.5472124,2.6016014,2.657803,2.712192,3.105605,3.4972048,3.8906176,4.2822175,4.6756306,4.2477713,3.8199122,3.392053,2.9641938,2.5381477,2.570781,2.6034143,2.6342347,2.666868,2.6995013,3.0149567,3.3304121,3.6458678,3.9595103,4.274966,4.115425,3.9558845,3.7945306,3.63499,3.4754493,1.5120108,1.5392052,1.5682126,1.5954071,1.6226015,1.649796,1.6280404,1.6044719,1.5827163,1.5591478,1.5373923,1.3597219,1.1820517,1.0043813,0.82671094,0.6508536,0.52032024,0.38978696,0.25925365,0.13053331,0.0,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,0.28826106,0.3245203,0.36259252,0.40066472,0.43692398,2.382233,4.327542,6.2728505,8.21816,10.161655,8.600695,7.037921,5.475147,3.9123733,2.3495996,2.3677292,2.3858588,2.4021754,2.420305,2.4366217,2.08672,1.7368182,1.3869164,1.0370146,0.6871128,1.651609,2.617918,3.5824142,4.5469103,5.5132194,4.7155156,3.917812,3.1201086,2.322405,1.5247015,3.919625,6.3145485,8.709473,11.104396,13.499319,12.279196,11.060884,9.840761,8.620637,7.400513,7.4494634,7.500226,7.549176,7.5999393,7.650702,6.630004,5.6093063,4.590421,3.5697234,2.5508385,2.079468,1.6099107,1.1403534,0.67079616,0.19942589,0.19217403,0.18492219,0.17767033,0.17041849,0.16316663,0.37165734,0.581961,0.79226464,1.0025684,1.2128719,1.1222239,1.0333886,0.94274056,0.8520924,0.76325727,1.0533313,1.3415923,1.6316663,1.9217403,2.2118144,2.0595255,1.9072367,1.7549478,1.6026589,1.4503701,1.4757515,1.49932,1.5247015,1.550083,1.5754645,1.7205015,1.8655385,2.0105755,2.1556125,2.3006494,3.2597067,4.220577,5.179634,6.1405044,7.0995617,6.9146395,6.7297173,6.544795,6.359873,6.1749506,5.955582,5.7344007,5.5150323,5.295664,5.0744824,4.361988,3.6494937,2.9369993,2.2245052,1.5120108,1.5881553,1.6624867,1.7368182,1.8129625,1.887294,1.6606737,1.4322405,1.2056202,0.97718686,0.7505665,0.85934424,0.969935,1.0805258,1.1893034,1.2998942,2.2571385,3.2143826,4.17344,5.130684,6.0879283,5.237649,4.3873696,3.53709,2.6868105,1.8383441,2.1592383,2.4819458,2.8046532,3.1273603,3.4500678,2.9369993,2.4257438,1.9126755,1.3996071,0.8883517,0.79226464,0.6979906,0.60190356,0.5076295,0.41335547,0.38978696,0.3680314,0.3444629,0.32270733,0.2991388,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.7995165,1.550083,2.3006494,3.049403,3.7999697,3.049403,2.3006494,1.550083,0.7995165,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.17041849,0.23931105,0.3100166,0.38072214,0.44961473,0.78319985,1.114972,1.4467441,1.7803292,2.1121013,2.084907,2.0577126,2.030518,2.0033236,1.9743162,2.1483607,2.3205922,2.4928236,2.665055,2.8372865,2.327844,1.8184015,1.3071461,0.79770356,0.28826106,0.23931105,0.19217403,0.14503701,0.09789998,0.05076295,0.5148814,0.9808127,1.4449311,1.9108626,2.374981,2.1900587,2.0051367,1.8202144,1.6352923,1.4503701,1.209246,0.969935,0.7306239,0.4894999,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07070554,0.13959812,0.21030366,0.27919623,0.34990177,1.3452182,2.3405347,3.3358512,4.329355,5.3246713,5.5531044,5.7797246,6.008158,6.2347784,6.4632115,7.059676,7.6579537,8.254418,8.852696,9.449161,8.564435,7.6797094,6.794984,5.910258,5.0255322,6.2384043,7.4494634,8.662335,9.875207,11.088079,10.919474,10.752681,10.585889,10.417283,10.25049,10.130835,10.009366,9.88971,9.770056,9.6504,9.742861,9.835322,9.927783,10.020245,10.112705,10.560507,11.008308,11.454298,11.9021,12.349901,11.622903,10.8959055,10.167094,9.440096,8.713099,7.895452,7.077806,6.26016,5.4425135,4.6248674,4.8134155,5.0001507,5.186886,5.375434,5.562169,5.614745,5.667321,5.719897,5.772473,5.825049,5.139749,4.454449,3.7691493,3.0856624,2.4003625,2.5290828,2.659616,2.7901495,2.9206827,3.049403,2.8880494,2.7248828,2.561716,2.4003625,2.2371957,1.9543737,1.6733645,1.3905423,1.1077201,0.824898,0.69436467,0.5656443,0.43511102,0.3045777,0.17585737,0.26287958,0.34990177,0.43692398,0.52575916,0.61278135,0.59283876,0.5728962,0.5529536,0.533011,0.51306844,0.67986095,0.8466535,1.015259,1.1820517,1.3506571,1.3923552,1.4358664,1.4775645,1.5192627,1.5627737,1.4268016,1.2926424,1.1566701,1.0225109,0.8883517,1.1530442,1.4177368,1.6824293,1.9471219,2.2118144,2.5018883,2.7919624,3.0820365,3.3721104,3.6621845,3.386614,3.1128569,2.8372865,2.561716,2.2879589,2.1447346,2.0033236,1.8600996,1.7168756,1.5754645,1.647983,1.7205015,1.79302,1.8655385,1.938057,2.0522738,2.1683033,2.2825198,2.3967366,2.5127661,2.9279346,3.343103,3.7582715,4.171627,4.5867953,4.0302157,3.4718235,2.9152439,2.3568513,1.8002719,1.8600996,1.9199274,1.9797552,2.039583,2.0994108,2.3441606,2.5907235,2.8354735,3.0802233,3.3249733,3.4083695,3.489953,3.5733492,3.6549325,3.738329,1.8746033,1.9126755,1.9507477,1.987007,2.0250793,2.0631514,2.0250793,1.987007,1.9507477,1.9126755,1.8746033,1.6624867,1.4503701,1.2382535,1.0243238,0.8122072,0.6508536,0.48768693,0.3245203,0.16316663,0.0,0.06164073,0.12509441,0.18673515,0.25018883,0.31182957,0.25018883,0.18673515,0.12509441,0.06164073,0.0,0.099712946,0.19942589,0.2991388,0.40066472,0.50037766,0.40066472,0.2991388,0.19942589,0.099712946,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.3506571,2.6995013,4.0501585,5.4008155,6.7496595,5.6999545,4.650249,3.6005437,2.5508385,1.49932,4.574105,7.650702,10.725487,13.800271,16.875055,15.350354,13.825653,12.299138,10.774437,9.249735,9.313189,9.374829,9.438283,9.499924,9.563377,8.287052,7.0125394,5.7380266,4.461701,3.1871881,2.5997884,2.0123885,1.4249886,0.8375887,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,1.49932,2.9369993,4.3746786,5.812358,7.250037,7.1992745,7.1503243,7.0995617,7.0506115,6.9998484,6.7623506,6.5248523,6.2873545,6.049856,5.812358,4.8623657,3.9123733,2.962381,2.0123885,1.062396,1.1874905,1.3125849,1.4376793,1.5627737,1.6878681,1.4503701,1.2128719,0.97537386,0.73787576,0.50037766,0.46230546,0.42423326,0.387974,0.34990177,0.31182957,1.7241274,3.1382382,4.550536,5.962834,7.3751316,6.300045,5.224958,4.1498713,3.0747845,1.9996977,2.3006494,2.5997884,2.9007401,3.199879,3.5008307,2.8499773,2.1991236,1.550083,0.89922947,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,1.0007553,1.938057,2.8753586,3.8126602,4.749962,3.8126602,2.8753586,1.938057,1.0007553,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.19942589,0.2755703,0.34990177,0.42423326,0.50037766,0.87566096,1.2491312,1.6244144,1.9996977,2.374981,2.2118144,2.0504606,1.887294,1.7241274,1.5627737,1.7495089,1.938057,2.124792,2.3133402,2.5000753,2.0631514,1.6244144,1.1874905,0.7505665,0.31182957,0.26287958,0.21211663,0.16316663,0.11240368,0.06164073,0.37528324,0.6871128,1.0007553,1.3125849,1.6244144,1.6624867,1.7005589,1.7368182,1.7748904,1.8129625,1.5120108,1.2128719,0.9119202,0.61278135,0.31182957,0.25018883,0.18673515,0.12509441,0.06164073,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,1.2255627,2.1991236,3.1744974,4.1498713,5.125245,5.487838,5.8504305,6.2130227,6.5756154,6.9382076,7.5256076,8.113008,8.700407,9.287807,9.875207,8.700407,7.5256076,6.350808,5.1741953,3.9993954,5.674573,7.3497505,9.024928,10.700105,12.375282,12.199425,12.025381,11.849524,11.675479,11.499621,11.349146,11.200482,11.050007,10.899531,10.750868,10.7871275,10.825199,10.863272,10.899531,10.937603,11.213174,11.486931,11.762501,12.038072,12.311829,11.849524,11.3872175,10.924912,10.462607,10.000301,9.012237,8.024173,7.037921,6.049856,5.0617914,5.087173,5.1125546,5.137936,5.163317,5.186886,5.125245,5.0617914,5.0001507,4.936697,4.8750563,3.9504454,3.0258346,2.0994108,1.1747998,0.25018883,0.5873999,0.9246109,1.261822,1.6008459,1.938057,2.08672,2.2371957,2.3876717,2.5381477,2.6868105,2.3495996,2.0123885,1.6751775,1.3379664,1.0007553,0.8375887,0.6744221,0.51306844,0.34990177,0.18673515,0.22480737,0.26287958,0.2991388,0.33721104,0.37528324,0.33721104,0.2991388,0.26287958,0.22480737,0.18673515,0.44961473,0.7124943,0.97537386,1.2382535,1.49932,1.5373923,1.5754645,1.6117238,1.649796,1.6878681,1.4757515,1.261822,1.0497054,0.8375887,0.62547207,0.8883517,1.1494182,1.4122978,1.6751775,1.938057,2.2879589,2.6378605,2.9877625,3.3376641,3.6875658,3.48814,3.2869012,3.0874753,2.8880494,2.6868105,2.4366217,2.1882458,1.938057,1.6878681,1.4376793,1.4376793,1.4376793,1.4376793,1.4376793,1.4376793,1.6117238,1.7875811,1.9616255,2.137483,2.3133402,2.7502642,3.1871881,3.6241121,4.062849,4.499773,3.8126602,3.1255474,2.4366217,1.7495089,1.062396,1.1494182,1.2382535,1.3252757,1.4122978,1.49932,1.6751775,1.8492218,2.0250793,2.1991236,2.374981,2.6995013,3.0258346,3.350355,3.6748753,3.9993954,1.6117238,1.6824293,1.7531348,1.8220274,1.892733,1.9616255,1.9906329,2.0178273,2.0450218,2.0722163,2.0994108,1.9054236,1.7096237,1.5156367,1.3198367,1.1258497,0.9318628,0.73968875,0.5475147,0.35534066,0.16316663,0.23205921,0.30276474,0.37165734,0.44236287,0.51306844,0.40972954,0.30820364,0.20486477,0.10333887,0.0,0.07977036,0.15954071,0.23931105,0.3208944,0.40066472,0.3444629,0.29007402,0.23568514,0.1794833,0.12509441,0.36984438,0.61459434,0.85934424,1.1059072,1.3506571,1.3125849,1.2745126,1.2382535,1.2001812,1.162109,2.030518,2.8971143,3.7655232,4.632119,5.5005283,4.7155156,3.930503,3.1454902,2.3604772,1.5754645,4.227829,6.880193,9.5325575,12.184921,14.837286,13.3506565,11.862214,10.375585,8.887142,7.400513,7.4494634,7.500226,7.549176,7.5999393,7.650702,6.6608243,5.669134,4.6792564,3.6893787,2.6995013,2.2027495,1.7041848,1.2074331,0.7106813,0.21211663,0.17223145,0.13234627,0.092461094,0.052575916,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.072518505,0.14503701,0.21755551,0.29007402,0.36259252,0.3770962,0.3934129,0.40791658,0.4224203,0.43692398,0.36440548,0.291887,0.21936847,0.14684997,0.07433146,1.2201238,2.3641033,3.5098956,4.655688,5.7996674,5.7597823,5.719897,5.6800117,5.6401267,5.600241,5.411693,5.224958,5.038223,4.8496747,4.6629395,4.2006345,3.738329,3.2742105,2.811905,2.3495996,2.47832,2.6052272,2.7321346,2.8608549,2.9877625,2.9478772,2.907992,2.8681068,2.8282216,2.7883365,2.5580902,2.327844,2.0975976,1.8673514,1.6371052,2.7557032,3.872488,4.989273,6.107871,7.224656,6.104245,4.985647,3.8652363,2.7448254,1.6244144,1.8600996,2.0957847,2.3296568,2.565342,2.7992141,2.280707,1.7603867,1.2400664,0.7197462,0.19942589,0.15954071,0.11965553,0.07977036,0.03988518,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.16679256,0.28463513,0.40247768,0.52032024,0.63816285,0.95180535,1.2672608,1.5827163,1.8981718,2.2118144,2.2426348,2.2734551,2.3024626,2.333283,2.3622901,2.6233568,2.8826106,3.141864,3.4029307,3.6621845,3.1799364,2.6976883,2.2154403,1.7331922,1.2491312,1.0098201,0.7705091,0.5293851,0.29007402,0.05076295,0.047137026,0.045324065,0.04169814,0.03988518,0.038072214,0.08520924,0.13234627,0.1794833,0.22662032,0.2755703,0.36077955,0.44417584,0.5293851,0.61459434,0.69980353,0.58014804,0.4604925,0.34083697,0.21936847,0.099712946,0.099712946,0.099712946,0.099712946,0.099712946,0.099712946,0.83940166,1.5790904,2.3205922,3.0602808,3.7999697,3.049403,2.3006494,1.550083,0.7995165,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.027194439,0.054388877,0.08339628,0.11059072,0.13778515,0.25562772,0.37165734,0.4894999,0.6073425,0.72518504,1.0279498,1.3307146,1.6316663,1.9344311,2.2371957,2.0957847,1.9525607,1.8093367,1.6679256,1.5247015,1.9579996,2.3894846,2.8227828,3.254268,3.6875658,3.007705,2.327844,1.647983,0.968122,0.28826106,0.26469254,0.24293698,0.21936847,0.19761293,0.17585737,0.48224804,0.7904517,1.0968424,1.405046,1.7132497,1.7150626,1.7168756,1.7205015,1.7223145,1.7241274,1.551896,1.3796645,1.2074331,1.0352017,0.8629702,0.7306239,0.5982776,0.46411842,0.33177215,0.19942589,0.15954071,0.11965553,0.07977036,0.03988518,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.25018883,0.50037766,0.7505665,1.0007553,1.2491312,2.0142014,2.7792716,3.5443418,4.309412,5.0744824,5.5095935,5.9447045,6.379815,6.814926,7.250037,7.931711,8.615198,9.296872,9.980359,10.662033,9.980359,9.296872,8.615198,7.931711,7.250037,8.482852,9.715667,10.948481,12.179482,13.412297,12.928236,12.442362,11.958302,11.472427,10.988366,11.392657,11.7969475,12.203052,12.607342,13.013446,12.589212,12.166792,11.744371,11.321951,10.899531,10.854207,10.810696,10.765372,10.720048,10.674724,10.4045925,10.13446,9.864329,9.594198,9.325879,8.582565,7.83925,7.0977483,6.354434,5.612932,6.1205616,6.628191,7.135821,7.6416373,8.149267,7.6833353,7.215591,6.7478466,6.2801023,5.812358,4.947575,4.082792,3.2180085,2.3532255,1.4866294,1.647983,1.8075237,1.9670644,2.126605,2.2879589,2.7683938,3.247016,3.727451,4.207886,4.688321,4.2477713,3.8072214,3.3666716,2.9279346,2.4873846,2.1900587,1.892733,1.5954071,1.2980812,1.0007553,0.86478317,0.7306239,0.5946517,0.4604925,0.3245203,0.33539808,0.3444629,0.35534066,0.36440548,0.37528324,0.58921283,0.80495536,1.020698,1.2346275,1.4503701,1.4576219,1.4648738,1.4721256,1.4793775,1.4866294,1.305333,1.1222239,0.93911463,0.75781834,0.5747091,0.8430276,1.1095331,1.3778516,1.6443571,1.9126755,2.1773682,2.4420607,2.7067533,2.9732587,3.2379513,3.149116,3.0620937,2.9750717,2.8880494,2.7992141,2.610666,2.420305,2.229944,2.039583,1.8492218,1.7857682,1.7205015,1.6552348,1.5899682,1.5247015,1.6769904,1.8292793,1.983381,2.13567,2.2879589,2.5979755,2.907992,3.2180085,3.5280252,3.8380418,3.2869012,2.7375734,2.1882458,1.6371052,1.0877775,1.1548572,1.2219368,1.2908293,1.357909,1.4249886,1.6153497,1.8057107,1.9942589,2.18462,2.374981,2.5798457,2.7847104,2.9895754,3.1944401,3.3993049,1.3506571,1.452183,1.5555218,1.6570477,1.7603867,1.8619126,1.9543737,2.0468347,2.1392958,2.231757,2.324218,2.1483607,1.9706904,1.79302,1.6153497,1.4376793,1.214685,0.9916905,0.7705091,0.5475147,0.3245203,0.40247768,0.48043507,0.55839247,0.6345369,0.7124943,0.56927025,0.42785916,0.28463513,0.14322405,0.0,0.059827764,0.11965553,0.1794833,0.23931105,0.2991388,0.29007402,0.27919623,0.27013144,0.25925365,0.25018883,0.73968875,1.2291887,1.7205015,2.2100015,2.6995013,2.6251698,2.5508385,2.474694,2.4003625,2.324218,2.7103791,3.094727,3.4808881,3.8652363,4.249584,3.729264,3.2107568,2.6904364,2.1701162,1.649796,3.87974,6.109684,8.339628,10.5695715,12.799516,11.349146,9.900589,8.450218,6.9998484,5.5494785,5.5875506,5.6256227,5.661882,5.6999545,5.7380266,5.032784,4.327542,3.6222992,2.9170568,2.2118144,1.8057107,1.3977941,0.9898776,0.581961,0.17585737,0.14503701,0.11421664,0.08520924,0.054388877,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14503701,0.29007402,0.43511102,0.58014804,0.72518504,0.7541924,0.7850128,0.81583315,0.8448406,0.87566096,0.7179332,0.56020546,0.40247768,0.24474995,0.0870222,0.93911463,1.79302,2.6451125,3.4972048,4.349297,4.3202896,4.2894692,4.2604623,4.229642,4.2006345,4.062849,3.925064,3.787279,3.6494937,3.5117085,3.53709,3.5624714,3.587853,3.6132345,3.636803,3.7673361,3.8978696,4.028403,4.157123,4.2876563,4.445384,4.603112,4.76084,4.9167547,5.0744824,4.652062,4.229642,3.8072214,3.3848011,2.962381,3.785466,4.606738,5.429823,6.2529078,7.07418,5.910258,4.744523,3.5806012,2.4148662,1.2491312,1.4195497,1.5899682,1.7603867,1.9308052,2.0994108,1.7096237,1.3198367,0.9300498,0.5402629,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.27194437,0.5076295,0.7433147,0.97718686,1.2128719,1.8546607,2.4982624,3.1400511,3.7818398,4.4254417,4.4852695,4.5450974,4.604925,4.664753,4.7245803,5.2449007,5.765221,6.285541,6.8058615,7.324369,6.359873,5.3953767,4.4308805,3.4645715,2.5000753,2.0196402,1.5392052,1.0605831,0.58014804,0.099712946,0.09427405,0.09064813,0.08520924,0.07977036,0.07433146,0.17041849,0.26469254,0.36077955,0.4550536,0.5493277,0.7197462,0.8901646,1.0605831,1.2291887,1.3996071,1.1602961,0.91917205,0.67986095,0.4405499,0.19942589,0.18673515,0.17585737,0.16316663,0.15047589,0.13778515,0.67986095,1.2219368,1.7658255,2.3079014,2.8499773,2.2879589,1.7241274,1.162109,0.6000906,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.3100166,0.46955732,0.630911,0.7904517,0.9499924,1.1802386,1.4104849,1.6407311,1.8691645,2.0994108,1.9779422,1.8546607,1.7331922,1.6099107,1.4866294,2.1646774,2.8427253,3.5207734,4.1970086,4.8750563,3.9522583,3.0294604,2.1066625,1.1856775,0.26287958,0.26831847,0.27194437,0.27738327,0.28282216,0.28826106,0.58921283,0.8919776,1.1947423,1.4975071,1.8002719,1.7676386,1.7350051,1.7023718,1.6697385,1.6371052,1.5917811,1.54827,1.502946,1.4576219,1.4122978,1.209246,1.0080072,0.80495536,0.60190356,0.40066472,0.3208944,0.23931105,0.15954071,0.07977036,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.44961473,0.89922947,1.3506571,1.8002719,2.2498865,2.8046532,3.3594196,3.9141862,4.4707656,5.0255322,5.5331616,6.0407915,6.548421,7.0542374,7.5618668,8.339628,9.117389,9.89515,10.672911,11.450671,11.26031,11.069949,10.879588,10.689227,10.500679,11.289318,12.07977,12.870221,13.660673,14.449312,13.655234,12.859344,12.065266,11.269376,10.475298,11.434355,12.395226,13.354282,14.315152,15.27421,14.39311,13.510198,12.627284,11.744371,10.863272,10.497053,10.1326475,9.768243,9.402024,9.037619,8.9596615,8.881703,8.805559,8.727602,8.649645,8.152893,7.654328,7.157576,6.6608243,6.16226,7.1521373,8.1420145,9.131892,10.12177,11.111648,10.239613,9.367578,8.495543,7.6216946,6.7496595,5.9447045,5.139749,4.3347936,3.529838,2.7248828,2.7067533,2.6904364,2.6723068,2.6541772,2.6378605,3.4482548,4.256836,5.06723,5.8776245,6.688019,6.14413,5.6020546,5.0599785,4.517903,3.975827,3.5425289,3.1092308,2.6777458,2.2444477,1.8129625,1.504759,1.1983683,0.8901646,0.581961,0.2755703,0.33177215,0.38978696,0.44780177,0.5058166,0.5620184,0.7306239,0.8974165,1.064209,1.2328146,1.3996071,1.3778516,1.3542831,1.3325275,1.310772,1.2872034,1.1349145,0.9826257,0.83033687,0.678048,0.52575916,0.79770356,1.0696479,1.3434052,1.6153497,1.887294,2.0667772,2.2480736,2.427557,2.6070402,2.7883365,2.811905,2.8372865,2.8626678,2.8880494,2.911618,2.7828975,2.6523643,2.521831,2.3931105,2.2625773,2.132044,2.0033236,1.8727903,1.742257,1.6117238,1.742257,1.8727903,2.0033236,2.132044,2.2625773,2.4456866,2.6269827,2.810092,2.9932013,3.1744974,2.762955,2.3495996,1.938057,1.5247015,1.1131591,1.1602961,1.2074331,1.2545701,1.3017071,1.3506571,1.5555218,1.7603867,1.9652514,2.1701162,2.374981,2.4601903,2.5453994,2.6306088,2.715818,2.7992141,1.0877775,1.2219368,1.357909,1.4920682,1.6280404,1.7621996,1.9199274,2.077655,2.2353828,2.3931105,2.5508385,2.3894846,2.229944,2.0704033,1.9108626,1.7495089,1.4975071,1.2455053,0.9916905,0.73968875,0.48768693,0.5728962,0.65810543,0.7433147,0.82671094,0.9119202,0.7306239,0.5475147,0.36440548,0.18310922,0.0,0.03988518,0.07977036,0.11965553,0.15954071,0.19942589,0.23568514,0.27013144,0.3045777,0.34083697,0.37528324,1.1095331,1.845596,2.5798457,3.3159087,4.0501585,3.9377546,3.825351,3.7129474,3.6005437,3.48814,3.39024,3.29234,3.1944401,3.0983531,3.000453,2.7448254,2.4891977,2.2353828,1.9797552,1.7241274,3.531651,5.3391747,7.1466985,8.954222,10.761745,9.349448,7.93715,6.5248523,5.1125546,3.7002566,3.7256382,3.7492065,3.774588,3.7999697,3.825351,3.4047437,2.9841363,2.565342,2.1447346,1.7241274,1.4068589,1.0895905,0.77232206,0.4550536,0.13778515,0.11784257,0.09789998,0.07795739,0.058014803,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.21755551,0.43511102,0.6526665,0.87022203,1.0877775,1.1331016,1.1766127,1.2219368,1.2672608,1.3125849,1.0696479,0.82671094,0.5855869,0.34264994,0.099712946,0.65991837,1.2201238,1.7803292,2.3405347,2.9007401,2.8807976,2.8608549,2.8409123,2.819157,2.7992141,2.712192,2.6251698,2.5381477,2.4493124,2.3622901,2.8753586,3.386614,3.8996825,4.4127507,4.9258194,5.0581656,5.1905117,5.3228583,5.4552045,5.5875506,5.942891,6.298232,6.6517596,7.0071006,7.362441,6.7478466,6.1332526,5.516845,4.902251,4.2876563,4.8152285,5.3428006,5.870373,6.397945,6.925517,5.714458,4.505212,3.294153,2.084907,0.87566096,0.9808127,1.0841516,1.1893034,1.2944553,1.3996071,1.1403534,0.8792868,0.6200332,0.36077955,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.3770962,0.7306239,1.0823387,1.4358664,1.7875811,2.7575161,3.727451,4.6973863,5.667321,6.637256,6.7279043,6.816739,6.9073873,6.9980354,7.0868707,7.8682575,8.647832,9.427405,10.20698,10.988366,9.539809,8.093065,6.644508,5.197764,3.7492065,3.0294604,2.3097143,1.5899682,0.87022203,0.15047589,0.14322405,0.13415924,0.12690738,0.11965553,0.11240368,0.25562772,0.39703882,0.5402629,0.68167394,0.824898,1.0805258,1.3343405,1.5899682,1.845596,2.0994108,1.7404441,1.3796645,1.020698,0.65991837,0.2991388,0.2755703,0.25018883,0.22480737,0.19942589,0.17585737,0.52032024,0.86478317,1.209246,1.5555218,1.8999848,1.5247015,1.1494182,0.774135,0.40066472,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.032633327,0.065266654,0.09789998,0.13053331,0.16316663,0.36440548,0.56745726,0.7705091,0.97174793,1.1747998,1.3325275,1.4902552,1.647983,1.8057107,1.9616255,1.8600996,1.7567607,1.6552348,1.551896,1.4503701,2.373168,3.294153,4.216951,5.139749,6.0625467,4.896812,3.73289,2.5671551,1.403233,0.2374981,0.27013144,0.30276474,0.33539808,0.3680314,0.40066472,0.6979906,0.99531645,1.2926424,1.5899682,1.887294,1.8202144,1.7531348,1.6842422,1.6171626,1.550083,1.6316663,1.7150626,1.7966459,1.8800422,1.9616255,1.6896812,1.4177368,1.1457924,0.872035,0.6000906,0.48043507,0.36077955,0.23931105,0.11965553,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.6508536,1.2998942,1.9507477,2.5997884,3.2506418,3.5951047,3.9395678,4.2858434,4.6303062,4.974769,5.5549173,6.1350656,6.7152133,7.2953615,7.8755093,8.747544,9.619579,10.493427,11.365462,12.237497,12.540262,12.843027,13.145792,13.446743,13.749508,14.097597,14.445685,14.791962,15.140051,15.488139,14.382232,13.278138,12.172231,11.068136,9.96223,11.477866,12.99169,14.507326,16.022963,17.536787,16.195194,14.851789,13.510198,12.166792,10.825199,10.139899,9.4546,8.7693,8.0858135,7.400513,7.51473,7.6307597,7.744976,7.859193,7.9752226,7.723221,7.4694057,7.217404,6.965402,6.7134004,8.185526,9.657652,11.129777,12.601903,14.075842,12.797703,11.519565,10.243238,8.9651,7.686961,6.9418335,6.1967063,5.4515786,4.708264,3.9631362,3.7673361,3.5733492,3.3775494,3.1817493,2.9877625,4.1281157,5.2666564,6.4070096,7.5473633,8.6877165,8.042302,7.3968873,6.7532854,6.107871,5.462456,4.894999,4.327542,3.7600844,3.1926272,2.6251698,2.1447346,1.6642996,1.1856775,0.70524246,0.22480737,0.32995918,0.43511102,0.5402629,0.64541465,0.7505665,0.87022203,0.9898776,1.1095331,1.2291887,1.3506571,1.2980812,1.2455053,1.1929294,1.1403534,1.0877775,0.9644961,0.8430276,0.7197462,0.5982776,0.4749962,0.7523795,1.0297627,1.3071461,1.5845293,1.8619126,1.9579996,2.0522738,2.1483607,2.2426348,2.3369088,2.474694,2.612479,2.7502642,2.8880494,3.0258346,2.955129,2.8844235,2.8155308,2.7448254,2.6741197,2.4801328,2.2843328,2.0903459,1.8945459,1.7005589,1.8075237,1.9144884,2.0232663,2.1302311,2.2371957,2.2933977,2.3477864,2.4021754,2.4583774,2.5127661,2.2371957,1.9616255,1.6878681,1.4122978,1.1367276,1.1657349,1.1929294,1.2201238,1.2473183,1.2745126,1.4956942,1.7150626,1.9344311,2.1556125,2.374981,2.3405347,2.3042755,2.269829,2.2353828,2.1991236,0.824898,0.9916905,1.1602961,1.3270886,1.4956942,1.6624867,1.8854811,2.1066625,2.3296568,2.5526514,2.7756457,2.6324217,2.4891977,2.3477864,2.2045624,2.0631514,1.7803292,1.4975071,1.214685,0.9318628,0.6508536,0.7433147,0.83577573,0.92823684,1.020698,1.1131591,0.8901646,0.6671702,0.44417584,0.2229944,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.1794833,0.25925365,0.34083697,0.42060733,0.50037766,1.4793775,2.4601903,3.43919,4.420003,5.4008155,5.2503395,5.0998635,4.949388,4.800725,4.650249,4.070101,3.489953,2.909805,2.3296568,1.7495089,1.7603867,1.7694515,1.7803292,1.789394,1.8002719,3.1853752,4.5704784,5.955582,7.3406854,8.725789,7.3497505,5.975525,4.599486,3.2252605,1.8492218,1.8619126,1.8746033,1.887294,1.8999848,1.9126755,1.7767034,1.6425442,1.5083848,1.3724127,1.2382535,1.0098201,0.78319985,0.55476654,0.32814622,0.099712946,0.09064813,0.07977036,0.07070554,0.059827764,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.29007402,0.58014804,0.87022203,1.1602961,1.4503701,1.5101979,1.5700256,1.6298534,1.6896812,1.7495089,1.4231756,1.0950294,0.7668832,0.4405499,0.11240368,0.38072214,0.64722764,0.9155461,1.1820517,1.4503701,1.4394923,1.4304274,1.4195497,1.4104849,1.3996071,1.3633479,1.3252757,1.2872034,1.2491312,1.2128719,2.2118144,3.2125697,4.213325,5.2122674,6.2130227,6.347182,6.4831543,6.6173134,6.7532854,6.887445,7.440398,7.993352,8.544493,9.097446,9.6504,8.841819,8.03505,7.228282,6.4197006,5.612932,5.844991,6.0770507,6.3091097,6.542982,6.775041,5.520471,4.265901,3.009518,1.7549478,0.50037766,0.5402629,0.58014804,0.6200332,0.65991837,0.69980353,0.56927025,0.4405499,0.3100166,0.1794833,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.48224804,0.95180535,1.4231756,1.892733,2.3622901,3.6603715,4.95664,6.2547207,7.552802,8.8508835,8.970539,9.090195,9.20985,9.329506,9.449161,10.489801,11.530442,12.569269,13.60991,14.650551,12.719746,10.790753,8.859948,6.929143,5.0001507,4.0392804,3.0802233,2.1193533,1.1602961,0.19942589,0.19036107,0.1794833,0.17041849,0.15954071,0.15047589,0.34083697,0.5293851,0.7197462,0.9101072,1.1004683,1.4394923,1.7803292,2.1193533,2.4601903,2.7992141,2.3205922,1.840157,1.3597219,0.8792868,0.40066472,0.36259252,0.3245203,0.28826106,0.25018883,0.21211663,0.36077955,0.5076295,0.6544795,0.8031424,0.9499924,0.76325727,0.5747091,0.387974,0.19942589,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.034446288,0.07070554,0.10515183,0.13959812,0.17585737,0.42060733,0.6653573,0.9101072,1.1548572,1.3996071,1.4848163,1.5700256,1.6552348,1.7404441,1.8256533,1.742257,1.6606737,1.5772774,1.4956942,1.4122978,2.5798457,3.7473936,4.914942,6.0824895,7.250037,5.8431783,4.4345064,3.0276475,1.6207886,0.21211663,0.27194437,0.33177215,0.39159992,0.45324063,0.51306844,0.80495536,1.0968424,1.3905423,1.6824293,1.9743162,1.8727903,1.7694515,1.6679256,1.5645868,1.4630609,1.6733645,1.8818551,2.0921588,2.3024626,2.5127661,2.1701162,1.8274662,1.4848163,1.1421664,0.7995165,0.6399758,0.48043507,0.3208944,0.15954071,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.85027945,1.7005589,2.5508385,3.3993049,4.249584,4.3855567,4.519716,4.655688,4.7898474,4.9258194,5.576673,6.2293396,6.882006,7.5346723,8.187339,9.155461,10.12177,11.089892,12.058014,13.024323,13.820213,14.614291,15.410182,16.20426,17.00015,16.905876,16.80979,16.715515,16.619429,16.525154,15.10923,13.695119,12.279196,10.865085,9.449161,11.519565,13.589968,15.660371,17.730774,19.799364,17.99728,16.195194,14.39311,12.589212,10.7871275,9.782746,8.778365,7.7721705,6.7677894,5.7615952,6.069799,6.378002,6.684393,6.9925966,7.3008003,7.2917356,7.2844834,7.2772317,7.26998,7.262728,9.217102,11.173288,13.127662,15.082036,17.038223,15.355793,13.673364,11.989121,10.308505,8.624263,7.9407763,7.2554765,6.5701766,5.8848767,5.199577,4.8279195,4.454449,4.082792,3.7093215,3.3376641,4.8079767,6.2782893,7.746789,9.217102,10.687414,9.940474,9.19172,8.444779,7.6978393,6.9508986,6.247469,5.5458527,4.842423,4.1408067,3.437377,2.7847104,2.132044,1.4793775,0.82671094,0.17585737,0.32814622,0.48043507,0.6327239,0.7850128,0.93730164,1.0098201,1.0823387,1.1548572,1.2273756,1.2998942,1.2183108,1.1349145,1.0533313,0.969935,0.8883517,0.79589057,0.7016165,0.6091554,0.5166943,0.42423326,0.7070554,0.9898776,1.2726997,1.5555218,1.8383441,1.8474089,1.8582866,1.8673514,1.8782293,1.887294,2.137483,2.3876717,2.6378605,2.8880494,3.1382382,3.1273603,3.1182957,3.1074178,3.0983531,3.0874753,2.8282216,2.5671551,2.3079014,2.0468347,1.7875811,1.8727903,1.9579996,2.0432088,2.126605,2.2118144,2.1392958,2.0667772,1.9942589,1.9217403,1.8492218,1.7132497,1.5754645,1.4376793,1.2998942,1.162109,1.1693609,1.1766127,1.1856775,1.1929294,1.2001812,1.4358664,1.6697385,1.9054236,2.1392958,2.374981,2.220879,2.0649643,1.9108626,1.7549478,1.6008459,0.5620184,0.76325727,0.96268314,1.162109,1.3633479,1.5627737,1.8492218,2.137483,2.4257438,2.712192,3.000453,2.8753586,2.7502642,2.6251698,2.5000753,2.374981,2.0631514,1.7495089,1.4376793,1.1258497,0.8122072,0.9119202,1.0116332,1.1131591,1.2128719,1.3125849,1.0497054,0.7868258,0.52575916,0.26287958,0.0,0.0,0.0,0.0,0.0,0.0,0.12509441,0.25018883,0.37528324,0.50037766,0.62547207,1.8492218,3.0747845,4.3003473,5.52591,6.7496595,6.5629244,6.3743763,6.187641,5.999093,5.812358,4.749962,3.6875658,2.6251698,1.5627737,0.50037766,0.774135,1.0497054,1.3252757,1.6008459,1.8746033,2.8372865,3.7999697,4.762653,5.7253356,6.688019,5.3500524,4.0120864,2.6741197,1.3379664,0.0,0.0,0.0,0.0,0.0,0.0,0.15047589,0.2991388,0.44961473,0.6000906,0.7505665,0.61278135,0.4749962,0.33721104,0.19942589,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.36259252,0.72518504,1.0877775,1.4503701,1.8129625,1.887294,1.9616255,2.03777,2.1121013,2.1882458,1.7748904,1.3633479,0.9499924,0.53663695,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,1.550083,3.0367124,4.5251546,6.011784,7.500226,7.6380115,7.7757964,7.911769,8.049554,8.187339,8.937905,9.686659,10.437225,11.187792,11.938358,10.937603,9.936848,8.937905,7.93715,6.9382076,6.874754,6.813113,6.7496595,6.688019,6.624565,5.3246713,4.024777,2.7248828,1.4249886,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.5873999,1.1747998,1.7621996,2.3495996,2.9369993,4.5632267,6.187641,7.8120556,9.438283,11.062697,11.213174,11.361836,11.512312,11.662788,11.813264,13.113158,14.413053,15.712947,17.01284,18.312735,15.899682,13.488441,11.075388,8.662335,6.249282,5.050914,3.8507326,2.6505513,1.4503701,0.25018883,0.2374981,0.22480737,0.21211663,0.19942589,0.18673515,0.42423326,0.66173136,0.89922947,1.1367276,1.3742256,1.8002719,2.2245052,2.6505513,3.0747845,3.5008307,2.9007401,2.3006494,1.7005589,1.1004683,0.50037766,0.44961473,0.40066472,0.34990177,0.2991388,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.4749962,0.76325727,1.0497054,1.3379664,1.6244144,1.6371052,1.649796,1.6624867,1.6751775,1.6878681,1.6244144,1.5627737,1.49932,1.4376793,1.3742256,2.7883365,4.2006345,5.612932,7.02523,8.437528,6.787732,5.137936,3.48814,1.8383441,0.18673515,0.2755703,0.36259252,0.44961473,0.53663695,0.62547207,0.9119202,1.2001812,1.4866294,1.7748904,2.0631514,1.9253663,1.7875811,1.649796,1.5120108,1.3742256,1.7132497,2.0504606,2.3876717,2.7248828,3.0620937,2.6505513,2.2371957,1.8256533,1.4122978,1.0007553,0.7995165,0.6000906,0.40066472,0.19942589,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.0497054,2.0994108,3.150929,4.2006345,5.2503395,5.1741953,5.0998635,5.0255322,4.949388,4.8750563,5.600241,6.3254266,7.0506115,7.7757964,8.499168,9.563377,10.625773,11.6881695,12.750566,13.812962,15.100165,16.38737,17.674572,18.961775,20.250792,19.712341,19.175705,18.637255,18.100618,17.562168,15.838041,14.112101,12.387974,10.662033,8.937905,11.563075,14.188245,16.813416,19.436771,22.061941,19.799364,17.536787,15.27421,13.011633,10.750868,9.425592,8.100317,6.775041,5.4497657,4.12449,4.6248674,5.125245,5.6256227,6.1241875,6.624565,6.8620634,7.0995617,7.3370595,7.574558,7.8120556,10.25049,12.687112,15.125546,17.562168,20.000603,17.912071,15.825351,13.736817,11.650098,9.563377,8.937905,8.312433,7.686961,7.063302,6.43783,5.8866897,5.337362,4.788034,4.2368937,3.6875658,5.487838,7.28811,9.088382,10.88684,12.687112,11.836833,10.988366,10.138086,9.287807,8.437528,7.5999393,6.7623506,5.924762,5.087173,4.249584,3.4246864,2.5997884,1.7748904,0.9499924,0.12509441,0.3245203,0.52575916,0.72518504,0.9246109,1.1258497,1.1494182,1.1747998,1.2001812,1.2255627,1.2491312,1.1367276,1.0243238,0.9119202,0.7995165,0.6871128,0.62547207,0.5620184,0.50037766,0.43692398,0.37528324,0.66173136,0.9499924,1.2382535,1.5247015,1.8129625,1.7368182,1.6624867,1.5881553,1.5120108,1.4376793,1.8002719,2.1628644,2.525457,2.8880494,3.2506418,3.299592,3.350355,3.3993049,3.4500678,3.5008307,3.1744974,2.8499773,2.525457,2.1991236,1.8746033,1.938057,1.9996977,2.0631514,2.124792,2.1882458,1.987007,1.7875811,1.5881553,1.3869164,1.1874905,1.1874905,1.1874905,1.1874905,1.1874905,1.1874905,1.1747998,1.162109,1.1494182,1.1367276,1.1258497,1.3742256,1.6244144,1.8746033,2.124792,2.374981,2.0994108,1.8256533,1.550083,1.2745126,1.0007553,0.48768693,0.67079616,0.8520924,1.0352017,1.2183108,1.3996071,1.6570477,1.9144884,2.1719291,2.42937,2.6868105,2.5744069,2.4620032,2.3495996,2.2371957,2.124792,1.8347181,1.5446441,1.2545701,0.9644961,0.6744221,0.7668832,0.85934424,0.95180535,1.0442665,1.1367276,0.922798,0.7070554,0.49312583,0.27738327,0.06164073,0.065266654,0.06707962,0.07070554,0.072518505,0.07433146,0.15954071,0.24474995,0.32995918,0.41516843,0.50037766,1.54827,2.5943494,3.6422417,4.690134,5.7380266,5.5875506,5.4370747,5.2865987,5.137936,4.98746,4.0954823,3.2016919,2.3097143,1.4177368,0.52575916,0.7868258,1.0497054,1.3125849,1.5754645,1.8383441,2.561716,3.2869012,4.0120864,4.7372713,5.462456,4.6266804,3.7927177,2.956942,2.1229792,1.2872034,1.064209,0.8430276,0.6200332,0.39703882,0.17585737,0.41516843,0.6544795,0.89560354,1.1349145,1.3742256,1.1421664,0.9101072,0.678048,0.44417584,0.21211663,0.18310922,0.15228885,0.12328146,0.092461094,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.29007402,0.58014804,0.87022203,1.1602961,1.4503701,1.5101979,1.5700256,1.6298534,1.6896812,1.7495089,1.4195497,1.0895905,0.75963134,0.42967212,0.099712946,0.0870222,0.07433146,0.06164073,0.05076295,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.22480737,0.26287958,0.2991388,0.33721104,0.37528324,0.41335547,1.7295663,3.04759,4.365614,5.6818247,6.9998484,7.17208,7.344311,7.518356,7.690587,7.8628187,8.339628,8.81825,9.295059,9.771869,10.25049,9.407463,8.564435,7.723221,6.880193,6.037165,5.8921285,5.7470913,5.6020546,5.4570174,5.3119802,4.269527,3.2270734,2.18462,1.1421664,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.5094425,0.969935,1.4304274,1.889107,2.3495996,3.6494937,4.949388,6.249282,7.549176,8.849071,8.970539,9.090195,9.20985,9.329506,9.449161,10.489801,11.530442,12.569269,13.60991,14.650551,12.732436,10.8143215,8.898021,6.979906,5.0617914,4.122677,3.1817493,2.2426348,1.3017071,0.36259252,0.34083697,0.31726846,0.2955129,0.27194437,0.25018883,0.4405499,0.629098,0.8194591,1.0098201,1.2001812,1.5228885,1.845596,2.1683033,2.4891977,2.811905,2.3296568,1.8474089,1.3651608,0.88291276,0.40066472,0.36077955,0.3208944,0.27919623,0.23931105,0.19942589,0.15954071,0.11965553,0.07977036,0.03988518,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.059827764,0.11965553,0.1794833,0.23931105,0.2991388,0.50037766,0.69980353,0.89922947,1.1004683,1.2998942,1.3923552,1.4848163,1.5772774,1.6697385,1.7621996,1.7368182,1.7132497,1.6878681,1.6624867,1.6371052,2.8282216,4.017525,5.2068286,6.397945,7.5872483,6.1006193,4.612177,3.1255474,1.6371052,0.15047589,0.26287958,0.37528324,0.48768693,0.6000906,0.7124943,0.922798,1.1331016,1.3434052,1.551896,1.7621996,1.6842422,1.6080978,1.5301404,1.452183,1.3742256,1.6117238,1.8492218,2.08672,2.324218,2.561716,2.2553256,1.9471219,1.6407311,1.3325275,1.0243238,0.86478317,0.70524246,0.54570174,0.38434806,0.22480737,0.18310922,0.13959812,0.09789998,0.054388877,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.90466833,1.7966459,2.6904364,3.5824142,4.4743915,4.501586,4.5305934,4.557788,4.5849824,4.612177,5.4407005,6.2674117,7.0941224,7.9226465,8.749357,9.637709,10.524248,11.4126,12.299138,13.1874895,14.110288,15.033086,15.955884,16.87687,17.799667,17.484211,17.170568,16.855114,16.539658,16.224201,15.636803,15.049402,14.462003,13.874602,13.287203,14.336908,15.386614,16.438131,17.487837,18.537542,17.534973,16.532406,15.529838,14.527269,13.524701,12.018129,10.509744,9.003172,7.494787,5.9882154,6.200332,6.412449,6.624565,6.836682,7.0506115,7.5056653,7.9607186,8.415772,8.870826,9.325879,11.300196,13.274512,15.250641,17.224958,19.199274,17.27572,15.350354,13.424988,11.499621,9.574255,8.943344,8.31062,7.6778965,7.0451727,6.412449,6.281915,6.153195,6.0226617,5.8921285,5.763408,7.309865,8.858135,10.4045925,11.952863,13.499319,12.897416,12.295512,11.691795,11.089892,10.487988,9.200785,7.911769,6.624565,5.337362,4.0501585,3.3376641,2.6251698,1.9126755,1.2001812,0.48768693,0.73424983,0.9826257,1.2291887,1.4775645,1.7241274,2.0649643,2.4058013,2.7448254,3.0856624,3.4246864,2.962381,2.5000753,2.03777,1.5754645,1.1131591,0.969935,0.82671094,0.6852999,0.5420758,0.40066472,0.69436467,0.9898776,1.2853905,1.5790904,1.8746033,1.794833,1.7150626,1.6352923,1.5555218,1.4757515,1.7767034,2.079468,2.382233,2.6849976,2.9877625,3.005892,3.0222087,3.0403383,3.056655,3.0747845,2.7883365,2.5000753,2.2118144,1.9253663,1.6371052,1.6806163,1.7223145,1.7658255,1.8075237,1.8492218,1.7132497,1.5754645,1.4376793,1.2998942,1.162109,1.1548572,1.1476053,1.1403534,1.1331016,1.1258497,1.0968424,1.0696479,1.0424535,1.015259,0.9880646,1.1893034,1.3923552,1.5954071,1.7966459,1.9996977,1.7748904,1.550083,1.3252757,1.1004683,0.87566096,0.41335547,0.57833505,0.7433147,0.90829426,1.0732739,1.2382535,1.4648738,1.693307,1.9199274,2.1483607,2.374981,2.275268,2.175555,2.0758421,1.9743162,1.8746033,1.6080978,1.3397794,1.0732739,0.80495536,0.53663695,0.62184614,0.7070554,0.79226464,0.8774739,0.96268314,0.79589057,0.62728506,0.4604925,0.291887,0.12509441,0.13053331,0.13415924,0.13959812,0.14503701,0.15047589,0.19579996,0.23931105,0.28463513,0.32995918,0.37528324,1.2455053,2.1157274,2.9841363,3.8543584,4.7245803,4.612177,4.499773,4.3873696,4.274966,4.162562,3.43919,2.7176309,1.9942589,1.2726997,0.5493277,0.7995165,1.0497054,1.2998942,1.550083,1.8002719,2.2879589,2.7756457,3.2633326,3.7492065,4.2368937,3.9051213,3.5733492,3.2397642,2.907992,2.5744069,2.1302311,1.6842422,1.2400664,0.79589057,0.34990177,0.67986095,1.0098201,1.3397794,1.6697385,1.9996977,1.6733645,1.3452182,1.017072,0.69073874,0.36259252,0.30276474,0.24293698,0.18310922,0.12328146,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.21755551,0.43511102,0.6526665,0.87022203,1.0877775,1.1331016,1.1766127,1.2219368,1.2672608,1.3125849,1.064209,0.81764615,0.56927025,0.32270733,0.07433146,0.07433146,0.07433146,0.07433146,0.07433146,0.07433146,0.15047589,0.22480737,0.2991388,0.37528324,0.44961473,0.51306844,0.5747091,0.63816285,0.69980353,0.76325727,1.9108626,3.056655,4.2042603,5.351866,6.4994707,6.7079616,6.9146395,7.12313,7.3298078,7.5382986,7.743163,7.948028,8.152893,8.357758,8.562622,7.877322,7.192023,6.506723,5.823236,5.137936,4.9095025,4.6828823,4.454449,4.227829,3.9993954,3.2143826,2.42937,1.6443571,0.85934424,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.43329805,0.7650702,1.0968424,1.4304274,1.7621996,2.7375734,3.7129474,4.688321,5.661882,6.637256,6.7279043,6.816739,6.9073873,6.9980354,7.0868707,7.8682575,8.647832,9.427405,10.20698,10.988366,9.56519,8.1420145,6.720652,5.297477,3.874301,3.1944401,2.514579,1.8347181,1.1548572,0.4749962,0.44236287,0.40972954,0.3770962,0.3444629,0.31182957,0.4550536,0.5982776,0.73968875,0.88291276,1.0243238,1.2455053,1.4648738,1.6842422,1.9054236,2.124792,1.7603867,1.3941683,1.0297627,0.6653573,0.2991388,0.27013144,0.23931105,0.21030366,0.1794833,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08339628,0.16497959,0.24837588,0.32995918,0.41335547,0.52575916,0.63816285,0.7505665,0.8629702,0.97537386,1.1476053,1.3198367,1.4920682,1.6642996,1.8383441,1.8492218,1.8619126,1.8746033,1.887294,1.8999848,2.8681068,3.834416,4.802538,5.77066,6.736969,5.411693,4.0882306,2.762955,1.4376793,0.11240368,0.25018883,0.387974,0.52575916,0.66173136,0.7995165,0.9318628,1.064209,1.1983683,1.3307146,1.4630609,1.4449311,1.4268016,1.4104849,1.3923552,1.3742256,1.5120108,1.649796,1.7875811,1.9253663,2.0631514,1.8600996,1.6570477,1.455809,1.2527572,1.0497054,0.9300498,0.8103943,0.69073874,0.56927025,0.44961473,0.36440548,0.27919623,0.19579996,0.11059072,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.75963134,1.4956942,2.229944,2.9641938,3.7002566,3.83079,3.9595103,4.0900435,4.220577,4.349297,5.279347,6.209397,7.1394467,8.069496,8.999546,9.712041,10.424535,11.137029,11.849524,12.562017,13.12041,13.67699,14.235382,14.791962,15.350354,15.257894,15.165432,15.072971,14.98051,14.888049,15.437376,15.986704,16.537846,17.087172,17.638313,17.112555,16.586794,16.062849,15.537089,15.013144,15.270584,15.528025,15.785465,16.042906,16.300346,14.610665,12.919171,11.22949,9.539809,7.850128,7.7757964,7.699652,7.6253204,7.549176,7.474845,8.147454,8.820063,9.492672,10.165281,10.837891,12.349901,13.861912,15.375735,16.887747,18.399757,16.637558,14.875358,13.113158,11.350959,9.5869465,8.94697,8.306994,7.667019,7.027043,6.3870673,6.677141,6.967215,7.2572894,7.5473633,7.837437,9.131892,10.428161,11.722616,13.017072,14.313339,13.957999,13.602658,13.247317,12.891977,12.536636,10.799818,9.063,7.324369,5.5875506,3.8507326,3.2506418,2.6505513,2.0504606,1.4503701,0.85027945,1.1457924,1.4394923,1.7350051,2.030518,2.324218,2.9805105,3.63499,4.2894692,4.945762,5.600241,4.788034,3.975827,3.1618068,2.3495996,1.5373923,1.3143979,1.0932164,0.87022203,0.64722764,0.42423326,0.726998,1.0297627,1.3325275,1.6352923,1.938057,1.8528478,1.7676386,1.6824293,1.5972201,1.5120108,1.7549478,1.9978848,2.2408218,2.4819458,2.7248828,2.7103791,2.6958754,2.6795588,2.665055,2.6505513,2.4003625,2.1501737,1.8999848,1.649796,1.3996071,1.4231756,1.4449311,1.4666867,1.4902552,1.5120108,1.4376793,1.3633479,1.2872034,1.2128719,1.1367276,1.1222239,1.1077201,1.0932164,1.0768998,1.062396,1.020698,0.97718686,0.9354887,0.8919776,0.85027945,1.0043813,1.1602961,1.3143979,1.4703126,1.6244144,1.4503701,1.2745126,1.1004683,0.9246109,0.7505665,0.33721104,0.48587397,0.6327239,0.7795739,0.92823684,1.0750868,1.2726997,1.4703126,1.6679256,1.8655385,2.0631514,1.9743162,1.887294,1.8002719,1.7132497,1.6244144,1.3796645,1.1349145,0.8901646,0.64541465,0.40066472,0.47680917,0.55476654,0.6327239,0.7106813,0.7868258,0.6671702,0.5475147,0.42785916,0.30820364,0.18673515,0.19579996,0.2030518,0.21030366,0.21755551,0.22480737,0.23024625,0.23568514,0.23931105,0.24474995,0.25018883,0.94274056,1.6352923,2.327844,3.0203958,3.7129474,3.636803,3.5624714,3.48814,3.4119956,3.3376641,2.7847104,2.231757,1.6806163,1.1276628,0.5747091,0.8122072,1.0497054,1.2872034,1.5247015,1.7621996,2.0123885,2.2625773,2.5127661,2.762955,3.0131438,3.1817493,3.3521678,3.5225863,3.6930048,3.8616104,3.1944401,2.5272698,1.8600996,1.1929294,0.52575916,0.9445535,1.3651608,1.7857682,2.2045624,2.6251698,2.2027495,1.7803292,1.357909,0.9354887,0.51306844,0.4224203,0.33177215,0.24293698,0.15228885,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14503701,0.29007402,0.43511102,0.58014804,0.72518504,0.7541924,0.7850128,0.81583315,0.8448406,0.87566096,0.7106813,0.54570174,0.38072214,0.21574254,0.05076295,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.22480737,0.33721104,0.44961473,0.5620184,0.6744221,0.76325727,0.85027945,0.93730164,1.0243238,1.1131591,2.0903459,3.0675328,4.0447197,5.0219064,6.000906,6.24203,6.484967,6.7279043,6.970841,7.211965,7.1448855,7.077806,7.0107265,6.9418335,6.874754,6.347182,5.81961,5.292038,4.764466,4.2368937,3.926877,3.6168604,3.3068438,2.9968271,2.6868105,2.1592383,1.6316663,1.1040943,0.57833505,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.35534066,0.56020546,0.7650702,0.969935,1.1747998,1.8256533,2.474694,3.1255474,3.774588,4.4254417,4.4852695,4.5450974,4.604925,4.664753,4.7245803,5.2449007,5.765221,6.285541,6.8058615,7.324369,6.397945,5.469708,4.5432844,3.6150475,2.6868105,2.268016,1.8474089,1.4268016,1.0080072,0.5873999,0.54570174,0.50219065,0.4604925,0.4169814,0.37528324,0.46955732,0.5656443,0.65991837,0.7541924,0.85027945,0.968122,1.0841516,1.2019942,1.3198367,1.4376793,1.1893034,0.94274056,0.69436467,0.44780177,0.19942589,0.1794833,0.15954071,0.13959812,0.11965553,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.10515183,0.21030366,0.3154555,0.42060733,0.52575916,0.5493277,0.5747091,0.6000906,0.62547207,0.6508536,0.90285534,1.1548572,1.4068589,1.6606737,1.9126755,1.9616255,2.0123885,2.0631514,2.1121013,2.1628644,2.907992,3.6531196,4.3982472,5.143375,5.8866897,4.7245803,3.5624714,2.4003625,1.2382535,0.07433146,0.2374981,0.40066472,0.5620184,0.72518504,0.8883517,0.94274056,0.99712944,1.0533313,1.1077201,1.162109,1.2056202,1.2473183,1.2908293,1.3325275,1.3742256,1.4122978,1.4503701,1.4866294,1.5247015,1.5627737,1.4648738,1.3669738,1.2708868,1.1729867,1.0750868,0.99531645,0.9155461,0.83577573,0.7541924,0.6744221,0.5475147,0.42060733,0.291887,0.16497959,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.61459434,1.1929294,1.7694515,2.3477864,2.9243085,3.1581807,3.39024,3.6222992,3.8543584,4.0882306,5.1198063,6.153195,7.1847706,8.21816,9.249735,9.788185,10.324821,10.863272,11.399909,11.938358,12.130532,12.322706,12.514881,12.707055,12.899229,13.029762,13.1602955,13.290829,13.419549,13.550082,15.23795,16.92582,18.611874,20.299742,21.98761,19.888199,17.786976,15.687565,13.588155,11.486931,13.00438,14.521831,16.03928,17.55673,19.074179,17.203201,15.330412,13.457622,11.584831,9.712041,9.349448,8.9868555,8.624263,8.26167,7.900891,8.789243,9.679407,10.5695715,11.459737,12.349901,13.399607,14.449312,15.50083,16.550535,17.60024,15.999394,14.400362,12.799516,11.200482,9.599637,8.952409,8.3051815,7.6579537,7.0107265,6.3616858,7.072367,7.783048,8.491917,9.202598,9.91328,10.955733,11.998186,13.04064,14.083094,15.125546,15.016769,14.909804,14.802839,14.695875,14.587097,12.400664,10.212419,8.024173,5.8377395,3.6494937,3.1618068,2.6741197,2.1882458,1.7005589,1.2128719,1.5555218,1.8981718,2.2408218,2.5816586,2.9243085,3.8942437,4.8641787,5.8341136,6.8040485,7.7757964,6.6118746,5.4497657,4.2876563,3.1255474,1.9616255,1.6606737,1.357909,1.0551442,0.7523795,0.44961473,0.75963134,1.0696479,1.3796645,1.6896812,1.9996977,1.9108626,1.8202144,1.7295663,1.6407311,1.550083,1.7331922,1.9144884,2.0975976,2.280707,2.4620032,2.4148662,2.3677292,2.3205922,2.2716422,2.2245052,2.0123885,1.8002719,1.5881553,1.3742256,1.162109,1.1657349,1.167548,1.1693609,1.1729867,1.1747998,1.162109,1.1494182,1.1367276,1.1258497,1.1131591,1.0895905,1.067835,1.0442665,1.0225109,1.0007553,0.94274056,0.88472575,0.82671094,0.7705091,0.7124943,0.8194591,0.92823684,1.0352017,1.1421664,1.2491312,1.1258497,1.0007553,0.87566096,0.7505665,0.62547207,0.26287958,0.39159992,0.52213323,0.6526665,0.78319985,0.9119202,1.0805258,1.2473183,1.4141108,1.5827163,1.7495089,1.6751775,1.6008459,1.5247015,1.4503701,1.3742256,1.1530442,0.9300498,0.7070554,0.48587397,0.26287958,0.33177215,0.40247768,0.47318324,0.5420758,0.61278135,0.5402629,0.46774435,0.39522585,0.32270733,0.25018883,0.25925365,0.27013144,0.27919623,0.29007402,0.2991388,0.26469254,0.23024625,0.19579996,0.15954071,0.12509441,0.6399758,1.1548572,1.6697385,2.18462,2.6995013,2.663242,2.6251698,2.5870976,2.5508385,2.5127661,2.1302311,1.7476959,1.3651608,0.9826257,0.6000906,0.824898,1.0497054,1.2745126,1.49932,1.7241274,1.7368182,1.7495089,1.7621996,1.7748904,1.7875811,2.4601903,3.1327994,3.8054085,4.478018,5.1506267,4.2604623,3.3702974,2.4801328,1.5899682,0.69980353,1.209246,1.7205015,2.229944,2.7393866,3.2506418,2.7321346,2.2154403,1.696933,1.1802386,0.66173136,0.5420758,0.4224203,0.30276474,0.18310922,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.072518505,0.14503701,0.21755551,0.29007402,0.36259252,0.3770962,0.39159992,0.40791658,0.4224203,0.43692398,0.35534066,0.27194437,0.19036107,0.10696479,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.15047589,0.2991388,0.44961473,0.6000906,0.7505665,0.89922947,1.0116332,1.1258497,1.2382535,1.3506571,1.4630609,2.269829,3.0765975,3.8851788,4.691947,5.5005283,5.7779117,6.055295,6.3326783,6.6100616,6.887445,6.546608,6.207584,5.866747,5.527723,5.186886,4.8170414,4.4471974,4.077353,3.7075086,3.3376641,2.9442513,2.5526514,2.1592383,1.7676386,1.3742256,1.1040943,0.83577573,0.5656443,0.2955129,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03988518,0.07977036,0.11965553,0.15954071,0.19942589,0.27738327,0.35534066,0.43329805,0.5094425,0.5873999,0.9119202,1.2382535,1.5627737,1.887294,2.2118144,2.2426348,2.2716422,2.3024626,2.333283,2.3622901,2.6233568,2.8826106,3.141864,3.4029307,3.6621845,3.2306993,2.7974012,2.3641033,1.9326181,1.49932,1.3397794,1.1802386,1.020698,0.85934424,0.69980353,0.64722764,0.5946517,0.5420758,0.4894999,0.43692398,0.48587397,0.533011,0.58014804,0.62728506,0.6744221,0.69073874,0.70524246,0.7197462,0.73424983,0.7505665,0.6200332,0.4894999,0.36077955,0.23024625,0.099712946,0.09064813,0.07977036,0.07070554,0.059827764,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.12690738,0.25562772,0.3825351,0.5094425,0.63816285,0.5747091,0.51306844,0.44961473,0.387974,0.3245203,0.65810543,0.9898776,1.3216497,1.6552348,1.987007,2.0758421,2.1628644,2.2498865,2.3369088,2.4257438,2.9478772,3.4700103,3.9921436,4.514277,5.038223,4.0374675,3.0367124,2.03777,1.0370146,0.038072214,0.22480737,0.41335547,0.6000906,0.7868258,0.97537386,0.95180535,0.9300498,0.90829426,0.88472575,0.8629702,0.9644961,1.067835,1.1693609,1.2726997,1.3742256,1.3125849,1.2491312,1.1874905,1.1258497,1.062396,1.0696479,1.0768998,1.0841516,1.0932164,1.1004683,1.0605831,1.020698,0.9808127,0.93911463,0.89922947,0.7306239,0.56020546,0.38978696,0.21936847,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.46955732,0.8901646,1.310772,1.7295663,2.1501737,2.4855716,2.819157,3.1545548,3.489953,3.825351,4.9602656,6.09518,7.230095,8.365009,9.499924,9.862516,10.225109,10.587702,10.950294,11.312886,11.1406555,10.966611,10.794379,10.622148,10.449916,10.801631,11.155159,11.506873,11.860401,12.212116,15.038525,17.863121,20.687716,23.512312,26.336908,22.662033,18.987158,15.312282,11.637406,7.9625316,10.73999,13.517449,16.294909,19.072367,21.849825,19.795738,17.73984,15.685752,13.629852,11.575767,10.924912,10.275872,9.625018,8.974165,8.325124,9.432844,10.540565,11.648285,12.754191,13.861912,14.449312,15.036712,15.625924,16.213324,16.800724,15.363045,13.925365,12.487686,11.050007,9.612328,8.957849,8.303369,7.647076,6.9925966,6.338117,7.4675927,8.597069,9.728357,10.857833,11.9873085,12.7777605,13.568212,14.356851,15.147303,15.937754,16.077353,16.21695,16.358362,16.49796,16.637558,13.999697,11.361836,8.725789,6.0879283,3.4500678,3.0747845,2.6995013,2.324218,1.9507477,1.5754645,1.9652514,2.3550384,2.7448254,3.1346123,3.5243993,4.8097897,6.09518,7.380571,8.664148,9.949538,8.437528,6.925517,5.411693,3.8996825,2.3876717,2.0051367,1.6226015,1.2400664,0.8575313,0.4749962,0.79226464,1.1095331,1.4268016,1.745883,2.0631514,1.9670644,1.8727903,1.7767034,1.6824293,1.5881553,1.7096237,1.8329052,1.9543737,2.077655,2.1991236,2.1193533,2.039583,1.9598125,1.8800422,1.8002719,1.6244144,1.4503701,1.2745126,1.1004683,0.9246109,0.90829426,0.8901646,0.872035,0.8557183,0.8375887,0.8883517,0.93730164,0.9880646,1.0370146,1.0877775,1.0569572,1.0279498,0.99712944,0.968122,0.93730164,0.86478317,0.79226464,0.7197462,0.64722764,0.5747091,0.6345369,0.69436467,0.7541924,0.81583315,0.87566096,0.7995165,0.72518504,0.6508536,0.5747091,0.50037766,0.18673515,0.2991388,0.41335547,0.52575916,0.63816285,0.7505665,0.8883517,1.0243238,1.162109,1.2998942,1.4376793,1.3742256,1.3125849,1.2491312,1.1874905,1.1258497,0.9246109,0.72518504,0.52575916,0.3245203,0.12509441,0.18673515,0.25018883,0.31182957,0.37528324,0.43692398,0.41335547,0.387974,0.36259252,0.33721104,0.31182957,0.3245203,0.33721104,0.34990177,0.36259252,0.37528324,0.2991388,0.22480737,0.15047589,0.07433146,0.0,0.33721104,0.6744221,1.0116332,1.3506571,1.6878681,1.6878681,1.6878681,1.6878681,1.6878681,1.6878681,1.4757515,1.261822,1.0497054,0.8375887,0.62547207,0.8375887,1.0497054,1.261822,1.4757515,1.6878681,1.4630609,1.2382535,1.0116332,0.7868258,0.5620184,1.7368182,2.911618,4.0882306,5.2630305,6.43783,5.3246713,4.213325,3.100166,1.987007,0.87566096,1.4757515,2.0758421,2.6741197,3.2742105,3.874301,3.2633326,2.6505513,2.03777,1.4249886,0.8122072,0.66173136,0.51306844,0.36259252,0.21211663,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.37528324,0.5620184,0.7505665,0.93730164,1.1258497,1.261822,1.3996071,1.5373923,1.6751775,1.8129625,2.4493124,3.0874753,3.7256382,4.361988,5.0001507,5.3119802,5.6256227,5.9374523,6.249282,6.5629244,5.9501433,5.337362,4.7245803,4.1117992,3.5008307,3.2869012,3.0747845,2.8626678,2.6505513,2.4366217,1.9616255,1.4866294,1.0116332,0.53663695,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06164073,0.12509441,0.18673515,0.25018883,0.31182957,0.41335547,0.51306844,0.61278135,0.7124943,0.8122072,0.7505665,0.6871128,0.62547207,0.5620184,0.50037766,0.50037766,0.50037766,0.50037766,0.50037766,0.50037766,0.41335547,0.3245203,0.2374981,0.15047589,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.15047589,0.2991388,0.44961473,0.6000906,0.7505665,0.6000906,0.44961473,0.2991388,0.15047589,0.0,0.41335547,0.824898,1.2382535,1.649796,2.0631514,2.1882458,2.3133402,2.4366217,2.561716,2.6868105,2.9877625,3.2869012,3.587853,3.8869917,4.1879435,3.350355,2.5127661,1.6751775,0.8375887,0.0,0.21211663,0.42423326,0.63816285,0.85027945,1.062396,0.96268314,0.8629702,0.76325727,0.66173136,0.5620184,0.72518504,0.8883517,1.0497054,1.2128719,1.3742256,1.2128719,1.0497054,0.8883517,0.72518504,0.5620184,0.6744221,0.7868258,0.89922947,1.0116332,1.1258497,1.1258497,1.1258497,1.1258497,1.1258497,1.1258497,0.9119202,0.69980353,0.48768693,0.2755703,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.3245203,0.5873999,0.85027945,1.1131591,1.3742256,1.8129625,2.2498865,2.6868105,3.1255474,3.5624714,4.800725,6.037165,7.2754188,8.511859,9.750113,9.936848,10.125396,10.312131,10.500679,10.687414,10.150778,9.612328,9.07569,8.537241,8.000604,8.575313,9.1500225,9.724731,10.29944,10.874149,14.837286,18.800423,22.761745,26.724882,30.688017,25.437677,20.187338,14.936998,9.686659,4.4381323,8.4756,12.513068,16.550535,20.588003,24.625471,22.386461,20.149265,17.912071,15.674874,13.437678,12.500377,11.563075,10.625773,9.686659,8.749357,10.074633,11.399909,12.725184,14.05046,15.375735,15.50083,15.624111,15.749206,15.8743,15.999394,14.724882,13.45037,12.175857,10.899531,9.625018,8.963287,8.299743,7.6380115,6.9744673,6.3127356,7.8628187,9.412902,10.962985,12.513068,14.06315,14.599788,15.138238,15.674874,16.213324,16.749962,17.137936,17.524096,17.912071,18.300045,18.688019,15.600543,12.513068,9.425592,6.338117,3.2506418,2.9877625,2.7248828,2.4620032,2.1991236,1.938057,2.374981,2.811905,3.2506418,3.6875658,4.12449,5.7253356,7.324369,8.925215,10.524248,12.125093,10.263181,8.399456,6.5375433,4.6756306,2.811905,2.3495996,1.887294,1.4249886,0.96268314,0.50037766,0.824898,1.1494182,1.4757515,1.8002719,2.124792,2.0250793,1.9253663,1.8256533,1.7241274,1.6244144,1.6878681,1.7495089,1.8129625,1.8746033,1.938057,1.8256533,1.7132497,1.6008459,1.4866294,1.3742256,1.2382535,1.1004683,0.96268314,0.824898,0.6871128,0.6508536,0.61278135,0.5747091,0.53663695,0.50037766,0.61278135,0.72518504,0.8375887,0.9499924,1.062396,1.0243238,0.9880646,0.9499924,0.9119202,0.87566096,0.7868258,0.69980353,0.61278135,0.52575916,0.43692398,0.44961473,0.46230546,0.4749962,0.48768693,0.50037766,0.4749962,0.44961473,0.42423326,0.40066472,0.37528324,0.15047589,0.23931105,0.32995918,0.42060733,0.5094425,0.6000906,0.7106813,0.8194591,0.9300498,1.0406405,1.1494182,1.1222239,1.0950294,1.067835,1.0406405,1.0116332,0.88472575,0.75781834,0.629098,0.50219065,0.37528324,0.36984438,0.36440548,0.36077955,0.35534066,0.34990177,0.32995918,0.3100166,0.29007402,0.27013144,0.25018883,0.25925365,0.27013144,0.27919623,0.29007402,0.2991388,0.23931105,0.1794833,0.11965553,0.059827764,0.0,0.27194437,0.54570174,0.81764615,1.0895905,1.3633479,1.3597219,1.357909,1.3542831,1.35247,1.3506571,1.1802386,1.0098201,0.83940166,0.67079616,0.50037766,0.6979906,0.89560354,1.0932164,1.2908293,1.4866294,1.3705997,1.2527572,1.1349145,1.017072,0.89922947,1.8655385,2.8300345,3.7945306,4.76084,5.7253356,4.784408,3.8452935,2.904366,1.9652514,1.0243238,1.4866294,1.9507477,2.4130533,2.8753586,3.3376641,3.0203958,2.7031271,2.3858588,2.0667772,1.7495089,1.7205015,1.6896812,1.6606737,1.6298534,1.6008459,1.3724127,1.1457924,0.91735905,0.69073874,0.46230546,0.36984438,0.27738327,0.18492219,0.092461094,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.2991388,0.44961473,0.6000906,0.7505665,0.89922947,1.0098201,1.1204109,1.2291887,1.3397794,1.4503701,1.9598125,2.469255,2.9805105,3.489953,3.9993954,4.249584,4.499773,4.749962,5.0001507,5.2503395,4.76084,4.269527,3.780027,3.290527,2.7992141,2.6306088,2.4601903,2.2897718,2.1193533,1.9507477,1.5827163,1.214685,0.8466535,0.48043507,0.11240368,0.09427405,0.07795739,0.059827764,0.04169814,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03988518,0.07977036,0.11965553,0.15954071,0.19942589,0.15954071,0.11965553,0.07977036,0.03988518,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,0.33539808,0.42060733,0.5058166,0.58921283,0.6744221,0.6399758,0.6055295,0.56927025,0.53482395,0.50037766,0.48587397,0.46955732,0.4550536,0.4405499,0.42423326,0.34990177,0.2755703,0.19942589,0.12509441,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.08339628,0.065266654,0.047137026,0.030820364,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.038072214,0.05076295,0.06164073,0.07433146,0.0870222,0.07070554,0.052575916,0.034446288,0.018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.11965553,0.23931105,0.36077955,0.48043507,0.6000906,0.48043507,0.36077955,0.23931105,0.11965553,0.0,0.32995918,0.65991837,0.9898776,1.3198367,1.649796,1.7694515,1.889107,2.0105755,2.1302311,2.2498865,2.4873846,2.7248828,2.962381,3.199879,3.437377,2.764768,2.0921588,1.4195497,0.7469406,0.07433146,0.27013144,0.46411842,0.65991837,0.8557183,1.0497054,0.9300498,0.8103943,0.69073874,0.56927025,0.44961473,0.59283876,0.73424983,0.8774739,1.020698,1.162109,1.020698,0.8774739,0.73424983,0.59283876,0.44961473,0.55476654,0.65991837,0.7650702,0.87022203,0.97537386,0.96087015,0.9445535,0.9300498,0.9155461,0.89922947,0.7306239,0.56020546,0.38978696,0.21936847,0.05076295,0.04169814,0.034446288,0.027194439,0.01994259,0.012690738,0.01994259,0.027194439,0.034446288,0.04169814,0.05076295,0.25925365,0.46955732,0.67986095,0.8901646,1.1004683,1.4757515,1.8492218,2.2245052,2.5997884,2.9750717,3.9957695,5.0146546,6.035352,7.0542374,8.074935,8.317872,8.560809,8.801933,9.04487,9.287807,9.099259,8.912524,8.725789,8.537241,8.350506,8.892582,9.434657,9.976733,10.520622,11.062697,14.273455,17.482399,20.693155,23.9021,27.112856,23.006495,18.901947,14.7974,10.692853,6.588306,10.047439,13.506571,16.967516,20.42665,23.887594,21.89515,19.902702,17.910257,15.917811,13.925365,12.594651,11.26575,9.935035,8.604321,7.2754188,9.115576,10.955733,12.79589,14.634234,16.474392,16.367426,16.260462,16.151684,16.04472,15.937754,14.400362,12.862969,11.325577,9.788185,8.2507925,8.194591,8.140202,8.0858135,8.029612,7.9752226,9.043057,10.109079,11.176914,12.244749,13.312584,13.827466,14.342347,14.857228,15.372109,15.8869915,16.445383,17.001963,17.560356,18.116936,18.675327,16.175253,13.675177,11.175101,8.675026,6.1749506,5.6455655,5.1143675,4.5849824,4.0555973,3.5243993,3.9105604,4.2949085,4.6792564,5.0654173,5.4497657,6.813113,8.174648,9.537996,10.899531,12.262879,10.48255,8.70222,6.921891,5.143375,3.3630457,2.7756457,2.1882458,1.6008459,1.0116332,0.42423326,0.69073874,0.9554313,1.2201238,1.4848163,1.7495089,1.696933,1.6443571,1.5917811,1.5392052,1.4866294,1.5881553,1.6878681,1.7875811,1.887294,1.987007,1.9054236,1.8220274,1.7404441,1.6570477,1.5754645,1.4141108,1.2545701,1.0950294,0.9354887,0.774135,0.7324369,0.69073874,0.64722764,0.6055295,0.5620184,0.64722764,0.7324369,0.81764615,0.90285534,0.9880646,0.9554313,0.922798,0.8901646,0.8575313,0.824898,0.7705091,0.71430725,0.65991837,0.6055295,0.5493277,0.5475147,0.54570174,0.5420758,0.5402629,0.53663695,0.52032024,0.50219065,0.48587397,0.46774435,0.44961473,0.11240368,0.1794833,0.24837588,0.3154555,0.3825351,0.44961473,0.533011,0.61459434,0.6979906,0.7795739,0.8629702,0.87022203,0.8774739,0.88472575,0.8919776,0.89922947,0.8448406,0.7904517,0.73424983,0.67986095,0.62547207,0.5529536,0.48043507,0.40791658,0.33539808,0.26287958,0.24837588,0.23205921,0.21755551,0.2030518,0.18673515,0.19579996,0.2030518,0.21030366,0.21755551,0.22480737,0.1794833,0.13415924,0.09064813,0.045324065,0.0,0.20667773,0.41516843,0.62184614,0.83033687,1.0370146,1.0333886,1.0279498,1.0225109,1.017072,1.0116332,0.88472575,0.75781834,0.629098,0.50219065,0.37528324,0.55839247,0.73968875,0.922798,1.1059072,1.2872034,1.2781386,1.2672608,1.258196,1.2473183,1.2382535,1.9924458,2.7466383,3.5026438,4.256836,5.0128417,4.2441454,3.4772623,2.7103791,1.9416829,1.1747998,1.49932,1.8256533,2.1501737,2.474694,2.7992141,2.7774587,2.7557032,2.7321346,2.7103791,2.6868105,2.7774587,2.8681068,2.956942,3.04759,3.1382382,2.6958754,2.2516994,1.8093367,1.3669738,0.9246109,0.73968875,0.55476654,0.36984438,0.18492219,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.22480737,0.33721104,0.44961473,0.5620184,0.6744221,0.75781834,0.83940166,0.922798,1.0043813,1.0877775,1.4703126,1.8528478,2.2353828,2.617918,3.000453,3.1871881,3.3757362,3.5624714,3.7492065,3.9377546,3.5697234,3.2016919,2.8354735,2.467442,2.0994108,1.9725033,1.845596,1.7168756,1.5899682,1.4630609,1.2019942,0.94274056,0.68167394,0.4224203,0.16316663,0.13959812,0.11784257,0.09427405,0.072518505,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.2574407,0.32814622,0.39703882,0.46774435,0.53663695,0.5293851,0.52213323,0.5148814,0.5076295,0.50037766,0.46955732,0.4405499,0.40972954,0.38072214,0.34990177,0.28826106,0.22480737,0.16316663,0.099712946,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03988518,0.07977036,0.11965553,0.15954071,0.19942589,0.16497959,0.13053331,0.09427405,0.059827764,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.07433146,0.099712946,0.12509441,0.15047589,0.17585737,0.13959812,0.10515183,0.07070554,0.034446288,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.09064813,0.1794833,0.27013144,0.36077955,0.44961473,0.36077955,0.27013144,0.1794833,0.09064813,0.0,0.24837588,0.4949388,0.7433147,0.9898776,1.2382535,1.35247,1.4666867,1.5827163,1.696933,1.8129625,1.987007,2.1628644,2.3369088,2.5127661,2.6868105,2.179181,1.6733645,1.1657349,0.65810543,0.15047589,0.32814622,0.5058166,0.68167394,0.85934424,1.0370146,0.8974165,0.75781834,0.61822027,0.47680917,0.33721104,0.4604925,0.581961,0.70524246,0.82671094,0.9499924,0.82671094,0.70524246,0.581961,0.4604925,0.33721104,0.43511102,0.533011,0.629098,0.726998,0.824898,0.79589057,0.7650702,0.73424983,0.70524246,0.6744221,0.5475147,0.42060733,0.291887,0.16497959,0.038072214,0.034446288,0.032633327,0.030820364,0.027194439,0.025381476,0.027194439,0.030820364,0.032633327,0.034446288,0.038072214,0.19579996,0.35171473,0.5094425,0.6671702,0.824898,1.1367276,1.4503701,1.7621996,2.0758421,2.3876717,3.1908143,3.9921436,4.795286,5.5966153,6.399758,6.697084,6.9944096,7.2917356,7.590874,7.8882003,8.049554,8.212721,8.375887,8.537241,8.700407,9.20985,9.719293,10.230548,10.73999,11.249433,13.70781,16.164375,18.622751,21.079315,23.537693,20.577126,17.61837,14.657803,11.697234,8.736667,11.62109,14.501887,17.384499,20.267109,23.14972,21.402023,19.654327,17.906631,16.160748,14.413053,12.690738,10.968424,9.244296,7.5219817,5.7996674,8.154706,10.509744,12.864782,15.219821,17.57486,17.235836,16.894999,16.554161,16.215137,15.8743,14.074029,12.27557,10.475298,8.675026,6.874754,7.4277077,7.9806614,8.531802,9.084756,9.637709,10.223296,10.80707,11.392657,11.978244,12.562017,13.055143,13.548269,14.039582,14.532708,15.025834,15.752831,16.47983,17.206827,17.935638,18.662638,16.749962,14.837286,12.92461,11.011934,9.099259,8.303369,7.5056653,6.7079616,5.910258,5.1125546,5.4443264,5.7779117,6.109684,6.4432693,6.775041,7.900891,9.024928,10.150778,11.274815,12.400664,10.701918,9.004985,7.308052,5.6093063,3.9123733,3.199879,2.4873846,1.7748904,1.062396,0.34990177,0.55476654,0.75963134,0.9644961,1.1693609,1.3742256,1.3705997,1.3651608,1.3597219,1.3542831,1.3506571,1.4866294,1.6244144,1.7621996,1.8999848,2.03777,1.9851941,1.9326181,1.8800422,1.8274662,1.7748904,1.5917811,1.4104849,1.2273756,1.0442665,0.8629702,0.81583315,0.7668832,0.7197462,0.6726091,0.62547207,0.68167394,0.73968875,0.79770356,0.8557183,0.9119202,0.88472575,0.8575313,0.83033687,0.8031424,0.774135,0.7523795,0.7306239,0.7070554,0.6852999,0.66173136,0.64541465,0.62728506,0.6091554,0.59283876,0.5747091,0.5656443,0.55476654,0.54570174,0.53482395,0.52575916,0.07433146,0.11965553,0.16497959,0.21030366,0.25562772,0.2991388,0.35534066,0.40972954,0.46411842,0.52032024,0.5747091,0.61822027,0.65991837,0.7016165,0.7451276,0.7868258,0.80495536,0.823085,0.83940166,0.8575313,0.87566096,0.73424983,0.5946517,0.4550536,0.3154555,0.17585737,0.16497959,0.15410182,0.14503701,0.13415924,0.12509441,0.13053331,0.13415924,0.13959812,0.14503701,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.14322405,0.28463513,0.42785916,0.56927025,0.7124943,0.70524246,0.6979906,0.69073874,0.68167394,0.6744221,0.58921283,0.5058166,0.42060733,0.33539808,0.25018883,0.4169814,0.5855869,0.7523795,0.91917205,1.0877775,1.1856775,1.2817645,1.3796645,1.4775645,1.5754645,2.1193533,2.665055,3.2107568,3.7546456,4.3003473,3.7056956,3.1092308,2.514579,1.9199274,1.3252757,1.5120108,1.7005589,1.887294,2.0758421,2.2625773,2.5345216,2.808279,3.0802233,3.3521678,3.6241121,3.834416,4.0447197,4.255023,4.465327,4.6756306,4.017525,3.3594196,2.7031271,2.0450218,1.3869164,1.1095331,0.8321498,0.55476654,0.27738327,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.15047589,0.22480737,0.2991388,0.37528324,0.44961473,0.5058166,0.56020546,0.61459434,0.67079616,0.72518504,0.9808127,1.2346275,1.4902552,1.745883,1.9996977,2.124792,2.2498865,2.374981,2.5000753,2.6251698,2.38042,2.13567,1.889107,1.6443571,1.3996071,1.3143979,1.2291887,1.1457924,1.0605831,0.97537386,0.823085,0.67079616,0.5166943,0.36440548,0.21211663,0.18492219,0.15772775,0.13053331,0.10333887,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.1794833,0.23568514,0.29007402,0.3444629,0.40066472,0.42060733,0.4405499,0.4604925,0.48043507,0.50037766,0.4550536,0.40972954,0.36440548,0.3208944,0.2755703,0.22480737,0.17585737,0.12509441,0.07433146,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.059827764,0.11965553,0.1794833,0.23931105,0.2991388,0.24837588,0.19579996,0.14322405,0.09064813,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.11240368,0.15047589,0.18673515,0.22480737,0.26287958,0.21030366,0.15772775,0.10515183,0.052575916,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.059827764,0.11965553,0.1794833,0.23931105,0.2991388,0.23931105,0.1794833,0.11965553,0.059827764,0.0,0.16497959,0.32995918,0.4949388,0.65991837,0.824898,0.9354887,1.0442665,1.1548572,1.2654479,1.3742256,1.4866294,1.6008459,1.7132497,1.8256533,1.938057,1.5954071,1.2527572,0.9101072,0.56745726,0.22480737,0.38434806,0.54570174,0.70524246,0.86478317,1.0243238,0.86478317,0.70524246,0.54570174,0.38434806,0.22480737,0.32814622,0.42967212,0.533011,0.6345369,0.73787576,0.6345369,0.533011,0.42967212,0.32814622,0.22480737,0.3154555,0.40429065,0.4949388,0.5855869,0.6744221,0.629098,0.5855869,0.5402629,0.4949388,0.44961473,0.36440548,0.27919623,0.19579996,0.11059072,0.025381476,0.027194439,0.030820364,0.032633327,0.034446288,0.038072214,0.034446288,0.032633327,0.030820364,0.027194439,0.025381476,0.13053331,0.23568514,0.34083697,0.44417584,0.5493277,0.7995165,1.0497054,1.2998942,1.550083,1.8002719,2.3858588,2.9696326,3.5552197,4.1408067,4.7245803,5.0781083,5.429823,5.7833505,6.1350656,6.48678,6.9998484,7.512917,8.024173,8.537241,9.050309,9.527119,10.00574,10.48255,10.959359,11.437981,13.142166,14.848164,16.55235,18.258347,19.96253,18.147755,16.33298,14.518205,12.701616,10.88684,13.192928,15.497204,17.803293,20.107569,22.411844,20.910711,19.407764,17.904818,16.401873,14.90074,12.785012,10.669285,8.55537,6.439643,4.325729,7.1956487,10.065568,12.935488,15.805408,18.675327,18.102432,17.529535,16.956638,16.385555,15.812659,13.749508,11.6881695,9.625018,7.5618668,5.5005283,6.6608243,7.819308,8.979604,10.139899,11.300196,11.401722,11.50506,11.608399,11.709926,11.813264,12.282822,12.752378,13.221936,13.693306,14.162864,15.06028,15.957697,16.855114,17.75253,18.649946,17.32467,15.999394,14.674119,13.3506565,12.025381,10.959359,9.89515,8.829127,7.764919,6.70071,6.979906,7.2591023,7.5401115,7.819308,8.100317,8.9868555,9.875207,10.761745,11.650098,12.536636,10.9230995,9.30775,7.6924005,6.0770507,4.461701,3.6241121,2.7865236,1.9507477,1.1131591,0.2755703,0.42060733,0.5656443,0.7106813,0.8557183,1.0007553,1.0424535,1.0841516,1.1276628,1.1693609,1.2128719,1.3869164,1.5627737,1.7368182,1.9126755,2.08672,2.0649643,2.0432088,2.0196402,1.9978848,1.9743162,1.7694515,1.5645868,1.3597219,1.1548572,0.9499924,0.8974165,0.8448406,0.79226464,0.73968875,0.6871128,0.7179332,0.7469406,0.7777609,0.80676836,0.8375887,0.81583315,0.79226464,0.7705091,0.7469406,0.72518504,0.73424983,0.7451276,0.7541924,0.7650702,0.774135,0.7433147,0.7106813,0.678048,0.64541465,0.61278135,0.6091554,0.6073425,0.6055295,0.60190356,0.6000906,0.038072214,0.059827764,0.08339628,0.10515183,0.12690738,0.15047589,0.17767033,0.20486477,0.23205921,0.25925365,0.28826106,0.36440548,0.44236287,0.52032024,0.5982776,0.6744221,0.7650702,0.8557183,0.9445535,1.0352017,1.1258497,0.91735905,0.7106813,0.50219065,0.2955129,0.0870222,0.08339628,0.07795739,0.072518505,0.06707962,0.06164073,0.065266654,0.06707962,0.07070554,0.072518505,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.07795739,0.15410182,0.23205921,0.3100166,0.387974,0.3770962,0.3680314,0.35715362,0.3480888,0.33721104,0.2955129,0.2520018,0.21030366,0.16679256,0.12509441,0.27738327,0.42967212,0.581961,0.73424983,0.8883517,1.0932164,1.2980812,1.502946,1.7078108,1.9126755,2.2480736,2.5816586,2.9170568,3.2524548,3.587853,3.1654327,2.7430124,2.3205922,1.8981718,1.4757515,1.5247015,1.5754645,1.6244144,1.6751775,1.7241274,2.2915847,2.8608549,3.4283123,3.9957695,4.5632267,4.893186,5.223145,5.5531044,5.883064,6.2130227,5.3391747,4.4671397,3.5951047,2.72307,1.8492218,1.4793775,1.1095331,0.73968875,0.36984438,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.22480737,0.2520018,0.27919623,0.30820364,0.33539808,0.36259252,0.4894999,0.61822027,0.7451276,0.872035,1.0007553,1.062396,1.1258497,1.1874905,1.2491312,1.3125849,1.1893034,1.067835,0.9445535,0.823085,0.69980353,0.65810543,0.61459434,0.5728962,0.5293851,0.48768693,0.44236287,0.39703882,0.35171473,0.30820364,0.26287958,0.23024625,0.19761293,0.16497959,0.13234627,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.10333887,0.14322405,0.18310922,0.2229944,0.26287958,0.3100166,0.35715362,0.40429065,0.45324063,0.50037766,0.4405499,0.38072214,0.3208944,0.25925365,0.19942589,0.16316663,0.12509441,0.0870222,0.05076295,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07977036,0.15954071,0.23931105,0.3208944,0.40066472,0.32995918,0.25925365,0.19036107,0.11965553,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.15047589,0.19942589,0.25018883,0.2991388,0.34990177,0.27919623,0.21030366,0.13959812,0.07070554,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.08339628,0.16497959,0.24837588,0.32995918,0.41335547,0.5166943,0.62184614,0.726998,0.8321498,0.93730164,0.9880646,1.0370146,1.0877775,1.1367276,1.1874905,1.0098201,0.8321498,0.6544795,0.47680917,0.2991388,0.44236287,0.5855869,0.726998,0.87022203,1.0116332,0.8321498,0.6526665,0.47318324,0.291887,0.11240368,0.19579996,0.27738327,0.36077955,0.44236287,0.52575916,0.44236287,0.36077955,0.27738327,0.19579996,0.11240368,0.19579996,0.27738327,0.36077955,0.44236287,0.52575916,0.46411842,0.40429065,0.3444629,0.28463513,0.22480737,0.18310922,0.13959812,0.09789998,0.054388877,0.012690738,0.01994259,0.027194439,0.034446288,0.04169814,0.05076295,0.04169814,0.034446288,0.027194439,0.01994259,0.012690738,0.065266654,0.11784257,0.17041849,0.2229944,0.2755703,0.46230546,0.6508536,0.8375887,1.0243238,1.2128719,1.5809034,1.9471219,2.3151531,2.6831846,3.049403,3.4573197,3.8652363,4.273153,4.6792564,5.087173,5.9501433,6.813113,7.6742706,8.537241,9.400211,9.844387,10.290376,10.734551,11.18054,11.624716,12.578335,13.53014,14.481945,15.435563,16.38737,15.716573,15.047589,14.376793,13.70781,13.037014,14.764768,16.492521,18.220274,19.948027,21.675781,20.417585,19.15939,17.903006,16.64481,15.386614,12.879286,10.371959,7.8646317,5.3573046,2.8499773,6.2347784,9.619579,13.00438,16.389181,19.775795,18.97084,18.165886,17.359118,16.554161,15.749206,13.424988,11.10077,8.774739,6.450521,4.12449,5.8921285,7.6597667,9.427405,11.195044,12.962683,12.581961,12.203052,11.822329,11.443419,11.062697,11.510499,11.958302,12.40429,12.852092,13.299893,14.367728,15.435563,16.503399,17.56942,18.637255,17.89938,17.163317,16.425442,15.687565,14.94969,13.617162,12.284635,10.952107,9.619579,8.287052,8.515485,8.7421055,8.970539,9.197159,9.425592,10.074633,10.725487,11.374527,12.025381,12.674421,11.142468,9.610515,8.076748,6.544795,5.0128417,4.0501585,3.0874753,2.124792,1.162109,0.19942589,0.28463513,0.36984438,0.4550536,0.5402629,0.62547207,0.71430725,0.80495536,0.89560354,0.98443866,1.0750868,1.2872034,1.49932,1.7132497,1.9253663,2.137483,2.1447346,2.1519866,2.1592383,2.1683033,2.175555,1.9471219,1.7205015,1.4920682,1.2654479,1.0370146,0.9808127,0.922798,0.86478317,0.80676836,0.7505665,0.7523795,0.7541924,0.75781834,0.75963134,0.76325727,0.7451276,0.726998,0.7106813,0.69255173,0.6744221,0.7179332,0.75963134,0.8031424,0.8448406,0.8883517,0.83940166,0.79226464,0.7451276,0.6979906,0.6508536,0.6544795,0.65991837,0.6653573,0.67079616,0.6744221,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.11240368,0.22480737,0.33721104,0.44961473,0.5620184,0.72518504,0.8883517,1.0497054,1.2128719,1.3742256,1.1004683,0.824898,0.5493277,0.2755703,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.13778515,0.2755703,0.41335547,0.5493277,0.6871128,1.0007553,1.3125849,1.6244144,1.938057,2.2498865,2.374981,2.5000753,2.6251698,2.7502642,2.8753586,2.6251698,2.374981,2.124792,1.8746033,1.6244144,1.5373923,1.4503701,1.3633479,1.2745126,1.1874905,2.0504606,2.911618,3.774588,4.6375585,5.5005283,5.9501433,6.399758,6.849373,7.3008003,7.750415,6.6626377,5.57486,4.4870825,3.3993049,2.3133402,1.8492218,1.3869164,0.9246109,0.46230546,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06164073,0.12509441,0.18673515,0.25018883,0.31182957,0.2755703,0.2374981,0.19942589,0.16316663,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.19942589,0.2755703,0.34990177,0.42423326,0.50037766,0.42423326,0.34990177,0.2755703,0.19942589,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.099712946,0.19942589,0.2991388,0.40066472,0.50037766,0.41335547,0.3245203,0.2374981,0.15047589,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.18673515,0.25018883,0.31182957,0.37528324,0.43692398,0.34990177,0.26287958,0.17585737,0.0870222,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.099712946,0.19942589,0.2991388,0.40066472,0.50037766,0.48768693,0.4749962,0.46230546,0.44961473,0.43692398,0.42423326,0.41335547,0.40066472,0.387974,0.37528324,0.50037766,0.62547207,0.7505665,0.87566096,1.0007553,0.7995165,0.6000906,0.40066472,0.19942589,0.0,0.06164073,0.12509441,0.18673515,0.25018883,0.31182957,0.25018883,0.18673515,0.12509441,0.06164073,0.0,0.07433146,0.15047589,0.22480737,0.2991388,0.37528324,0.2991388,0.22480737,0.15047589,0.07433146,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.12509441,0.25018883,0.37528324,0.50037766,0.62547207,0.774135,0.9246109,1.0750868,1.2255627,1.3742256,1.8383441,2.3006494,2.762955,3.2252605,3.6875658,4.900438,6.11331,7.324369,8.537241,9.750113,10.161655,10.57501,10.988366,11.399909,11.813264,12.012691,12.212116,12.413355,12.612781,12.812206,13.287203,13.762199,14.237195,14.712192,15.187187,16.338419,17.487837,18.637255,19.786674,20.937904,19.92446,18.912827,17.89938,16.887747,15.8743,12.975373,10.074633,7.175706,4.274966,1.3742256,5.275721,9.175404,13.075087,16.97477,20.87445,19.837437,18.800423,17.761595,16.72458,15.687565,13.100468,10.51337,7.9244595,5.337362,2.7502642,5.125245,7.500226,9.875207,12.250188,14.625169,13.762199,12.899229,12.038072,11.175101,10.312131,10.738177,11.162411,11.586644,12.012691,12.436923,13.675177,14.911617,16.14987,17.388124,18.624565,18.474089,18.325426,18.17495,18.024473,17.87581,16.274965,14.675932,13.075087,11.47424,9.875207,10.049252,10.225109,10.399154,10.57501,10.750868,11.162411,11.575767,11.9873085,12.400664,12.812206,11.361836,9.91328,8.46291,7.0125394,5.562169,4.4743915,3.386614,2.3006494,1.2128719,0.12509441,0.15047589,0.17585737,0.19942589,0.22480737,0.25018883,0.387974,0.52575916,0.66173136,0.7995165,0.93730164,1.1874905,1.4376793,1.6878681,1.938057,2.1882458,2.2245052,2.2625773,2.3006494,2.3369088,2.374981,2.124792,1.8746033,1.6244144,1.3742256,1.1258497,1.062396,1.0007553,0.93730164,0.87566096,0.8122072,0.7868258,0.76325727,0.73787576,0.7124943,0.6871128,0.6744221,0.66173136,0.6508536,0.63816285,0.62547207,0.69980353,0.774135,0.85027945,0.9246109,1.0007553,0.93730164,0.87566096,0.8122072,0.7505665,0.6871128,0.69980353,0.7124943,0.72518504,0.73787576,0.7505665,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.09064813,0.1794833,0.27013144,0.36077955,0.44961473,0.58014804,0.7106813,0.83940166,0.969935,1.1004683,0.8792868,0.65991837,0.4405499,0.21936847,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.07070554,0.065266654,0.059827764,0.054388877,0.05076295,0.047137026,0.045324065,0.04169814,0.03988518,0.038072214,0.21574254,0.39159992,0.56927025,0.7469406,0.9246109,1.1204109,1.3143979,1.5101979,1.7041848,1.8999848,1.9797552,2.0595255,2.1392958,2.220879,2.3006494,2.1030366,1.9054236,1.7078108,1.5101979,1.3125849,1.3325275,1.35247,1.3724127,1.3923552,1.4122978,2.034144,2.657803,3.2796493,3.9033084,4.5251546,5.23221,5.9392653,6.6481338,7.3551893,8.062244,7.6597667,7.2572894,6.8548117,6.452334,6.049856,5.9700856,5.8903155,5.810545,5.730775,5.6510043,4.5342193,3.4192474,2.3042755,1.1893034,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,0.21936847,0.19036107,0.15954071,0.13053331,0.099712946,0.08339628,0.065266654,0.047137026,0.030820364,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.05076295,0.06164073,0.07433146,0.0870222,0.099712946,0.17041849,0.23931105,0.3100166,0.38072214,0.44961473,0.46774435,0.48587397,0.50219065,0.52032024,0.53663695,0.48768693,0.43692398,0.387974,0.33721104,0.28826106,0.3045777,0.32270733,0.34083697,0.35715362,0.37528324,0.33539808,0.2955129,0.25562772,0.21574254,0.17585737,0.15410182,0.13415924,0.11421664,0.09427405,0.07433146,0.29007402,0.5058166,0.7197462,0.9354887,1.1494182,1.0333886,0.9155461,0.79770356,0.67986095,0.5620184,0.4604925,0.35715362,0.25562772,0.15228885,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.092461094,0.08520924,0.07795739,0.07070554,0.06164073,0.052575916,0.04169814,0.032633327,0.02175555,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.10515183,0.21030366,0.3154555,0.42060733,0.52575916,0.42060733,0.3154555,0.21030366,0.10515183,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.07977036,0.08520924,0.09064813,0.09427405,0.099712946,0.15047589,0.19942589,0.25018883,0.2991388,0.34990177,0.27919623,0.21030366,0.13959812,0.07070554,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.15954071,0.2955129,0.42967212,0.5656443,0.69980353,0.629098,0.56020546,0.4894999,0.42060733,0.34990177,0.37528324,0.40066472,0.42423326,0.44961473,0.4749962,0.5747091,0.6744221,0.774135,0.87566096,0.97537386,0.89922947,0.824898,0.7505665,0.6744221,0.6000906,0.6073425,0.61459434,0.62184614,0.630911,0.63816285,0.5094425,0.3825351,0.25562772,0.12690738,0.0,0.059827764,0.11965553,0.1794833,0.23931105,0.2991388,0.23931105,0.1794833,0.11965553,0.059827764,0.0,0.032633327,0.065266654,0.09789998,0.13053331,0.16316663,0.16679256,0.17223145,0.17767033,0.18310922,0.18673515,0.16497959,0.14322405,0.11965553,0.09789998,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.099712946,0.19942589,0.2991388,0.40066472,0.50037766,0.6327239,0.7650702,0.8974165,1.0297627,1.162109,1.6080978,2.0522738,2.4982624,2.9424384,3.386614,4.273153,5.1578784,6.0426044,6.92733,7.8120556,8.1420145,8.471974,8.801933,9.131892,9.461852,9.731983,10.002114,10.272246,10.542377,10.812509,11.704487,12.598277,13.490254,14.382232,15.27421,16.051971,16.829731,17.607492,18.385254,19.163015,18.280102,17.397188,16.514277,15.633177,14.750263,12.864782,10.979301,9.0956335,7.210152,5.3246713,7.723221,10.119957,12.516694,14.915243,17.31198,16.635744,15.957697,15.279649,14.601601,13.925365,11.862214,9.800876,7.7377243,5.674573,3.6132345,5.7833505,7.951654,10.12177,12.291886,14.462003,13.675177,12.888351,12.099712,11.312886,10.524248,10.990179,11.454298,11.920229,12.384347,12.850279,14.180993,15.509895,16.840609,18.169512,19.500225,18.79317,18.084301,17.377247,16.67019,15.963136,14.380419,12.797703,11.214987,9.63227,8.049554,8.39039,8.729415,9.070251,9.409276,9.750113,10.493427,11.234929,11.978244,12.719746,13.46306,12.164979,10.866898,9.570629,8.272549,6.9744673,5.732588,4.4907084,3.247016,2.0051367,0.76325727,0.6544795,0.5475147,0.4405499,0.33177215,0.22480737,0.3444629,0.46411842,0.5855869,0.70524246,0.824898,1.0605831,1.2944553,1.5301404,1.7658255,1.9996977,2.039583,2.079468,2.1193533,2.1592383,2.1991236,2.039583,1.8800422,1.7205015,1.5591478,1.3996071,1.305333,1.209246,1.114972,1.020698,0.9246109,0.90466833,0.88472575,0.86478317,0.8448406,0.824898,0.80495536,0.7850128,0.7650702,0.7451276,0.72518504,0.77232206,0.8194591,0.8665961,0.9155461,0.96268314,0.90829426,0.8520924,0.79770356,0.7433147,0.6871128,0.6979906,0.7070554,0.7179332,0.726998,0.73787576,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06707962,0.13415924,0.2030518,0.27013144,0.33721104,0.43511102,0.533011,0.629098,0.726998,0.824898,0.65991837,0.4949388,0.32995918,0.16497959,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.018129626,0.034446288,0.052575916,0.07070554,0.0870222,0.09064813,0.092461094,0.09427405,0.09789998,0.099712946,0.09427405,0.09064813,0.08520924,0.07977036,0.07433146,0.291887,0.5094425,0.726998,0.9445535,1.162109,1.2400664,1.3180238,1.3941683,1.4721256,1.550083,1.5845293,1.6207886,1.6552348,1.6896812,1.7241274,1.5809034,1.4358664,1.2908293,1.1457924,1.0007553,1.1276628,1.2545701,1.3832904,1.5101979,1.6371052,2.0196402,2.4021754,2.7847104,3.1672456,3.5497808,4.514277,5.480586,6.445082,7.409578,8.375887,8.656897,8.939718,9.222541,9.5053625,9.788185,10.089137,10.391902,10.694666,10.997431,11.300196,9.057561,6.814926,4.572292,2.3296568,0.0870222,0.07070554,0.052575916,0.034446288,0.018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.16497959,0.14322405,0.11965553,0.09789998,0.07433146,0.065266654,0.054388877,0.045324065,0.034446288,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.07433146,0.07433146,0.07433146,0.07433146,0.07433146,0.13959812,0.20486477,0.27013144,0.33539808,0.40066472,0.5094425,0.6200332,0.7306239,0.83940166,0.9499924,0.87566096,0.7995165,0.72518504,0.6508536,0.5747091,0.6091554,0.64541465,0.67986095,0.71430725,0.7505665,0.67079616,0.58921283,0.5094425,0.42967212,0.34990177,0.3100166,0.27013144,0.23024625,0.19036107,0.15047589,0.58014804,1.0098201,1.4394923,1.8691645,2.3006494,1.9652514,1.6298534,1.2944553,0.96087015,0.62547207,0.5076295,0.38978696,0.27194437,0.15410182,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.08520924,0.09427405,0.10515183,0.11421664,0.12509441,0.10515183,0.08520924,0.065266654,0.045324065,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.21030366,0.42060733,0.630911,0.83940166,1.0497054,0.83940166,0.630911,0.42060733,0.21030366,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.13415924,0.11965553,0.10515183,0.09064813,0.07433146,0.11240368,0.15047589,0.18673515,0.22480737,0.26287958,0.21030366,0.15772775,0.10515183,0.052575916,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.21936847,0.38978696,0.56020546,0.7306239,0.89922947,0.77232206,0.64541465,0.5166943,0.38978696,0.26287958,0.3245203,0.387974,0.44961473,0.51306844,0.5747091,0.6508536,0.72518504,0.7995165,0.87566096,0.9499924,1.0007553,1.0497054,1.1004683,1.1494182,1.2001812,1.1530442,1.1059072,1.0569572,1.0098201,0.96268314,0.7705091,0.57833505,0.38434806,0.19217403,0.0,0.045324065,0.09064813,0.13415924,0.1794833,0.22480737,0.1794833,0.13415924,0.09064813,0.045324065,0.0,0.065266654,0.13053331,0.19579996,0.25925365,0.3245203,0.32270733,0.3208944,0.31726846,0.3154555,0.31182957,0.27919623,0.24837588,0.21574254,0.18310922,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.07433146,0.15047589,0.22480737,0.2991388,0.37528324,0.4894999,0.6055295,0.7197462,0.83577573,0.9499924,1.3778516,1.8057107,2.231757,2.659616,3.0874753,3.6458678,4.2024474,4.76084,5.317419,5.8758116,6.1223745,6.3707504,6.6173134,6.8656893,7.112252,7.453089,7.7921133,8.13295,8.471974,8.812811,10.12177,11.432542,12.743314,14.052273,15.363045,15.767336,16.171627,16.57773,16.982021,17.388124,16.635744,15.883366,15.129172,14.376793,13.6244135,12.754191,11.885782,11.015561,10.145339,9.275117,10.17072,11.06451,11.9601145,12.855718,13.749508,13.43224,13.114971,12.797703,12.480434,12.163166,10.625773,9.088382,7.549176,6.011784,4.4743915,6.439643,8.404895,10.370146,12.335398,14.300649,13.588155,12.87566,12.163166,11.450671,10.738177,11.242181,11.747997,12.252001,12.757817,13.261822,14.684997,16.108173,17.529535,18.952711,20.375887,19.11044,17.84499,16.579542,15.3159075,14.05046,12.48406,10.919474,9.354887,7.7903004,6.2257137,6.7297173,7.2355337,7.7395372,8.245354,8.749357,9.822631,10.894093,11.967366,13.04064,14.112101,12.968122,11.822329,10.6783495,9.5325575,8.386765,6.9907837,5.5929894,4.195195,2.7974012,1.3996071,1.1602961,0.91917205,0.67986095,0.4405499,0.19942589,0.30276474,0.40429065,0.5076295,0.6091554,0.7124943,0.9318628,1.1530442,1.3724127,1.5917811,1.8129625,1.8546607,1.8981718,1.93987,1.983381,2.0250793,1.9543737,1.8854811,1.8147756,1.745883,1.6751775,1.54827,1.4195497,1.2926424,1.1657349,1.0370146,1.0225109,1.0080072,0.9916905,0.97718686,0.96268314,0.9354887,0.90829426,0.8792868,0.8520924,0.824898,0.8448406,0.86478317,0.88472575,0.90466833,0.9246109,0.8774739,0.83033687,0.78319985,0.73424983,0.6871128,0.69436467,0.7016165,0.7106813,0.7179332,0.72518504,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.045324065,0.09064813,0.13415924,0.1794833,0.22480737,0.29007402,0.35534066,0.42060733,0.48587397,0.5493277,0.4405499,0.32995918,0.21936847,0.11059072,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.11059072,0.11965553,0.13053331,0.13959812,0.15047589,0.14322405,0.13415924,0.12690738,0.11965553,0.11240368,0.36984438,0.62728506,0.88472575,1.1421664,1.3996071,1.3597219,1.3198367,1.2799516,1.2400664,1.2001812,1.1893034,1.1802386,1.1693609,1.1602961,1.1494182,1.0569572,0.9644961,0.872035,0.7795739,0.6871128,0.922798,1.1566701,1.3923552,1.6280404,1.8619126,2.0051367,2.1483607,2.2897718,2.4329958,2.5744069,3.7981565,5.0200934,6.24203,7.46578,8.6877165,9.655839,10.622148,11.59027,12.558392,13.524701,14.210001,14.895301,15.580601,16.264088,16.949387,13.580903,10.210606,6.8403077,3.4700103,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.11059072,0.09427405,0.07977036,0.065266654,0.05076295,0.047137026,0.045324065,0.04169814,0.03988518,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.05076295,0.11059072,0.17041849,0.23024625,0.29007402,0.34990177,0.5529536,0.7541924,0.9572442,1.1602961,1.3633479,1.261822,1.162109,1.062396,0.96268314,0.8629702,0.9155461,0.968122,1.020698,1.0732739,1.1258497,1.0043813,0.88472575,0.7650702,0.64541465,0.52575916,0.46411842,0.40429065,0.3444629,0.28463513,0.22480737,0.87022203,1.5156367,2.1592383,2.8046532,3.4500678,2.8971143,2.3441606,1.79302,1.2400664,0.6871128,0.55476654,0.4224203,0.29007402,0.15772775,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.07795739,0.10515183,0.13234627,0.15954071,0.18673515,0.15772775,0.12690738,0.09789998,0.06707962,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.3154555,0.629098,0.9445535,1.260009,1.5754645,1.260009,0.9445535,0.629098,0.3154555,0.0,0.045324065,0.09064813,0.13415924,0.1794833,0.22480737,0.19036107,0.15410182,0.11965553,0.08520924,0.05076295,0.07433146,0.099712946,0.12509441,0.15047589,0.17585737,0.13959812,0.10515183,0.07070554,0.034446288,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.27919623,0.48587397,0.69073874,0.89560354,1.1004683,0.9155461,0.7306239,0.54570174,0.36077955,0.17585737,0.2755703,0.37528324,0.4749962,0.5747091,0.6744221,0.72518504,0.774135,0.824898,0.87566096,0.9246109,1.1004683,1.2745126,1.4503701,1.6244144,1.8002719,1.696933,1.5954071,1.4920682,1.3905423,1.2872034,1.0297627,0.77232206,0.5148814,0.2574407,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.09789998,0.19579996,0.291887,0.38978696,0.48768693,0.47680917,0.46774435,0.45686656,0.44780177,0.43692398,0.39522585,0.35171473,0.3100166,0.26831847,0.22480737,0.1794833,0.13415924,0.09064813,0.045324065,0.0,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,0.3480888,0.44417584,0.5420758,0.6399758,0.73787576,1.1476053,1.5573349,1.9670644,2.3767939,2.7883365,3.0167696,3.247016,3.4772623,3.7075086,3.9377546,4.102734,4.267714,4.4326935,4.597673,4.762653,5.1723824,5.582112,5.9918413,6.4033837,6.813113,8.540867,10.266808,11.99456,13.722314,15.4500675,15.4827,15.515334,15.547967,15.580601,15.613234,14.989574,14.367728,13.745882,13.122223,12.500377,12.645414,12.790451,12.935488,13.080525,13.225562,12.618219,12.010877,11.401722,10.794379,10.1870365,10.230548,10.272246,10.315757,10.357455,10.399154,9.38752,8.375887,7.362441,6.350808,5.337362,7.0977483,8.858135,10.616709,12.377095,14.137483,13.499319,12.862969,12.224807,11.586644,10.950294,11.494183,12.039885,12.585587,13.129475,13.675177,15.190813,16.704638,18.220274,19.734098,21.249735,19.427708,17.60568,15.781839,13.959812,12.137785,10.589515,9.043057,7.494787,5.9483304,4.40006,5.0708566,5.7398396,6.4106355,7.079619,7.750415,9.151835,10.555068,11.958302,13.359721,14.762955,13.769451,12.7777605,11.784257,10.792566,9.800876,8.247167,6.695271,5.141562,3.589666,2.03777,1.6642996,1.2926424,0.91917205,0.5475147,0.17585737,0.25925365,0.3444629,0.42967212,0.5148814,0.6000906,0.80495536,1.0098201,1.214685,1.4195497,1.6244144,1.6697385,1.7150626,1.7603867,1.8057107,1.8492218,1.8691645,1.889107,1.9108626,1.9308052,1.9507477,1.789394,1.6298534,1.4703126,1.310772,1.1494182,1.1403534,1.1294757,1.1204109,1.1095331,1.1004683,1.064209,1.0297627,0.99531645,0.96087015,0.9246109,0.91735905,0.9101072,0.90285534,0.89560354,0.8883517,0.8466535,0.80676836,0.7668832,0.726998,0.6871128,0.69255173,0.6979906,0.7016165,0.7070554,0.7124943,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.14503701,0.17767033,0.21030366,0.24293698,0.2755703,0.21936847,0.16497959,0.11059072,0.054388877,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.13053331,0.14684997,0.16497959,0.18310922,0.19942589,0.19036107,0.1794833,0.17041849,0.15954071,0.15047589,0.44780177,0.7451276,1.0424535,1.3397794,1.6371052,1.4793775,1.3216497,1.1657349,1.0080072,0.85027945,0.79589057,0.73968875,0.6852999,0.629098,0.5747091,0.53482395,0.4949388,0.4550536,0.41516843,0.37528324,0.7179332,1.0605831,1.403233,1.745883,2.08672,1.9906329,1.892733,1.794833,1.696933,1.6008459,3.0802233,4.559601,6.0407915,7.520169,8.999546,10.652968,12.304577,13.957999,15.609608,17.26303,18.330864,19.396887,20.464722,21.532557,22.600391,18.102432,13.604471,9.106511,4.610364,0.11240368,0.09064813,0.06707962,0.045324065,0.02175555,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.054388877,0.047137026,0.03988518,0.032633327,0.025381476,0.030820364,0.034446288,0.03988518,0.045324065,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.07977036,0.13415924,0.19036107,0.24474995,0.2991388,0.5946517,0.8901646,1.1856775,1.4793775,1.7748904,1.649796,1.5247015,1.3996071,1.2745126,1.1494182,1.2201238,1.2908293,1.3597219,1.4304274,1.49932,1.3397794,1.1802386,1.020698,0.85934424,0.69980353,0.6200332,0.5402629,0.4604925,0.38072214,0.2991388,1.1602961,2.0196402,2.8807976,3.7401419,4.599486,3.83079,3.0602808,2.2897718,1.5192627,0.7505665,0.60190356,0.4550536,0.30820364,0.15954071,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.07070554,0.11421664,0.15954071,0.20486477,0.25018883,0.21030366,0.17041849,0.13053331,0.09064813,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.42060733,0.83940166,1.260009,1.6806163,2.0994108,1.6806163,1.260009,0.83940166,0.42060733,0.0,0.059827764,0.11965553,0.1794833,0.23931105,0.2991388,0.24474995,0.19036107,0.13415924,0.07977036,0.025381476,0.038072214,0.05076295,0.06164073,0.07433146,0.0870222,0.07070554,0.052575916,0.034446288,0.018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.34083697,0.58014804,0.8194591,1.0605831,1.2998942,1.0569572,0.81583315,0.5728962,0.32995918,0.0870222,0.22480737,0.36259252,0.50037766,0.63816285,0.774135,0.7995165,0.824898,0.85027945,0.87566096,0.89922947,1.2001812,1.49932,1.8002719,2.0994108,2.4003625,2.2426348,2.084907,1.9271792,1.7694515,1.6117238,1.2908293,0.968122,0.64541465,0.32270733,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.13053331,0.25925365,0.38978696,0.52032024,0.6508536,0.6327239,0.61459434,0.5982776,0.58014804,0.5620184,0.5094425,0.45686656,0.40429065,0.35171473,0.2991388,0.23931105,0.1794833,0.11965553,0.059827764,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.20486477,0.28463513,0.36440548,0.44417584,0.52575916,0.91735905,1.310772,1.7023718,2.0957847,2.4873846,2.3894846,2.2915847,2.1954978,2.0975976,1.9996977,2.0830941,2.1646774,2.2480736,2.3296568,2.4130533,2.8916752,3.3721104,3.8525455,4.3329806,4.8116026,6.9581504,9.102885,11.24762,13.392355,15.537089,15.198066,14.857228,14.518205,14.177367,13.838344,13.345218,12.852092,12.360779,11.867653,11.374527,12.534823,13.695119,14.855415,16.01571,17.174194,15.065719,12.955431,10.845142,8.734854,6.624565,7.027043,7.4295206,7.8319983,8.234476,8.636953,8.149267,7.663393,7.175706,6.688019,6.200332,7.755854,9.309563,10.865085,12.420607,13.974316,13.412297,12.850279,12.28826,11.724429,11.162411,11.747997,12.331772,12.917358,13.502945,14.0867195,15.694818,17.302916,18.9092,20.517298,22.125395,19.744976,17.364555,14.984136,12.605529,10.225109,8.694968,7.1648283,5.634688,4.1045475,2.5744069,3.4101827,4.2441454,5.0799212,5.915697,6.7496595,8.482852,10.2142315,11.947423,13.680615,15.411995,14.572594,13.7331915,12.891977,12.052575,11.213174,9.5053625,7.797552,6.089741,4.3819304,2.6741197,2.1701162,1.6642996,1.1602961,0.6544795,0.15047589,0.21755551,0.28463513,0.35171473,0.42060733,0.48768693,0.678048,0.8684091,1.0569572,1.2473183,1.4376793,1.4848163,1.5319533,1.5809034,1.6280404,1.6751775,1.7857682,1.8945459,2.0051367,2.1157274,2.2245052,2.032331,1.840157,1.647983,1.455809,1.261822,1.258196,1.2527572,1.2473183,1.2418793,1.2382535,1.1947423,1.1530442,1.1095331,1.067835,1.0243238,0.9898776,0.9554313,0.91917205,0.88472575,0.85027945,0.81764615,0.7850128,0.7523795,0.7197462,0.6871128,0.69073874,0.69255173,0.69436467,0.6979906,0.69980353,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.15047589,0.17585737,0.19942589,0.22480737,0.25018883,0.2374981,0.22480737,0.21211663,0.19942589,0.18673515,0.52575916,0.8629702,1.2001812,1.5373923,1.8746033,1.6008459,1.3252757,1.0497054,0.774135,0.50037766,0.40066472,0.2991388,0.19942589,0.099712946,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.51306844,0.96268314,1.4122978,1.8619126,2.3133402,1.9743162,1.6371052,1.2998942,0.96268314,0.62547207,2.3622901,4.099108,5.8377395,7.574558,9.313189,11.650098,13.987006,16.325727,18.662638,20.999546,22.449915,23.900286,25.350657,26.799213,28.249582,22.625772,17.00015,11.374527,5.750717,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,0.63816285,1.0243238,1.4122978,1.8002719,2.1882458,2.03777,1.887294,1.7368182,1.5881553,1.4376793,1.5247015,1.6117238,1.7005589,1.7875811,1.8746033,1.6751775,1.4757515,1.2745126,1.0750868,0.87566096,0.774135,0.6744221,0.5747091,0.4749962,0.37528324,1.4503701,2.525457,3.6005437,4.6756306,5.750717,4.762653,3.774588,2.7883365,1.8002719,0.8122072,0.6508536,0.48768693,0.3245203,0.16316663,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06164073,0.12509441,0.18673515,0.25018883,0.31182957,0.26287958,0.21211663,0.16316663,0.11240368,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.52575916,1.0497054,1.5754645,2.0994108,2.6251698,2.0994108,1.5754645,1.0497054,0.52575916,0.0,0.07433146,0.15047589,0.22480737,0.2991388,0.37528324,0.2991388,0.22480737,0.15047589,0.07433146,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.40066472,0.6744221,0.9499924,1.2255627,1.49932,1.2001812,0.89922947,0.6000906,0.2991388,0.0,0.17585737,0.34990177,0.52575916,0.69980353,0.87566096,0.87566096,0.87566096,0.87566096,0.87566096,0.87566096,1.2998942,1.7241274,2.1501737,2.5744069,3.000453,2.7883365,2.5744069,2.3622901,2.1501737,1.938057,1.550083,1.162109,0.774135,0.387974,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.16316663,0.3245203,0.48768693,0.6508536,0.8122072,0.7868258,0.76325727,0.73787576,0.7124943,0.6871128,0.62547207,0.5620184,0.50037766,0.43692398,0.37528324,0.2991388,0.22480737,0.15047589,0.07433146,0.0,0.0,0.0,0.0,0.0,0.0,0.06164073,0.12509441,0.18673515,0.25018883,0.31182957,0.6871128,1.062396,1.4376793,1.8129625,2.1882458,1.7621996,1.3379664,0.9119202,0.48768693,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.61278135,1.162109,1.7132497,2.2625773,2.811905,5.375434,7.93715,10.500679,13.062395,15.624111,14.911617,14.199123,13.486629,12.774135,12.06164,11.700861,11.338268,10.975676,10.613083,10.25049,12.4242325,14.599788,16.775343,18.950897,21.12464,17.511406,13.899984,10.28675,6.6753283,3.0620937,3.825351,4.5867953,5.3500524,6.11331,6.874754,6.9128265,6.9508986,6.987158,7.02523,7.063302,8.412147,9.762803,11.111648,12.462305,13.812962,13.325275,12.837588,12.349901,11.862214,11.374527,11.999999,12.625471,13.24913,13.874602,14.500074,16.200634,17.89938,19.59994,21.300497,22.999243,20.062244,17.125244,14.188245,11.249433,8.312433,6.8004227,5.2884116,3.774588,2.2625773,0.7505665,1.7495089,2.7502642,3.7492065,4.749962,5.750717,7.8120556,9.875207,11.938358,13.999697,16.062849,15.375735,14.68681,13.999697,13.312584,12.625471,10.761745,8.899834,7.037921,5.176008,3.3122826,2.6741197,2.03777,1.3996071,0.76325727,0.12509441,0.17585737,0.22480737,0.2755703,0.3245203,0.37528324,0.5493277,0.72518504,0.89922947,1.0750868,1.2491312,1.2998942,1.3506571,1.3996071,1.4503701,1.49932,1.7005589,1.8999848,2.0994108,2.3006494,2.5000753,2.275268,2.0504606,1.8256533,1.6008459,1.3742256,1.3742256,1.3742256,1.3742256,1.3742256,1.3742256,1.3252757,1.2745126,1.2255627,1.1747998,1.1258497,1.062396,1.0007553,0.93730164,0.87566096,0.8122072,0.7868258,0.76325727,0.73787576,0.7124943,0.6871128,0.6871128,0.6871128,0.6871128,0.6871128,0.6871128,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.15410182,0.21030366,0.26469254,0.3208944,0.37528324,0.35715362,0.34083697,0.32270733,0.3045777,0.28826106,0.5873999,0.8883517,1.1874905,1.4866294,1.7875811,1.5754645,1.3633479,1.1494182,0.93730164,0.72518504,0.62547207,0.52575916,0.42423326,0.3245203,0.22480737,0.20667773,0.19036107,0.17223145,0.15410182,0.13778515,0.6073425,1.0768998,1.54827,2.0178273,2.4873846,2.179181,1.8727903,1.5645868,1.258196,0.9499924,2.3296568,3.7093215,5.090799,6.4704633,7.850128,9.657652,11.465176,13.272699,15.080223,16.887747,18.029913,19.17208,20.314245,21.458225,22.600391,18.100618,13.600845,9.099259,4.599486,0.099712946,0.13053331,0.15954071,0.19036107,0.21936847,0.25018883,0.46955732,0.69073874,0.9101072,1.1294757,1.3506571,1.0968424,0.8448406,0.59283876,0.34083697,0.0870222,0.07070554,0.052575916,0.034446288,0.018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.03988518,0.07977036,0.11965553,0.15954071,0.19942589,0.5094425,0.8194591,1.1294757,1.4394923,1.7495089,1.6298534,1.5101979,1.3905423,1.2708868,1.1494182,1.2201238,1.2908293,1.3597219,1.4304274,1.49932,1.3397794,1.1802386,1.020698,0.85934424,0.69980353,0.62184614,0.54570174,0.46774435,0.38978696,0.31182957,1.1729867,2.032331,2.8916752,3.7528327,4.612177,3.825351,3.0367124,2.2498865,1.4630609,0.6744221,0.56927025,0.46411842,0.36077955,0.25562772,0.15047589,0.17767033,0.20486477,0.23205921,0.25925365,0.28826106,0.3770962,0.46774435,0.55839247,0.64722764,0.73787576,0.64722764,0.55839247,0.46774435,0.3770962,0.28826106,0.23931105,0.19217403,0.14503701,0.09789998,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.46411842,0.9300498,1.3941683,1.8600996,2.324218,1.889107,1.455809,1.020698,0.5855869,0.15047589,0.27738327,0.40429065,0.533011,0.65991837,0.7868258,0.6671702,0.5475147,0.42785916,0.30820364,0.18673515,0.15410182,0.12328146,0.09064813,0.058014803,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.11240368,0.16316663,0.21211663,0.26287958,0.31182957,0.27194437,0.23205921,0.19217403,0.15228885,0.11240368,0.34083697,0.56745726,0.79589057,1.0225109,1.2491312,1.0007553,0.7505665,0.50037766,0.25018883,0.0,0.13959812,0.27919623,0.42060733,0.56020546,0.69980353,0.7070554,0.71430725,0.72337204,0.7306239,0.73787576,1.0768998,1.4177368,1.7567607,2.0975976,2.4366217,2.3568513,2.277081,2.1973107,2.1175404,2.03777,1.693307,1.3470312,1.0025684,0.65810543,0.31182957,0.25925365,0.20667773,0.15410182,0.10333887,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.13053331,0.25925365,0.38978696,0.52032024,0.6508536,0.629098,0.6091554,0.58921283,0.56927025,0.5493277,0.50037766,0.44961473,0.40066472,0.34990177,0.2991388,0.23931105,0.1794833,0.11965553,0.059827764,0.0,0.0,0.0,0.0,0.0,0.0,0.059827764,0.11965553,0.1794833,0.23931105,0.2991388,0.6399758,0.9808127,1.3198367,1.6606737,1.9996977,1.6624867,1.3252757,0.9880646,0.6508536,0.31182957,0.25925365,0.20667773,0.15410182,0.10333887,0.05076295,0.4894999,0.9300498,1.3705997,1.8093367,2.2498865,4.795286,7.3406854,9.884272,12.429671,14.975071,14.054086,13.134913,12.215742,11.294757,10.375585,10.817947,11.26031,11.702674,12.145037,12.5873995,14.052273,15.517147,16.982021,18.446894,19.911768,16.697386,13.483003,10.266808,7.0524244,3.8380418,4.4798307,5.121619,5.765221,6.4070096,7.0506115,7.3896356,7.7304726,8.069496,8.410334,8.749357,9.644961,10.540565,11.434355,12.329959,13.225562,13.037014,12.850279,12.661731,12.474996,12.28826,12.817645,13.347031,13.878228,14.407614,14.936998,16.117237,17.297476,18.477715,19.657953,20.838192,18.17495,15.511708,12.850279,10.1870365,7.5256076,6.1731377,4.8206677,3.4681973,2.1157274,0.76325727,1.5627737,2.3622901,3.1618068,3.9631362,4.762653,6.8203654,8.8780775,10.93579,12.99169,15.049402,14.757515,14.465629,14.171928,13.880041,13.588155,11.787883,9.987611,8.187339,6.3870673,4.5867953,3.7727752,2.956942,2.1429217,1.3270886,0.51306844,0.48587397,0.45686656,0.42967212,0.40247768,0.37528324,0.5058166,0.6345369,0.7650702,0.89560354,1.0243238,1.114972,1.2056202,1.2944553,1.3851035,1.4757515,1.6244144,1.7748904,1.9253663,2.0758421,2.2245052,2.034144,1.845596,1.6552348,1.4648738,1.2745126,1.3252757,1.3742256,1.4249886,1.4757515,1.5247015,1.4594349,1.3941683,1.3307146,1.2654479,1.2001812,1.1566701,1.114972,1.0732739,1.0297627,0.9880646,0.9354887,0.88291276,0.83033687,0.7777609,0.72518504,0.7433147,0.75963134,0.7777609,0.79589057,0.8122072,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.15954071,0.24474995,0.32995918,0.41516843,0.50037766,0.47680917,0.4550536,0.43329805,0.40972954,0.387974,0.6508536,0.9119202,1.1747998,1.4376793,1.7005589,1.550083,1.3996071,1.2491312,1.1004683,0.9499924,0.85027945,0.7505665,0.6508536,0.5493277,0.44961473,0.40247768,0.35534066,0.30820364,0.25925365,0.21211663,0.7016165,1.1929294,1.6824293,2.1719291,2.663242,2.3858588,2.1066625,1.8292793,1.551896,1.2745126,2.2970235,3.3195345,4.3420453,5.3645563,6.3870673,7.665206,8.943344,10.21967,11.497808,12.774135,13.60991,14.445685,15.279649,16.115425,16.949387,13.575464,10.199727,6.8239913,3.4500678,0.07433146,0.15954071,0.24474995,0.32995918,0.41516843,0.50037766,0.93911463,1.3796645,1.8202144,2.2607644,2.6995013,2.1954978,1.6896812,1.1856775,0.67986095,0.17585737,0.13959812,0.10515183,0.07070554,0.034446288,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.09064813,0.06707962,0.045324065,0.02175555,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.3825351,0.61459434,0.8466535,1.0805258,1.3125849,1.2219368,1.1331016,1.0424535,0.95180535,0.8629702,0.9155461,0.968122,1.020698,1.0732739,1.1258497,1.0043813,0.88472575,0.7650702,0.64541465,0.52575916,0.46955732,0.41516843,0.36077955,0.3045777,0.25018883,0.89560354,1.5392052,2.18462,2.8300345,3.4754493,2.8880494,2.3006494,1.7132497,1.1258497,0.53663695,0.4894999,0.44236287,0.39522585,0.3480888,0.2991388,0.35534066,0.40972954,0.46411842,0.52032024,0.5747091,0.7541924,0.9354887,1.114972,1.2944553,1.4757515,1.2328146,0.9898776,0.7469406,0.5058166,0.26287958,0.21755551,0.17223145,0.12690738,0.08339628,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.40429065,0.8103943,1.214685,1.6207886,2.0250793,1.6806163,1.3343405,0.9898776,0.64541465,0.2991388,0.48043507,0.65991837,0.83940166,1.020698,1.2001812,1.0352017,0.87022203,0.70524246,0.5402629,0.37528324,0.3100166,0.24474995,0.1794833,0.11421664,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.22480737,0.3245203,0.42423326,0.52575916,0.62547207,0.52032024,0.41516843,0.3100166,0.20486477,0.099712946,0.27919623,0.4604925,0.6399758,0.8194591,1.0007553,0.7995165,0.6000906,0.40066472,0.19942589,0.0,0.10515183,0.21030366,0.3154555,0.42060733,0.52575916,0.5402629,0.55476654,0.56927025,0.5855869,0.6000906,0.8557183,1.1095331,1.3651608,1.6207886,1.8746033,1.9271792,1.9797552,2.032331,2.084907,2.137483,1.8347181,1.5319533,1.2291887,0.92823684,0.62547207,0.52032024,0.41516843,0.3100166,0.20486477,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.09789998,0.19579996,0.291887,0.38978696,0.48768693,0.47318324,0.45686656,0.44236287,0.42785916,0.41335547,0.37528324,0.33721104,0.2991388,0.26287958,0.22480737,0.1794833,0.13415924,0.09064813,0.045324065,0.0,0.0,0.0,0.0,0.0,0.0,0.058014803,0.11421664,0.17223145,0.23024625,0.28826106,0.59283876,0.8974165,1.2019942,1.5083848,1.8129625,1.5627737,1.3125849,1.062396,0.8122072,0.5620184,0.45686656,0.35171473,0.24837588,0.14322405,0.038072214,0.3680314,0.6979906,1.0279498,1.357909,1.6878681,4.215138,6.742408,9.269678,11.7969475,14.324218,13.196554,12.070704,10.943042,9.815379,8.6877165,9.935035,11.182353,12.429671,13.67699,14.924308,15.680313,16.434505,17.190512,17.944704,18.700708,15.881553,13.064208,10.246864,7.4295206,4.612177,5.1343102,5.658256,6.1803894,6.7025228,7.224656,7.8682575,8.510046,9.151835,9.795437,10.437225,10.877775,11.318325,11.757062,12.197612,12.638163,12.750566,12.862969,12.975373,13.087777,13.200181,13.635292,14.070402,14.505513,14.940624,15.375735,16.035654,16.695572,17.355492,18.01541,18.675327,16.287657,13.899984,11.512312,9.12464,6.736969,5.5440397,4.3529234,3.159994,1.9670644,0.774135,1.3742256,1.9743162,2.5744069,3.1744974,3.774588,5.826862,7.8791356,9.933222,11.985496,14.037769,14.139296,14.242634,14.34416,14.447499,14.5508375,12.812206,11.075388,9.336758,7.5999393,5.863121,4.8696175,3.877927,2.8844235,1.892733,0.89922947,0.79589057,0.69073874,0.5855869,0.48043507,0.37528324,0.4604925,0.54570174,0.629098,0.71430725,0.7995165,0.9300498,1.0605831,1.1893034,1.3198367,1.4503701,1.550083,1.649796,1.7495089,1.8492218,1.9507477,1.794833,1.6407311,1.4848163,1.3307146,1.1747998,1.2745126,1.3742256,1.4757515,1.5754645,1.6751775,1.5954071,1.5156367,1.4358664,1.3542831,1.2745126,1.2527572,1.2291887,1.2074331,1.1856775,1.162109,1.0823387,1.0025684,0.922798,0.8430276,0.76325727,0.79770356,0.8321498,0.8665961,0.90285534,0.93730164,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.16497959,0.27919623,0.39522585,0.5094425,0.62547207,0.5982776,0.56927025,0.5420758,0.5148814,0.48768693,0.7124943,0.93730164,1.162109,1.3869164,1.6117238,1.5247015,1.4376793,1.3506571,1.261822,1.1747998,1.0750868,0.97537386,0.87566096,0.774135,0.6744221,0.5982776,0.52032024,0.44236287,0.36440548,0.28826106,0.79770356,1.3071461,1.8184015,2.327844,2.8372865,2.5907235,2.3423476,2.0957847,1.8474089,1.6008459,2.2643902,2.9297476,3.5951047,4.2604623,4.9258194,5.67276,6.4197006,7.166641,7.915395,8.662335,9.189907,9.71748,10.245051,10.772624,11.300196,9.050309,6.8004227,4.550536,2.3006494,0.05076295,0.19036107,0.32995918,0.46955732,0.6091554,0.7505665,1.4104849,2.0704033,2.7303216,3.39024,4.0501585,3.29234,2.5345216,1.7767034,1.020698,0.26287958,0.21030366,0.15772775,0.10515183,0.052575916,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.25562772,0.40972954,0.5656443,0.7197462,0.87566096,0.81583315,0.7541924,0.69436467,0.6345369,0.5747091,0.6091554,0.64541465,0.67986095,0.71430725,0.7505665,0.67079616,0.58921283,0.5094425,0.42967212,0.34990177,0.31726846,0.28463513,0.2520018,0.21936847,0.18673515,0.61822027,1.0478923,1.4775645,1.9072367,2.3369088,1.9507477,1.5627737,1.1747998,0.7868258,0.40066472,0.40972954,0.42060733,0.42967212,0.4405499,0.44961473,0.533011,0.61459434,0.6979906,0.7795739,0.8629702,1.1331016,1.403233,1.6733645,1.9416829,2.2118144,1.8184015,1.4231756,1.0279498,0.6327239,0.2374981,0.19579996,0.15228885,0.11059072,0.06707962,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.3444629,0.69073874,1.0352017,1.3796645,1.7241274,1.4703126,1.214685,0.96087015,0.70524246,0.44961473,0.68167394,0.9155461,1.1476053,1.3796645,1.6117238,1.403233,1.1929294,0.9826257,0.77232206,0.5620184,0.46411842,0.3680314,0.27013144,0.17223145,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.33721104,0.48768693,0.63816285,0.7868258,0.93730164,0.7668832,0.5982776,0.42785916,0.2574407,0.0870222,0.21936847,0.35171473,0.48587397,0.61822027,0.7505665,0.6000906,0.44961473,0.2991388,0.15047589,0.0,0.07070554,0.13959812,0.21030366,0.27919623,0.34990177,0.37165734,0.39522585,0.4169814,0.4405499,0.46230546,0.6327239,0.8031424,0.97174793,1.1421664,1.3125849,1.4975071,1.6824293,1.8673514,2.0522738,2.2371957,1.9779422,1.7168756,1.4576219,1.1983683,0.93730164,0.7795739,0.62184614,0.46411842,0.30820364,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.065266654,0.13053331,0.19579996,0.25925365,0.3245203,0.3154555,0.3045777,0.2955129,0.28463513,0.2755703,0.25018883,0.22480737,0.19942589,0.17585737,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.0,0.0,0.0,0.0,0.0,0.054388877,0.11059072,0.16497959,0.21936847,0.2755703,0.54570174,0.81583315,1.0841516,1.3542831,1.6244144,1.4630609,1.2998942,1.1367276,0.97537386,0.8122072,0.6544795,0.49675176,0.34083697,0.18310922,0.025381476,0.24474995,0.46411842,0.6852999,0.90466833,1.1258497,3.63499,6.14413,8.655084,11.164224,13.675177,12.339024,11.004683,9.670342,8.334189,6.9998484,9.052122,11.104396,13.15667,15.210756,17.26303,17.308353,17.351866,17.397188,17.442513,17.487837,15.067532,12.647227,10.226922,7.8084297,5.388125,5.7906027,6.19308,6.5955577,6.9980354,7.400513,8.345067,9.28962,10.234174,11.18054,12.125093,12.11059,12.094274,12.07977,12.065266,12.050762,12.462305,12.87566,13.287203,13.700559,14.112101,14.452938,14.791962,15.132799,15.471823,15.812659,15.952258,16.091856,16.233267,16.372866,16.512463,14.400362,12.28826,10.174346,8.062244,5.9501433,4.9167547,3.8851788,2.8517902,1.8202144,0.7868258,1.1874905,1.5881553,1.987007,2.3876717,2.7883365,4.835171,6.882006,8.930654,10.9774885,13.024323,13.522888,14.01964,14.518205,15.014956,15.511708,13.836531,12.163166,10.487988,8.812811,7.137634,5.9682727,4.797099,3.6277382,2.4583774,1.2872034,1.1040943,0.922798,0.73968875,0.55839247,0.37528324,0.41516843,0.4550536,0.4949388,0.53482395,0.5747091,0.7451276,0.9155461,1.0841516,1.2545701,1.4249886,1.4757515,1.5247015,1.5754645,1.6244144,1.6751775,1.5555218,1.4358664,1.3143979,1.1947423,1.0750868,1.2255627,1.3742256,1.5247015,1.6751775,1.8256533,1.7295663,1.6352923,1.5392052,1.4449311,1.3506571,1.3470312,1.3452182,1.3434052,1.3397794,1.3379664,1.2291887,1.1222239,1.015259,0.90829426,0.7995165,0.8520924,0.90466833,0.9572442,1.0098201,1.062396,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.17041849,0.3154555,0.4604925,0.6055295,0.7505665,0.7179332,0.6852999,0.6526665,0.6200332,0.5873999,0.774135,0.96268314,1.1494182,1.3379664,1.5247015,1.49932,1.4757515,1.4503701,1.4249886,1.3996071,1.2998942,1.2001812,1.1004683,1.0007553,0.89922947,0.79226464,0.6852999,0.57833505,0.46955732,0.36259252,0.8919776,1.4231756,1.9525607,2.4819458,3.0131438,2.7955883,2.5780327,2.3604772,2.1429217,1.9253663,2.231757,2.5399606,2.8481643,3.1545548,3.4627585,3.680314,3.8978696,4.115425,4.3329806,4.550536,4.7699046,4.989273,5.2104545,5.429823,5.6491914,4.5251546,3.3993049,2.275268,1.1494182,0.025381476,0.21936847,0.41516843,0.6091554,0.80495536,1.0007553,1.8800422,2.759329,3.6404288,4.519716,5.4008155,4.3891826,3.3793623,2.3695421,1.3597219,0.34990177,0.27919623,0.21030366,0.13959812,0.07070554,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.12690738,0.20486477,0.28282216,0.36077955,0.43692398,0.40791658,0.3770962,0.3480888,0.31726846,0.28826106,0.3045777,0.32270733,0.34083697,0.35715362,0.37528324,0.33539808,0.2955129,0.25562772,0.21574254,0.17585737,0.16497959,0.15410182,0.14503701,0.13415924,0.12509441,0.34083697,0.55476654,0.7705091,0.98443866,1.2001812,1.0116332,0.824898,0.63816285,0.44961473,0.26287958,0.32995918,0.39703882,0.46411842,0.533011,0.6000906,0.7106813,0.8194591,0.9300498,1.0406405,1.1494182,1.5101979,1.8691645,2.229944,2.5907235,2.94969,2.4021754,1.8546607,1.3071461,0.75963134,0.21211663,0.17223145,0.13234627,0.092461094,0.052575916,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.28463513,0.56927025,0.8557183,1.1403534,1.4249886,1.260009,1.0950294,0.9300498,0.7650702,0.6000906,0.88472575,1.1693609,1.455809,1.7404441,2.0250793,1.7694515,1.5156367,1.260009,1.0043813,0.7505665,0.6200332,0.4894999,0.36077955,0.23024625,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,0.44961473,0.6508536,0.85027945,1.0497054,1.2491312,1.015259,0.7795739,0.54570174,0.3100166,0.07433146,0.15954071,0.24474995,0.32995918,0.41516843,0.50037766,0.40066472,0.2991388,0.19942589,0.099712946,0.0,0.034446288,0.07070554,0.10515183,0.13959812,0.17585737,0.20486477,0.23568514,0.26469254,0.2955129,0.3245203,0.40972954,0.4949388,0.58014804,0.6653573,0.7505665,1.067835,1.3851035,1.7023718,2.0196402,2.3369088,2.1193533,1.9017978,1.6842422,1.4666867,1.2491312,1.0406405,0.83033687,0.6200332,0.40972954,0.19942589,0.15954071,0.11965553,0.07977036,0.03988518,0.0,0.032633327,0.065266654,0.09789998,0.13053331,0.16316663,0.15772775,0.15228885,0.14684997,0.14322405,0.13778515,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.052575916,0.10515183,0.15772775,0.21030366,0.26287958,0.49675176,0.7324369,0.968122,1.2019942,1.4376793,1.3633479,1.2872034,1.2128719,1.1367276,1.062396,0.8520924,0.6417888,0.43329805,0.2229944,0.012690738,0.12328146,0.23205921,0.34264994,0.45324063,0.5620184,3.054842,5.5476656,8.040489,10.533313,13.024323,11.481492,9.940474,8.397643,6.8548117,5.3119802,8.171022,11.028252,13.885481,16.74271,19.59994,18.934582,18.269224,17.60568,16.940323,16.274965,14.2516985,12.230246,10.20698,8.185526,6.16226,6.445082,6.7279043,7.0107265,7.2917356,7.574558,8.821876,10.069194,11.318325,12.565643,13.812962,13.341592,12.872034,12.402477,11.9329195,11.463363,12.175857,12.888351,13.600845,14.313339,15.025834,15.270584,15.515334,15.760084,16.004833,16.249584,15.870674,15.489952,15.10923,14.730321,14.349599,12.513068,10.674724,8.838193,6.9998484,5.163317,4.2894692,3.4174345,2.5453994,1.6733645,0.7995165,1.0007553,1.2001812,1.3996071,1.6008459,1.8002719,3.8434806,5.8848767,7.9280853,9.969481,12.012691,12.904668,13.796645,14.690435,15.582414,16.474392,14.862667,13.24913,11.637406,10.025683,8.412147,7.065115,5.718084,4.36924,3.0222087,1.6751775,1.4141108,1.1548572,0.89560354,0.6345369,0.37528324,0.36984438,0.36440548,0.36077955,0.35534066,0.34990177,0.56020546,0.7705091,0.9808127,1.1893034,1.3996071,1.3996071,1.3996071,1.3996071,1.3996071,1.3996071,1.3143979,1.2291887,1.1457924,1.0605831,0.97537386,1.1747998,1.3742256,1.5754645,1.7748904,1.9743162,1.8655385,1.7549478,1.6443571,1.5355793,1.4249886,1.4431182,1.4594349,1.4775645,1.4956942,1.5120108,1.3778516,1.2418793,1.1077201,0.97174793,0.8375887,0.90829426,0.97718686,1.0478923,1.1167849,1.1874905,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.17585737,0.34990177,0.52575916,0.69980353,0.87566096,0.8375887,0.7995165,0.76325727,0.72518504,0.6871128,0.8375887,0.9880646,1.1367276,1.2872034,1.4376793,1.4757515,1.5120108,1.550083,1.5881553,1.6244144,1.5247015,1.4249886,1.3252757,1.2255627,1.1258497,0.9880646,0.85027945,0.7124943,0.5747091,0.43692398,0.9880646,1.5373923,2.08672,2.6378605,3.1871881,3.000453,2.811905,2.6251698,2.4366217,2.2498865,2.1991236,2.1501737,2.0994108,2.0504606,1.9996977,1.6878681,1.3742256,1.062396,0.7505665,0.43692398,0.34990177,0.26287958,0.17585737,0.0870222,0.0,0.0,0.0,0.0,0.0,0.0,0.25018883,0.50037766,0.7505665,1.0007553,1.2491312,2.3495996,3.4500678,4.550536,5.6491914,6.7496595,5.487838,4.2242026,2.962381,1.7005589,0.43692398,0.34990177,0.26287958,0.17585737,0.0870222,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.25018883,0.37528324,0.50037766,0.62547207,0.7505665,0.8883517,1.0243238,1.162109,1.2998942,1.4376793,1.887294,2.3369088,2.7883365,3.2379513,3.6875658,2.9877625,2.2879589,1.5881553,0.8883517,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06164073,0.12509441,0.18673515,0.25018883,0.31182957,0.25018883,0.18673515,0.12509441,0.06164073,0.0,0.22480737,0.44961473,0.6744221,0.89922947,1.1258497,1.0497054,0.97537386,0.89922947,0.824898,0.7505665,1.0877775,1.4249886,1.7621996,2.0994108,2.4366217,2.137483,1.8383441,1.5373923,1.2382535,0.93730164,0.774135,0.61278135,0.44961473,0.28826106,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06164073,0.12509441,0.18673515,0.25018883,0.31182957,0.5620184,0.8122072,1.062396,1.3125849,1.5627737,1.261822,0.96268314,0.66173136,0.36259252,0.06164073,0.099712946,0.13778515,0.17585737,0.21211663,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.0,0.0,0.0,0.0,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.18673515,0.18673515,0.18673515,0.18673515,0.18673515,0.63816285,1.0877775,1.5373923,1.987007,2.4366217,2.2625773,2.08672,1.9126755,1.7368182,1.5627737,1.2998942,1.0370146,0.774135,0.51306844,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,0.44961473,0.6508536,0.85027945,1.0497054,1.2491312,1.261822,1.2745126,1.2872034,1.2998942,1.3125849,1.0497054,0.7868258,0.52575916,0.26287958,0.0,0.0,0.0,0.0,0.0,0.0,2.474694,4.949388,7.4258947,9.900589,12.375282,10.625773,8.874452,7.124943,5.375434,3.6241121,7.28811,10.950294,14.612478,18.274662,21.936848,20.562622,19.188396,17.812357,16.438131,15.062093,13.437678,11.813264,10.1870365,8.562622,6.9382076,7.0995617,7.262728,7.4258947,7.5872483,7.750415,9.300498,10.850581,12.400664,13.9507475,15.50083,14.574407,13.649796,12.725184,11.800573,10.874149,11.887595,12.899229,13.912675,14.924308,15.937754,16.08823,16.236893,16.38737,16.537846,16.68832,15.787278,14.888049,13.987006,13.087777,12.186734,10.625773,9.063,7.500226,5.9374523,4.3746786,3.6621845,2.94969,2.2371957,1.5247015,0.8122072,0.8122072,0.8122072,0.8122072,0.8122072,0.8122072,2.8499773,4.8877473,6.925517,8.961474,10.999244,12.28826,13.575464,14.862667,16.14987,17.437075,15.8869915,14.336908,12.786825,11.236742,9.686659,8.161958,6.637256,5.1125546,3.587853,2.0631514,1.7241274,1.3869164,1.0497054,0.7124943,0.37528324,0.3245203,0.2755703,0.22480737,0.17585737,0.12509441,0.37528324,0.62547207,0.87566096,1.1258497,1.3742256,1.3252757,1.2745126,1.2255627,1.1747998,1.1258497,1.0750868,1.0243238,0.97537386,0.9246109,0.87566096,1.1258497,1.3742256,1.6244144,1.8746033,2.124792,1.9996977,1.8746033,1.7495089,1.6244144,1.49932,1.5373923,1.5754645,1.6117238,1.649796,1.6878681,1.5247015,1.3633479,1.2001812,1.0370146,0.87566096,0.96268314,1.0497054,1.1367276,1.2255627,1.3125849,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.034446288,0.058014803,0.07977036,0.10333887,0.12509441,0.24474995,0.36440548,0.48587397,0.6055295,0.72518504,0.73787576,0.7505665,0.76325727,0.774135,0.7868258,0.9445535,1.1022812,1.260009,1.4177368,1.5754645,1.7096237,1.845596,1.9797552,2.1157274,2.2498865,2.0069497,1.7658255,1.5228885,1.2799516,1.0370146,0.9246109,0.8122072,0.69980353,0.5873999,0.4749962,0.9300498,1.3851035,1.840157,2.2952106,2.7502642,2.6523643,2.5544643,2.4583774,2.3604772,2.2625773,2.2154403,2.1683033,2.1193533,2.0722163,2.0250793,1.7277533,1.4304274,1.1331016,0.83577573,0.53663695,0.43511102,0.33177215,0.23024625,0.12690738,0.025381476,0.02175555,0.01994259,0.018129626,0.014503701,0.012690738,0.21030366,0.40791658,0.6055295,0.8031424,1.0007553,1.8800422,2.759329,3.6404288,4.519716,5.4008155,4.3891826,3.3793623,2.3695421,1.3597219,0.34990177,0.27919623,0.21030366,0.13959812,0.07070554,0.0,0.032633327,0.065266654,0.09789998,0.13053331,0.16316663,0.13415924,0.10696479,0.07977036,0.052575916,0.025381476,0.12690738,0.23024625,0.33177215,0.43511102,0.53663695,0.5293851,0.52213323,0.5148814,0.5076295,0.50037766,0.40972954,0.3208944,0.23024625,0.13959812,0.05076295,0.04169814,0.034446288,0.027194439,0.01994259,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.01994259,0.027194439,0.034446288,0.04169814,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.059827764,0.07070554,0.07977036,0.09064813,0.099712946,0.19942589,0.2991388,0.40066472,0.50037766,0.6000906,0.7124943,0.824898,0.93730164,1.0497054,1.162109,1.5319533,1.9017978,2.2716422,2.6432993,3.0131438,2.5526514,2.0921588,1.6316663,1.1729867,0.7124943,0.56927025,0.42785916,0.28463513,0.14322405,0.0,0.0,0.0,0.0,0.0,0.0,0.07070554,0.13959812,0.21030366,0.27919623,0.34990177,0.40972954,0.46955732,0.5293851,0.58921283,0.6508536,0.6852999,0.7197462,0.7541924,0.7904517,0.824898,0.8774739,0.9300498,0.9826257,1.0352017,1.0877775,1.0025684,0.91735905,0.8321498,0.7469406,0.66173136,0.922798,1.1820517,1.4431182,1.7023718,1.9616255,1.7223145,1.4830034,1.2418793,1.0025684,0.76325727,0.629098,0.49675176,0.36440548,0.23205921,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.032633327,0.065266654,0.09789998,0.13053331,0.16316663,0.26831847,0.37165734,0.47680917,0.581961,0.6871128,1.0116332,1.3379664,1.6624867,1.987007,2.3133402,1.8600996,1.4068589,0.9554313,0.50219065,0.05076295,0.08520924,0.11965553,0.15410182,0.19036107,0.22480737,0.1794833,0.13415924,0.09064813,0.045324065,0.0,0.0,0.0,0.0,0.0,0.0,0.034446288,0.07070554,0.10515183,0.13959812,0.17585737,0.19036107,0.20486477,0.21936847,0.23568514,0.25018883,0.59283876,0.9354887,1.2781386,1.6207886,1.9616255,2.030518,2.0975976,2.1646774,2.231757,2.3006494,1.9181144,1.5355793,1.1530442,0.7705091,0.387974,0.35715362,0.32814622,0.29732585,0.26831847,0.2374981,0.19036107,0.14322405,0.09427405,0.047137026,0.0,0.07795739,0.15410182,0.23205921,0.3100166,0.387974,0.32270733,0.2574407,0.19217403,0.12690738,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.11059072,0.21936847,0.32995918,0.4405499,0.5493277,0.6526665,0.7541924,0.8575313,0.96087015,1.062396,1.1204109,1.1766127,1.2346275,1.2926424,1.3506571,1.1095331,0.87022203,0.629098,0.38978696,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,2.0160143,4.0302157,6.0444174,8.0604315,10.074633,8.887142,7.699652,6.5121617,5.3246713,4.137181,6.8529987,9.567003,12.282822,14.996826,17.712645,16.697386,15.682126,14.666867,13.651608,12.638163,11.563075,10.487988,9.412902,8.337815,7.262728,7.0904965,6.9182653,6.7442207,6.5719895,6.399758,7.795739,9.189907,10.585889,11.980057,13.374225,13.05333,12.730623,12.407916,12.085209,11.762501,12.215742,12.66717,13.12041,13.571837,14.025079,14.347786,14.670493,14.9932,15.314095,15.636803,14.7974,13.957999,13.116784,12.277383,11.437981,10.197914,8.957849,7.7177815,6.4777155,5.237649,4.572292,3.9069343,3.24339,2.5780327,1.9126755,1.7368182,1.5627737,1.3869164,1.2128719,1.0370146,2.9478772,4.856927,6.7677894,8.676839,10.587702,11.947423,13.307145,14.666867,16.026588,17.388124,16.091856,14.7974,13.502945,12.20849,10.912222,9.293246,7.6724577,6.051669,4.4326935,2.811905,2.4474995,2.0830941,1.7168756,1.35247,0.9880646,0.8321498,0.678048,0.52213323,0.3680314,0.21211663,0.43692398,0.66173136,0.8883517,1.1131591,1.3379664,1.2944553,1.2527572,1.209246,1.167548,1.1258497,1.0823387,1.0406405,0.99712944,0.9554313,0.9119202,1.162109,1.4122978,1.6624867,1.9126755,2.1628644,2.0667772,1.9725033,1.8782293,1.7821422,1.6878681,1.6697385,1.651609,1.6352923,1.6171626,1.6008459,1.4775645,1.3542831,1.2328146,1.1095331,0.9880646,1.0569572,1.1276628,1.1983683,1.2672608,1.3379664,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.07070554,0.11421664,0.15954071,0.20486477,0.25018883,0.3154555,0.38072214,0.44417584,0.5094425,0.5747091,0.63816285,0.69980353,0.76325727,0.824898,0.8883517,1.0533313,1.2183108,1.3832904,1.54827,1.7132497,1.9453088,2.1773682,2.4094272,2.6432993,2.8753586,2.4891977,2.1048496,1.7205015,1.3343405,0.9499924,0.8629702,0.774135,0.6871128,0.6000906,0.51306844,0.872035,1.2328146,1.5917811,1.9525607,2.3133402,2.3042755,2.2970235,2.2897718,2.2825198,2.275268,2.229944,2.18462,2.1392958,2.0957847,2.0504606,1.7676386,1.4848163,1.2019942,0.91917205,0.63816285,0.52032024,0.40247768,0.28463513,0.16679256,0.05076295,0.045324065,0.03988518,0.034446288,0.030820364,0.025381476,0.17041849,0.3154555,0.4604925,0.6055295,0.7505665,1.4104849,2.0704033,2.7303216,3.39024,4.0501585,3.29234,2.5345216,1.7767034,1.020698,0.26287958,0.21030366,0.15772775,0.10515183,0.052575916,0.0,0.065266654,0.13053331,0.19579996,0.25925365,0.3245203,0.27013144,0.21574254,0.15954071,0.10515183,0.05076295,0.25562772,0.4604925,0.6653573,0.87022203,1.0750868,1.0605831,1.0442665,1.0297627,1.015259,1.0007553,0.8194591,0.6399758,0.4604925,0.27919623,0.099712946,0.08520924,0.07070554,0.054388877,0.03988518,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.027194439,0.030820364,0.032633327,0.034446288,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.045324065,0.052575916,0.059827764,0.06707962,0.07433146,0.15047589,0.22480737,0.2991388,0.37528324,0.44961473,0.53663695,0.62547207,0.7124943,0.7995165,0.8883517,1.1766127,1.4666867,1.7567607,2.0468347,2.3369088,2.1175404,1.8981718,1.6769904,1.4576219,1.2382535,0.9898776,0.7433147,0.4949388,0.24837588,0.0,0.0,0.0,0.0,0.0,0.0,0.13959812,0.27919623,0.42060733,0.56020546,0.69980353,0.75781834,0.81583315,0.872035,0.9300498,0.9880646,1.1204109,1.2527572,1.3851035,1.5174497,1.649796,1.5301404,1.4104849,1.2908293,1.1693609,1.0497054,0.9554313,0.85934424,0.7650702,0.67079616,0.5747091,0.75781834,0.93911463,1.1222239,1.305333,1.4866294,1.3071461,1.1276628,0.9481794,0.7668832,0.5873999,0.48587397,0.3825351,0.27919623,0.17767033,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.065266654,0.13053331,0.19579996,0.25925365,0.3245203,0.47318324,0.6200332,0.7668832,0.9155461,1.062396,1.4630609,1.8619126,2.2625773,2.663242,3.0620937,2.4565642,1.8528478,1.2473183,0.6417888,0.038072214,0.07070554,0.10333887,0.13415924,0.16679256,0.19942589,0.15954071,0.11965553,0.07977036,0.03988518,0.0,0.0,0.0,0.0,0.0,0.0,0.032633327,0.065266654,0.09789998,0.13053331,0.16316663,0.19217403,0.2229944,0.2520018,0.28282216,0.31182957,0.5475147,0.78319985,1.017072,1.2527572,1.4866294,1.7966459,2.1066625,2.4166791,2.7266958,3.0367124,2.5345216,2.032331,1.5301404,1.0279498,0.52575916,0.5148814,0.5058166,0.4949388,0.48587397,0.4749962,0.38072214,0.28463513,0.19036107,0.09427405,0.0,0.15591478,0.3100166,0.46411842,0.6200332,0.774135,0.64541465,0.5148814,0.38434806,0.25562772,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.17041849,0.34083697,0.5094425,0.67986095,0.85027945,0.8557183,0.85934424,0.86478317,0.87022203,0.87566096,0.97718686,1.0805258,1.1820517,1.2853905,1.3869164,1.1693609,0.95180535,0.73424983,0.5166943,0.2991388,0.23931105,0.1794833,0.11965553,0.059827764,0.0,1.5555218,3.1092308,4.664753,6.2202744,7.7757964,7.1503243,6.5248523,5.89938,5.275721,4.650249,6.4178877,8.185526,9.953164,11.720803,13.486629,12.8321495,12.17767,11.5231905,10.866898,10.212419,9.686659,9.162713,8.636953,8.113008,7.5872483,7.079619,6.5719895,6.0643597,5.5567303,5.049101,6.2891674,7.5292335,8.7693,10.009366,11.249433,11.530442,11.809638,12.090648,12.3698435,12.650853,12.542075,12.43511,12.328146,12.219368,12.112403,12.607342,13.102281,13.597219,14.092158,14.587097,13.807523,13.027949,12.248375,11.466989,10.687414,9.770056,8.852696,7.935337,7.017978,6.1006193,5.482399,4.8641787,4.2477713,3.6295512,3.0131438,2.663242,2.3133402,1.9616255,1.6117238,1.261822,3.045777,4.8279195,6.6100616,8.392203,10.174346,11.608399,13.04064,14.47288,15.905121,17.33736,16.29672,15.257894,14.217253,13.178425,12.137785,10.422722,8.70766,6.9925966,5.277534,3.5624714,3.1708715,2.7774587,2.3858588,1.9924458,1.6008459,1.3397794,1.0805258,0.8194591,0.56020546,0.2991388,0.50037766,0.69980353,0.89922947,1.1004683,1.2998942,1.2654479,1.2291887,1.1947423,1.1602961,1.1258497,1.0895905,1.0551442,1.020698,0.98443866,0.9499924,1.2001812,1.4503701,1.7005589,1.9507477,2.1991236,2.13567,2.0704033,2.0051367,1.93987,1.8746033,1.8020848,1.7295663,1.6570477,1.5845293,1.5120108,1.4304274,1.3470312,1.2654479,1.1820517,1.1004683,1.1530442,1.2056202,1.258196,1.310772,1.3633479,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.10515183,0.17223145,0.23931105,0.30820364,0.37528324,0.38434806,0.39522585,0.40429065,0.41516843,0.42423326,0.53663695,0.6508536,0.76325727,0.87566096,0.9880646,1.1602961,1.3325275,1.504759,1.6769904,1.8492218,2.179181,2.5091403,2.8409123,3.1708715,3.5008307,2.9732587,2.4456866,1.9181144,1.3905423,0.8629702,0.7995165,0.73787576,0.6744221,0.61278135,0.5493277,0.81583315,1.0805258,1.3452182,1.6099107,1.8746033,1.9579996,2.039583,2.1229792,2.2045624,2.2879589,2.2444477,2.2027495,2.1592383,2.1175404,2.0758421,1.8075237,1.5392052,1.2726997,1.0043813,0.73787576,0.6055295,0.47318324,0.34083697,0.20667773,0.07433146,0.06707962,0.059827764,0.052575916,0.045324065,0.038072214,0.13053331,0.2229944,0.3154555,0.40791658,0.50037766,0.93911463,1.3796645,1.8202144,2.2607644,2.6995013,2.1954978,1.6896812,1.1856775,0.67986095,0.17585737,0.13959812,0.10515183,0.07070554,0.034446288,0.0,0.09789998,0.19579996,0.291887,0.38978696,0.48768693,0.40429065,0.32270733,0.23931105,0.15772775,0.07433146,0.3825351,0.69073874,0.99712944,1.305333,1.6117238,1.5899682,1.5682126,1.5446441,1.5228885,1.49932,1.2291887,0.96087015,0.69073874,0.42060733,0.15047589,0.12690738,0.10515183,0.08339628,0.059827764,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.045324065,0.09064813,0.13415924,0.1794833,0.22480737,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.034446288,0.032633327,0.030820364,0.027194439,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.030820364,0.034446288,0.03988518,0.045324065,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,0.2991388,0.36259252,0.42423326,0.48768693,0.5493277,0.61278135,0.823085,1.0333886,1.2418793,1.452183,1.6624867,1.6824293,1.7023718,1.7223145,1.742257,1.7621996,1.4104849,1.0569572,0.70524246,0.35171473,0.0,0.0,0.0,0.0,0.0,0.0,0.21030366,0.42060733,0.630911,0.83940166,1.0497054,1.1040943,1.1602961,1.214685,1.2708868,1.3252757,1.5555218,1.7857682,2.0142014,2.2444477,2.474694,2.182807,1.889107,1.5972201,1.305333,1.0116332,0.90829426,0.8031424,0.6979906,0.59283876,0.48768693,0.59283876,0.6979906,0.8031424,0.90829426,1.0116332,0.8919776,0.77232206,0.6526665,0.533011,0.41335547,0.34083697,0.26831847,0.19579996,0.12328146,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.09789998,0.19579996,0.291887,0.38978696,0.48768693,0.678048,0.8665961,1.0569572,1.2473183,1.4376793,1.9126755,2.3876717,2.8626678,3.3376641,3.8126602,3.054842,2.2970235,1.5392052,0.78319985,0.025381476,0.054388877,0.08520924,0.11421664,0.14503701,0.17585737,0.13959812,0.10515183,0.07070554,0.034446288,0.0,0.0,0.0,0.0,0.0,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.19579996,0.23931105,0.28463513,0.32995918,0.37528324,0.50219065,0.629098,0.75781834,0.88472575,1.0116332,1.5645868,2.1175404,2.6704938,3.2216346,3.774588,3.152742,2.5308957,1.9072367,1.2853905,0.66173136,0.6726091,0.68167394,0.69255173,0.7016165,0.7124943,0.56927025,0.42785916,0.28463513,0.14322405,0.0,0.23205921,0.46411842,0.6979906,0.9300498,1.162109,0.968122,0.77232206,0.57833505,0.3825351,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.0,0.0,0.0,0.0,0.0,0.23024625,0.4604925,0.69073874,0.91917205,1.1494182,1.0569572,0.9644961,0.872035,0.7795739,0.6871128,0.83577573,0.9826257,1.1294757,1.2781386,1.4249886,1.2291887,1.0352017,0.83940166,0.64541465,0.44961473,0.36077955,0.27013144,0.1794833,0.09064813,0.0,1.0950294,2.1900587,3.2850883,4.3801174,5.475147,5.411693,5.3500524,5.2865987,5.224958,5.163317,5.9827766,6.8022356,7.6216946,8.442966,9.262425,8.966913,8.673213,8.3777,8.082188,7.7866745,7.8120556,7.837437,7.8628187,7.8882003,7.911769,7.0705543,6.2275267,5.384499,4.5432844,3.7002566,4.784408,5.870373,6.9545245,8.040489,9.12464,10.007553,10.890467,11.773379,12.654479,13.537392,12.870221,12.203052,11.535881,10.866898,10.199727,10.866898,11.535881,12.203052,12.870221,13.537392,12.817645,12.097899,11.378153,10.658407,9.936848,9.342196,8.747544,8.152893,7.558241,6.9617763,6.392506,5.823236,5.2521524,4.6828823,4.1117992,3.587853,3.0620937,2.5381477,2.0123885,1.4866294,3.141864,4.797099,6.452334,8.107569,9.762803,11.267563,12.772322,14.277081,15.781839,17.286598,16.501585,15.716573,14.9333725,14.14836,13.363347,11.552197,9.742861,7.931711,6.1223745,4.313038,3.8924308,3.4718235,3.053029,2.6324217,2.2118144,1.8474089,1.4830034,1.1167849,0.7523795,0.387974,0.5620184,0.73787576,0.9119202,1.0877775,1.261822,1.2346275,1.2074331,1.1802386,1.1530442,1.1258497,1.0968424,1.0696479,1.0424535,1.015259,0.9880646,1.2382535,1.4866294,1.7368182,1.987007,2.2371957,2.2027495,2.1683033,2.132044,2.0975976,2.0631514,1.9344311,1.8075237,1.6806163,1.551896,1.4249886,1.3832904,1.3397794,1.2980812,1.2545701,1.2128719,1.2473183,1.2817645,1.3180238,1.35247,1.3869164,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.13959812,0.23024625,0.3208944,0.40972954,0.50037766,0.4550536,0.40972954,0.36440548,0.3208944,0.2755703,0.43692398,0.6000906,0.76325727,0.9246109,1.0877775,1.2672608,1.4467441,1.6280404,1.8075237,1.987007,2.4148662,2.8427253,3.2705846,3.6966307,4.12449,3.4555066,2.7847104,2.1157274,1.4449311,0.774135,0.73787576,0.69980353,0.66173136,0.62547207,0.5873999,0.75781834,0.92823684,1.0968424,1.2672608,1.4376793,1.6099107,1.7821422,1.9543737,2.126605,2.3006494,2.2607644,2.220879,2.179181,2.1392958,2.0994108,1.8474089,1.5954071,1.3415923,1.0895905,0.8375887,0.69073874,0.5420758,0.39522585,0.24837588,0.099712946,0.09064813,0.07977036,0.07070554,0.059827764,0.05076295,0.09064813,0.13053331,0.17041849,0.21030366,0.25018883,0.46955732,0.69073874,0.9101072,1.1294757,1.3506571,1.0968424,0.8448406,0.59283876,0.34083697,0.0870222,0.07070554,0.052575916,0.034446288,0.018129626,0.0,0.13053331,0.25925365,0.38978696,0.52032024,0.6508536,0.5402629,0.42967212,0.3208944,0.21030366,0.099712946,0.5094425,0.91917205,1.3307146,1.7404441,2.1501737,2.1193533,2.0903459,2.0595255,2.030518,1.9996977,1.6407311,1.2799516,0.91917205,0.56020546,0.19942589,0.17041849,0.13959812,0.11059072,0.07977036,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.059827764,0.11965553,0.1794833,0.23931105,0.2991388,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.04169814,0.034446288,0.027194439,0.01994259,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.014503701,0.018129626,0.01994259,0.02175555,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.15047589,0.18673515,0.22480737,0.26287958,0.2991388,0.33721104,0.46774435,0.5982776,0.726998,0.8575313,0.9880646,1.2473183,1.5083848,1.7676386,2.0268922,2.2879589,1.8292793,1.3724127,0.9155461,0.45686656,0.0,0.0,0.0,0.0,0.0,0.0,0.27919623,0.56020546,0.83940166,1.1204109,1.3996071,1.452183,1.504759,1.5573349,1.6099107,1.6624867,1.9906329,2.3169663,2.6451125,2.9732587,3.299592,2.8354735,2.3695421,1.9054236,1.4394923,0.97537386,0.85934424,0.7451276,0.629098,0.5148814,0.40066472,0.42785916,0.4550536,0.48224804,0.5094425,0.53663695,0.47680917,0.4169814,0.35715362,0.29732585,0.2374981,0.19579996,0.15228885,0.11059072,0.06707962,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13053331,0.25925365,0.38978696,0.52032024,0.6508536,0.88291276,1.114972,1.3470312,1.5809034,1.8129625,2.3622901,2.911618,3.4627585,4.0120864,4.5632267,3.6531196,2.7430124,1.8329052,0.922798,0.012690738,0.03988518,0.06707962,0.09427405,0.12328146,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.0,0.0,0.0,0.0,0.0,0.027194439,0.054388877,0.08339628,0.11059072,0.13778515,0.19761293,0.2574407,0.31726846,0.3770962,0.43692398,0.45686656,0.47680917,0.49675176,0.5166943,0.53663695,1.3325275,2.126605,2.9224956,3.7183862,4.512464,3.7691493,3.0276475,2.2843328,1.5428312,0.7995165,0.83033687,0.85934424,0.8901646,0.91917205,0.9499924,0.75963134,0.56927025,0.38072214,0.19036107,0.0,0.3100166,0.6200332,0.9300498,1.2400664,1.550083,1.2908293,1.0297627,0.7705091,0.5094425,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.0,0.0,0.0,0.0,0.0,0.29007402,0.58014804,0.87022203,1.1602961,1.4503701,1.260009,1.0696479,0.8792868,0.69073874,0.50037766,0.69255173,0.88472575,1.0768998,1.2708868,1.4630609,1.2908293,1.1167849,0.9445535,0.77232206,0.6000906,0.48043507,0.36077955,0.23931105,0.11965553,0.0,0.6345369,1.2690738,1.9054236,2.5399606,3.1744974,3.6748753,4.175253,4.6756306,5.1741953,5.674573,5.5476656,5.4207582,5.292038,5.1651306,5.038223,5.101677,5.1669436,5.23221,5.297477,5.3627434,5.9374523,6.5121617,7.0868707,7.66158,8.238102,7.059676,5.883064,4.704638,3.5280252,2.3495996,3.2796493,4.209699,5.139749,6.069799,6.9998484,8.484665,9.969481,11.454298,12.939114,14.425743,13.196554,11.969179,10.741803,9.514427,8.287052,9.128266,9.967669,10.80707,11.648285,12.487686,11.827768,11.16785,10.507931,9.848013,9.188094,8.914337,8.642392,8.370448,8.096691,7.8247466,7.3026133,6.78048,6.258347,5.7344007,5.2122674,4.512464,3.8126602,3.1128569,2.4130533,1.7132497,3.2397642,4.7680917,6.294606,7.8229337,9.349448,10.926725,12.5058155,14.083094,15.660371,17.237648,16.708263,16.177065,15.64768,15.118295,14.587097,12.681673,10.778063,8.872639,6.967215,5.0617914,4.615803,4.168001,3.720199,3.2723975,2.8245957,2.3550384,1.8854811,1.4141108,0.9445535,0.4749962,0.62547207,0.774135,0.9246109,1.0750868,1.2255627,1.2056202,1.1856775,1.1657349,1.1457924,1.1258497,1.1040943,1.0841516,1.064209,1.0442665,1.0243238,1.2745126,1.5247015,1.7748904,2.0250793,2.275268,2.269829,2.2643902,2.2607644,2.2553256,2.2498865,2.0667772,1.8854811,1.7023718,1.5192627,1.3379664,1.3343405,1.3325275,1.3307146,1.3270886,1.3252757,1.3434052,1.3597219,1.3778516,1.3941683,1.4122978,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.17585737,0.28826106,0.40066472,0.51306844,0.62547207,0.52575916,0.42423326,0.3245203,0.22480737,0.12509441,0.33721104,0.5493277,0.76325727,0.97537386,1.1874905,1.3742256,1.5627737,1.7495089,1.938057,2.124792,2.6505513,3.1744974,3.7002566,4.2242026,4.749962,3.9377546,3.1255474,2.3133402,1.49932,0.6871128,0.6744221,0.66173136,0.6508536,0.63816285,0.62547207,0.69980353,0.774135,0.85027945,0.9246109,1.0007553,1.261822,1.5247015,1.7875811,2.0504606,2.3133402,2.275268,2.2371957,2.1991236,2.1628644,2.124792,1.887294,1.649796,1.4122978,1.1747998,0.93730164,0.774135,0.61278135,0.44961473,0.28826106,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.16316663,0.3245203,0.48768693,0.6508536,0.8122072,0.6744221,0.53663695,0.40066472,0.26287958,0.12509441,0.63816285,1.1494182,1.6624867,2.175555,2.6868105,2.6505513,2.612479,2.5744069,2.5381477,2.5000753,2.0504606,1.6008459,1.1494182,0.69980353,0.25018883,0.21211663,0.17585737,0.13778515,0.099712946,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07433146,0.15047589,0.22480737,0.2991388,0.37528324,0.31182957,0.25018883,0.18673515,0.12509441,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.11240368,0.16316663,0.21211663,0.26287958,0.31182957,0.8122072,1.3125849,1.8129625,2.3133402,2.811905,2.2498865,1.6878681,1.1258497,0.5620184,0.0,0.0,0.0,0.0,0.0,0.0,0.34990177,0.69980353,1.0497054,1.3996071,1.7495089,1.8002719,1.8492218,1.8999848,1.9507477,1.9996977,2.4257438,2.8499773,3.2742105,3.7002566,4.12449,3.48814,2.8499773,2.2118144,1.5754645,0.93730164,0.8122072,0.6871128,0.5620184,0.43692398,0.31182957,0.26287958,0.21211663,0.16316663,0.11240368,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.16316663,0.3245203,0.48768693,0.6508536,0.8122072,1.0877775,1.3633479,1.6371052,1.9126755,2.1882458,2.811905,3.437377,4.062849,4.688321,5.3119802,4.249584,3.1871881,2.124792,1.062396,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.19942589,0.2755703,0.34990177,0.42423326,0.50037766,0.41335547,0.3245203,0.2374981,0.15047589,0.06164073,1.1004683,2.137483,3.1744974,4.213325,5.2503395,4.3873696,3.5243993,2.663242,1.8002719,0.93730164,0.9880646,1.0370146,1.0877775,1.1367276,1.1874905,0.9499924,0.7124943,0.4749962,0.2374981,0.0,0.387974,0.774135,1.162109,1.550083,1.938057,1.6117238,1.2872034,0.96268314,0.63816285,0.31182957,0.25018883,0.18673515,0.12509441,0.06164073,0.0,0.0,0.0,0.0,0.0,0.0,0.34990177,0.69980353,1.0497054,1.3996071,1.7495089,1.4630609,1.1747998,0.8883517,0.6000906,0.31182957,0.5493277,0.7868258,1.0243238,1.261822,1.49932,1.3506571,1.2001812,1.0497054,0.89922947,0.7505665,0.6000906,0.44961473,0.2991388,0.15047589,0.0,0.17585737,0.34990177,0.52575916,0.69980353,0.87566096,1.938057,3.000453,4.062849,5.125245,6.187641,5.1125546,4.0374675,2.962381,1.887294,0.8122072,1.2382535,1.6624867,2.08672,2.5127661,2.9369993,4.062849,5.186886,6.3127356,7.4367723,8.562622,7.0506115,5.5367875,4.024777,2.5127661,1.0007553,1.7748904,2.5508385,3.3249733,4.099108,4.8750563,6.9617763,9.050309,11.137029,13.225562,15.312282,13.524701,11.73712,9.949538,8.161958,6.3743763,7.3878226,8.399456,9.412902,10.424535,11.437981,10.837891,10.2378,9.637709,9.037619,8.437528,8.488291,8.537241,8.588004,8.636953,8.6877165,8.212721,7.7377243,7.262728,6.787732,6.3127356,5.4370747,4.5632267,3.6875658,2.811905,1.938057,3.3376641,4.7372713,6.1368785,7.5382986,8.937905,10.587702,12.237497,13.887294,15.537089,17.186886,16.913128,16.637558,16.361988,16.08823,15.812659,13.812962,11.811451,9.811753,7.8120556,5.812358,5.337362,4.8623657,4.3873696,3.9123733,3.437377,2.8626678,2.2879589,1.7132497,1.1367276,0.5620184,0.6871128,0.8122072,0.93730164,1.062396,1.1874905,1.1747998,1.162109,1.1494182,1.1367276,1.1258497,1.1131591,1.1004683,1.0877775,1.0750868,1.062396,1.3125849,1.5627737,1.8129625,2.0631514,2.3133402,2.3369088,2.3622901,2.3876717,2.4130533,2.4366217,2.1991236,1.9616255,1.7241274,1.4866294,1.2491312,1.2872034,1.3252757,1.3633479,1.3996071,1.4376793,1.4376793,1.4376793,1.4376793,1.4376793,1.4376793,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.14684997,0.24474995,0.34264994,0.4405499,0.53663695,0.5148814,0.49312583,0.46955732,0.44780177,0.42423326,0.63816285,0.85027945,1.062396,1.2745126,1.4866294,1.6824293,1.8782293,2.0722163,2.268016,2.4620032,2.8028402,3.141864,3.482701,3.8217251,4.162562,3.4772623,2.7919624,2.1066625,1.4231756,0.73787576,0.78319985,0.82671094,0.872035,0.91735905,0.96268314,1.0768998,1.1929294,1.3071461,1.4231756,1.5373923,1.7748904,2.0123885,2.2498865,2.4873846,2.7248828,2.6432993,2.5599031,2.47832,2.3949237,2.3133402,2.0432088,1.7730774,1.502946,1.2328146,0.96268314,0.81764615,0.6726091,0.5275721,0.3825351,0.2374981,0.2030518,0.16679256,0.13234627,0.09789998,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.44236287,0.88472575,1.3270886,1.7694515,2.2118144,2.0051367,1.7966459,1.5899682,1.3832904,1.1747998,1.452183,1.7295663,2.0069497,2.2843328,2.561716,2.6976883,2.8318477,2.9678197,3.101979,3.2379513,2.6324217,2.0268922,1.4231756,0.81764615,0.21211663,0.1794833,0.14684997,0.11421664,0.08339628,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.10515183,0.11059072,0.11421664,0.11965553,0.12509441,0.15047589,0.17585737,0.19942589,0.22480737,0.25018883,0.28282216,0.3154555,0.3480888,0.38072214,0.41335547,0.36259252,0.31182957,0.26287958,0.21211663,0.16316663,0.17223145,0.18310922,0.19217403,0.2030518,0.21211663,0.21211663,0.21211663,0.21211663,0.21211663,0.21211663,0.19942589,0.18673515,0.17585737,0.16316663,0.15047589,0.22662032,0.3045777,0.3825351,0.4604925,0.53663695,0.44236287,0.3480888,0.2520018,0.15772775,0.06164073,0.099712946,0.13778515,0.17585737,0.21211663,0.25018883,0.20486477,0.15954071,0.11421664,0.07070554,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.047137026,0.09427405,0.14322405,0.19036107,0.2374981,0.19942589,0.16316663,0.12509441,0.0870222,0.05076295,0.09064813,0.13053331,0.17041849,0.21030366,0.25018883,0.6508536,1.0497054,1.4503701,1.8492218,2.2498865,1.8002719,1.3506571,0.89922947,0.44961473,0.0,0.12509441,0.25018883,0.37528324,0.50037766,0.62547207,0.83940166,1.0551442,1.2708868,1.4848163,1.7005589,1.6896812,1.6806163,1.6697385,1.6606737,1.649796,2.3622901,3.0747845,3.787279,4.499773,5.2122674,4.4870825,3.7618973,3.0367124,2.3133402,1.5881553,1.3452182,1.1022812,0.85934424,0.61822027,0.37528324,0.50037766,0.62547207,0.7505665,0.87566096,1.0007553,1.0823387,1.1657349,1.2473183,1.3307146,1.4122978,1.1294757,0.8466535,0.5656443,0.28282216,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.054388877,0.11059072,0.16497959,0.21936847,0.2755703,0.49312583,0.7106813,0.92823684,1.1457924,1.3633479,1.6099107,1.8582866,2.1048496,2.3532255,2.5997884,3.2524548,3.9051213,4.557788,5.2104545,5.863121,4.762653,3.6621845,2.561716,1.4630609,0.36259252,0.37528324,0.387974,0.40066472,0.41335547,0.42423326,0.38434806,0.3444629,0.3045777,0.26469254,0.22480737,0.20486477,0.18492219,0.16497959,0.14503701,0.12509441,0.12690738,0.13053331,0.13234627,0.13415924,0.13778515,0.20667773,0.27738327,0.3480888,0.4169814,0.48768693,0.68167394,0.8774739,1.0732739,1.2672608,1.4630609,2.277081,3.092914,3.9069343,4.7227674,5.5367875,4.744523,3.9522583,3.159994,2.3677292,1.5754645,1.4956942,1.4141108,1.3343405,1.2545701,1.1747998,0.9481794,0.7197462,0.49312583,0.26469254,0.038072214,0.37528324,0.7124943,1.0497054,1.3869164,1.7241274,1.4304274,1.1349145,0.83940166,0.54570174,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.0,0.0,0.0,0.0,0.0,0.27919623,0.56020546,0.83940166,1.1204109,1.3996071,1.1693609,0.93911463,0.7106813,0.48043507,0.25018883,0.4405499,0.629098,0.8194591,1.0098201,1.2001812,1.0805258,0.96087015,0.83940166,0.7197462,0.6000906,0.5148814,0.42967212,0.3444629,0.25925365,0.17585737,0.3154555,0.4550536,0.5946517,0.73424983,0.87566096,2.0432088,3.2107568,4.3783045,5.5458527,6.7134004,6.1278133,5.542227,4.95664,4.3728657,3.787279,4.004834,4.2223897,4.439945,4.6575007,4.8750563,5.4044414,5.9356394,6.4650245,6.9944096,7.5256076,6.4668374,5.40988,4.3529234,3.295966,2.2371957,2.9877625,3.738329,4.4870825,5.237649,5.9882154,7.567306,9.14821,10.7273,12.308203,13.887294,12.594651,11.302009,10.009366,8.716724,7.4258947,8.258044,9.090195,9.922344,10.754494,11.586644,11.445232,11.302009,11.160598,11.017374,10.874149,10.839704,10.805257,10.770811,10.734551,10.700105,9.655839,8.609759,7.5654926,6.5194135,5.475147,4.7354584,3.9957695,3.254268,2.514579,1.7748904,3.0403383,4.305786,5.569421,6.834869,8.100317,9.557939,11.015561,12.473183,13.928991,15.386614,15.422873,15.457319,15.491765,15.528025,15.56247,13.898171,12.232059,10.567759,8.90346,7.2373466,7.0995617,6.9617763,6.825804,6.688019,6.550234,6.1169357,5.6854506,5.2521524,4.8206677,4.3873696,4.220577,4.0519714,3.8851788,3.7183862,3.5497808,3.1346123,2.7194438,2.3042755,1.8909199,1.4757515,1.7567607,2.039583,2.322405,2.6052272,2.8880494,3.053029,3.2180085,3.3829882,3.5479677,3.7129474,3.4645715,3.2180085,2.9696326,2.72307,2.474694,2.2879589,2.0994108,1.9126755,1.7241274,1.5373923,1.5355793,1.5319533,1.5301404,1.5283275,1.5247015,1.5083848,1.4902552,1.4721256,1.455809,1.4376793,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.11965553,0.2030518,0.28463513,0.3680314,0.44961473,0.5058166,0.56020546,0.61459434,0.67079616,0.72518504,0.93730164,1.1494182,1.3633479,1.5754645,1.7875811,1.9906329,2.1918716,2.3949237,2.5979755,2.7992141,2.955129,3.1092308,3.2651455,3.4192474,3.5751622,3.0167696,2.4601903,1.9017978,1.3452182,0.7868258,0.8901646,0.9916905,1.0950294,1.1983683,1.2998942,1.455809,1.6099107,1.7658255,1.9199274,2.0758421,2.2879589,2.5000753,2.712192,2.9243085,3.1382382,3.009518,2.8826106,2.7557032,2.6269827,2.5000753,2.1973107,1.8945459,1.5917811,1.2908293,0.9880646,0.85934424,0.7324369,0.6055295,0.47680917,0.34990177,0.291887,0.23568514,0.17767033,0.11965553,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.72337204,1.4449311,2.1683033,2.8898623,3.6132345,3.3358512,3.056655,2.7792716,2.5018883,2.2245052,2.268016,2.3097143,2.3532255,2.3949237,2.4366217,2.7448254,3.053029,3.3594196,3.6676233,3.975827,3.2143826,2.4547513,1.69512,0.9354887,0.17585737,0.14684997,0.11965553,0.092461094,0.065266654,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.11059072,0.14503701,0.1794833,0.21574254,0.25018883,0.2991388,0.34990177,0.40066472,0.44961473,0.50037766,0.5656443,0.629098,0.69436467,0.75963134,0.824898,0.72518504,0.62547207,0.52575916,0.42423326,0.3245203,0.3444629,0.36440548,0.38434806,0.40429065,0.42423326,0.42423326,0.42423326,0.42423326,0.42423326,0.42423326,0.40066472,0.37528324,0.34990177,0.3245203,0.2991388,0.38072214,0.4604925,0.5402629,0.6200332,0.69980353,0.5728962,0.44417584,0.31726846,0.19036107,0.06164073,0.15047589,0.2374981,0.3245203,0.41335547,0.50037766,0.40972954,0.3208944,0.23024625,0.13959812,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.09427405,0.19036107,0.28463513,0.38072214,0.4749962,0.387974,0.2991388,0.21211663,0.12509441,0.038072214,0.06707962,0.09789998,0.12690738,0.15772775,0.18673515,0.48768693,0.7868258,1.0877775,1.3869164,1.6878681,1.3506571,1.0116332,0.6744221,0.33721104,0.0,0.25018883,0.50037766,0.7505665,1.0007553,1.2491312,1.3307146,1.4104849,1.4902552,1.5700256,1.649796,1.5809034,1.5101979,1.4394923,1.3705997,1.2998942,2.3006494,3.299592,4.3003473,5.2992897,6.300045,5.487838,4.6756306,3.8616104,3.049403,2.2371957,1.8782293,1.5174497,1.1566701,0.79770356,0.43692398,0.73787576,1.0370146,1.3379664,1.6371052,1.938057,2.1030366,2.268016,2.4329958,2.5979755,2.762955,2.2100015,1.6570477,1.1040943,0.5529536,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.11059072,0.21936847,0.32995918,0.4405499,0.5493277,0.823085,1.0950294,1.3669738,1.6407311,1.9126755,2.132044,2.3532255,2.572594,2.7919624,3.0131438,3.6930048,4.3728657,5.0527267,5.732588,6.412449,5.275721,4.137181,3.000453,1.8619126,0.72518504,0.72518504,0.72518504,0.72518504,0.72518504,0.72518504,0.67079616,0.61459434,0.56020546,0.5058166,0.44961473,0.40972954,0.36984438,0.32995918,0.29007402,0.25018883,0.23024625,0.21030366,0.19036107,0.17041849,0.15047589,0.21574254,0.27919623,0.3444629,0.40972954,0.4749962,0.95180535,1.4304274,1.9072367,2.3858588,2.8626678,3.4555066,4.0483456,4.6393714,5.23221,5.825049,5.101677,4.3801174,3.6567454,2.9351864,2.2118144,2.0033236,1.79302,1.5827163,1.3724127,1.162109,0.9445535,0.726998,0.5094425,0.291887,0.07433146,0.36259252,0.6508536,0.93730164,1.2255627,1.5120108,1.2473183,0.9826257,0.7179332,0.45324063,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.0,0.0,0.0,0.0,0.0,0.21030366,0.42060733,0.630911,0.83940166,1.0497054,0.8774739,0.70524246,0.533011,0.36077955,0.18673515,0.32995918,0.47318324,0.61459434,0.75781834,0.89922947,0.8103943,0.7197462,0.629098,0.5402629,0.44961473,0.42967212,0.40972954,0.38978696,0.36984438,0.34990177,0.4550536,0.56020546,0.6653573,0.7705091,0.87566096,2.1483607,3.4192474,4.691947,5.964647,7.2373466,7.1430726,7.0469856,6.9527116,6.8566246,6.7623506,6.773228,6.782293,6.793171,6.8022356,6.813113,6.7478466,6.68258,6.6173134,6.552047,6.48678,5.8848767,5.282973,4.6792564,4.077353,3.4754493,4.2006345,4.9258194,5.6491914,6.3743763,7.0995617,8.172835,9.244296,10.31757,11.389031,12.462305,11.664601,10.866898,10.069194,9.273304,8.4756,9.128266,9.77912,10.431787,11.084454,11.73712,12.052575,12.368031,12.681673,12.9971285,13.312584,13.192928,13.073273,12.951805,12.8321495,12.712494,11.097144,9.481794,7.8682575,6.2529078,4.6375585,4.0320287,3.4283123,2.8227828,2.2172532,1.6117238,2.7430124,3.872488,5.0019636,6.1332526,7.262728,8.528176,9.791811,11.057259,12.322706,13.588155,13.932617,14.277081,14.623356,14.967819,15.312282,13.981567,12.652666,11.321951,9.99305,8.662335,8.861761,9.063,9.262425,9.461852,9.663091,9.373016,9.082943,8.792869,8.502794,8.212721,7.752228,7.2917356,6.833056,6.3725634,5.9120708,5.0944247,4.2767787,3.4591327,2.6432993,1.8256533,2.4021754,2.9805105,3.5570326,4.135368,4.7118897,4.7916603,4.8732433,4.953014,5.032784,5.1125546,4.592234,4.071914,3.5515938,3.0330863,2.5127661,2.374981,2.2371957,2.0994108,1.9616255,1.8256533,1.7821422,1.7404441,1.696933,1.6552348,1.6117238,1.5772774,1.5428312,1.5083848,1.4721256,1.4376793,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.092461094,0.15954071,0.22662032,0.2955129,0.36259252,0.4949388,0.62728506,0.75963134,0.8919776,1.0243238,1.2382535,1.4503701,1.6624867,1.8746033,2.08672,2.2970235,2.5073273,2.7176309,2.9279346,3.1382382,3.1074178,3.0765975,3.04759,3.0167696,2.9877625,2.5580902,2.128418,1.696933,1.2672608,0.8375887,0.99712944,1.1566701,1.3180238,1.4775645,1.6371052,1.8329052,2.0268922,2.222692,2.4166791,2.612479,2.7992141,2.9877625,3.1744974,3.3630457,3.5497808,3.3775494,3.2053177,3.0330863,2.8608549,2.6868105,2.3532255,2.0178273,1.6824293,1.3470312,1.0116332,0.90285534,0.79226464,0.68167394,0.5728962,0.46230546,0.3825351,0.30276474,0.2229944,0.14322405,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.0025684,2.0051367,3.007705,4.0102735,5.0128417,4.664753,4.3166637,3.9703882,3.6222992,3.2742105,3.0820365,2.8898623,2.6976883,2.5055144,2.3133402,2.7919624,3.2723975,3.7528327,4.233268,4.7118897,3.7981565,2.8826106,1.9670644,1.0533313,0.13778515,0.11421664,0.092461094,0.07070554,0.047137026,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.11421664,0.1794833,0.24474995,0.3100166,0.37528324,0.44961473,0.52575916,0.6000906,0.6744221,0.7505665,0.8466535,0.9445535,1.0424535,1.1403534,1.2382535,1.0877775,0.93730164,0.7868258,0.63816285,0.48768693,0.5166943,0.5475147,0.57833505,0.6073425,0.63816285,0.63816285,0.63816285,0.63816285,0.63816285,0.63816285,0.6000906,0.5620184,0.52575916,0.48768693,0.44961473,0.533011,0.61459434,0.6979906,0.7795739,0.8629702,0.7016165,0.5420758,0.3825351,0.2229944,0.06164073,0.19942589,0.33721104,0.4749962,0.61278135,0.7505665,0.61459434,0.48043507,0.3444629,0.21030366,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.14322405,0.28463513,0.42785916,0.56927025,0.7124943,0.5747091,0.43692398,0.2991388,0.16316663,0.025381476,0.045324065,0.065266654,0.08520924,0.10515183,0.12509441,0.3245203,0.52575916,0.72518504,0.9246109,1.1258497,0.89922947,0.6744221,0.44961473,0.22480737,0.0,0.37528324,0.7505665,1.1258497,1.49932,1.8746033,1.8202144,1.7658255,1.7096237,1.6552348,1.6008459,1.4703126,1.3397794,1.209246,1.0805258,0.9499924,2.2371957,3.5243993,4.8134155,6.1006193,7.3878226,6.48678,5.5875506,4.688321,3.787279,2.8880494,2.4094272,1.9326181,1.455809,0.97718686,0.50037766,0.97537386,1.4503701,1.9253663,2.4003625,2.8753586,3.1219215,3.3702974,3.6168604,3.8652363,4.1117992,3.290527,2.467442,1.6443571,0.823085,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.16497959,0.32995918,0.4949388,0.65991837,0.824898,1.1530442,1.4793775,1.8075237,2.13567,2.4620032,2.6541772,2.8481643,3.0403383,3.2325122,3.4246864,4.1317415,4.84061,5.5476656,6.2547207,6.9617763,5.7869763,4.612177,3.437377,2.2625773,1.0877775,1.0750868,1.062396,1.0497054,1.0370146,1.0243238,0.9554313,0.88472575,0.81583315,0.7451276,0.6744221,0.61459434,0.55476654,0.4949388,0.43511102,0.37528324,0.33177215,0.29007402,0.24837588,0.20486477,0.16316663,0.2229944,0.28282216,0.34264994,0.40247768,0.46230546,1.2219368,1.9815681,2.7430124,3.5026438,4.262275,4.632119,5.0019636,5.371808,5.7416525,6.11331,5.4606433,4.8079767,4.15531,3.5026438,2.8499773,2.5091403,2.1701162,1.8292793,1.4902552,1.1494182,0.94274056,0.73424983,0.5275721,0.3208944,0.11240368,0.34990177,0.5873999,0.824898,1.062396,1.2998942,1.064209,0.83033687,0.5946517,0.36077955,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.13959812,0.27919623,0.42060733,0.56020546,0.69980353,0.5855869,0.46955732,0.35534066,0.23931105,0.12509441,0.21936847,0.3154555,0.40972954,0.5058166,0.6000906,0.5402629,0.48043507,0.42060733,0.36077955,0.2991388,0.3444629,0.38978696,0.43511102,0.48043507,0.52575916,0.5946517,0.6653573,0.73424983,0.80495536,0.87566096,2.2516994,3.6295512,5.0074024,6.3852544,7.763106,8.158332,8.551744,8.94697,9.342196,9.737422,9.539809,9.342196,9.144584,8.94697,8.749357,8.089439,7.4295206,6.7696023,6.109684,5.4497657,5.3029156,5.1542525,5.0074024,4.860553,4.7118897,5.411693,6.11331,6.813113,7.512917,8.212721,8.778365,9.342196,9.907841,10.471672,11.037316,10.734551,10.431787,10.130835,9.82807,9.525306,9.9966755,10.469859,10.943042,11.4144125,11.887595,12.659918,13.43224,14.204562,14.976884,15.749206,15.544341,15.339477,15.134612,14.929747,14.724882,12.540262,10.355642,8.1692095,5.9845896,3.7999697,3.3304121,2.8608549,2.3894846,1.9199274,1.4503701,2.4456866,3.43919,4.4345064,5.429823,6.4251394,7.498413,8.569874,9.643148,10.714609,11.787883,12.442362,13.096842,13.753134,14.407614,15.062093,14.066776,13.073273,12.077957,11.082641,10.087324,10.625773,11.162411,11.700861,12.237497,12.774135,12.627284,12.480434,12.331772,12.184921,12.038072,11.285692,10.5315,9.77912,9.026741,8.274362,7.0542374,5.8341136,4.615803,3.395679,2.175555,3.04759,3.919625,4.7916603,5.6655083,6.5375433,6.532104,6.526665,6.5230393,6.5176005,6.5121617,5.719897,4.9276323,4.135368,3.343103,2.5508385,2.4620032,2.374981,2.2879589,2.1991236,2.1121013,2.030518,1.9471219,1.8655385,1.7821422,1.7005589,1.647983,1.5954071,1.5428312,1.4902552,1.4376793,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.065266654,0.11784257,0.17041849,0.2229944,0.2755703,0.48587397,0.69436467,0.90466833,1.114972,1.3252757,1.5373923,1.7495089,1.9616255,2.175555,2.3876717,2.6052272,2.8227828,3.0403383,3.2578938,3.4754493,3.2597067,3.045777,2.8300345,2.6142921,2.4003625,2.0975976,1.794833,1.4920682,1.1893034,0.8883517,1.1040943,1.3216497,1.5392052,1.7567607,1.9743162,2.2100015,2.4456866,2.6795588,2.9152439,3.149116,3.3122826,3.4754493,3.636803,3.7999697,3.9631362,3.7455807,3.5280252,3.3104696,3.092914,2.8753586,2.5073273,2.1392958,1.7730774,1.405046,1.0370146,0.9445535,0.8520924,0.75963134,0.6671702,0.5747091,0.47318324,0.36984438,0.26831847,0.16497959,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.2817645,2.565342,3.8471067,5.130684,6.412449,5.995467,5.576673,5.1596913,4.74271,4.325729,3.8978696,3.4700103,3.0421512,2.6142921,2.1882458,2.8390994,3.491766,4.1444325,4.797099,5.4497657,4.3801174,3.3104696,2.2408218,1.1693609,0.099712946,0.08339628,0.065266654,0.047137026,0.030820364,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.11965553,0.21574254,0.3100166,0.40429065,0.50037766,0.6000906,0.69980353,0.7995165,0.89922947,1.0007553,1.1294757,1.260009,1.3905423,1.5192627,1.649796,1.4503701,1.2491312,1.0497054,0.85027945,0.6508536,0.69073874,0.7306239,0.7705091,0.8103943,0.85027945,0.85027945,0.85027945,0.85027945,0.85027945,0.85027945,0.7995165,0.7505665,0.69980353,0.6508536,0.6000906,0.6852999,0.7705091,0.8557183,0.93911463,1.0243238,0.8321498,0.6399758,0.44780177,0.25562772,0.06164073,0.25018883,0.43692398,0.62547207,0.8122072,1.0007553,0.8194591,0.6399758,0.4604925,0.27919623,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.19036107,0.38072214,0.56927025,0.75963134,0.9499924,0.76325727,0.5747091,0.387974,0.19942589,0.012690738,0.02175555,0.032633327,0.04169814,0.052575916,0.06164073,0.16316663,0.26287958,0.36259252,0.46230546,0.5620184,0.44961473,0.33721104,0.22480737,0.11240368,0.0,0.50037766,1.0007553,1.49932,1.9996977,2.5000753,2.3097143,2.1193533,1.9308052,1.7404441,1.550083,1.3597219,1.1693609,0.9808127,0.7904517,0.6000906,2.175555,3.7492065,5.3246713,6.9001355,8.4756,7.4875355,6.4994707,5.5132194,4.5251546,3.53709,2.9424384,2.3477864,1.7531348,1.1566701,0.5620184,1.2128719,1.8619126,2.5127661,3.1618068,3.8126602,4.1426196,4.4725785,4.802538,5.132497,5.462456,4.36924,3.2778363,2.18462,1.0932164,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.21936847,0.4405499,0.65991837,0.8792868,1.1004683,1.4830034,1.8655385,2.2480736,2.6306088,3.0131438,3.1781235,3.343103,3.5080826,3.673062,3.8380418,4.572292,5.3083544,6.0426044,6.776854,7.512917,6.300045,5.087173,3.874301,2.663242,1.4503701,1.4249886,1.3996071,1.3742256,1.3506571,1.3252757,1.2400664,1.1548572,1.0696479,0.98443866,0.89922947,0.8194591,0.73968875,0.65991837,0.58014804,0.50037766,0.43511102,0.36984438,0.3045777,0.23931105,0.17585737,0.23024625,0.28463513,0.34083697,0.39522585,0.44961473,1.4920682,2.5345216,3.576975,4.6194286,5.661882,5.810545,5.957395,6.104245,6.2529078,6.399758,5.8177967,5.235836,4.652062,4.070101,3.48814,3.0167696,2.5472124,2.077655,1.6080978,1.1367276,0.93911463,0.7433147,0.54570174,0.3480888,0.15047589,0.33721104,0.52575916,0.7124943,0.89922947,1.0877775,0.88291276,0.678048,0.47318324,0.26831847,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.07070554,0.13959812,0.21030366,0.27919623,0.34990177,0.291887,0.23568514,0.17767033,0.11965553,0.06164073,0.11059072,0.15772775,0.20486477,0.2520018,0.2991388,0.27013144,0.23931105,0.21030366,0.1794833,0.15047589,0.25925365,0.36984438,0.48043507,0.58921283,0.69980353,0.73424983,0.7705091,0.80495536,0.83940166,0.87566096,2.3568513,3.8398547,5.3228583,6.8058615,8.287052,9.171778,10.058316,10.943042,11.827768,12.712494,12.308203,11.9021,11.497808,11.091705,10.687414,9.432844,8.178274,6.921891,5.667321,4.4127507,4.7191415,5.027345,5.335549,5.6419396,5.9501433,6.624565,7.3008003,7.9752226,8.649645,9.325879,9.382081,9.440096,9.498111,9.554313,9.612328,9.804502,9.9966755,10.190662,10.382836,10.57501,10.866898,11.160598,11.452485,11.744371,12.038072,13.267261,14.498261,15.72745,16.956638,18.187641,17.897566,17.607492,17.31742,17.027344,16.73727,13.981567,11.227677,8.471974,5.718084,2.962381,2.6269827,2.2933977,1.9579996,1.6226015,1.2872034,2.1483607,3.007705,3.8670492,4.7282066,5.5875506,6.4668374,7.3479376,8.227224,9.108324,9.987611,10.952107,11.918416,12.882912,13.847408,14.811904,14.151986,13.492067,12.8321495,12.172231,11.512312,12.387974,13.261822,14.137483,15.013144,15.8869915,15.883366,15.877926,15.872487,15.867048,15.863422,14.817343,13.773077,12.726997,11.682731,10.636651,9.01405,7.3914485,5.77066,4.1480584,2.525457,3.6930048,4.860553,6.0281005,7.1956487,8.363196,8.272549,8.1819,8.093065,8.002417,7.911769,6.8475595,5.7815375,4.7173285,3.6531196,2.5870976,2.5508385,2.5127661,2.474694,2.4366217,2.4003625,2.277081,2.1556125,2.032331,1.9108626,1.7875811,1.7168756,1.647983,1.5772774,1.5083848,1.4376793,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.4749962,0.76325727,1.0497054,1.3379664,1.6244144,1.8383441,2.0504606,2.2625773,2.474694,2.6868105,2.911618,3.1382382,3.3630457,3.587853,3.8126602,3.4119956,3.0131438,2.612479,2.2118144,1.8129625,1.6371052,1.4630609,1.2872034,1.1131591,0.93730164,1.2128719,1.4866294,1.7621996,2.03777,2.3133402,2.5870976,2.8626678,3.1382382,3.4119956,3.6875658,3.825351,3.9631362,4.099108,4.2368937,4.3746786,4.1117992,3.8507326,3.587853,3.3249733,3.0620937,2.663242,2.2625773,1.8619126,1.4630609,1.062396,0.9880646,0.9119202,0.8375887,0.76325727,0.6871128,0.5620184,0.43692398,0.31182957,0.18673515,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.5627737,3.1255474,4.688321,6.249282,7.8120556,7.324369,6.836682,6.350808,5.863121,5.375434,4.7118897,4.0501585,3.386614,2.7248828,2.0631514,2.8880494,3.7129474,4.537845,5.3627434,6.187641,4.9620786,3.738329,2.5127661,1.2872034,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.12509441,0.25018883,0.37528324,0.50037766,0.62547207,0.7505665,0.87566096,1.0007553,1.1258497,1.2491312,1.4122978,1.5754645,1.7368182,1.8999848,2.0631514,1.8129625,1.5627737,1.3125849,1.062396,0.8122072,0.8629702,0.9119202,0.96268314,1.0116332,1.062396,1.062396,1.062396,1.062396,1.062396,1.062396,1.0007553,0.93730164,0.87566096,0.8122072,0.7505665,0.8375887,0.9246109,1.0116332,1.1004683,1.1874905,0.96268314,0.73787576,0.51306844,0.28826106,0.06164073,0.2991388,0.53663695,0.774135,1.0116332,1.2491312,1.0243238,0.7995165,0.5747091,0.34990177,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.2374981,0.4749962,0.7124943,0.9499924,1.1874905,0.9499924,0.7124943,0.4749962,0.2374981,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.62547207,1.2491312,1.8746033,2.5000753,3.1255474,2.7992141,2.474694,2.1501737,1.8256533,1.49932,1.2491312,1.0007553,0.7505665,0.50037766,0.25018883,2.1121013,3.975827,5.8377395,7.699652,9.563377,8.488291,7.413204,6.338117,5.2630305,4.1879435,3.4754493,2.762955,2.0504606,1.3379664,0.62547207,1.4503701,2.275268,3.100166,3.925064,4.749962,5.163317,5.57486,5.9882154,6.399758,6.813113,5.4497657,4.0882306,2.7248828,1.3633479,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.2755703,0.5493277,0.824898,1.1004683,1.3742256,1.8129625,2.2498865,2.6868105,3.1255474,3.5624714,3.7002566,3.8380418,3.975827,4.1117992,4.249584,5.0128417,5.774286,6.5375433,7.3008003,8.062244,6.813113,5.562169,4.313038,3.0620937,1.8129625,1.7748904,1.7368182,1.7005589,1.6624867,1.6244144,1.5247015,1.4249886,1.3252757,1.2255627,1.1258497,1.0243238,0.9246109,0.824898,0.72518504,0.62547207,0.53663695,0.44961473,0.36259252,0.2755703,0.18673515,0.2374981,0.28826106,0.33721104,0.387974,0.43692398,1.7621996,3.0874753,4.4127507,5.7380266,7.063302,6.987158,6.9128265,6.836682,6.7623506,6.688019,6.1749506,5.661882,5.1506267,4.6375585,4.12449,3.5243993,2.9243085,2.324218,1.7241274,1.1258497,0.93730164,0.7505665,0.5620184,0.37528324,0.18673515,0.3245203,0.46230546,0.6000906,0.73787576,0.87566096,0.69980353,0.52575916,0.34990177,0.17585737,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.17585737,0.34990177,0.52575916,0.69980353,0.87566096,0.87566096,0.87566096,0.87566096,0.87566096,0.87566096,2.4620032,4.0501585,5.638314,7.224656,8.812811,10.1870365,11.563075,12.937301,14.313339,15.687565,15.074784,14.462003,13.849221,13.238253,12.625471,10.774437,8.925215,7.07418,5.224958,3.3757362,4.137181,4.900438,5.661882,6.4251394,7.1883965,7.837437,8.488291,9.137331,9.788185,10.437225,9.987611,9.537996,9.088382,8.636953,8.187339,8.874452,9.563377,10.25049,10.937603,11.624716,11.73712,11.849524,11.961927,12.07433,12.186734,13.874602,15.56247,17.25034,18.938208,20.624262,20.250792,19.87551,19.500225,19.124943,18.749659,15.4246855,12.099712,8.774739,5.4497657,2.124792,1.9253663,1.7241274,1.5247015,1.3252757,1.1258497,1.8492218,2.5744069,3.299592,4.024777,4.749962,5.4370747,6.1241875,6.813113,7.500226,8.187339,9.461852,10.738177,12.012691,13.287203,14.561715,14.237195,13.912675,13.588155,13.261822,12.937301,14.150173,15.363045,16.575916,17.786976,18.999847,19.137632,19.275417,19.413204,19.549175,19.68696,18.350807,17.01284,15.674874,14.336908,13.000754,10.975676,8.950596,6.925517,4.900438,2.8753586,4.3384194,5.7996674,7.262728,8.725789,10.1870365,10.012992,9.837135,9.663091,9.487233,9.313189,7.9752226,6.637256,5.2992897,3.9631362,2.6251698,2.6378605,2.6505513,2.663242,2.6741197,2.6868105,2.525457,2.3622901,2.1991236,2.03777,1.8746033,1.7875811,1.7005589,1.6117238,1.5247015,1.4376793,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.38072214,0.6091554,0.83940166,1.0696479,1.2998942,1.4920682,1.6842422,1.8782293,2.0704033,2.2625773,2.5290828,2.7974012,3.0657198,3.3322253,3.6005437,3.2778363,2.955129,2.6324217,2.3097143,1.987007,1.794833,1.6026589,1.4104849,1.2183108,1.0243238,1.214685,1.405046,1.5954071,1.7857682,1.9743162,2.222692,2.469255,2.7176309,2.9641938,3.2125697,3.3648586,3.5171473,3.6694362,3.8217251,3.975827,3.6766882,3.3793623,3.0820365,2.7847104,2.4873846,2.1701162,1.8528478,1.5355793,1.2183108,0.89922947,0.8466535,0.79589057,0.7433147,0.69073874,0.63816285,0.52032024,0.40247768,0.28463513,0.16679256,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.2491312,2.5000753,3.7492065,5.0001507,6.249282,5.859495,5.469708,5.0799212,4.690134,4.3003473,3.785466,3.2705846,2.7557032,2.2408218,1.7241274,2.3695421,3.0149567,3.6603715,4.305786,4.949388,4.1081734,3.2651455,2.422118,1.5790904,0.73787576,1.017072,1.2980812,1.5772774,1.8582866,2.137483,1.789394,1.4431182,1.0950294,0.7469406,0.40066472,0.3208944,0.23931105,0.15954071,0.07977036,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.099712946,0.19942589,0.2991388,0.40066472,0.50037766,0.63816285,0.774135,0.9119202,1.0497054,1.1874905,1.3270886,1.4666867,1.6080978,1.7476959,1.887294,1.7476959,1.6080978,1.4666867,1.3270886,1.1874905,1.3742256,1.5627737,1.7495089,1.938057,2.124792,2.229944,2.335096,2.4402475,2.5453994,2.6505513,2.3006494,1.9507477,1.6008459,1.2491312,0.89922947,0.9101072,0.91917205,0.9300498,0.93911463,0.9499924,0.78319985,0.61459434,0.44780177,0.27919623,0.11240368,0.29007402,0.46774435,0.64541465,0.823085,1.0007553,0.8194591,0.6399758,0.4604925,0.27919623,0.099712946,0.0870222,0.07433146,0.06164073,0.05076295,0.038072214,0.21936847,0.40247768,0.5855869,0.7668832,0.9499924,0.75963134,0.56927025,0.38072214,0.19036107,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.047137026,0.08339628,0.11784257,0.15228885,0.18673515,0.27013144,0.35171473,0.43511102,0.5166943,0.6000906,1.0732739,1.5446441,2.0178273,2.4891977,2.962381,2.6469254,2.333283,2.0178273,1.7023718,1.3869164,1.2980812,1.2074331,1.1167849,1.0279498,0.93730164,2.9369993,4.936697,6.9382076,8.937905,10.937603,9.514427,8.093065,6.6698895,5.2467136,3.825351,3.1799364,2.5345216,1.889107,1.2455053,0.6000906,1.4666867,2.335096,3.2016919,4.070101,4.936697,5.040036,5.143375,5.2449007,5.3482394,5.4497657,4.360175,3.2705846,2.179181,1.0895905,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.3208944,0.5148814,0.7106813,0.90466833,1.1004683,1.6407311,2.179181,2.7194438,3.2597067,3.7999697,4.004834,4.209699,4.4145637,4.6194286,4.8242936,5.315606,5.805106,6.294606,6.784106,7.2754188,6.301858,5.33011,4.358362,3.3848011,2.4130533,2.2897718,2.1683033,2.0450218,1.9217403,1.8002719,1.6207886,1.4394923,1.260009,1.0805258,0.89922947,0.8194591,0.73968875,0.65991837,0.58014804,0.50037766,0.42967212,0.36077955,0.29007402,0.21936847,0.15047589,0.2030518,0.25562772,0.30820364,0.36077955,0.41335547,1.6008459,2.7883365,3.975827,5.163317,6.350808,6.5756154,6.8004227,7.02523,7.250037,7.474845,6.985345,6.495845,6.004532,5.5150323,5.0255322,4.2604623,3.4953918,2.7303216,1.9652514,1.2001812,0.99712944,0.79589057,0.59283876,0.38978696,0.18673515,0.29732585,0.40791658,0.5166943,0.62728506,0.73787576,0.58921283,0.44236287,0.2955129,0.14684997,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.11784257,0.23568514,0.35171473,0.46955732,0.5873999,0.61278135,0.63816285,0.66173136,0.6871128,0.7124943,0.7451276,0.7777609,0.8103943,0.8430276,0.87566096,2.275268,3.6748753,5.0744824,6.4759026,7.8755093,9.079316,10.284937,11.490557,12.694364,13.899984,13.406858,12.915545,12.42242,11.929294,11.437981,10.239613,9.043057,7.844689,6.6481338,5.4497657,5.810545,6.169512,6.530291,6.889258,7.250037,7.8229337,8.39583,8.966913,9.539809,10.112705,9.527119,8.943344,8.357758,7.7721705,7.1865835,7.6851482,8.1819,8.680465,9.177217,9.675781,10.025683,10.375585,10.725487,11.075388,11.42529,13.055143,14.684997,16.31485,17.944704,19.574556,19.17933,18.784105,18.390692,17.995466,17.60024,14.614291,11.630155,8.644206,5.660069,2.6741197,2.3550384,2.034144,1.7150626,1.3941683,1.0750868,1.987007,2.9007401,3.8126602,4.7245803,5.638314,6.247469,6.8566246,7.4675927,8.076748,8.6877165,9.735609,10.783502,11.829581,12.877473,13.925365,13.544643,13.165734,12.785012,12.40429,12.025381,13.274512,14.525456,15.774588,17.025532,18.274662,18.305483,18.33449,18.36531,18.394318,18.425138,17.112555,15.799969,14.487384,13.174799,11.862214,10.323009,8.781991,7.2427855,5.7017674,4.162562,5.0980506,6.0317264,6.967215,7.902704,8.838193,8.892582,8.94697,9.003172,9.057561,9.11195,7.7903004,6.4668374,5.145188,3.8217251,2.5000753,2.6378605,2.7756457,2.911618,3.049403,3.1871881,3.045777,2.902553,2.759329,2.617918,2.474694,2.2607644,2.0450218,1.8292793,1.6153497,1.3996071,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.28463513,0.45686656,0.629098,0.8031424,0.97537386,1.1476053,1.3198367,1.4920682,1.6642996,1.8383441,2.1483607,2.4583774,2.7683938,3.0765975,3.386614,3.141864,2.8971143,2.6523643,2.4076142,2.1628644,1.9525607,1.742257,1.5319533,1.3216497,1.1131591,1.2183108,1.3216497,1.4268016,1.5319533,1.6371052,1.8582866,2.077655,2.2970235,2.518205,2.7375734,2.904366,3.0729716,3.2397642,3.4083695,3.5751622,3.24339,2.909805,2.5780327,2.2444477,1.9126755,1.6769904,1.4431182,1.2074331,0.97174793,0.73787576,0.7070554,0.678048,0.64722764,0.61822027,0.5873999,0.47680917,0.3680314,0.2574407,0.14684997,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.93730164,1.8746033,2.811905,3.7492065,4.688321,4.3946214,4.102734,3.8108473,3.5171473,3.2252605,2.857229,2.4891977,2.1229792,1.7549478,1.3869164,1.8528478,2.3169663,2.7828975,3.247016,3.7129474,3.2524548,2.7919624,2.333283,1.8727903,1.4122978,1.9851941,2.5580902,3.1291735,3.7020695,4.274966,3.5806012,2.8844235,2.1900587,1.4956942,0.7995165,0.6399758,0.48043507,0.3208944,0.15954071,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07433146,0.15047589,0.22480737,0.2991388,0.37528324,0.52575916,0.6744221,0.824898,0.97537386,1.1258497,1.2418793,1.3597219,1.4775645,1.5954071,1.7132497,1.6824293,1.651609,1.6226015,1.5917811,1.5627737,1.887294,2.2118144,2.5381477,2.8626678,3.1871881,3.397492,3.6077955,3.8180993,4.028403,4.2368937,3.6005437,2.962381,2.324218,1.6878681,1.0497054,0.9826257,0.9155461,0.8466535,0.7795739,0.7124943,0.60190356,0.49312583,0.3825351,0.27194437,0.16316663,0.27919623,0.39703882,0.5148814,0.6327239,0.7505665,0.61459434,0.48043507,0.3444629,0.21030366,0.07433146,0.07433146,0.07433146,0.07433146,0.07433146,0.07433146,0.2030518,0.32995918,0.45686656,0.5855869,0.7124943,0.56927025,0.42785916,0.28463513,0.14322405,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.09427405,0.16497959,0.23568514,0.3045777,0.37528324,0.5402629,0.70524246,0.87022203,1.0352017,1.2001812,1.5192627,1.840157,2.1592383,2.4801328,2.7992141,2.4946365,2.1900587,1.8854811,1.5790904,1.2745126,1.3452182,1.4141108,1.4848163,1.5555218,1.6244144,3.7618973,5.89938,8.036863,10.174346,12.311829,10.542377,8.772926,7.0016613,5.23221,3.4627585,2.8844235,2.3079014,1.7295663,1.1530442,0.5747091,1.4848163,2.3949237,3.3050308,4.215138,5.125245,4.9167547,4.710077,4.501586,4.2949085,4.0882306,3.2705846,2.4529383,1.6352923,0.81764615,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,0.36440548,0.48043507,0.5946517,0.7106813,0.824898,1.4666867,2.1102884,2.752077,3.395679,4.0374675,4.309412,4.5831695,4.855114,5.127058,5.4008155,5.618371,5.8341136,6.051669,6.2692246,6.48678,5.7924156,5.0980506,4.401873,3.7075086,3.0131438,2.8046532,2.5979755,2.3894846,2.182807,1.9743162,1.7150626,1.455809,1.1947423,0.9354887,0.6744221,0.61459434,0.55476654,0.4949388,0.43511102,0.37528324,0.32270733,0.27013144,0.21755551,0.16497959,0.11240368,0.16679256,0.2229944,0.27738327,0.33177215,0.387974,1.4376793,2.4873846,3.53709,4.5867953,5.638314,6.16226,6.688019,7.211965,7.7377243,8.26167,7.795739,7.327995,6.8602505,6.392506,5.924762,4.994712,4.064662,3.1346123,2.2045624,1.2745126,1.0569572,0.83940166,0.62184614,0.40429065,0.18673515,0.27013144,0.35171473,0.43511102,0.5166943,0.6000906,0.48043507,0.36077955,0.23931105,0.11965553,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.23568514,0.46955732,0.70524246,0.93911463,1.1747998,1.0497054,0.9246109,0.7995165,0.6744221,0.5493277,0.61459434,0.67986095,0.7451276,0.8103943,0.87566096,2.08672,3.299592,4.512464,5.7253356,6.9382076,7.9734097,9.006798,10.042,11.077202,12.112403,11.740746,11.367275,10.995618,10.622148,10.25049,9.704789,9.1609,8.615198,8.069496,7.5256076,7.4820967,7.440398,7.3968873,7.3551893,7.311678,7.8084297,8.303369,8.798307,9.293246,9.788185,9.066626,8.34688,7.6271334,6.9073873,6.187641,6.495845,6.8022356,7.1104393,7.41683,7.7250338,8.312433,8.899834,9.487233,10.074633,10.662033,12.235684,13.807523,15.379361,16.953012,18.52485,18.109684,17.694515,17.279346,16.864178,16.450823,13.80571,11.160598,8.515485,5.870373,3.2252605,2.7847104,2.3441606,1.9054236,1.4648738,1.0243238,2.124792,3.2252605,4.325729,5.424384,6.5248523,7.057863,7.590874,8.122072,8.655084,9.188094,10.007553,10.827013,11.648285,12.467744,13.287203,12.852092,12.416981,11.98187,11.546759,11.111648,12.400664,13.687867,14.975071,16.262274,17.549479,17.473333,17.395376,17.31742,17.239462,17.163317,15.8743,14.587097,13.299893,12.012691,10.725487,9.670342,8.615198,7.560054,6.5049095,5.4497657,5.857682,6.265599,6.6717024,7.079619,7.4875355,7.7721705,8.056806,8.343254,8.627889,8.912524,7.605378,6.298232,4.989273,3.682127,2.374981,2.6378605,2.9007401,3.1618068,3.4246864,3.6875658,3.5642843,3.442816,3.3195345,3.198066,3.0747845,2.7321346,2.3894846,2.0468347,1.7041848,1.3633479,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.07433146,0.07433146,0.07433146,0.07433146,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.19036107,0.3045777,0.42060733,0.53482395,0.6508536,0.8031424,0.9554313,1.1077201,1.260009,1.4122978,1.7658255,2.1175404,2.469255,2.8227828,3.1744974,3.007705,2.8390994,2.6723068,2.5055144,2.3369088,2.1102884,1.8818551,1.6552348,1.4268016,1.2001812,1.2201238,1.2400664,1.260009,1.2799516,1.2998942,1.4920682,1.6842422,1.8782293,2.0704033,2.2625773,2.4456866,2.6269827,2.810092,2.9932013,3.1744974,2.808279,2.4402475,2.0722163,1.7041848,1.3379664,1.1856775,1.0333886,0.8792868,0.726998,0.5747091,0.56745726,0.56020546,0.5529536,0.54570174,0.53663695,0.43511102,0.33177215,0.23024625,0.12690738,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.62547207,1.2491312,1.8746033,2.5000753,3.1255474,2.9297476,2.7357605,2.5399606,2.3441606,2.1501737,1.9308052,1.7096237,1.4902552,1.2708868,1.0497054,1.3343405,1.6207886,1.9054236,2.1900587,2.474694,2.3967366,2.3205922,2.2426348,2.1646774,2.08672,2.953316,3.8180993,4.6828823,5.5476656,6.412449,5.369995,4.327542,3.2850883,2.2426348,1.2001812,0.96087015,0.7197462,0.48043507,0.23931105,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,0.41335547,0.5747091,0.73787576,0.89922947,1.062396,1.1566701,1.2527572,1.3470312,1.4431182,1.5373923,1.6171626,1.696933,1.7767034,1.8582866,1.938057,2.4003625,2.8626678,3.3249733,3.787279,4.249584,4.5650396,4.880495,5.1941376,5.5095935,5.825049,4.900438,3.975827,3.049403,2.124792,1.2001812,1.0551442,0.9101072,0.7650702,0.6200332,0.4749962,0.4224203,0.36984438,0.31726846,0.26469254,0.21211663,0.27013144,0.32814622,0.38434806,0.44236287,0.50037766,0.40972954,0.3208944,0.23024625,0.13959812,0.05076295,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.18492219,0.2574407,0.32995918,0.40247768,0.4749962,0.38072214,0.28463513,0.19036107,0.09427405,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.14322405,0.24837588,0.35171473,0.45686656,0.5620184,0.8103943,1.0569572,1.305333,1.551896,1.8002719,1.9670644,2.13567,2.3024626,2.469255,2.6378605,2.3423476,2.0468347,1.7531348,1.4576219,1.162109,1.3923552,1.6226015,1.8528478,2.0830941,2.3133402,4.5867953,6.8620634,9.137331,11.4126,13.687867,11.570327,9.452786,7.3352466,5.217706,3.100166,2.5907235,2.079468,1.5700256,1.0605831,0.5493277,1.502946,2.4547513,3.4083695,4.360175,5.3119802,4.795286,4.2767787,3.7600844,3.24339,2.7248828,2.179181,1.6352923,1.0895905,0.54570174,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07433146,0.15047589,0.22480737,0.2991388,0.37528324,0.40972954,0.44417584,0.48043507,0.5148814,0.5493277,1.2944553,2.039583,2.7847104,3.529838,4.274966,4.615803,4.954827,5.295664,5.634688,5.975525,5.919323,5.864934,5.810545,5.754343,5.6999545,5.282973,4.8641787,4.4471974,4.0302157,3.6132345,3.3195345,3.0276475,2.7357605,2.4420607,2.1501737,1.8093367,1.4703126,1.1294757,0.7904517,0.44961473,0.40972954,0.36984438,0.32995918,0.29007402,0.25018883,0.21574254,0.1794833,0.14503701,0.11059072,0.07433146,0.13234627,0.19036107,0.24837588,0.3045777,0.36259252,1.2745126,2.1882458,3.100166,4.0120864,4.9258194,5.750717,6.5756154,7.400513,8.225411,9.050309,8.604321,8.160145,7.7141557,7.26998,6.825804,5.730775,4.6357455,3.540716,2.4456866,1.3506571,1.1167849,0.88472575,0.6526665,0.42060733,0.18673515,0.24293698,0.29732585,0.35171473,0.40791658,0.46230546,0.36984438,0.27738327,0.18492219,0.092461094,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.35171473,0.70524246,1.0569572,1.4104849,1.7621996,1.4866294,1.2128719,0.93730164,0.66173136,0.387974,0.48587397,0.581961,0.67986095,0.7777609,0.87566096,1.8999848,2.9243085,3.9504454,4.974769,6.000906,6.8656893,7.7304726,8.595256,9.460039,10.324821,10.07282,9.820818,9.567003,9.3150015,9.063,9.169965,9.27693,9.385707,9.492672,9.599637,9.155461,8.709473,8.265296,7.819308,7.3751316,7.7921133,8.209095,8.627889,9.04487,9.461852,8.607946,7.752228,6.8983226,6.0426044,5.186886,5.3047285,5.422571,5.540414,5.658256,5.774286,6.599184,7.424082,8.2507925,9.07569,9.900589,11.4144125,12.930049,14.445685,15.95951,17.475147,17.040035,16.604925,16.169813,15.734702,15.299591,12.995316,10.689227,8.384952,6.0806766,3.774588,3.2143826,2.6541772,2.0957847,1.5355793,0.97537386,2.2625773,3.5497808,4.836984,6.1241875,7.413204,7.8682575,8.323311,8.778365,9.231606,9.686659,10.279498,10.872336,11.465176,12.058014,12.650853,12.15954,11.67004,11.18054,10.689227,10.199727,11.525003,12.850279,14.175554,15.50083,16.824293,16.63937,16.454449,16.269526,16.084604,15.899682,14.63786,13.374225,12.112403,10.850581,9.5869465,9.017676,8.446592,7.877322,7.308052,6.736969,6.6173134,6.497658,6.378002,6.258347,6.1368785,6.6517596,7.168454,7.6833353,8.198216,8.713099,7.420456,6.1278133,4.835171,3.5425289,2.2498865,2.6378605,3.0258346,3.4119956,3.7999697,4.1879435,4.0846047,3.9830787,3.87974,3.778214,3.6748753,3.2053177,2.7357605,2.2643902,1.794833,1.3252757,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.099712946,0.099712946,0.099712946,0.099712946,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.09427405,0.15228885,0.21030366,0.26831847,0.3245203,0.45686656,0.58921283,0.72337204,0.8557183,0.9880646,1.3832904,1.7767034,2.1719291,2.5671551,2.962381,2.8717327,2.7828975,2.6922495,2.6016014,2.5127661,2.268016,2.0232663,1.7767034,1.5319533,1.2872034,1.2219368,1.1566701,1.0932164,1.0279498,0.96268314,1.1276628,1.2926424,1.4576219,1.6226015,1.7875811,1.9851941,2.182807,2.38042,2.5780327,2.7756457,2.373168,1.9706904,1.5682126,1.1657349,0.76325727,0.69255173,0.62184614,0.5529536,0.48224804,0.41335547,0.42785916,0.44236287,0.45686656,0.47318324,0.48768693,0.39159992,0.29732585,0.2030518,0.10696479,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.31182957,0.62547207,0.93730164,1.2491312,1.5627737,1.4648738,1.3669738,1.2690738,1.1729867,1.0750868,1.0025684,0.9300498,0.8575313,0.7850128,0.7124943,0.81764615,0.922798,1.0279498,1.1331016,1.2382535,1.5428312,1.8474089,2.1519866,2.4583774,2.762955,3.919625,5.0781083,6.2347784,7.3932614,8.549932,7.159389,5.77066,4.3801174,2.9895754,1.6008459,1.2799516,0.96087015,0.6399758,0.3208944,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.2991388,0.4749962,0.6508536,0.824898,1.0007553,1.0732739,1.1457924,1.2183108,1.2908293,1.3633479,1.551896,1.742257,1.9326181,2.1229792,2.3133402,2.911618,3.5117085,4.1117992,4.7118897,5.3119802,5.732588,6.153195,6.5719895,6.9925966,7.413204,6.200332,4.98746,3.774588,2.561716,1.3506571,1.1276628,0.90466833,0.68167394,0.4604925,0.2374981,0.24293698,0.24837588,0.2520018,0.2574407,0.26287958,0.25925365,0.2574407,0.25562772,0.2520018,0.25018883,0.20486477,0.15954071,0.11421664,0.07070554,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.15047589,0.16679256,0.18492219,0.2030518,0.21936847,0.2374981,0.19036107,0.14322405,0.09427405,0.047137026,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.19036107,0.32995918,0.46955732,0.6091554,0.7505665,1.0805258,1.4104849,1.7404441,2.0704033,2.4003625,2.4148662,2.42937,2.4456866,2.4601903,2.474694,2.1900587,1.9054236,1.6207886,1.3343405,1.0497054,1.4394923,1.8292793,2.220879,2.610666,3.000453,5.411693,7.8247466,10.2378,12.650853,15.062093,12.598277,10.1326475,7.667019,5.2032027,2.7375734,2.2952106,1.8528478,1.4104849,0.968122,0.52575916,1.5192627,2.514579,3.5098956,4.505212,5.5005283,4.6720047,3.8452935,3.0167696,2.1900587,1.3633479,1.0895905,0.81764615,0.54570174,0.27194437,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.099712946,0.19942589,0.2991388,0.40066472,0.50037766,0.4550536,0.40972954,0.36440548,0.3208944,0.2755703,1.1222239,1.9706904,2.817344,3.6658103,4.512464,4.9203806,5.328297,5.7344007,6.1423173,6.550234,6.2220874,5.8957543,5.567608,5.239462,4.9131284,4.7717175,4.632119,4.4925213,4.3529234,4.213325,3.834416,3.4573197,3.0802233,2.7031271,2.324218,1.9054236,1.4848163,1.064209,0.64541465,0.22480737,0.20486477,0.18492219,0.16497959,0.14503701,0.12509441,0.10696479,0.09064813,0.072518505,0.054388877,0.038072214,0.09789998,0.15772775,0.21755551,0.27738327,0.33721104,1.1131591,1.887294,2.663242,3.437377,4.213325,5.337362,6.4632115,7.5872483,8.713099,9.837135,9.414715,8.992294,8.569874,8.147454,7.7250338,6.4650245,5.2050157,3.9450066,2.6849976,1.4249886,1.1766127,0.9300498,0.68167394,0.43511102,0.18673515,0.21574254,0.24293698,0.27013144,0.29732585,0.3245203,0.25925365,0.19579996,0.13053331,0.065266654,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.46955732,0.93911463,1.4104849,1.8800422,2.3495996,1.9253663,1.49932,1.0750868,0.6508536,0.22480737,0.35534066,0.48587397,0.61459434,0.7451276,0.87566096,1.7132497,2.5508385,3.386614,4.2242026,5.0617914,5.7579694,6.452334,7.1466985,7.842876,8.537241,8.404895,8.272549,8.140202,8.007855,7.8755093,8.63514,9.394773,10.154404,10.915848,11.675479,10.827013,9.980359,9.131892,8.285239,7.4367723,7.7776093,8.116633,8.457471,8.798307,9.137331,8.147454,7.157576,6.167699,5.177821,4.1879435,4.115425,4.0429068,3.9703882,3.8978696,3.825351,4.8877473,5.9501433,7.0125394,8.074935,9.137331,10.594954,12.052575,13.510198,14.967819,16.425442,15.970387,15.515334,15.06028,14.6052265,14.150173,12.184921,10.21967,8.254418,6.2909803,4.325729,3.6458678,2.9641938,2.2843328,1.6044719,0.9246109,2.4003625,3.874301,5.3500524,6.825804,8.299743,8.676839,9.055748,9.432844,9.80994,10.1870365,10.553255,10.917661,11.282066,11.648285,12.012691,11.466989,10.9230995,10.377398,9.8316965,9.287807,10.649343,12.012691,13.374225,14.737573,16.099108,15.80722,15.515334,15.221634,14.929747,14.63786,13.399607,12.163166,10.924912,9.686659,8.450218,8.365009,8.2798,8.194591,8.109382,8.024173,7.3769445,6.7297173,6.0824895,5.4352617,4.788034,5.5331616,6.2782893,7.023417,7.7667317,8.511859,7.2355337,5.957395,4.6792564,3.4029307,2.124792,2.6378605,3.150929,3.6621845,4.175253,4.688321,4.604925,4.5233417,4.439945,4.358362,4.274966,3.6766882,3.0802233,2.4819458,1.8854811,1.2872034,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.11240368,0.22480737,0.33721104,0.44961473,0.5620184,1.0007553,1.4376793,1.8746033,2.3133402,2.7502642,2.7375734,2.7248828,2.712192,2.6995013,2.6868105,2.4257438,2.1628644,1.8999848,1.6371052,1.3742256,1.2255627,1.0750868,0.9246109,0.774135,0.62547207,0.76325727,0.89922947,1.0370146,1.1747998,1.3125849,1.5247015,1.7368182,1.9507477,2.1628644,2.374981,1.938057,1.49932,1.062396,0.62547207,0.18673515,0.19942589,0.21211663,0.22480737,0.2374981,0.25018883,0.28826106,0.3245203,0.36259252,0.40066472,0.43692398,0.34990177,0.26287958,0.17585737,0.0870222,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07433146,0.15047589,0.22480737,0.2991388,0.37528324,0.2991388,0.22480737,0.15047589,0.07433146,0.0,0.6871128,1.3742256,2.0631514,2.7502642,3.437377,4.8877473,6.338117,7.7866745,9.237044,10.687414,8.950596,7.211965,5.475147,3.738329,1.9996977,1.6008459,1.2001812,0.7995165,0.40066472,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.18673515,0.37528324,0.5620184,0.7505665,0.93730164,0.9880646,1.0370146,1.0877775,1.1367276,1.1874905,1.4866294,1.7875811,2.08672,2.3876717,2.6868105,3.4246864,4.162562,4.900438,5.638314,6.3743763,6.9001355,7.424082,7.949841,8.4756,8.999546,7.500226,6.000906,4.499773,3.000453,1.49932,1.2001812,0.89922947,0.6000906,0.2991388,0.0,0.06164073,0.12509441,0.18673515,0.25018883,0.31182957,0.25018883,0.18673515,0.12509441,0.06164073,0.0,0.0,0.0,0.0,0.0,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.2374981,0.41335547,0.5873999,0.76325727,0.93730164,1.3506571,1.7621996,2.175555,2.5870976,3.000453,2.8626678,2.7248828,2.5870976,2.4493124,2.3133402,2.03777,1.7621996,1.4866294,1.2128719,0.93730164,1.4866294,2.03777,2.5870976,3.1382382,3.6875658,6.2365913,8.78743,11.338268,13.887294,16.438131,13.6244135,10.812509,8.000604,5.186886,2.374981,1.9996977,1.6244144,1.2491312,0.87566096,0.50037766,1.5373923,2.5744069,3.6132345,4.650249,5.6872635,4.550536,3.4119956,2.275268,1.1367276,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.12509441,0.25018883,0.37528324,0.50037766,0.62547207,0.50037766,0.37528324,0.25018883,0.12509441,0.0,0.9499924,1.8999848,2.8499773,3.7999697,4.749962,5.224958,5.6999545,6.1749506,6.6499467,7.124943,6.5248523,5.924762,5.3246713,4.7245803,4.12449,4.262275,4.40006,4.537845,4.6756306,4.8116026,4.349297,3.8869917,3.4246864,2.962381,2.5000753,1.9996977,1.49932,1.0007553,0.50037766,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06164073,0.12509441,0.18673515,0.25018883,0.31182957,0.9499924,1.5881553,2.2245052,2.8626678,3.5008307,4.9258194,6.350808,7.7757964,9.200785,10.625773,10.225109,9.824444,9.425592,9.024928,8.624263,7.1992745,5.774286,4.349297,2.9243085,1.49932,1.2382535,0.97537386,0.7124943,0.44961473,0.18673515,0.18673515,0.18673515,0.18673515,0.18673515,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.5873999,1.1747998,1.7621996,2.3495996,2.9369993,2.3622901,1.7875811,1.2128719,0.63816285,0.06164073,0.22480737,0.387974,0.5493277,0.7124943,0.87566096,1.5247015,2.175555,2.8245957,3.4754493,4.12449,4.650249,5.1741953,5.6999545,6.2257137,6.7496595,6.736969,6.7242785,6.7134004,6.70071,6.688019,8.100317,9.512614,10.924912,12.337211,13.749508,12.500377,11.249433,10.000301,8.749357,7.500226,7.763106,8.024173,8.287052,8.549932,8.812811,7.686961,6.5629244,5.4370747,4.313038,3.1871881,2.9243085,2.663242,2.4003625,2.137483,1.8746033,3.1744974,4.4743915,5.774286,7.07418,8.375887,9.775495,11.175101,12.574709,13.974316,15.375735,14.90074,14.425743,13.9507475,13.475751,13.000754,11.374527,9.750113,8.125698,6.4994707,4.8750563,4.07554,3.2742105,2.474694,1.6751775,0.87566096,2.5381477,4.2006345,5.863121,7.5256076,9.188094,9.487233,9.788185,10.087324,10.388275,10.687414,10.825199,10.962985,11.10077,11.236742,11.374527,10.774437,10.174346,9.574255,8.974165,8.375887,9.775495,11.175101,12.574709,13.974316,15.375735,14.975071,14.574407,14.175554,13.77489,13.374225,12.163166,10.950294,9.737422,8.52455,7.311678,7.7123427,8.113008,8.511859,8.912524,9.313189,8.136576,6.9617763,5.7869763,4.612177,3.437377,4.4127507,5.388125,6.3616858,7.3370595,8.312433,7.0506115,5.7869763,4.5251546,3.2633326,1.9996977,2.6378605,3.2742105,3.9123733,4.550536,5.186886,5.125245,5.0617914,5.0001507,4.936697,4.8750563,4.1498713,3.4246864,2.6995013,1.9743162,1.2491312,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.099712946,0.099712946,0.099712946,0.099712946,0.099712946,0.08339628,0.065266654,0.047137026,0.030820364,0.012690738,0.018129626,0.02175555,0.027194439,0.032633327,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.09064813,0.1794833,0.27013144,0.36077955,0.44961473,0.7995165,1.1494182,1.49932,1.8492218,2.1991236,2.2027495,2.2045624,2.2081885,2.2100015,2.2118144,2.0903459,1.9670644,1.845596,1.7223145,1.6008459,1.4304274,1.260009,1.0895905,0.91917205,0.7505665,0.872035,0.99531645,1.1167849,1.2400664,1.3633479,1.4920682,1.6226015,1.7531348,1.8818551,2.0123885,1.6733645,1.3325275,0.9916905,0.6526665,0.31182957,0.291887,0.27194437,0.2520018,0.23205921,0.21211663,0.24293698,0.27194437,0.30276474,0.33177215,0.36259252,0.29007402,0.21755551,0.14503701,0.072518505,0.0,0.018129626,0.034446288,0.052575916,0.07070554,0.0870222,0.24293698,0.39703882,0.5529536,0.7070554,0.8629702,0.70524246,0.5475147,0.38978696,0.23205921,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.10333887,0.20486477,0.30820364,0.40972954,0.51306844,0.533011,0.5529536,0.5728962,0.59283876,0.61278135,1.0406405,1.4666867,1.8945459,2.322405,2.7502642,3.9105604,5.069043,6.2293396,7.3896356,8.549932,7.159389,5.77066,4.3801174,2.9895754,1.6008459,1.2799516,0.96087015,0.6399758,0.3208944,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.17767033,0.34264994,0.5076295,0.6726091,0.8375887,0.8665961,0.8974165,0.92823684,0.9572442,0.9880646,1.2745126,1.5627737,1.8492218,2.137483,2.4257438,2.9950142,3.5642843,4.135368,4.704638,5.275721,5.674573,6.0752378,6.474089,6.874754,7.2754188,6.069799,4.8641787,3.6603715,2.4547513,1.2491312,1.0007553,0.7505665,0.50037766,0.25018883,0.0,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.0,0.0,0.0,0.0,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.2030518,0.35534066,0.5076295,0.65991837,0.8122072,1.1494182,1.4866294,1.8256533,2.1628644,2.5000753,2.514579,2.5308957,2.5453994,2.5599031,2.5744069,2.275268,1.9743162,1.6751775,1.3742256,1.0750868,1.4956942,1.9144884,2.335096,2.7557032,3.1744974,5.1705694,7.1648283,9.1609,11.155159,13.149418,10.899531,8.649645,6.399758,4.1498713,1.8999848,1.6008459,1.2998942,1.0007553,0.69980353,0.40066472,1.2291887,2.0595255,2.8898623,3.720199,4.550536,3.6404288,2.7303216,1.8202144,0.9101072,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.12690738,0.23024625,0.33177215,0.43511102,0.53663695,0.4604925,0.3825351,0.3045777,0.22662032,0.15047589,0.9880646,1.8256533,2.663242,3.5008307,4.3366065,4.655688,4.972956,5.290225,5.6074934,5.924762,5.4026284,4.880495,4.358362,3.834416,3.3122826,3.4246864,3.53709,3.6494937,3.7618973,3.874301,3.5280252,3.1799364,2.8318477,2.4855716,2.137483,1.7132497,1.2872034,0.8629702,0.43692398,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,0.9119202,1.5754645,2.2371957,2.9007401,3.5624714,5.328297,7.0923095,8.858135,10.622148,12.387974,12.021755,11.65735,11.292944,10.926725,10.56232,8.7421055,6.921891,5.101677,3.2832751,1.4630609,1.3397794,1.2183108,1.0950294,0.97174793,0.85027945,0.75963134,0.67079616,0.58014804,0.4894999,0.40066472,0.3208944,0.23931105,0.15954071,0.07977036,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.49675176,0.969935,1.4431182,1.9144884,2.3876717,1.9815681,1.5772774,1.1729867,0.7668832,0.36259252,0.5094425,0.65810543,0.80495536,0.95180535,1.1004683,1.7621996,2.4257438,3.0874753,3.7492065,4.4127507,4.8079767,5.2032027,5.5966153,5.9918413,6.3870673,6.590119,6.793171,6.9944096,7.1974616,7.400513,8.46291,9.525306,10.587702,11.650098,12.712494,11.856775,11.00287,10.147152,9.293246,8.437528,8.629702,8.821876,9.015862,9.208037,9.400211,8.345067,7.2899227,6.2347784,5.179634,4.12449,3.8833659,3.6404288,3.397492,3.1545548,2.911618,3.9522583,4.992899,6.0317264,7.072367,8.113008,9.402024,10.692853,11.98187,13.272699,14.561715,14.157425,13.753134,13.347031,12.9427395,12.536636,11.035503,9.5325575,8.029612,6.528478,5.0255322,4.2894692,3.5552197,2.819157,2.084907,1.3506571,2.7847104,4.220577,5.65463,7.0904965,8.52455,9.128266,9.73017,10.332074,10.93579,11.537694,11.709926,11.882156,12.054388,12.22662,12.400664,11.985496,11.570327,11.155159,10.73999,10.324821,11.399909,12.474996,13.550082,14.625169,15.700256,15.245202,14.790149,14.335095,13.880041,13.424988,12.197612,10.970237,9.742861,8.515485,7.28811,7.6380115,7.987913,8.337815,8.6877165,9.037619,7.915395,6.793171,5.669134,4.5469103,3.4246864,4.349297,5.275721,6.200332,7.124943,8.049554,6.8076744,5.563982,4.322103,3.0802233,1.8383441,2.3949237,2.953316,3.5098956,4.068288,4.6248674,4.699199,4.7753434,4.8496747,4.9258194,5.0001507,4.3819304,3.7655232,3.147303,2.5308957,1.9126755,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.07433146,0.07433146,0.07433146,0.07433146,0.07433146,0.065266654,0.054388877,0.045324065,0.034446288,0.025381476,0.034446288,0.045324065,0.054388877,0.065266654,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06707962,0.13415924,0.2030518,0.27013144,0.33721104,0.6000906,0.8629702,1.1258497,1.3869164,1.649796,1.6679256,1.6842422,1.7023718,1.7205015,1.7368182,1.7549478,1.7730774,1.789394,1.8075237,1.8256533,1.6352923,1.4449311,1.2545701,1.064209,0.87566096,0.9826257,1.0895905,1.1983683,1.305333,1.4122978,1.4594349,1.5083848,1.5555218,1.6026589,1.649796,1.4068589,1.1657349,0.922798,0.67986095,0.43692398,0.38434806,0.33177215,0.27919623,0.22662032,0.17585737,0.19761293,0.21936847,0.24293698,0.26469254,0.28826106,0.23024625,0.17223145,0.11421664,0.058014803,0.0,0.034446288,0.07070554,0.10515183,0.13959812,0.17585737,0.48587397,0.79589057,1.1059072,1.4141108,1.7241274,1.4104849,1.0950294,0.7795739,0.46411842,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13053331,0.25925365,0.38978696,0.52032024,0.6508536,0.7650702,0.8792868,0.99531645,1.1095331,1.2255627,1.3923552,1.5591478,1.7277533,1.8945459,2.0631514,2.9333735,3.8017826,4.6720047,5.542227,6.412449,5.369995,4.327542,3.2850883,2.2426348,1.2001812,0.96087015,0.7197462,0.48043507,0.23931105,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.16679256,0.3100166,0.45324063,0.5946517,0.73787576,0.7469406,0.75781834,0.7668832,0.7777609,0.7868258,1.062396,1.3379664,1.6117238,1.887294,2.1628644,2.565342,2.9678197,3.3702974,3.7727752,4.175253,4.4508233,4.7245803,5.0001507,5.275721,5.5494785,4.6393714,3.729264,2.819157,1.9108626,1.0007553,0.7995165,0.6000906,0.40066472,0.19942589,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.0,0.0,0.0,0.0,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.09064813,0.06707962,0.045324065,0.02175555,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.16679256,0.29732585,0.42785916,0.55839247,0.6871128,0.9499924,1.2128719,1.4757515,1.7368182,1.9996977,2.1683033,2.335096,2.5018883,2.6704938,2.8372865,2.5127661,2.1882458,1.8619126,1.5373923,1.2128719,1.502946,1.79302,2.0830941,2.373168,2.663242,4.102734,5.542227,6.981719,8.423024,9.862516,8.174648,6.48678,4.800725,3.1128569,1.4249886,1.2001812,0.97537386,0.7505665,0.52575916,0.2991388,0.922798,1.5446441,2.1683033,2.7901495,3.4119956,2.7303216,2.0468347,1.3651608,0.68167394,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.13053331,0.21030366,0.29007402,0.36984438,0.44961473,0.42060733,0.38978696,0.36077955,0.32995918,0.2991388,1.0243238,1.7495089,2.474694,3.199879,3.925064,4.0846047,4.2441454,4.405499,4.5650396,4.7245803,4.2804046,3.834416,3.39024,2.9442513,2.5000753,2.5870976,2.6741197,2.762955,2.8499773,2.9369993,2.70494,2.472881,2.2408218,2.0069497,1.7748904,1.4249886,1.0750868,0.72518504,0.37528324,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.87566096,1.5627737,2.2498865,2.9369993,3.6241121,5.730775,7.835624,9.940474,12.045323,14.150173,13.820213,13.490254,13.1602955,12.830337,12.500377,10.284937,8.069496,5.8540564,3.6404288,1.4249886,1.4431182,1.4594349,1.4775645,1.4956942,1.5120108,1.3325275,1.1530442,0.97174793,0.79226464,0.61278135,0.4894999,0.3680314,0.24474995,0.12328146,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.40791658,0.7650702,1.1222239,1.4793775,1.8383441,1.6026589,1.3669738,1.1331016,0.8974165,0.66173136,0.79589057,0.92823684,1.0605831,1.1929294,1.3252757,1.9996977,2.6741197,3.350355,4.024777,4.699199,4.9657044,5.230397,5.4950895,5.7597823,6.0244746,6.4432693,6.8602505,7.2772317,7.6942134,8.113008,8.825501,9.537996,10.25049,10.962985,11.675479,11.214987,10.754494,10.2958145,9.835322,9.374829,9.498111,9.619579,9.742861,9.864329,9.987611,9.003172,8.01692,7.0324817,6.0480433,5.0617914,4.84061,4.6176157,4.3946214,4.171627,3.9504454,4.7300196,5.5095935,6.2891674,7.0705543,7.850128,9.030367,10.210606,11.390844,12.569269,13.749508,13.41411,13.080525,12.745127,12.409729,12.07433,10.694666,9.3150015,7.935337,6.5556726,5.1741953,4.505212,3.834416,3.1654327,2.4946365,1.8256533,3.0330863,4.2405195,5.4479527,6.6553855,7.8628187,8.767487,9.672155,10.576823,11.483305,12.387974,12.594651,12.803142,13.009819,13.21831,13.424988,13.194741,12.964496,12.734249,12.5058155,12.27557,13.024323,13.77489,14.525456,15.27421,16.024776,15.515334,15.004078,14.494636,13.985193,13.475751,12.232059,10.990179,9.7483,8.504607,7.262728,7.5618668,7.8628187,8.161958,8.46291,8.762048,7.6924005,6.622752,5.5531044,4.4834566,3.4119956,4.2876563,5.163317,6.037165,6.9128265,7.7866745,6.5647373,5.3428006,4.120864,2.8971143,1.6751775,2.1519866,2.6306088,3.1074178,3.584227,4.062849,4.274966,4.4870825,4.699199,4.9131284,5.125245,4.615803,4.1045475,3.5951047,3.0856624,2.5744069,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.047137026,0.045324065,0.04169814,0.03988518,0.038072214,0.052575916,0.06707962,0.08339628,0.09789998,0.11240368,0.09064813,0.06707962,0.045324065,0.02175555,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.045324065,0.09064813,0.13415924,0.1794833,0.22480737,0.40066472,0.5747091,0.7505665,0.9246109,1.1004683,1.1331016,1.1657349,1.1983683,1.2291887,1.261822,1.4195497,1.5772774,1.7350051,1.892733,2.0504606,1.840157,1.6298534,1.4195497,1.209246,1.0007553,1.0932164,1.1856775,1.2781386,1.3705997,1.4630609,1.4268016,1.3923552,1.357909,1.3216497,1.2872034,1.1421664,0.99712944,0.8520924,0.7070554,0.5620184,0.47680917,0.39159992,0.30820364,0.2229944,0.13778515,0.15228885,0.16679256,0.18310922,0.19761293,0.21211663,0.17041849,0.12690738,0.08520924,0.04169814,0.0,0.052575916,0.10515183,0.15772775,0.21030366,0.26287958,0.726998,1.1929294,1.6570477,2.1229792,2.5870976,2.1157274,1.6425442,1.1693609,0.6979906,0.22480737,0.1794833,0.13415924,0.09064813,0.045324065,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.15772775,0.3154555,0.47318324,0.629098,0.7868258,0.99712944,1.2074331,1.4177368,1.6280404,1.8383441,1.745883,1.651609,1.5591478,1.4666867,1.3742256,1.9543737,2.5345216,3.1146698,3.6948178,4.274966,3.5806012,2.8844235,2.1900587,1.4956942,0.7995165,0.6399758,0.48043507,0.3208944,0.15954071,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.15772775,0.27738327,0.39703882,0.5166943,0.63816285,0.62728506,0.61822027,0.6073425,0.5982776,0.5873999,0.85027945,1.1131591,1.3742256,1.6371052,1.8999848,2.13567,2.3695421,2.6052272,2.8409123,3.0747845,3.2252605,3.3757362,3.5243993,3.6748753,3.825351,3.2107568,2.5943494,1.9797552,1.3651608,0.7505665,0.6000906,0.44961473,0.2991388,0.15047589,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.13234627,0.23931105,0.3480888,0.4550536,0.5620184,0.7505665,0.93730164,1.1258497,1.3125849,1.49932,1.8202144,2.1392958,2.4601903,2.7792716,3.100166,2.7502642,2.4003625,2.0504606,1.7005589,1.3506571,1.5101979,1.6697385,1.8292793,1.9906329,2.1501737,3.0348995,3.919625,4.804351,5.6908894,6.5756154,5.4497657,4.325729,3.199879,2.0758421,0.9499924,0.7995165,0.6508536,0.50037766,0.34990177,0.19942589,0.61459434,1.0297627,1.4449311,1.8600996,2.275268,1.8202144,1.3651608,0.9101072,0.4550536,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.13234627,0.19036107,0.24837588,0.3045777,0.36259252,0.38072214,0.39703882,0.41516843,0.43329805,0.44961473,1.062396,1.6751775,2.2879589,2.9007401,3.5117085,3.5153344,3.5171473,3.5207734,3.5225863,3.5243993,3.1581807,2.7901495,2.422118,2.0558996,1.6878681,1.7495089,1.8129625,1.8746033,1.938057,1.9996977,1.8818551,1.7658255,1.647983,1.5301404,1.4122978,1.1367276,0.8629702,0.5873999,0.31182957,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.8375887,1.550083,2.2625773,2.9750717,3.6875658,6.1332526,8.577126,11.022813,13.466686,15.912373,15.616859,15.32316,15.027647,14.732134,14.436621,11.827768,9.217102,6.6082487,3.9975824,1.3869164,1.5446441,1.7023718,1.8600996,2.0178273,2.175555,1.9054236,1.6352923,1.3651608,1.0950294,0.824898,0.65991837,0.4949388,0.32995918,0.16497959,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.31726846,0.56020546,0.8031424,1.0442665,1.2872034,1.2219368,1.1566701,1.0932164,1.0279498,0.96268314,1.0805258,1.1983683,1.3143979,1.4322405,1.550083,2.2371957,2.9243085,3.6132345,4.3003473,4.98746,5.121619,5.2575917,5.391751,5.527723,5.661882,6.294606,6.92733,7.560054,8.192778,8.825501,9.188094,9.550687,9.91328,10.275872,10.636651,10.573197,10.507931,10.442664,10.377398,10.312131,10.364707,10.417283,10.469859,10.522435,10.57501,9.659465,8.745731,7.8301854,6.9146395,5.999093,5.7978544,5.5948024,5.391751,5.1905117,4.98746,5.5077806,6.0281005,6.546608,7.066928,7.5872483,8.656897,9.728357,10.798005,11.867653,12.937301,12.672608,12.407916,12.143224,11.876718,11.612025,10.355642,9.097446,7.83925,6.582867,5.3246713,4.7191415,4.115425,3.5098956,2.904366,2.3006494,3.2796493,4.2604623,5.239462,6.2202744,7.1992745,8.406708,9.6141405,10.823386,12.03082,13.238253,13.479377,13.722314,13.965251,14.208188,14.449312,14.405801,14.3604765,14.315152,14.269829,14.224504,14.650551,15.074784,15.50083,15.925063,16.349297,15.785465,15.219821,14.654177,14.090345,13.524701,12.268318,11.010121,9.751925,8.495543,7.2373466,7.4875355,7.7377243,7.987913,8.238102,8.488291,7.4694057,6.452334,5.4352617,4.41819,3.3993049,4.2242026,5.050914,5.8758116,6.70071,7.5256076,6.3218007,5.1198063,3.917812,2.715818,1.5120108,1.9108626,2.3079014,2.70494,3.101979,3.5008307,3.8507326,4.2006345,4.550536,4.900438,5.2503395,4.847862,4.445384,4.0429068,3.6404288,3.2379513,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.030820364,0.034446288,0.03988518,0.045324065,0.05076295,0.07070554,0.09064813,0.11059072,0.13053331,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.19942589,0.28826106,0.37528324,0.46230546,0.5493277,0.5982776,0.64541465,0.69255173,0.73968875,0.7868258,1.0841516,1.3832904,1.6806163,1.9779422,2.275268,2.0450218,1.8147756,1.5845293,1.3542831,1.1258497,1.2019942,1.2799516,1.357909,1.4358664,1.5120108,1.3941683,1.2781386,1.1602961,1.0424535,0.9246109,0.8774739,0.83033687,0.78319985,0.73424983,0.6871128,0.56927025,0.45324063,0.33539808,0.21755551,0.099712946,0.10696479,0.11421664,0.12328146,0.13053331,0.13778515,0.11059072,0.08339628,0.054388877,0.027194439,0.0,0.07070554,0.13959812,0.21030366,0.27919623,0.34990177,0.969935,1.5899682,2.2100015,2.8300345,3.4500678,2.819157,2.1900587,1.5591478,0.9300498,0.2991388,0.23931105,0.1794833,0.11965553,0.059827764,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.18492219,0.36984438,0.55476654,0.73968875,0.9246109,1.2291887,1.5355793,1.840157,2.1447346,2.4493124,2.0975976,1.745883,1.3923552,1.0406405,0.6871128,0.97718686,1.2672608,1.5573349,1.8474089,2.137483,1.789394,1.4431182,1.0950294,0.7469406,0.40066472,0.3208944,0.23931105,0.15954071,0.07977036,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.14684997,0.24474995,0.34264994,0.4405499,0.53663695,0.5076295,0.47680917,0.44780177,0.4169814,0.387974,0.63816285,0.8883517,1.1367276,1.3869164,1.6371052,1.7041848,1.7730774,1.840157,1.9072367,1.9743162,1.9996977,2.0250793,2.0504606,2.0758421,2.0994108,1.7803292,1.4594349,1.1403534,0.8194591,0.50037766,0.40066472,0.2991388,0.19942589,0.099712946,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.09789998,0.18310922,0.26831847,0.35171473,0.43692398,0.5493277,0.66173136,0.774135,0.8883517,1.0007553,1.4721256,1.9453088,2.4166791,2.8898623,3.3630457,2.9877625,2.612479,2.2371957,1.8619126,1.4866294,1.5174497,1.54827,1.5772774,1.6080978,1.6371052,1.9670644,2.2970235,2.6269827,2.956942,3.2869012,2.7248828,2.1628644,1.6008459,1.0370146,0.4749962,0.40066472,0.3245203,0.25018883,0.17585737,0.099712946,0.30820364,0.5148814,0.72337204,0.9300498,1.1367276,0.9101072,0.68167394,0.4550536,0.22662032,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.13415924,0.17041849,0.20486477,0.23931105,0.2755703,0.34083697,0.40429065,0.46955732,0.53482395,0.6000906,1.1004683,1.6008459,2.0994108,2.5997884,3.100166,2.9442513,2.7901495,2.6342347,2.4801328,2.324218,2.034144,1.745883,1.455809,1.1657349,0.87566096,0.9119202,0.9499924,0.9880646,1.0243238,1.062396,1.0605831,1.0569572,1.0551442,1.0533313,1.0497054,0.85027945,0.6508536,0.44961473,0.25018883,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.7995165,1.5373923,2.275268,3.0131438,3.7492065,6.53573,9.32044,12.105151,14.889862,17.674572,17.41532,17.154251,16.894999,16.635744,16.374678,13.370599,10.364707,7.360628,4.3547363,1.3506571,1.647983,1.9453088,2.2426348,2.5399606,2.8372865,2.47832,2.1175404,1.7567607,1.3977941,1.0370146,0.83033687,0.62184614,0.41516843,0.20667773,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.22662032,0.35534066,0.48224804,0.6091554,0.73787576,0.8430276,0.9481794,1.0533313,1.1566701,1.261822,1.3651608,1.4666867,1.5700256,1.6733645,1.7748904,2.474694,3.1744974,3.874301,4.5759177,5.275721,5.279347,5.2847857,5.290225,5.295664,5.2992897,6.147756,6.9944096,7.842876,8.689529,9.537996,9.550687,9.563377,9.574255,9.5869465,9.599637,9.929596,10.259555,10.589515,10.919474,11.249433,11.233116,11.214987,11.1968565,11.18054,11.162411,10.31757,9.47273,8.627889,7.783048,6.9382076,6.755099,6.5719895,6.390693,6.207584,6.0244746,6.285541,6.544795,6.8058615,7.065115,7.324369,8.285239,9.244296,10.205167,11.164224,12.125093,11.929294,11.735307,11.539507,11.34552,11.14972,10.014805,8.87989,7.744976,6.6100616,5.475147,4.934884,4.3946214,3.8543584,3.3159087,2.7756457,3.5280252,4.2804046,5.032784,5.7851634,6.5375433,8.047741,9.557939,11.068136,12.576522,14.0867195,14.365915,14.643299,14.920682,15.198066,15.475449,15.6150465,15.754644,15.894243,16.035654,16.175253,16.274965,16.374678,16.474392,16.574104,16.67563,16.055597,15.435563,14.81553,14.195497,13.575464,12.302764,11.030065,9.757364,8.484665,7.211965,7.413204,7.61263,7.8120556,8.013294,8.212721,7.2482243,6.281915,5.317419,4.3529234,3.386614,4.162562,4.936697,5.712645,6.48678,7.262728,6.0806766,4.896812,3.7147603,2.5327086,1.3506571,1.6679256,1.9851941,2.3024626,2.619731,2.9369993,3.4246864,3.9123733,4.40006,4.8877473,5.375434,5.0799212,4.784408,4.4907084,4.195195,3.8996825,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.0870222,0.11240368,0.13778515,0.16316663,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06164073,0.12509441,0.18673515,0.25018883,0.31182957,0.7505665,1.1874905,1.6244144,2.0631514,2.5000753,2.2498865,1.9996977,1.7495089,1.49932,1.2491312,1.3125849,1.3742256,1.4376793,1.49932,1.5627737,1.3633479,1.162109,0.96268314,0.76325727,0.5620184,0.61278135,0.66173136,0.7124943,0.76325727,0.8122072,0.66173136,0.51306844,0.36259252,0.21211663,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0870222,0.17585737,0.26287958,0.34990177,0.43692398,1.2128719,1.987007,2.762955,3.53709,4.313038,3.5243993,2.7375734,1.9507477,1.162109,0.37528324,0.2991388,0.22480737,0.15047589,0.07433146,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.21211663,0.42423326,0.63816285,0.85027945,1.062396,1.4630609,1.8619126,2.2625773,2.663242,3.0620937,2.4493124,1.8383441,1.2255627,0.61278135,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.13778515,0.21211663,0.28826106,0.36259252,0.43692398,0.387974,0.33721104,0.28826106,0.2374981,0.18673515,0.42423326,0.66173136,0.89922947,1.1367276,1.3742256,1.2745126,1.1747998,1.0750868,0.97537386,0.87566096,0.774135,0.6744221,0.5747091,0.4749962,0.37528324,0.34990177,0.3245203,0.2991388,0.2755703,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06164073,0.12509441,0.18673515,0.25018883,0.31182957,0.34990177,0.387974,0.42423326,0.46230546,0.50037766,1.1258497,1.7495089,2.374981,3.000453,3.6241121,3.2252605,2.8245957,2.4257438,2.0250793,1.6244144,1.5247015,1.4249886,1.3252757,1.2255627,1.1258497,0.89922947,0.6744221,0.44961473,0.22480737,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.13778515,0.15047589,0.16316663,0.17585737,0.18673515,0.2991388,0.41335547,0.52575916,0.63816285,0.7505665,1.1367276,1.5247015,1.9126755,2.3006494,2.6868105,2.374981,2.0631514,1.7495089,1.4376793,1.1258497,0.9119202,0.69980353,0.48768693,0.2755703,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.2374981,0.34990177,0.46230546,0.5747091,0.6871128,0.5620184,0.43692398,0.31182957,0.18673515,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.76325727,1.5247015,2.2879589,3.049403,3.8126602,6.9382076,10.061942,13.1874895,16.313038,19.436771,19.211964,18.987158,18.76235,18.537542,18.312735,14.911617,11.512312,8.113008,4.7118897,1.3125849,1.7495089,2.1882458,2.6251698,3.0620937,3.5008307,3.049403,2.5997884,2.1501737,1.7005589,1.2491312,1.0007553,0.7505665,0.50037766,0.25018883,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.13778515,0.15047589,0.16316663,0.17585737,0.18673515,0.46230546,0.73787576,1.0116332,1.2872034,1.5627737,1.649796,1.7368182,1.8256533,1.9126755,1.9996977,2.712192,3.4246864,4.137181,4.8496747,5.562169,5.4370747,5.3119802,5.186886,5.0617914,4.936697,6.000906,7.063302,8.125698,9.188094,10.25049,9.91328,9.574255,9.237044,8.899834,8.562622,9.287807,10.012992,10.738177,11.463363,12.186734,12.099712,12.012691,11.925668,11.836833,11.74981,10.975676,10.199727,9.425592,8.649645,7.8755093,7.7123427,7.549176,7.3878226,7.224656,7.063302,7.063302,7.063302,7.063302,7.063302,7.063302,7.911769,8.762048,9.612328,10.462607,11.312886,11.187792,11.062697,10.937603,10.812509,10.687414,9.675781,8.662335,7.650702,6.637256,5.6256227,5.1506267,4.6756306,4.2006345,3.7256382,3.2506418,3.774588,4.3003473,4.8242936,5.3500524,5.8758116,7.686961,9.499924,11.312886,13.124036,14.936998,15.250641,15.56247,15.8743,16.187943,16.499773,16.824293,17.150625,17.475147,17.799667,18.124187,17.89938,17.674572,17.449764,17.224958,17.00015,16.325727,15.649493,14.975071,14.300649,13.6244135,12.337211,11.050007,9.762803,8.4756,7.1883965,7.3370595,7.4875355,7.6380115,7.7866745,7.93715,7.02523,6.111497,5.199577,4.2876563,3.3757362,4.100921,4.8242936,5.5494785,6.2746634,6.9998484,5.8377395,4.6756306,3.5117085,2.3495996,1.1874905,1.4249886,1.6624867,1.8999848,2.137483,2.374981,3.000453,3.625925,4.249584,4.8750563,5.5005283,5.3119802,5.125245,4.936697,4.749962,4.5632267,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.11784257,0.15954071,0.2030518,0.24474995,0.28826106,0.2374981,0.18673515,0.13778515,0.0870222,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,0.6000906,0.9499924,1.2998942,1.649796,1.9996977,1.8147756,1.6298534,1.4449311,1.260009,1.0750868,1.1530442,1.2291887,1.3071461,1.3851035,1.4630609,1.3125849,1.162109,1.0116332,0.8629702,0.7124943,0.7124943,0.7124943,0.7124943,0.7124943,0.7124943,0.58014804,0.44780177,0.3154555,0.18310922,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.07977036,0.15954071,0.23931105,0.3208944,0.40066472,1.1004683,1.8002719,2.5000753,3.199879,3.8996825,3.198066,2.4946365,1.79302,1.0895905,0.387974,0.31182957,0.2374981,0.16316663,0.0870222,0.012690738,0.014503701,0.018129626,0.01994259,0.02175555,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.17041849,0.34083697,0.5094425,0.67986095,0.85027945,1.1693609,1.4902552,1.8093367,2.1302311,2.4493124,1.9598125,1.4703126,0.9808127,0.4894999,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.052575916,0.10515183,0.15772775,0.21030366,0.26287958,0.27919623,0.29732585,0.3154555,0.33177215,0.34990177,0.54570174,0.73968875,0.9354887,1.1294757,1.3252757,1.3125849,1.2998942,1.2872034,1.2745126,1.261822,1.1530442,1.0424535,0.9318628,0.823085,0.7124943,0.63816285,0.5620184,0.48768693,0.41335547,0.33721104,0.31182957,0.28826106,0.26287958,0.2374981,0.21211663,0.17041849,0.12690738,0.08520924,0.04169814,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,0.27919623,0.3100166,0.34083697,0.36984438,0.40066472,0.89922947,1.3996071,1.8999848,2.4003625,2.9007401,2.5798457,2.2607644,1.93987,1.6207886,1.2998942,1.2201238,1.1403534,1.0605831,0.9808127,0.89922947,0.7197462,0.5402629,0.36077955,0.1794833,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.13234627,0.16497959,0.19761293,0.23024625,0.26287958,0.34083697,0.4169814,0.4949388,0.5728962,0.6508536,0.95180535,1.2545701,1.5573349,1.8600996,2.1628644,1.9108626,1.6570477,1.405046,1.1530442,0.89922947,0.7306239,0.56020546,0.38978696,0.21936847,0.05076295,0.059827764,0.07070554,0.07977036,0.09064813,0.099712946,0.19036107,0.27919623,0.36984438,0.4604925,0.5493277,0.5076295,0.46411842,0.4224203,0.38072214,0.33721104,0.27013144,0.2030518,0.13415924,0.06707962,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.6091554,1.2201238,1.8292793,2.4402475,3.049403,5.844991,8.640579,11.434355,14.229943,17.025532,17.94289,18.86025,19.777609,20.694967,21.612328,17.660069,13.70781,9.755551,5.803293,1.8492218,2.2970235,2.7448254,3.1926272,3.6404288,4.0882306,3.7909048,3.491766,3.1944401,2.8971143,2.5997884,2.0830941,1.5645868,1.0478923,0.5293851,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.32814622,0.6544795,0.9826257,1.310772,1.6371052,1.6733645,1.7078108,1.742257,1.7767034,1.8129625,1.7404441,1.6679256,1.5954071,1.5228885,1.4503701,1.5809034,1.7096237,1.840157,1.9706904,2.0994108,2.7357605,3.3702974,4.004834,4.6393714,5.275721,5.2648435,5.2557783,5.2449007,5.235836,5.224958,6.008158,6.789545,7.572745,8.354132,9.137331,8.943344,8.747544,8.551744,8.357758,8.161958,9.055748,9.947725,10.839704,11.731681,12.625471,12.456866,12.290073,12.123281,11.954676,11.787883,11.10077,10.411844,9.724731,9.037619,8.350506,8.3777,8.404895,8.432089,8.459284,8.488291,8.3051815,8.122072,7.9407763,7.757667,7.574558,8.172835,8.7693,9.367578,9.965856,10.56232,10.377398,10.192475,10.007553,9.822631,9.637709,8.680465,7.723221,6.7641635,5.806919,4.8496747,4.5342193,4.220577,3.9051213,3.589666,3.2742105,3.7655232,4.255023,4.744523,5.235836,5.7253356,7.28811,8.849071,10.411844,11.974618,13.537392,13.918114,14.297023,14.677745,15.056654,15.437376,15.620485,15.801782,15.984891,16.168001,16.349297,16.41819,16.48527,16.55235,16.619429,16.68832,16.091856,15.497204,14.902553,14.3079,13.713249,12.8321495,11.952863,11.071762,10.192475,9.313189,8.785617,8.258044,7.7304726,7.2029004,6.6753283,5.903006,5.130684,4.358362,3.584227,2.811905,3.3721104,3.9323158,4.4925213,5.0527267,5.612932,4.7390842,3.8670492,2.9950142,2.1229792,1.2491312,1.4068589,1.5645868,1.7223145,1.8800422,2.03777,2.561716,3.0874753,3.6132345,4.137181,4.6629395,4.632119,4.603112,4.572292,4.5432844,4.512464,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.018129626,0.034446288,0.052575916,0.07070554,0.0870222,0.14684997,0.20667773,0.26831847,0.32814622,0.387974,0.3245203,0.26287958,0.19942589,0.13778515,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.44961473,0.7124943,0.97537386,1.2382535,1.49932,1.3796645,1.260009,1.1403534,1.020698,0.89922947,0.9916905,1.0841516,1.1766127,1.2708868,1.3633479,1.261822,1.162109,1.062396,0.96268314,0.8629702,0.8122072,0.76325727,0.7124943,0.66173136,0.61278135,0.49675176,0.3825351,0.26831847,0.15228885,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.072518505,0.14503701,0.21755551,0.29007402,0.36259252,0.9880646,1.6117238,2.2371957,2.8626678,3.48814,2.8699198,2.2516994,1.6352923,1.017072,0.40066472,0.3245203,0.25018883,0.17585737,0.099712946,0.025381476,0.030820364,0.034446288,0.03988518,0.045324065,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.12690738,0.25562772,0.3825351,0.5094425,0.63816285,0.8774739,1.1167849,1.357909,1.5972201,1.8383441,1.4703126,1.1022812,0.73424983,0.3680314,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.092461094,0.18492219,0.27738327,0.36984438,0.46230546,0.4224203,0.3825351,0.34264994,0.30276474,0.26287958,0.7016165,1.1421664,1.5827163,2.0232663,2.4620032,2.1991236,1.938057,1.6751775,1.4122978,1.1494182,1.0297627,0.9101072,0.7904517,0.67079616,0.5493277,0.50037766,0.44961473,0.40066472,0.34990177,0.2991388,0.2755703,0.25018883,0.22480737,0.19942589,0.17585737,0.13959812,0.10515183,0.07070554,0.034446288,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.21030366,0.23205921,0.25562772,0.27738327,0.2991388,0.6744221,1.0497054,1.4249886,1.8002719,2.175555,1.9344311,1.69512,1.455809,1.214685,0.97537386,0.9155461,0.8557183,0.79589057,0.73424983,0.6744221,0.5402629,0.40429065,0.27013144,0.13415924,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.12690738,0.1794833,0.23205921,0.28463513,0.33721104,0.38072214,0.4224203,0.46411842,0.5076295,0.5493277,0.7668832,0.98443866,1.2019942,1.4195497,1.6371052,1.4449311,1.2527572,1.0605831,0.8665961,0.6744221,0.5475147,0.42060733,0.291887,0.16497959,0.038072214,0.045324065,0.052575916,0.059827764,0.06707962,0.07433146,0.14322405,0.21030366,0.27738327,0.3444629,0.41335547,0.45324063,0.49312583,0.533011,0.5728962,0.61278135,0.4894999,0.3680314,0.24474995,0.12328146,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.45686656,0.9155461,1.3724127,1.8292793,2.2879589,4.751775,7.217404,9.683033,12.14685,14.612478,16.672005,18.733343,20.792868,22.852394,24.911919,20.406708,15.903308,11.398096,6.892884,2.3876717,2.8445382,3.303218,3.7600844,4.216951,4.6756306,4.5305934,4.3855567,4.2405195,4.0954823,3.9504454,3.1654327,2.38042,1.5954071,0.8103943,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.630911,1.260009,1.8909199,2.520018,3.149116,3.207131,3.2651455,3.3231604,3.3793623,3.437377,3.0167696,2.5979755,2.1773682,1.7567607,1.3379664,1.5101979,1.6824293,1.8546607,2.0268922,2.1991236,2.7575161,3.3140955,3.872488,4.4308805,4.98746,5.092612,5.197764,5.3029156,5.408067,5.5132194,6.01541,6.5176005,7.019791,7.5219817,8.024173,7.9715962,7.9208336,7.8682575,7.8156815,7.763106,8.821876,9.882459,10.943042,12.001812,13.062395,12.815832,12.567456,12.320893,12.072517,11.8241415,11.225864,10.625773,10.025683,9.425592,8.825501,9.043057,9.2606125,9.4781685,9.695724,9.91328,9.547061,9.182655,8.81825,8.452031,8.087626,8.432089,8.778365,9.122828,9.467291,9.811753,9.567003,9.322253,9.077503,8.832754,8.588004,7.6851482,6.782293,5.8794374,4.9783955,4.07554,3.919625,3.7655232,3.6096084,3.4555066,3.299592,3.7546456,4.209699,4.664753,5.1198063,5.57486,6.887445,8.200029,9.512614,10.825199,12.137785,12.585587,13.033388,13.479377,13.927178,14.37498,14.4148655,14.454751,14.494636,14.534521,14.574407,14.935185,15.294152,15.654932,16.01571,16.374678,15.859797,15.344915,14.830034,14.315152,13.800271,13.327088,12.855718,12.382534,11.909351,11.437981,10.232361,9.026741,7.8229337,6.6173134,5.411693,4.780782,4.1480584,3.5153344,2.8826106,2.2498865,2.6451125,3.0403383,3.435564,3.83079,4.2242026,3.6422417,3.0602808,2.47832,1.8945459,1.3125849,1.3905423,1.4666867,1.5446441,1.6226015,1.7005589,2.124792,2.5508385,2.9750717,3.3993049,3.825351,3.9522583,4.079166,4.207886,4.3347936,4.461701,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.17767033,0.25562772,0.33177215,0.40972954,0.48768693,0.41335547,0.33721104,0.26287958,0.18673515,0.11240368,0.09064813,0.06707962,0.045324065,0.02175555,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.2991388,0.4749962,0.6508536,0.824898,1.0007553,0.9445535,0.8901646,0.83577573,0.7795739,0.72518504,0.8321498,0.93911463,1.0478923,1.1548572,1.261822,1.2128719,1.162109,1.1131591,1.062396,1.0116332,0.9119202,0.8122072,0.7124943,0.61278135,0.51306844,0.41516843,0.31726846,0.21936847,0.12328146,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.065266654,0.13053331,0.19579996,0.25925365,0.3245203,0.87566096,1.4249886,1.9743162,2.525457,3.0747845,2.5417736,2.0105755,1.4775645,0.9445535,0.41335547,0.33721104,0.26287958,0.18673515,0.11240368,0.038072214,0.045324065,0.052575916,0.059827764,0.06707962,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.08520924,0.17041849,0.25562772,0.34083697,0.42423326,0.5855869,0.7451276,0.90466833,1.064209,1.2255627,0.9808127,0.73424983,0.4894999,0.24474995,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13234627,0.26469254,0.39703882,0.5293851,0.66173136,0.5656443,0.46774435,0.36984438,0.27194437,0.17585737,0.85934424,1.5446441,2.229944,2.9152439,3.6005437,3.0874753,2.5744069,2.0631514,1.550083,1.0370146,0.90829426,0.7777609,0.64722764,0.5166943,0.387974,0.36259252,0.33721104,0.31182957,0.28826106,0.26287958,0.2374981,0.21211663,0.18673515,0.16316663,0.13778515,0.11059072,0.08339628,0.054388877,0.027194439,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.13959812,0.15410182,0.17041849,0.18492219,0.19942589,0.44961473,0.69980353,0.9499924,1.2001812,1.4503701,1.2908293,1.1294757,0.969935,0.8103943,0.6508536,0.6091554,0.56927025,0.5293851,0.4894999,0.44961473,0.36077955,0.27013144,0.1794833,0.09064813,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.12328146,0.19579996,0.26831847,0.34083697,0.41335547,0.42060733,0.42785916,0.43511102,0.44236287,0.44961473,0.581961,0.71430725,0.8466535,0.9808127,1.1131591,0.9808127,0.8466535,0.71430725,0.581961,0.44961473,0.36440548,0.27919623,0.19579996,0.11059072,0.025381476,0.030820364,0.034446288,0.03988518,0.045324065,0.05076295,0.09427405,0.13959812,0.18492219,0.23024625,0.2755703,0.39703882,0.52032024,0.6417888,0.7650702,0.8883517,0.7106813,0.533011,0.35534066,0.17767033,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.3045777,0.6091554,0.9155461,1.2201238,1.5247015,3.6603715,5.7942286,7.9298983,10.065568,12.199425,15.40293,18.604622,21.808126,25.009819,28.213324,23.155159,18.096992,13.04064,7.9824743,2.9243085,3.392053,3.8597972,4.327542,4.795286,5.2630305,5.2702823,5.277534,5.2847857,5.292038,5.2992897,4.2477713,3.1944401,2.1429217,1.0895905,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.9318628,1.8655385,2.7974012,3.729264,4.6629395,4.74271,4.8224807,4.902251,4.9820213,5.0617914,4.2949085,3.5280252,2.759329,1.9924458,1.2255627,1.4394923,1.6552348,1.8691645,2.084907,2.3006494,2.7792716,3.2597067,3.7401419,4.220577,4.699199,4.9203806,5.139749,5.3591175,5.580299,5.7996674,6.0226617,6.245656,6.4668374,6.6898317,6.9128265,7.0016613,7.0923095,7.1829576,7.271793,7.362441,8.589817,9.817192,11.044568,12.271944,13.499319,13.172986,12.84484,12.516694,12.19036,11.862214,11.349146,10.837891,10.324821,9.811753,9.300498,9.708415,10.114518,10.522435,10.930351,11.338268,10.790753,10.243238,9.695724,9.14821,8.600695,8.693155,8.785617,8.8780775,8.970539,9.063,8.756609,8.452031,8.147454,7.842876,7.5382986,6.6898317,5.8431783,4.994712,4.1480584,3.299592,3.3050308,3.3104696,3.3159087,3.3195345,3.3249733,3.7455807,4.164375,4.5849824,5.0055895,5.424384,6.48678,7.549176,8.613385,9.675781,10.738177,11.253058,11.7679405,12.282822,12.797703,13.312584,13.209246,13.107719,13.00438,12.902855,12.799516,13.452183,14.104849,14.757515,15.410182,16.062849,15.627737,15.192626,14.757515,14.322405,13.887294,13.822026,13.75676,13.693306,13.628039,13.562773,11.679105,9.79725,7.915395,6.0317264,4.1498713,3.6567454,3.1654327,2.6723068,2.179181,1.6878681,1.9181144,2.1483607,2.3767939,2.6070402,2.8372865,2.5453994,2.2516994,1.9598125,1.6679256,1.3742256,1.3724127,1.3705997,1.3669738,1.3651608,1.3633479,1.6878681,2.0123885,2.3369088,2.663242,2.9877625,3.2723975,3.5570326,3.8416677,4.1281157,4.4127507,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.20667773,0.30276474,0.39703882,0.49312583,0.5873999,0.50037766,0.41335547,0.3245203,0.2374981,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.15047589,0.2374981,0.3245203,0.41335547,0.50037766,0.5094425,0.52032024,0.5293851,0.5402629,0.5493277,0.6726091,0.79589057,0.91735905,1.0406405,1.162109,1.162109,1.162109,1.162109,1.162109,1.162109,1.0116332,0.8629702,0.7124943,0.5620184,0.41335547,0.33177215,0.2520018,0.17223145,0.092461094,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.058014803,0.11421664,0.17223145,0.23024625,0.28826106,0.76325727,1.2382535,1.7132497,2.1882458,2.663242,2.2154403,1.7676386,1.3198367,0.872035,0.42423326,0.34990177,0.2755703,0.19942589,0.12509441,0.05076295,0.059827764,0.07070554,0.07977036,0.09064813,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.04169814,0.08520924,0.12690738,0.17041849,0.21211663,0.291887,0.37165734,0.45324063,0.533011,0.61278135,0.4894999,0.3680314,0.24474995,0.12328146,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.17223145,0.3444629,0.5166943,0.69073874,0.8629702,0.7070554,0.5529536,0.39703882,0.24293698,0.0870222,1.017072,1.9471219,2.8771715,3.8072214,4.7372713,3.975827,3.2125697,2.4493124,1.6878681,0.9246109,0.7850128,0.64541465,0.5058166,0.36440548,0.22480737,0.22480737,0.22480737,0.22480737,0.22480737,0.22480737,0.19942589,0.17585737,0.15047589,0.12509441,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.07070554,0.07795739,0.08520924,0.092461094,0.099712946,0.22480737,0.34990177,0.4749962,0.6000906,0.72518504,0.64541465,0.5656443,0.48587397,0.40429065,0.3245203,0.3045777,0.28463513,0.26469254,0.24474995,0.22480737,0.1794833,0.13415924,0.09064813,0.045324065,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.11784257,0.21030366,0.30276474,0.39522585,0.48768693,0.4604925,0.43329805,0.40429065,0.3770962,0.34990177,0.39703882,0.44417584,0.49312583,0.5402629,0.5873999,0.5148814,0.44236287,0.36984438,0.29732585,0.22480737,0.18310922,0.13959812,0.09789998,0.054388877,0.012690738,0.014503701,0.018129626,0.01994259,0.02175555,0.025381476,0.047137026,0.07070554,0.092461094,0.11421664,0.13778515,0.34264994,0.5475147,0.7523795,0.9572442,1.162109,0.9300498,0.6979906,0.46411842,0.23205921,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.15228885,0.3045777,0.45686656,0.6091554,0.76325727,2.5671551,4.3728657,6.1767635,7.9824743,9.788185,14.132043,18.477715,22.823385,27.167244,31.512915,25.901796,20.29249,14.683184,9.072064,3.4627585,3.9395678,4.41819,4.894999,5.371808,5.8504305,6.009971,6.169512,6.3308654,6.490406,6.6499467,5.33011,4.0102735,2.6904364,1.3705997,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.2346275,2.469255,3.7056956,4.940323,6.1749506,6.2782893,6.379815,6.4831543,6.58468,6.688019,5.573047,4.458075,3.343103,2.228131,1.1131591,1.3705997,1.6280404,1.8854811,2.1429217,2.4003625,2.8028402,3.2053177,3.6077955,4.0102735,4.4127507,4.748149,5.081734,5.4171324,5.75253,6.0879283,6.0299134,5.9718986,5.915697,5.857682,5.7996674,6.0317264,6.265599,6.497658,6.7297173,6.9617763,8.357758,9.751925,11.147907,12.542075,13.938056,13.53014,13.122223,12.714307,12.308203,11.900287,11.47424,11.050007,10.625773,10.199727,9.775495,10.371959,10.970237,11.566701,12.164979,12.763257,12.032633,11.302009,10.573197,9.842574,9.11195,8.952409,8.792869,8.6333275,8.471974,8.312433,7.948028,7.5818095,7.217404,6.8529987,6.48678,5.6945157,4.902251,4.1099863,3.3177216,2.525457,2.6904364,2.855416,3.0203958,3.1853752,3.350355,3.7347028,4.120864,4.505212,4.88956,5.275721,6.0879283,6.9001355,7.7123427,8.52455,9.336758,9.920531,10.502492,11.084454,11.668227,12.250188,12.005438,11.760688,11.514126,11.269376,11.024626,11.969179,12.915545,13.860099,14.804652,15.749206,15.3956785,15.040338,14.684997,14.329657,13.974316,14.316965,14.6596155,15.002265,15.344915,15.687565,13.127662,10.567759,8.007855,5.4479527,2.8880494,2.5345216,2.182807,1.8292793,1.4775645,1.1258497,1.1893034,1.2545701,1.3198367,1.3851035,1.4503701,1.4467441,1.4449311,1.4431182,1.4394923,1.4376793,1.3542831,1.2726997,1.1893034,1.1077201,1.0243238,1.2491312,1.4757515,1.7005589,1.9253663,2.1501737,2.5925364,3.0348995,3.4772623,3.919625,4.361988,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.2374981,0.34990177,0.46230546,0.5747091,0.6871128,0.5873999,0.48768693,0.387974,0.28826106,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07433146,0.15047589,0.22480737,0.2991388,0.37528324,0.51306844,0.6508536,0.7868258,0.9246109,1.062396,1.1131591,1.162109,1.2128719,1.261822,1.3125849,1.1131591,0.9119202,0.7124943,0.51306844,0.31182957,0.25018883,0.18673515,0.12509441,0.06164073,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,0.6508536,1.0497054,1.4503701,1.8492218,2.2498865,1.887294,1.5247015,1.162109,0.7995165,0.43692398,0.36259252,0.28826106,0.21211663,0.13778515,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.21211663,0.42423326,0.63816285,0.85027945,1.062396,0.85027945,0.63816285,0.42423326,0.21211663,0.0,1.1747998,2.3495996,3.5243993,4.699199,5.8758116,4.8623657,3.8507326,2.8372865,1.8256533,0.8122072,0.66173136,0.51306844,0.36259252,0.21211663,0.06164073,0.0870222,0.11240368,0.13778515,0.16316663,0.18673515,0.16316663,0.13778515,0.11240368,0.0870222,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.11240368,0.22480737,0.33721104,0.44961473,0.5620184,0.50037766,0.43692398,0.37528324,0.31182957,0.25018883,0.21211663,0.17585737,0.13778515,0.099712946,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.28826106,0.5747091,0.8629702,1.1494182,1.4376793,1.1494182,0.8629702,0.5747091,0.28826106,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.4757515,2.94969,4.4254417,5.89938,7.3751316,12.862969,18.348995,23.836832,29.324669,34.812508,28.650248,22.487988,16.323915,10.161655,3.9993954,4.4870825,4.974769,5.462456,5.9501433,6.43783,6.7496595,7.063302,7.3751316,7.686961,8.000604,6.412449,4.8242936,3.2379513,1.649796,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.5373923,3.0747845,4.612177,6.149569,7.686961,7.8120556,7.93715,8.062244,8.187339,8.312433,6.849373,5.388125,3.925064,2.4620032,1.0007553,1.2998942,1.6008459,1.8999848,2.1991236,2.5000753,2.8245957,3.149116,3.4754493,3.7999697,4.12449,4.5759177,5.0255322,5.475147,5.924762,6.3743763,6.037165,5.6999545,5.3627434,5.0255322,4.688321,5.0617914,5.4370747,5.812358,6.187641,6.5629244,8.125698,9.686659,11.249433,12.812206,14.37498,13.887294,13.399607,12.91192,12.4242325,11.938358,11.599335,11.262123,10.924912,10.587702,10.25049,11.037316,11.8241415,12.612781,13.399607,14.188245,13.274512,12.362592,11.450671,10.536939,9.625018,9.211663,8.80012,8.386765,7.9752226,7.5618668,7.137634,6.7134004,6.2873545,5.863121,5.4370747,4.699199,3.9631362,3.2252605,2.4873846,1.7495089,2.0758421,2.4003625,2.7248828,3.049403,3.3757362,3.7256382,4.07554,4.4254417,4.7753434,5.125245,5.6872635,6.249282,6.813113,7.3751316,7.93715,8.588004,9.237044,9.8878975,10.536939,11.187792,10.799818,10.411844,10.025683,9.637709,9.249735,10.487988,11.724429,12.962683,14.199123,15.437376,15.161806,14.888049,14.612478,14.336908,14.06315,14.811904,15.56247,16.313038,17.06179,17.812357,14.574407,11.336455,8.100317,4.8623657,1.6244144,1.4122978,1.2001812,0.9880646,0.774135,0.5620184,0.46230546,0.36259252,0.26287958,0.16316663,0.06164073,0.34990177,0.63816285,0.9246109,1.2128719,1.49932,1.3379664,1.1747998,1.0116332,0.85027945,0.6871128,0.8122072,0.93730164,1.062396,1.1874905,1.3125849,1.9126755,2.5127661,3.1128569,3.7129474,4.313038,0.5747091,0.5094425,0.44417584,0.38072214,0.3154555,0.25018883,0.23568514,0.21936847,0.20486477,0.19036107,0.17585737,0.1794833,0.18492219,0.19036107,0.19579996,0.19942589,0.3100166,0.42060733,0.5293851,0.6399758,0.7505665,0.629098,0.5094425,0.38978696,0.27013144,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.06707962,0.072518505,0.07795739,0.08339628,0.0870222,0.099712946,0.11240368,0.12509441,0.13778515,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.059827764,0.11965553,0.1794833,0.23931105,0.2991388,0.40972954,0.52032024,0.629098,0.73968875,0.85027945,0.90829426,0.9644961,1.0225109,1.0805258,1.1367276,0.968122,0.79770356,0.62728506,0.45686656,0.28826106,0.23568514,0.18310922,0.13053331,0.07795739,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.03988518,0.07977036,0.11965553,0.15954071,0.19942589,0.53482395,0.87022203,1.2056202,1.5392052,1.8746033,1.5809034,1.2853905,0.9898776,0.69436467,0.40066472,0.34083697,0.27919623,0.21936847,0.15954071,0.099712946,0.18492219,0.27013144,0.35534066,0.4405499,0.52575916,0.42423326,0.3245203,0.22480737,0.12509441,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.018129626,0.034446288,0.052575916,0.07070554,0.0870222,0.10696479,0.12690738,0.14684997,0.16679256,0.18673515,0.34083697,0.49312583,0.64541465,0.79770356,0.9499924,0.823085,0.69436467,0.56745726,0.4405499,0.31182957,1.3869164,2.4620032,3.53709,4.612177,5.6872635,4.6792564,3.673062,2.665055,1.6570477,0.6508536,0.533011,0.41516843,0.29732585,0.1794833,0.06164073,0.08520924,0.10696479,0.13053331,0.15228885,0.17585737,0.17767033,0.1794833,0.18310922,0.18492219,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08339628,0.16497959,0.24837588,0.32995918,0.41335547,0.32995918,0.24837588,0.16497959,0.08339628,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.032633327,0.027194439,0.02175555,0.018129626,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.018129626,0.034446288,0.052575916,0.07070554,0.0870222,0.07070554,0.052575916,0.034446288,0.018129626,0.0,0.12509441,0.25018883,0.37528324,0.50037766,0.62547207,0.7306239,0.83577573,0.93911463,1.0442665,1.1494182,1.0352017,0.91917205,0.80495536,0.69073874,0.5747091,0.4604925,0.3444629,0.23024625,0.11421664,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.23024625,0.4604925,0.69073874,0.91917205,1.1494182,0.91917205,0.69073874,0.4604925,0.23024625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,1.2056202,2.3967366,3.589666,4.782595,5.975525,10.662033,15.350354,20.036863,24.725183,29.411692,25.24913,21.08838,16.924006,12.763257,8.600695,8.074935,7.549176,7.02523,6.4994707,5.975525,6.156821,6.33993,6.5230393,6.7043357,6.887445,5.8903155,4.893186,3.8942437,2.8971143,1.8999848,1.5192627,1.1403534,0.75963134,0.38072214,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.260009,2.520018,3.780027,5.040036,6.300045,6.6118746,6.925517,7.2373466,7.549176,7.8628187,6.7641635,5.667321,4.5704784,3.4718235,2.374981,2.3441606,2.3151531,2.2843328,2.2553256,2.2245052,2.6269827,3.0294604,3.4319382,3.834416,4.2368937,4.599486,4.9620786,5.3246713,5.6872635,6.049856,5.6945157,5.3391747,4.985647,4.6303062,4.274966,4.6756306,5.0744824,5.475147,5.8758116,6.2746634,7.6833353,9.090195,10.497053,11.9057255,13.312584,13.062395,12.812206,12.562017,12.311829,12.06164,11.722616,11.381779,11.042755,10.701918,10.362894,11.104396,11.847711,12.589212,13.332527,14.075842,13.142166,12.210303,11.276628,10.344765,9.412902,9.003172,8.59163,8.1819,7.7721705,7.362441,6.8004227,6.2384043,5.674573,5.1125546,4.550536,4.062849,3.5751622,3.0874753,2.5997884,2.1121013,2.4583774,2.8028402,3.147303,3.491766,3.8380418,4.169814,4.503399,4.835171,5.1669436,5.5005283,5.979151,6.4595857,6.9400206,7.420456,7.900891,8.548119,9.195346,9.842574,10.489801,11.137029,10.823386,10.507931,10.192475,9.87702,9.563377,10.681975,11.802386,12.922797,14.043208,15.161806,14.947877,14.732134,14.518205,14.302462,14.0867195,14.755702,15.422873,16.090042,16.757214,17.424383,14.597975,11.769753,8.941531,6.115123,3.2869012,2.7774587,2.268016,1.7567607,1.2473183,0.73787576,0.60190356,0.46774435,0.33177215,0.19761293,0.06164073,0.29732585,0.533011,0.7668832,1.0025684,1.2382535,1.1022812,0.968122,0.8321498,0.6979906,0.5620184,0.6852999,0.80676836,0.9300498,1.0533313,1.1747998,1.7005589,2.2245052,2.7502642,3.2742105,3.7999697,1.1494182,1.020698,0.8901646,0.75963134,0.629098,0.50037766,0.46955732,0.4405499,0.40972954,0.38072214,0.34990177,0.33539808,0.3208944,0.3045777,0.29007402,0.2755703,0.3825351,0.4894999,0.5982776,0.70524246,0.8122072,0.6726091,0.533011,0.39159992,0.2520018,0.11240368,0.09064813,0.06707962,0.045324065,0.02175555,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.08520924,0.10696479,0.13053331,0.15228885,0.17585737,0.19942589,0.22480737,0.25018883,0.2755703,0.2991388,0.23931105,0.1794833,0.11965553,0.059827764,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.045324065,0.09064813,0.13415924,0.1794833,0.22480737,0.30820364,0.38978696,0.47318324,0.55476654,0.63816285,0.7016165,0.7668832,0.8321498,0.8974165,0.96268314,0.823085,0.68167394,0.5420758,0.40247768,0.26287958,0.21936847,0.17767033,0.13415924,0.092461094,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.42060733,0.69073874,0.96087015,1.2291887,1.49932,1.2726997,1.0442665,0.81764615,0.58921283,0.36259252,0.31726846,0.27194437,0.22662032,0.18310922,0.13778515,0.2955129,0.45324063,0.6091554,0.7668832,0.9246109,0.7505665,0.5747091,0.40066472,0.22480737,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.034446288,0.07070554,0.10515183,0.13959812,0.17585737,0.21574254,0.25562772,0.2955129,0.33539808,0.37528324,0.46774435,0.56020546,0.6526665,0.7451276,0.8375887,0.79589057,0.7523795,0.7106813,0.6671702,0.62547207,1.6008459,2.5744069,3.5497808,4.5251546,5.5005283,4.49796,3.4953918,2.4928236,1.4902552,0.48768693,0.40247768,0.31726846,0.23205921,0.14684997,0.06164073,0.08339628,0.10333887,0.12328146,0.14322405,0.16316663,0.19217403,0.2229944,0.2520018,0.28282216,0.31182957,0.25018883,0.18673515,0.12509441,0.06164073,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.16497959,0.32995918,0.4949388,0.65991837,0.824898,0.65991837,0.4949388,0.32995918,0.16497959,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03988518,0.07977036,0.11965553,0.15954071,0.19942589,0.15954071,0.11965553,0.07977036,0.03988518,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.065266654,0.054388877,0.045324065,0.034446288,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.034446288,0.07070554,0.10515183,0.13959812,0.17585737,0.13959812,0.10515183,0.07070554,0.034446288,0.0,0.13778515,0.2755703,0.41335547,0.5493277,0.6871128,0.96087015,1.2328146,1.504759,1.7767034,2.0504606,1.8582866,1.6642996,1.4721256,1.2799516,1.0877775,0.87022203,0.6526665,0.43511102,0.21755551,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.17223145,0.3444629,0.5166943,0.69073874,0.8629702,0.69073874,0.5166943,0.3444629,0.17223145,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.9354887,1.845596,2.7557032,3.6658103,4.574105,8.46291,12.349901,16.236893,20.125698,24.01269,21.849825,19.68696,17.524096,15.363045,13.200181,11.662788,10.125396,8.588004,7.0506115,5.5132194,5.565795,5.618371,5.669134,5.7217097,5.774286,5.368182,4.9602656,4.552349,4.1444325,3.738329,2.9895754,2.2426348,1.4956942,0.7469406,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.9826257,1.9652514,2.9478772,3.930503,4.9131284,5.411693,5.9120708,6.412449,6.9128265,7.413204,6.680767,5.9483304,5.2140803,4.4816437,3.7492065,3.39024,3.0294604,2.6704938,2.3097143,1.9507477,2.42937,2.909805,3.39024,3.870675,4.349297,4.6248674,4.900438,5.1741953,5.4497657,5.7253356,5.351866,4.9802084,4.606738,4.2350807,3.8616104,4.2876563,4.7118897,5.137936,5.562169,5.9882154,7.2409725,8.491917,9.744674,10.997431,12.250188,12.237497,12.224807,12.212116,12.199425,12.186734,11.844085,11.503247,11.160598,10.817947,10.475298,11.173288,11.869466,12.567456,13.265448,13.961625,13.009819,12.058014,11.104396,10.152591,9.200785,8.792869,8.384952,7.9770355,7.569119,7.1630154,6.4632115,5.763408,5.0617914,4.361988,3.6621845,3.4246864,3.1871881,2.94969,2.712192,2.474694,2.8409123,3.2053177,3.5697234,3.9341288,4.3003473,4.615803,4.9294453,5.2449007,5.560356,5.8758116,6.2728505,6.6698895,7.066928,7.46578,7.8628187,8.508233,9.151835,9.79725,10.442664,11.088079,10.845142,10.602205,10.359268,10.118144,9.875207,10.877775,11.880343,12.882912,13.885481,14.888049,14.732134,14.5780325,14.422117,14.268016,14.112101,14.697688,15.283275,15.867048,16.452635,17.038223,14.61973,12.203052,9.784559,7.36788,4.949388,4.1426196,3.3340383,2.5272698,1.7205015,0.9119202,0.7433147,0.5728962,0.40247768,0.23205921,0.06164073,0.24474995,0.42785916,0.6091554,0.79226464,0.97537386,0.8665961,0.75963134,0.6526665,0.54570174,0.43692398,0.55839247,0.678048,0.79770356,0.91735905,1.0370146,1.4866294,1.938057,2.3876717,2.8372865,3.2869012,1.7241274,1.5301404,1.3343405,1.1403534,0.9445535,0.7505665,0.70524246,0.65991837,0.61459434,0.56927025,0.52575916,0.4894999,0.4550536,0.42060733,0.38434806,0.34990177,0.4550536,0.56020546,0.6653573,0.7705091,0.87566096,0.71430725,0.55476654,0.39522585,0.23568514,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.10333887,0.14322405,0.18310922,0.2229944,0.26287958,0.2991388,0.33721104,0.37528324,0.41335547,0.44961473,0.36077955,0.27013144,0.1794833,0.09064813,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.20486477,0.25925365,0.3154555,0.36984438,0.42423326,0.49675176,0.56927025,0.6417888,0.71430725,0.7868258,0.678048,0.56745726,0.45686656,0.3480888,0.2374981,0.20486477,0.17223145,0.13959812,0.10696479,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.3045777,0.5094425,0.71430725,0.91917205,1.1258497,0.9644961,0.80495536,0.64541465,0.48587397,0.3245203,0.2955129,0.26469254,0.23568514,0.20486477,0.17585737,0.40429065,0.6345369,0.86478317,1.0950294,1.3252757,1.0750868,0.824898,0.5747091,0.3245203,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.052575916,0.10515183,0.15772775,0.21030366,0.26287958,0.32270733,0.3825351,0.44236287,0.50219065,0.5620184,0.5946517,0.62728506,0.65991837,0.69255173,0.72518504,0.7668832,0.8103943,0.8520924,0.89560354,0.93730164,1.8129625,2.6868105,3.5624714,4.4381323,5.3119802,4.314851,3.3177216,2.3205922,1.3216497,0.3245203,0.27194437,0.21936847,0.16679256,0.11421664,0.06164073,0.07977036,0.09789998,0.11421664,0.13234627,0.15047589,0.20667773,0.26469254,0.32270733,0.38072214,0.43692398,0.34990177,0.26287958,0.17585737,0.0870222,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.24837588,0.4949388,0.7433147,0.9898776,1.2382535,0.9898776,0.7433147,0.4949388,0.24837588,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.059827764,0.11965553,0.1794833,0.23931105,0.2991388,0.23931105,0.1794833,0.11965553,0.059827764,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.09789998,0.08339628,0.06707962,0.052575916,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.052575916,0.10515183,0.15772775,0.21030366,0.26287958,0.21030366,0.15772775,0.10515183,0.052575916,0.0,0.15047589,0.2991388,0.44961473,0.6000906,0.7505665,1.1893034,1.6298534,2.0704033,2.5091403,2.94969,2.6795588,2.4094272,2.1392958,1.8691645,1.6008459,1.2799516,0.96087015,0.6399758,0.3208944,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.11421664,0.23024625,0.3444629,0.4604925,0.5747091,0.4604925,0.3444629,0.23024625,0.11421664,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.6653573,1.2926424,1.9199274,2.5472124,3.1744974,6.261973,9.349448,12.436923,15.524399,18.611874,18.45052,18.287354,18.124187,17.962833,17.799667,15.250641,12.699803,10.150778,7.5999393,5.049101,4.972956,4.894999,4.8170414,4.740897,4.6629395,4.844236,5.027345,5.2104545,5.391751,5.57486,4.459888,3.3449159,2.229944,1.114972,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.70524246,1.4104849,2.1157274,2.819157,3.5243993,4.213325,4.900438,5.5875506,6.2746634,6.9617763,6.5955577,6.2275267,5.859495,5.4932766,5.125245,4.4345064,3.7455807,3.054842,2.3641033,1.6751775,2.231757,2.7901495,3.346729,3.9051213,4.461701,4.650249,4.836984,5.0255322,5.2122674,5.4008155,5.009216,4.6194286,4.229642,3.8398547,3.4500678,3.8996825,4.349297,4.800725,5.2503395,5.6999545,6.796797,7.895452,8.992294,10.089137,11.187792,11.4126,11.637406,11.862214,12.087022,12.311829,11.967366,11.622903,11.276628,10.932164,10.587702,11.240368,11.893035,12.545701,13.198368,13.849221,12.877473,11.9057255,10.932164,9.960417,8.9868555,8.582565,8.178274,7.7721705,7.36788,6.9617763,6.1241875,5.2884116,4.4508233,3.6132345,2.7756457,2.7883365,2.7992141,2.811905,2.8245957,2.8372865,3.2216346,3.6077955,3.9921436,4.3783045,4.762653,5.0599785,5.3573046,5.65463,5.9519563,6.249282,6.5647373,6.880193,7.1956487,7.509291,7.8247466,8.4683485,9.110137,9.751925,10.395528,11.037316,10.866898,10.698292,10.527874,10.357455,10.1870365,11.071762,11.958302,12.843027,13.727753,14.612478,14.518205,14.422117,14.327844,14.231756,14.137483,14.639673,15.141864,15.645867,16.148058,16.650248,14.641486,12.634536,10.627586,8.620637,6.6118746,5.5077806,4.401873,3.2977788,2.1918716,1.0877775,0.88291276,0.678048,0.47318324,0.26831847,0.06164073,0.19217403,0.32270733,0.45324063,0.581961,0.7124943,0.6327239,0.5529536,0.47318324,0.39159992,0.31182957,0.42967212,0.5475147,0.6653573,0.78319985,0.89922947,1.2745126,1.649796,2.0250793,2.4003625,2.7756457,2.3006494,2.039583,1.7803292,1.5192627,1.260009,1.0007553,0.93911463,0.8792868,0.8194591,0.75963134,0.69980353,0.64541465,0.58921283,0.53482395,0.48043507,0.42423326,0.5275721,0.629098,0.7324369,0.83577573,0.93730164,0.75781834,0.57833505,0.39703882,0.21755551,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.11965553,0.17767033,0.23568514,0.291887,0.34990177,0.40066472,0.44961473,0.50037766,0.5493277,0.6000906,0.48043507,0.36077955,0.23931105,0.11965553,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.10333887,0.13053331,0.15772775,0.18492219,0.21211663,0.291887,0.37165734,0.45324063,0.533011,0.61278135,0.533011,0.45324063,0.37165734,0.291887,0.21211663,0.19036107,0.16679256,0.14503701,0.12328146,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.19036107,0.32995918,0.46955732,0.6091554,0.7505665,0.65810543,0.5656443,0.47318324,0.38072214,0.28826106,0.27194437,0.2574407,0.24293698,0.22662032,0.21211663,0.5148814,0.81764615,1.1204109,1.4231756,1.7241274,1.3996071,1.0750868,0.7505665,0.42423326,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07070554,0.13959812,0.21030366,0.27919623,0.34990177,0.42967212,0.5094425,0.58921283,0.67079616,0.7505665,0.72337204,0.69436467,0.6671702,0.6399758,0.61278135,0.73968875,0.8665961,0.99531645,1.1222239,1.2491312,2.0250793,2.7992141,3.5751622,4.349297,5.125245,4.1317415,3.1400511,2.1483607,1.1548572,0.16316663,0.14322405,0.12328146,0.10333887,0.08339628,0.06164073,0.07795739,0.092461094,0.10696479,0.12328146,0.13778515,0.2229944,0.30820364,0.39159992,0.47680917,0.5620184,0.44961473,0.33721104,0.22480737,0.11240368,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.32995918,0.65991837,0.9898776,1.3198367,1.649796,1.3198367,0.9898776,0.65991837,0.32995918,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07977036,0.15954071,0.23931105,0.3208944,0.40066472,0.3208944,0.23931105,0.15954071,0.07977036,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.13053331,0.11059072,0.09064813,0.07070554,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07070554,0.13959812,0.21030366,0.27919623,0.34990177,0.27919623,0.21030366,0.13959812,0.07070554,0.0,0.16316663,0.3245203,0.48768693,0.6508536,0.8122072,1.4195497,2.0268922,2.6342347,3.24339,3.8507326,3.5026438,3.1545548,2.808279,2.4601903,2.1121013,1.6896812,1.2672608,0.8448406,0.4224203,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.058014803,0.11421664,0.17223145,0.23024625,0.28826106,0.23024625,0.17223145,0.11421664,0.058014803,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.39522585,0.73968875,1.0841516,1.4304274,1.7748904,4.062849,6.3489947,8.636953,10.924912,13.212872,15.049402,16.887747,18.724277,20.562622,22.400965,18.836681,15.276023,11.711739,8.149267,4.5867953,4.3801174,4.171627,3.9649491,3.7582715,3.5497808,4.322103,5.0944247,5.866747,6.640882,7.413204,5.9302006,4.4471974,2.9641938,1.4830034,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.42785916,0.8557183,1.2817645,1.7096237,2.137483,3.0131438,3.8869917,4.762653,5.638314,6.5121617,6.510349,6.506723,6.5049095,6.5030966,6.4994707,5.480586,4.459888,3.43919,2.420305,1.3996071,2.034144,2.6704938,3.3050308,3.9395678,4.574105,4.6756306,4.7753434,4.8750563,4.974769,5.0744824,4.666566,4.2604623,3.8525455,3.444629,3.0367124,3.5117085,3.9867048,4.461701,4.936697,5.411693,6.354434,7.2971745,8.239915,9.182655,10.125396,10.587702,11.050007,11.512312,11.974618,12.436923,12.090648,11.7425585,11.39447,11.048194,10.700105,11.307447,11.91479,12.522133,13.129475,13.736817,12.745127,11.751623,10.7599325,9.768243,8.774739,8.372261,7.9697833,7.567306,7.1648283,6.7623506,5.7869763,4.8134155,3.8380418,2.8626678,1.887294,2.1501737,2.4130533,2.6741197,2.9369993,3.199879,3.6041696,4.0102735,4.4145637,4.8206677,5.224958,5.504154,5.7851634,6.0643597,6.345369,6.624565,6.8566246,7.0904965,7.322556,7.554615,7.7866745,8.42665,9.068439,9.708415,10.346578,10.988366,10.890467,10.792566,10.694666,10.596766,10.500679,11.267563,12.034446,12.803142,13.5700245,14.336908,14.302462,14.268016,14.231756,14.19731,14.162864,14.581658,15.002265,15.422873,15.841667,16.262274,14.665054,13.067834,11.470614,9.873394,8.274362,6.872941,5.469708,4.068288,2.665055,1.261822,1.0225109,0.78319985,0.5420758,0.30276474,0.06164073,0.13959812,0.21755551,0.2955129,0.37165734,0.44961473,0.39703882,0.3444629,0.291887,0.23931105,0.18673515,0.30276474,0.4169814,0.533011,0.64722764,0.76325727,1.062396,1.3633479,1.6624867,1.9616255,2.2625773,2.8753586,2.5508385,2.2245052,1.8999848,1.5754645,1.2491312,1.1747998,1.1004683,1.0243238,0.9499924,0.87566096,0.7995165,0.72518504,0.6508536,0.5747091,0.50037766,0.6000906,0.69980353,0.7995165,0.89922947,1.0007553,0.7995165,0.6000906,0.40066472,0.19942589,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.13778515,0.21211663,0.28826106,0.36259252,0.43692398,0.50037766,0.5620184,0.62547207,0.6871128,0.7505665,0.6000906,0.44961473,0.2991388,0.15047589,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0870222,0.17585737,0.26287958,0.34990177,0.43692398,0.387974,0.33721104,0.28826106,0.2374981,0.18673515,0.17585737,0.16316663,0.15047589,0.13778515,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07433146,0.15047589,0.22480737,0.2991388,0.37528324,0.34990177,0.3245203,0.2991388,0.2755703,0.25018883,0.25018883,0.25018883,0.25018883,0.25018883,0.25018883,0.62547207,1.0007553,1.3742256,1.7495089,2.124792,1.7241274,1.3252757,0.9246109,0.52575916,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0870222,0.17585737,0.26287958,0.34990177,0.43692398,0.53663695,0.63816285,0.73787576,0.8375887,0.93730164,0.85027945,0.76325727,0.6744221,0.5873999,0.50037766,0.7124943,0.9246109,1.1367276,1.3506571,1.5627737,2.2371957,2.911618,3.587853,4.262275,4.936697,3.9504454,2.962381,1.9743162,0.9880646,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.2374981,0.34990177,0.46230546,0.5747091,0.6871128,0.5493277,0.41335547,0.2755703,0.13778515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.41335547,0.824898,1.2382535,1.649796,2.0631514,1.649796,1.2382535,0.824898,0.41335547,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.099712946,0.19942589,0.2991388,0.40066472,0.50037766,0.40066472,0.2991388,0.19942589,0.099712946,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.16316663,0.13778515,0.11240368,0.0870222,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0870222,0.17585737,0.26287958,0.34990177,0.43692398,0.34990177,0.26287958,0.17585737,0.0870222,0.0,0.17585737,0.34990177,0.52575916,0.69980353,0.87566096,1.649796,2.4257438,3.199879,3.975827,4.749962,4.325729,3.8996825,3.4754493,3.049403,2.6251698,2.0994108,1.5754645,1.0497054,0.52575916,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.12509441,0.18673515,0.25018883,0.31182957,0.37528324,1.8619126,3.350355,4.836984,6.3254266,7.8120556,11.650098,15.488139,19.324368,23.16241,27.000452,22.424534,17.85043,13.274512,8.700407,4.12449,3.787279,3.4500678,3.1128569,2.7756457,2.4366217,3.7999697,5.163317,6.5248523,7.8882003,9.249735,7.400513,5.5494785,3.7002566,1.8492218,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.15047589,0.2991388,0.44961473,0.6000906,0.7505665,1.8129625,2.8753586,3.9377546,5.0001507,6.0625467,6.4251394,6.787732,7.1503243,7.512917,7.8755093,6.5248523,5.1741953,3.825351,2.474694,1.1258497,1.8383441,2.5508385,3.2633326,3.975827,4.688321,4.699199,4.7118897,4.7245803,4.7372713,4.749962,4.325729,3.8996825,3.4754493,3.049403,2.6251698,3.1255474,3.6241121,4.12449,4.6248674,5.125245,5.9120708,6.70071,7.4875355,8.274362,9.063,9.762803,10.462607,11.162411,11.862214,12.562017,12.212116,11.862214,11.512312,11.162411,10.812509,11.374527,11.938358,12.500377,13.062395,13.6244135,12.612781,11.599335,10.587702,9.574255,8.562622,8.161958,7.763106,7.362441,6.9617763,6.5629244,5.4497657,4.3384194,3.2252605,2.1121013,1.0007553,1.5120108,2.0250793,2.5381477,3.049403,3.5624714,3.9867048,4.4127507,4.836984,5.2630305,5.6872635,5.9501433,6.2130227,6.4759026,6.736969,6.9998484,7.1503243,7.3008003,7.4494634,7.5999393,7.750415,8.386765,9.024928,9.663091,10.29944,10.937603,10.912222,10.88684,10.863272,10.837891,10.812509,11.463363,12.112403,12.763257,13.412297,14.06315,14.0867195,14.112101,14.137483,14.162864,14.188245,14.525456,14.862667,15.199879,15.537089,15.8743,14.68681,13.499319,12.311829,11.124338,9.936848,8.238102,6.5375433,4.836984,3.1382382,1.4376793,1.162109,0.8883517,0.61278135,0.33721104,0.06164073,0.0870222,0.11240368,0.13778515,0.16316663,0.18673515,0.16316663,0.13778515,0.11240368,0.0870222,0.06164073,0.17585737,0.28826106,0.40066472,0.51306844,0.62547207,0.85027945,1.0750868,1.2998942,1.5247015,1.7495089,3.636803,3.1871881,2.7375734,2.2879589,1.8383441,1.3869164,1.4576219,1.5283275,1.5972201,1.6679256,1.7368182,1.7041848,1.6733645,1.6407311,1.6080978,1.5754645,1.5881553,1.6008459,1.6117238,1.6244144,1.6371052,1.3343405,1.0333886,0.7306239,0.42785916,0.12509441,0.2229944,0.3208944,0.4169814,0.5148814,0.61278135,0.5148814,0.4169814,0.3208944,0.2229944,0.12509441,0.18673515,0.25018883,0.31182957,0.37528324,0.43692398,0.5058166,0.5728962,0.6399758,0.7070554,0.774135,0.6508536,0.52575916,0.40066472,0.2755703,0.15047589,0.13234627,0.11421664,0.09789998,0.07977036,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07070554,0.13959812,0.21030366,0.27919623,0.34990177,0.3100166,0.27013144,0.23024625,0.19036107,0.15047589,0.14322405,0.13415924,0.12690738,0.11965553,0.11240368,0.09064813,0.06707962,0.045324065,0.02175555,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.059827764,0.11965553,0.1794833,0.23931105,0.2991388,0.27919623,0.25925365,0.23931105,0.21936847,0.19942589,0.19942589,0.19942589,0.19942589,0.19942589,0.19942589,0.51306844,0.824898,1.1367276,1.4503701,1.7621996,1.4304274,1.0968424,0.7650702,0.43329805,0.099712946,0.08520924,0.07070554,0.054388877,0.03988518,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.15047589,1.0116332,1.8746033,2.7375734,3.6005437,4.461701,4.004834,3.5479677,3.0892882,2.6324217,2.175555,1.7531348,1.3307146,0.90829426,0.48587397,0.06164073,0.07070554,0.07795739,0.08520924,0.092461094,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.05076295,0.0870222,0.12509441,0.16316663,0.19942589,0.15954071,0.11965553,0.07977036,0.03988518,0.0,0.07070554,0.13959812,0.21030366,0.27919623,0.34990177,0.42967212,0.5094425,0.58921283,0.67079616,0.7505665,0.67986095,0.6091554,0.5402629,0.46955732,0.40066472,0.5728962,0.7451276,0.91735905,1.0895905,1.261822,1.8075237,2.3532255,2.8971143,3.442816,3.9867048,3.2198215,2.4529383,1.6842422,0.91735905,0.15047589,0.30276474,0.4550536,0.6073425,0.75963134,0.9119202,0.7650702,0.61822027,0.46955732,0.32270733,0.17585737,0.29007402,0.40429065,0.52032024,0.6345369,0.7505665,0.6055295,0.4604925,0.3154555,0.17041849,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.32995918,0.65991837,0.9898776,1.3198367,1.649796,1.3198367,0.9898776,0.65991837,0.32995918,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07977036,0.15954071,0.23931105,0.3208944,0.40066472,0.3208944,0.23931105,0.15954071,0.07977036,0.0,0.12509441,0.25018883,0.37528324,0.50037766,0.62547207,0.62728506,0.630911,0.6327239,0.6345369,0.63816285,0.5094425,0.3825351,0.25562772,0.12690738,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.030820364,0.034446288,0.03988518,0.045324065,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.13415924,0.11965553,0.10515183,0.09064813,0.07433146,0.08339628,0.09064813,0.09789998,0.10515183,0.11240368,0.11784257,0.12328146,0.12690738,0.13234627,0.13778515,0.11240368,0.0870222,0.06164073,0.038072214,0.012690738,0.047137026,0.08339628,0.11784257,0.15228885,0.18673515,0.15954071,0.13234627,0.10515183,0.07795739,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0870222,0.17585737,0.26287958,0.34990177,0.43692398,0.36440548,0.291887,0.21936847,0.14684997,0.07433146,0.19942589,0.3245203,0.44961473,0.5747091,0.69980353,1.3506571,1.9996977,2.6505513,3.299592,3.9504454,3.729264,3.5098956,3.290527,3.0693457,2.8499773,2.3006494,1.7495089,1.2001812,0.6508536,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,0.2991388,1.7150626,3.1291735,4.5450974,5.959208,7.3751316,10.469859,13.564586,16.659313,19.755854,22.85058,19.072367,15.294152,11.517752,7.7395372,3.9631362,3.7256382,3.48814,3.2506418,3.0131438,2.7756457,3.9830787,5.1905117,6.397945,7.605378,8.812811,7.066928,5.3228583,3.576975,1.8329052,0.0870222,0.07070554,0.052575916,0.034446288,0.018129626,0.0,0.018129626,0.034446288,0.052575916,0.07070554,0.0870222,0.13778515,0.18673515,0.2374981,0.28826106,0.33721104,0.41516843,0.49312583,0.56927025,0.64722764,0.72518504,1.8528478,2.9805105,4.1081734,5.235836,6.3616858,6.773228,7.1829576,7.592687,8.002417,8.412147,7.3751316,6.338117,5.2992897,4.262275,3.2252605,3.444629,3.6658103,3.8851788,4.1045475,4.325729,4.25321,4.1806917,4.1081734,4.0356545,3.9631362,3.5932918,3.2216346,2.8517902,2.4819458,2.1121013,2.521831,2.9333735,3.343103,3.7528327,4.162562,4.784408,5.408067,6.0299134,6.6517596,7.2754188,7.8483152,8.419398,8.992294,9.56519,10.138086,9.857078,9.577881,9.296872,9.017676,8.736667,9.583321,10.428161,11.273002,12.117842,12.962683,12.427858,11.893035,11.358211,10.823386,10.28675,9.570629,8.852696,8.134763,7.41683,6.70071,5.6401267,4.5795436,3.5207734,2.4601903,1.3996071,1.7223145,2.0450218,2.3677292,2.6904364,3.0131438,3.3576066,3.7020695,4.0483456,4.3928084,4.7372713,5.3971896,6.057108,6.717026,7.3769445,8.036863,7.8755093,7.7123427,7.549176,7.3878226,7.224656,7.703278,8.180087,8.656897,9.135518,9.612328,9.944099,10.277685,10.609457,10.943042,11.274815,11.543133,11.809638,12.077957,12.344462,12.612781,12.951805,13.292642,13.631665,13.972503,14.313339,14.757515,15.201692,15.64768,16.091856,16.537846,15.607795,14.677745,13.747695,12.817645,11.887595,10.29944,8.713099,7.124943,5.5367875,3.9504454,3.4500678,2.94969,2.4493124,1.9507477,1.4503701,1.2328146,1.015259,0.79770356,0.58014804,0.36259252,0.32814622,0.291887,0.2574407,0.2229944,0.18673515,0.27738327,0.3680314,0.45686656,0.5475147,0.63816285,0.8031424,0.968122,1.1331016,1.2980812,1.4630609,4.40006,3.825351,3.2506418,2.6741197,2.0994108,1.5247015,1.7404441,1.9543737,2.1701162,2.3858588,2.5997884,2.610666,2.619731,2.6306088,2.6396735,2.6505513,2.5744069,2.5000753,2.4257438,2.3495996,2.275268,1.8691645,1.4648738,1.0605831,0.6544795,0.25018883,0.44417584,0.6399758,0.83577573,1.0297627,1.2255627,1.017072,0.8103943,0.60190356,0.39522585,0.18673515,0.2374981,0.28826106,0.33721104,0.387974,0.43692398,0.5094425,0.581961,0.6544795,0.726998,0.7995165,0.69980353,0.6000906,0.50037766,0.40066472,0.2991388,0.26469254,0.23024625,0.19579996,0.15954071,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.052575916,0.10515183,0.15772775,0.21030366,0.26287958,0.23205921,0.2030518,0.17223145,0.14322405,0.11240368,0.11059072,0.10696479,0.10515183,0.10333887,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.045324065,0.09064813,0.13415924,0.1794833,0.22480737,0.21030366,0.19579996,0.1794833,0.16497959,0.15047589,0.15047589,0.15047589,0.15047589,0.15047589,0.15047589,0.40066472,0.6508536,0.89922947,1.1494182,1.3996071,1.1349145,0.87022203,0.6055295,0.34083697,0.07433146,0.07070554,0.065266654,0.059827764,0.054388877,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,0.2991388,2.0250793,3.7492065,5.475147,7.1992745,8.925215,8.009668,7.0959353,6.1803894,5.2648435,4.349297,3.5044568,2.659616,1.8147756,0.969935,0.12509441,0.11421664,0.10515183,0.09427405,0.08520924,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.099712946,0.17585737,0.25018883,0.3245203,0.40066472,0.3208944,0.23931105,0.15954071,0.07977036,0.0,0.052575916,0.10515183,0.15772775,0.21030366,0.26287958,0.32270733,0.3825351,0.44236287,0.50219065,0.5620184,0.5094425,0.45686656,0.40429065,0.35171473,0.2991388,0.43329805,0.5656443,0.6979906,0.83033687,0.96268314,1.3778516,1.79302,2.2081885,2.6233568,3.0367124,2.4891977,1.9416829,1.3941683,0.8466535,0.2991388,0.59283876,0.88472575,1.1766127,1.4703126,1.7621996,1.455809,1.1476053,0.83940166,0.533011,0.22480737,0.34264994,0.4604925,0.57833505,0.69436467,0.8122072,0.65991837,0.5076295,0.35534066,0.2030518,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.24837588,0.4949388,0.7433147,0.9898776,1.2382535,0.9898776,0.7433147,0.4949388,0.24837588,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.059827764,0.11965553,0.1794833,0.23931105,0.2991388,0.23931105,0.1794833,0.11965553,0.059827764,0.0,0.25018883,0.50037766,0.7505665,1.0007553,1.2491312,1.2545701,1.260009,1.2654479,1.2708868,1.2745126,1.020698,0.7650702,0.5094425,0.25562772,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.059827764,0.07070554,0.07977036,0.09064813,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.059827764,0.11965553,0.1794833,0.23931105,0.2991388,0.27013144,0.23931105,0.21030366,0.1794833,0.15047589,0.16497959,0.1794833,0.19579996,0.21030366,0.22480737,0.23568514,0.24474995,0.25562772,0.26469254,0.2755703,0.22480737,0.17585737,0.12509441,0.07433146,0.025381476,0.058014803,0.09064813,0.12328146,0.15410182,0.18673515,0.15772775,0.12690738,0.09789998,0.06707962,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0870222,0.17585737,0.26287958,0.34990177,0.43692398,0.38072214,0.32270733,0.26469254,0.20667773,0.15047589,0.22480737,0.2991388,0.37528324,0.44961473,0.52575916,1.0497054,1.5754645,2.0994108,2.6251698,3.149116,3.1346123,3.1201086,3.105605,3.0892882,3.0747845,2.5000753,1.9253663,1.3506571,0.774135,0.19942589,0.15954071,0.11965553,0.07977036,0.03988518,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.22480737,1.5682126,2.909805,4.25321,5.5948024,6.9382076,9.28962,11.642846,13.994258,16.347483,18.700708,15.720199,12.739688,9.759177,6.78048,3.7999697,3.6621845,3.5243993,3.386614,3.2506418,3.1128569,4.164375,5.217706,6.2692246,7.322556,8.375887,6.735156,5.0944247,3.4555066,1.8147756,0.17585737,0.13959812,0.10515183,0.07070554,0.034446288,0.0,0.034446288,0.07070554,0.10515183,0.13959812,0.17585737,0.2755703,0.37528324,0.4749962,0.5747091,0.6744221,0.67986095,0.6852999,0.69073874,0.69436467,0.69980353,1.892733,3.0856624,4.2767787,5.469708,6.6626377,7.119504,7.5781837,8.03505,8.491917,8.950596,8.225411,7.500226,6.775041,6.049856,5.3246713,5.0527267,4.780782,4.507025,4.2350807,3.9631362,3.8054085,3.6476808,3.489953,3.3322253,3.1744974,2.8608549,2.5453994,2.229944,1.9144884,1.6008459,1.9199274,2.2408218,2.5599031,2.8807976,3.199879,3.6567454,4.115425,4.572292,5.029158,5.487838,5.9320135,6.378002,6.8221784,7.268167,7.7123427,7.502039,7.2917356,7.083245,6.872941,6.6626377,7.7903004,8.917963,10.045626,11.173288,12.299138,12.242936,12.184921,12.126906,12.070704,12.012691,10.9774885,9.9422865,8.907085,7.8718834,6.836682,5.8304877,4.8224807,3.8144734,2.808279,1.8002719,1.9326181,2.0649643,2.1973107,2.3296568,2.4620032,2.7266958,2.9932013,3.2578938,3.5225863,3.787279,4.844236,5.903006,6.9599633,8.01692,9.07569,8.600695,8.125698,7.650702,7.175706,6.70071,7.017978,7.3352466,7.652515,7.9697833,8.287052,8.977791,9.666717,10.357455,11.048194,11.73712,11.622903,11.506873,11.392657,11.276628,11.162411,11.81689,12.473183,13.127662,13.782142,14.436621,14.989574,15.542528,16.095482,16.646622,17.199575,16.526966,15.854358,15.181748,14.510953,13.838344,12.362592,10.88684,9.412902,7.93715,6.4632115,5.7380266,5.0128417,4.2876563,3.5624714,2.8372865,2.3767939,1.9181144,1.4576219,0.99712944,0.53663695,0.49312583,0.44780177,0.40247768,0.35715362,0.31182957,0.38072214,0.44780177,0.5148814,0.581961,0.6508536,0.7541924,0.85934424,0.9644961,1.0696479,1.1747998,5.163317,4.461701,3.7618973,3.0620937,2.3622901,1.6624867,2.0232663,2.382233,2.7430124,3.101979,3.4627585,3.5153344,3.5679104,3.6204863,3.673062,3.7256382,3.5624714,3.3993049,3.2379513,3.0747845,2.911618,2.4058013,1.8981718,1.3905423,0.88291276,0.37528324,0.6671702,0.96087015,1.2527572,1.5446441,1.8383441,1.5192627,1.2019942,0.88472575,0.56745726,0.25018883,0.28826106,0.3245203,0.36259252,0.40066472,0.43692398,0.5148814,0.59283876,0.67079616,0.7469406,0.824898,0.7505665,0.6744221,0.6000906,0.52575916,0.44961473,0.39703882,0.3444629,0.291887,0.23931105,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.034446288,0.07070554,0.10515183,0.13959812,0.17585737,0.15410182,0.13415924,0.11421664,0.09427405,0.07433146,0.07795739,0.07977036,0.08339628,0.08520924,0.0870222,0.07070554,0.052575916,0.034446288,0.018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.13959812,0.13053331,0.11965553,0.11059072,0.099712946,0.099712946,0.099712946,0.099712946,0.099712946,0.099712946,0.28826106,0.4749962,0.66173136,0.85027945,1.0370146,0.83940166,0.6417888,0.44417584,0.24837588,0.05076295,0.054388877,0.059827764,0.065266654,0.07070554,0.07433146,0.15047589,0.22480737,0.2991388,0.37528324,0.44961473,3.0367124,5.6256227,8.212721,10.799818,13.386916,12.0145035,10.642091,9.269678,7.897265,6.5248523,5.2575917,3.9903307,2.72307,1.455809,0.18673515,0.15954071,0.13234627,0.10515183,0.07795739,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.15047589,0.26287958,0.37528324,0.48768693,0.6000906,0.48043507,0.36077955,0.23931105,0.11965553,0.0,0.034446288,0.07070554,0.10515183,0.13959812,0.17585737,0.21574254,0.25562772,0.2955129,0.33539808,0.37528324,0.34083697,0.3045777,0.27013144,0.23568514,0.19942589,0.291887,0.38434806,0.47680917,0.56927025,0.66173136,0.9481794,1.2328146,1.5174497,1.8020848,2.08672,1.7603867,1.4322405,1.1040943,0.7777609,0.44961473,0.88291276,1.3143979,1.7476959,2.179181,2.612479,2.1447346,1.6769904,1.209246,0.7433147,0.2755703,0.39522585,0.5148814,0.6345369,0.7541924,0.87566096,0.71430725,0.55476654,0.39522585,0.23568514,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.16497959,0.32995918,0.4949388,0.65991837,0.824898,0.65991837,0.4949388,0.32995918,0.16497959,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03988518,0.07977036,0.11965553,0.15954071,0.19942589,0.15954071,0.11965553,0.07977036,0.03988518,0.0,0.37528324,0.7505665,1.1258497,1.49932,1.8746033,1.8818551,1.889107,1.8981718,1.9054236,1.9126755,1.5301404,1.1476053,0.7650702,0.3825351,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.09064813,0.10515183,0.11965553,0.13415924,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.09064813,0.1794833,0.27013144,0.36077955,0.44961473,0.40429065,0.36077955,0.3154555,0.27013144,0.22480737,0.24837588,0.27013144,0.291887,0.3154555,0.33721104,0.35171473,0.3680314,0.3825351,0.39703882,0.41335547,0.33721104,0.26287958,0.18673515,0.11240368,0.038072214,0.06707962,0.09789998,0.12690738,0.15772775,0.18673515,0.15410182,0.12328146,0.09064813,0.058014803,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0870222,0.17585737,0.26287958,0.34990177,0.43692398,0.39522585,0.35171473,0.3100166,0.26831847,0.22480737,0.25018883,0.2755703,0.2991388,0.3245203,0.34990177,0.7505665,1.1494182,1.550083,1.9507477,2.3495996,2.5399606,2.7303216,2.9206827,3.1092308,3.299592,2.6995013,2.0994108,1.49932,0.89922947,0.2991388,0.23931105,0.1794833,0.11965553,0.059827764,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.15047589,1.4195497,2.6904364,3.9595103,5.230397,6.4994707,8.109382,9.719293,11.329204,12.940927,14.5508375,12.368031,10.185224,8.002417,5.81961,3.636803,3.6005437,3.5624714,3.5243993,3.48814,3.4500678,4.347484,5.2449007,6.1423173,7.039734,7.93715,6.401571,4.8678045,3.3322253,1.7966459,0.26287958,0.21030366,0.15772775,0.10515183,0.052575916,0.0,0.052575916,0.10515183,0.15772775,0.21030366,0.26287958,0.41335547,0.5620184,0.7124943,0.8629702,1.0116332,0.9445535,0.8774739,0.8103943,0.7433147,0.6744221,1.9326181,3.1908143,4.4471974,5.7053933,6.9617763,7.4675927,7.9715962,8.477413,8.98323,9.487233,9.07569,8.662335,8.2507925,7.837437,7.424082,6.6608243,5.8957543,5.130684,4.365614,3.6005437,3.3576066,3.1146698,2.8717327,2.6306088,2.3876717,2.126605,1.8673514,1.6080978,1.3470312,1.0877775,1.3180238,1.54827,1.7767034,2.0069497,2.2371957,2.5308957,2.8227828,3.1146698,3.4083695,3.7002566,4.017525,4.3347936,4.652062,4.9693303,5.2884116,5.147001,5.0074024,4.8678045,4.7282066,4.5867953,5.99728,7.407765,8.81825,10.226922,11.637406,12.058014,12.476809,12.897416,13.318023,13.736817,12.384347,11.0318775,9.679407,8.326937,6.9744673,6.019036,5.0654173,4.1099863,3.1545548,2.1991236,2.1429217,2.084907,2.0268922,1.9706904,1.9126755,2.0975976,2.2825198,2.467442,2.6523643,2.8372865,4.2930956,5.7470913,7.2029004,8.656897,10.112705,9.324066,8.537241,7.750415,6.9617763,6.1749506,6.3326783,6.490406,6.6481338,6.8058615,6.9617763,8.009668,9.057561,10.1054535,11.151533,12.199425,11.702674,11.204109,10.707357,10.210606,9.712041,10.681975,11.651911,12.621845,13.591781,14.561715,15.221634,15.883366,16.543283,17.203201,17.863121,17.447952,17.032784,16.617615,16.202446,15.787278,14.425743,13.062395,11.699047,10.337513,8.974165,8.024173,7.07418,6.1241875,5.1741953,4.2242026,3.5225863,2.819157,2.1175404,1.4159238,0.7124943,0.65810543,0.60190356,0.5475147,0.49312583,0.43692398,0.48224804,0.5275721,0.5728962,0.61822027,0.66173136,0.7070554,0.7523795,0.79770356,0.8430276,0.8883517,5.924762,5.0998635,4.274966,3.4500678,2.6251698,1.8002719,2.3042755,2.810092,3.3159087,3.8199122,4.325729,4.420003,4.514277,4.610364,4.704638,4.800725,4.550536,4.3003473,4.0501585,3.7999697,3.5497808,2.9406252,2.3296568,1.7205015,1.1095331,0.50037766,0.8901646,1.2799516,1.6697385,2.0595255,2.4493124,2.0232663,1.5954071,1.167548,0.73968875,0.31182957,0.33721104,0.36259252,0.387974,0.41335547,0.43692398,0.52032024,0.60190356,0.6852999,0.7668832,0.85027945,0.7995165,0.7505665,0.69980353,0.6508536,0.6000906,0.5293851,0.4604925,0.38978696,0.3208944,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.018129626,0.034446288,0.052575916,0.07070554,0.0870222,0.07795739,0.06707962,0.058014803,0.047137026,0.038072214,0.045324065,0.052575916,0.059827764,0.06707962,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.07070554,0.065266654,0.059827764,0.054388877,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.17585737,0.2991388,0.42423326,0.5493277,0.6744221,0.54570174,0.41516843,0.28463513,0.15410182,0.025381476,0.03988518,0.054388877,0.07070554,0.08520924,0.099712946,0.19942589,0.2991388,0.40066472,0.50037766,0.6000906,4.0501585,7.500226,10.950294,14.400362,17.85043,16.019337,14.190058,12.360779,10.529687,8.700407,7.0107265,5.319232,3.6295512,1.93987,0.25018883,0.20486477,0.15954071,0.11421664,0.07070554,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.19942589,0.34990177,0.50037766,0.6508536,0.7995165,0.6399758,0.48043507,0.3208944,0.15954071,0.0,0.018129626,0.034446288,0.052575916,0.07070554,0.0870222,0.10696479,0.12690738,0.14684997,0.16679256,0.18673515,0.17041849,0.15228885,0.13415924,0.11784257,0.099712946,0.15228885,0.20486477,0.2574407,0.3100166,0.36259252,0.5166943,0.6726091,0.82671094,0.9826257,1.1367276,1.0297627,0.922798,0.81583315,0.7070554,0.6000906,1.1729867,1.745883,2.3169663,2.8898623,3.4627585,2.8354735,2.2081885,1.5790904,0.95180535,0.3245203,0.44780177,0.56927025,0.69255173,0.81583315,0.93730164,0.7705091,0.60190356,0.43511102,0.26831847,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0,0.0,0.0,0.0,0.0,0.08339628,0.16497959,0.24837588,0.32995918,0.41335547,0.32995918,0.24837588,0.16497959,0.08339628,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.50037766,1.0007553,1.49932,1.9996977,2.5000753,2.5091403,2.520018,2.5308957,2.5399606,2.5508385,2.039583,1.5301404,1.020698,0.5094425,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.11965553,0.13959812,0.15954071,0.1794833,0.19942589,0.15954071,0.11965553,0.07977036,0.03988518,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.11965553,0.23931105,0.36077955,0.48043507,0.6000906,0.5402629,0.48043507,0.42060733,0.36077955,0.2991388,0.32995918,0.36077955,0.38978696,0.42060733,0.44961473,0.46955732,0.4894999,0.5094425,0.5293851,0.5493277,0.44961473,0.34990177,0.25018883,0.15047589,0.05076295,0.07795739,0.10515183,0.13234627,0.15954071,0.18673515,0.15228885,0.11784257,0.08339628,0.047137026,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0870222,0.17585737,0.26287958,0.34990177,0.43692398,0.40972954,0.3825351,0.35534066,0.32814622,0.2991388,0.2755703,0.25018883,0.22480737,0.19942589,0.17585737,0.44961473,0.72518504,1.0007553,1.2745126,1.550083,1.9453088,2.3405347,2.7357605,3.1291735,3.5243993,2.9007401,2.275268,1.649796,1.0243238,0.40066472,0.3208944,0.23931105,0.15954071,0.07977036,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.07433146,1.2726997,2.469255,3.6676233,4.8641787,6.0625467,6.929143,7.797552,8.664148,9.5325575,10.399154,9.01405,7.6307597,6.245656,4.860553,3.4754493,3.53709,3.6005437,3.6621845,3.7256382,3.787279,4.5305934,5.272095,6.01541,6.7569118,7.500226,6.069799,4.6393714,3.2107568,1.7803292,0.34990177,0.27919623,0.21030366,0.13959812,0.07070554,0.0,0.07070554,0.13959812,0.21030366,0.27919623,0.34990177,0.5493277,0.7505665,0.9499924,1.1494182,1.3506571,1.209246,1.0696479,0.9300498,0.7904517,0.6508536,1.9725033,3.294153,4.6176157,5.9392653,7.262728,7.8156815,8.366822,8.919776,9.47273,10.025683,9.924157,9.824444,9.724731,9.625018,9.525306,8.267109,7.0107265,5.75253,4.494334,3.2379513,2.909805,2.5816586,2.2553256,1.9271792,1.6008459,1.3941683,1.1893034,0.98443866,0.7795739,0.5747091,0.71430725,0.8557183,0.99531645,1.1349145,1.2745126,1.403233,1.5301404,1.6570477,1.7857682,1.9126755,2.1030366,2.2915847,2.4819458,2.6723068,2.8626678,2.7919624,2.72307,2.6523643,2.5816586,2.5127661,4.2042603,5.8975673,7.590874,9.282369,10.975676,11.873092,12.770509,13.667925,14.565341,15.462758,13.793019,12.123281,10.451729,8.781991,7.112252,6.209397,5.3083544,4.405499,3.5026438,2.5997884,2.3532255,2.1048496,1.8582866,1.6099107,1.3633479,1.4666867,1.5718386,1.6769904,1.7821422,1.887294,3.7401419,5.5929894,7.4458375,9.296872,11.14972,10.049252,8.950596,7.850128,6.7496595,5.6491914,5.6473784,5.6455655,5.6419396,5.6401267,5.638314,7.0433598,8.448405,9.851639,11.256684,12.661731,11.782444,10.903157,10.022058,9.142771,8.26167,9.547061,10.832452,12.117842,13.403233,14.68681,15.455506,16.22239,16.989273,17.757969,18.52485,18.367125,18.209396,18.051668,17.895754,17.738026,16.487082,15.23795,13.987006,12.737875,11.486931,10.312131,9.137331,7.9625316,6.787732,5.612932,4.666566,3.7220123,2.7774587,1.8329052,0.8883517,0.823085,0.75781834,0.69255173,0.62728506,0.5620184,0.5855869,0.6073425,0.629098,0.6526665,0.6744221,0.65991837,0.64541465,0.629098,0.61459434,0.6000906,6.688019,5.7380266,4.788034,3.8380418,2.8880494,1.938057,2.5870976,3.2379513,3.8869917,4.537845,5.186886,5.3246713,5.462456,5.600241,5.7380266,5.8758116,5.5367875,5.199577,4.8623657,4.5251546,4.1879435,3.4754493,2.762955,2.0504606,1.3379664,0.62547207,1.1131591,1.6008459,2.08672,2.5744069,3.0620937,2.525457,1.987007,1.4503701,0.9119202,0.37528324,0.387974,0.40066472,0.41335547,0.42423326,0.43692398,0.52575916,0.61278135,0.69980353,0.7868258,0.87566096,0.85027945,0.824898,0.7995165,0.774135,0.7505665,0.66173136,0.5747091,0.48768693,0.40066472,0.31182957,0.25018883,0.18673515,0.12509441,0.06164073,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06164073,0.12509441,0.18673515,0.25018883,0.31182957,0.25018883,0.18673515,0.12509441,0.06164073,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.25018883,0.37528324,0.50037766,0.62547207,0.7505665,5.0617914,9.374829,13.687867,18.000906,22.31213,20.024172,17.738026,15.4500675,13.162108,10.874149,8.762048,6.6499467,4.537845,2.4257438,0.31182957,0.25018883,0.18673515,0.12509441,0.06164073,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.25018883,0.43692398,0.62547207,0.8122072,1.0007553,0.7995165,0.6000906,0.40066472,0.19942589,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.0870222,0.11240368,0.13778515,0.16316663,0.18673515,0.2991388,0.41335547,0.52575916,0.63816285,0.7505665,1.4630609,2.175555,2.8880494,3.6005437,4.313038,3.5243993,2.7375734,1.9507477,1.162109,0.37528324,0.50037766,0.62547207,0.7505665,0.87566096,1.0007553,0.824898,0.6508536,0.4749962,0.2991388,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.62547207,1.2491312,1.8746033,2.5000753,3.1255474,3.1382382,3.149116,3.1618068,3.1744974,3.1871881,2.5508385,1.9126755,1.2745126,0.63816285,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.15047589,0.17585737,0.19942589,0.22480737,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.15047589,0.2991388,0.44961473,0.6000906,0.7505665,0.6744221,0.6000906,0.52575916,0.44961473,0.37528324,0.41335547,0.44961473,0.48768693,0.52575916,0.5620184,0.5873999,0.61278135,0.63816285,0.66173136,0.6871128,0.5620184,0.43692398,0.31182957,0.18673515,0.06164073,0.0870222,0.11240368,0.13778515,0.16316663,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0870222,0.17585737,0.26287958,0.34990177,0.43692398,0.42423326,0.41335547,0.40066472,0.387974,0.37528324,0.2991388,0.22480737,0.15047589,0.07433146,0.0,0.15047589,0.2991388,0.44961473,0.6000906,0.7505665,1.3506571,1.9507477,2.5508385,3.149116,3.7492065,3.100166,2.4493124,1.8002719,1.1494182,0.50037766,0.40066472,0.2991388,0.19942589,0.099712946,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.1258497,2.2498865,3.3757362,4.499773,5.6256227,5.750717,5.8758116,6.000906,6.1241875,6.249282,5.661882,5.0744824,4.4870825,3.8996825,3.3122826,3.4754493,3.636803,3.7999697,3.9631362,4.12449,4.7118897,5.2992897,5.8866897,6.4759026,7.063302,5.7380266,4.4127507,3.0874753,1.7621996,0.43692398,0.34990177,0.26287958,0.17585737,0.0870222,0.0,0.0870222,0.17585737,0.26287958,0.34990177,0.43692398,0.6871128,0.93730164,1.1874905,1.4376793,1.6878681,1.4757515,1.261822,1.0497054,0.8375887,0.62547207,2.0123885,3.3993049,4.788034,6.1749506,7.5618668,8.161958,8.762048,9.362139,9.96223,10.56232,10.774437,10.988366,11.200482,11.4126,11.624716,9.875207,8.125698,6.3743763,4.6248674,2.8753586,2.4620032,2.0504606,1.6371052,1.2255627,0.8122072,0.66173136,0.51306844,0.36259252,0.21211663,0.06164073,0.11240368,0.16316663,0.21211663,0.26287958,0.31182957,0.2755703,0.2374981,0.19942589,0.16316663,0.12509441,0.18673515,0.25018883,0.31182957,0.37528324,0.43692398,0.43692398,0.43692398,0.43692398,0.43692398,0.43692398,2.4130533,4.3873696,6.3616858,8.337815,10.312131,11.6881695,13.062395,14.438434,15.812659,17.186886,15.199879,13.212872,11.224051,9.237044,7.250037,6.399758,5.5494785,4.699199,3.8507326,3.000453,2.561716,2.124792,1.6878681,1.2491312,0.8122072,0.8375887,0.8629702,0.8883517,0.9119202,0.93730164,3.1871881,5.4370747,7.686961,9.936848,12.186734,10.774437,9.362139,7.949841,6.5375433,5.125245,4.9620786,4.800725,4.6375585,4.4743915,4.313038,6.0752378,7.837437,9.599637,11.361836,13.125849,11.862214,10.600392,9.336758,8.074935,6.813113,8.412147,10.012992,11.612025,13.212872,14.811904,15.687565,16.563227,17.437075,18.312735,19.188396,19.288109,19.387821,19.487535,19.587248,19.68696,18.550234,17.411694,16.274965,15.138238,13.999697,12.60009,11.200482,9.799063,8.399456,6.9998484,5.812358,4.6248674,3.437377,2.2498865,1.062396,0.9880646,0.9119202,0.8375887,0.76325727,0.6871128,0.6871128,0.6871128,0.6871128,0.6871128,0.6871128,0.61278135,0.53663695,0.46230546,0.387974,0.31182957,7.3370595,6.68258,6.0281005,5.371808,4.7173285,4.062849,4.2405195,4.41819,4.59586,4.7717175,4.949388,4.994712,5.040036,5.08536,5.130684,5.1741953,4.9203806,4.664753,4.409125,4.15531,3.8996825,3.245203,2.5907235,1.9344311,1.2799516,0.62547207,1.0098201,1.3941683,1.7803292,2.1646774,2.5508385,2.137483,1.7241274,1.3125849,0.89922947,0.48768693,0.58921283,0.69255173,0.79589057,0.8974165,1.0007553,0.9554313,0.9101072,0.86478317,0.8194591,0.774135,0.7433147,0.7106813,0.678048,0.64541465,0.61278135,0.5493277,0.48768693,0.42423326,0.36259252,0.2991388,0.24474995,0.19036107,0.13415924,0.07977036,0.025381476,0.02175555,0.01994259,0.018129626,0.014503701,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.06707962,0.13415924,0.2030518,0.27013144,0.33721104,0.27919623,0.2229944,0.16497959,0.10696479,0.05076295,0.09064813,0.13053331,0.17041849,0.21030366,0.25018883,0.33721104,0.42423326,0.51306844,0.6000906,0.6871128,4.119051,7.552802,10.98474,14.416678,17.85043,16.019337,14.190058,12.360779,10.529687,8.700407,7.0107265,5.319232,3.6295512,1.93987,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.17585737,0.34990177,0.52575916,0.69980353,0.87566096,0.71430725,0.55476654,0.39522585,0.23568514,0.07433146,0.21936847,0.36440548,0.5094425,0.6544795,0.7995165,0.6653573,0.5293851,0.39522585,0.25925365,0.12509441,0.16679256,0.21030366,0.2520018,0.2955129,0.33721104,0.3100166,0.28282216,0.25562772,0.22662032,0.19942589,0.22480737,0.25018883,0.2755703,0.2991388,0.3245203,0.27013144,0.21574254,0.15954071,0.10515183,0.05076295,0.0870222,0.12509441,0.16316663,0.19942589,0.2374981,0.72337204,1.2074331,1.693307,2.1773682,2.663242,2.8227828,2.9823234,3.141864,3.303218,3.4627585,2.8318477,2.2027495,1.5718386,0.94274056,0.31182957,0.42060733,0.5275721,0.6345369,0.7433147,0.85027945,0.79589057,0.73968875,0.6852999,0.630911,0.5747091,0.4749962,0.37528324,0.2755703,0.17585737,0.07433146,0.06707962,0.059827764,0.052575916,0.045324065,0.038072214,0.059827764,0.08339628,0.10515183,0.12690738,0.15047589,0.15228885,0.15410182,0.15772775,0.15954071,0.16316663,0.14503701,0.12690738,0.11059072,0.092461094,0.07433146,0.09064813,0.10515183,0.11965553,0.13415924,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.0,0.0,0.0,0.0,0.0,0.50037766,1.0007553,1.49932,1.9996977,2.5000753,2.5091403,2.520018,2.5290828,2.5399606,2.5508385,2.039583,1.5301404,1.020698,0.5094425,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.13778515,0.17585737,0.21211663,0.25018883,0.28826106,0.23024625,0.17223145,0.11421664,0.058014803,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.065266654,0.13053331,0.19579996,0.25925365,0.3245203,0.52032024,0.71430725,0.9101072,1.1059072,1.2998942,1.1204109,0.93911463,0.75963134,0.58014804,0.40066472,0.4224203,0.44417584,0.46774435,0.4894999,0.51306844,0.5275721,0.5420758,0.55839247,0.5728962,0.5873999,0.50219065,0.4169814,0.33177215,0.24837588,0.16316663,0.17223145,0.18310922,0.19217403,0.2030518,0.21211663,0.19036107,0.16679256,0.14503701,0.12328146,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.2030518,0.40429065,0.6073425,0.8103943,1.0116332,0.88291276,0.7523795,0.62184614,0.49312583,0.36259252,0.291887,0.2229944,0.15228885,0.08339628,0.012690738,0.17041849,0.32814622,0.48587397,0.6417888,0.7995165,1.35247,1.9054236,2.4583774,3.009518,3.5624714,2.9297476,2.2970235,1.6642996,1.0333886,0.40066472,0.3208944,0.23931105,0.15954071,0.07977036,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.968122,1.9344311,2.902553,3.870675,4.836984,5.1198063,5.4026284,5.6854506,5.9682727,6.249282,5.8758116,5.5005283,5.125245,4.749962,4.3746786,4.220577,4.064662,3.9105604,3.7546456,3.6005437,4.0157123,4.4290676,4.844236,5.2594047,5.674573,4.655688,3.63499,2.6142921,1.5954071,0.5747091,0.5058166,0.43511102,0.36440548,0.2955129,0.22480737,0.2955129,0.36440548,0.43511102,0.5058166,0.5747091,0.7306239,0.88472575,1.0406405,1.1947423,1.3506571,1.305333,1.260009,1.214685,1.1693609,1.1258497,2.1773682,3.2306993,4.2822175,5.335549,6.3870673,7.3008003,8.212721,9.12464,10.038374,10.950294,10.966611,10.98474,11.00287,11.019187,11.037316,9.412902,7.7866745,6.16226,4.537845,2.911618,2.518205,2.1229792,1.7277533,1.3325275,0.93730164,0.8194591,0.7016165,0.5855869,0.46774435,0.34990177,0.3770962,0.40429065,0.43329805,0.4604925,0.48768693,0.43329805,0.3770962,0.32270733,0.26831847,0.21211663,0.24293698,0.27194437,0.30276474,0.33177215,0.36259252,0.45324063,0.5420758,0.6327239,0.72337204,0.8122072,2.6432993,4.4725785,6.301858,8.13295,9.96223,11.227677,12.493125,13.75676,15.022208,16.287657,14.777458,13.267261,11.757062,10.246864,8.736667,8.392203,8.047741,7.703278,7.3570023,7.0125394,6.644508,6.2782893,5.910258,5.542227,5.1741953,4.4272547,3.680314,2.9333735,2.18462,1.4376793,3.1618068,4.8877473,6.6118746,8.337815,10.061942,9.300498,8.537241,7.7757964,7.0125394,6.249282,5.9718986,5.6945157,5.4171324,5.139749,4.8623657,6.58468,8.306994,10.029309,11.751623,13.475751,12.23931,11.004683,9.770056,8.535428,7.3008003,8.934279,10.5695715,12.2048645,13.840157,15.475449,16.189756,16.905876,17.620184,18.33449,19.050611,19.066927,19.085056,19.103188,19.119503,19.137632,18.116936,17.09805,16.077353,15.058467,14.037769,12.890164,11.7425585,10.594954,9.447348,8.299743,7.440398,6.5792413,5.719897,4.860553,3.9993954,3.4156215,2.8300345,2.2444477,1.6606737,1.0750868,1.0080072,0.93911463,0.872035,0.80495536,0.73787576,0.6526665,0.56745726,0.48224804,0.39703882,0.31182957,7.987913,7.6271334,7.268167,6.9073873,6.546608,6.187641,5.8921285,5.5966153,5.3029156,5.0074024,4.7118897,4.664753,4.6176157,4.5704784,4.5233417,4.4743915,4.3021603,4.1299286,3.9576974,3.785466,3.6132345,3.0149567,2.4166791,1.8202144,1.2219368,0.62547207,0.90829426,1.1893034,1.4721256,1.7549478,2.03777,1.7495089,1.4630609,1.1747998,0.8883517,0.6000906,0.79226464,0.98443866,1.1766127,1.3705997,1.5627737,1.3851035,1.2074331,1.0297627,0.8520924,0.6744221,0.6345369,0.5946517,0.55476654,0.5148814,0.4749962,0.43692398,0.40066472,0.36259252,0.3245203,0.28826106,0.23931105,0.19217403,0.14503701,0.09789998,0.05076295,0.045324065,0.03988518,0.034446288,0.030820364,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.072518505,0.14503701,0.21755551,0.29007402,0.36259252,0.3100166,0.2574407,0.20486477,0.15228885,0.099712946,0.15410182,0.21030366,0.26469254,0.3208944,0.37528324,0.42423326,0.4749962,0.52575916,0.5747091,0.62547207,3.1781235,5.730775,8.283426,10.834265,13.386916,12.0145035,10.642091,9.269678,7.897265,6.5248523,5.2575917,3.9903307,2.72307,1.455809,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.34990177,0.69980353,1.0497054,1.3996071,1.7495089,1.4177368,1.0841516,0.7523795,0.42060733,0.0870222,0.19036107,0.291887,0.39522585,0.49675176,0.6000906,0.5293851,0.4604925,0.38978696,0.3208944,0.25018883,0.33539808,0.42060733,0.5058166,0.58921283,0.6744221,0.6200332,0.5656443,0.5094425,0.4550536,0.40066472,0.44961473,0.50037766,0.5493277,0.6000906,0.6508536,0.5275721,0.40429065,0.28282216,0.15954071,0.038072214,0.0870222,0.13778515,0.18673515,0.2374981,0.28826106,1.1457924,2.0033236,2.8608549,3.7183862,4.5759177,4.1825047,3.7909048,3.397492,3.005892,2.612479,2.1392958,1.6679256,1.1947423,0.72337204,0.25018883,0.34083697,0.42967212,0.52032024,0.6091554,0.69980353,0.7650702,0.83033687,0.89560354,0.96087015,1.0243238,0.85027945,0.6744221,0.50037766,0.3245203,0.15047589,0.13415924,0.11965553,0.10515183,0.09064813,0.07433146,0.11965553,0.16497959,0.21030366,0.25562772,0.2991388,0.3045777,0.3100166,0.3154555,0.3208944,0.3245203,0.29007402,0.25562772,0.21936847,0.18492219,0.15047589,0.1794833,0.21030366,0.23931105,0.27013144,0.2991388,0.23931105,0.1794833,0.11965553,0.059827764,0.0,0.0,0.0,0.0,0.0,0.0,0.37528324,0.7505665,1.1258497,1.49932,1.8746033,1.8818551,1.889107,1.8981718,1.9054236,1.9126755,1.5301404,1.1476053,0.7650702,0.3825351,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.12509441,0.17585737,0.22480737,0.2755703,0.3245203,0.25925365,0.19579996,0.13053331,0.065266654,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13053331,0.25925365,0.38978696,0.52032024,0.6508536,0.8901646,1.1294757,1.3705997,1.6099107,1.8492218,1.5645868,1.2799516,0.99531645,0.7106813,0.42423326,0.43329805,0.4405499,0.44780177,0.4550536,0.46230546,0.46774435,0.47318324,0.47680917,0.48224804,0.48768693,0.44236287,0.39703882,0.35171473,0.30820364,0.26287958,0.2574407,0.2520018,0.24837588,0.24293698,0.2374981,0.23024625,0.2229944,0.21574254,0.20667773,0.19942589,0.15954071,0.11965553,0.07977036,0.03988518,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.31726846,0.6345369,0.95180535,1.2708868,1.5881553,1.3397794,1.0932164,0.8448406,0.5982776,0.34990177,0.28463513,0.21936847,0.15410182,0.09064813,0.025381476,0.19036107,0.35534066,0.52032024,0.6852999,0.85027945,1.3542831,1.8600996,2.3659163,2.8699198,3.3757362,2.759329,2.1447346,1.5301404,0.9155461,0.2991388,0.23931105,0.1794833,0.11965553,0.059827764,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.8103943,1.6207886,2.42937,3.2397642,4.0501585,4.4907084,4.9294453,5.369995,5.810545,6.249282,6.0879283,5.924762,5.7615952,5.600241,5.4370747,4.9657044,4.4925213,4.019338,3.5479677,3.0747845,3.3177216,3.5606585,3.8017826,4.0447197,4.2876563,3.5733492,2.857229,2.1429217,1.4268016,0.7124943,0.65991837,0.6073425,0.55476654,0.50219065,0.44961473,0.50219065,0.55476654,0.6073425,0.65991837,0.7124943,0.77232206,0.8321498,0.8919776,0.95180535,1.0116332,1.1349145,1.258196,1.3796645,1.502946,1.6244144,2.3423476,3.0602808,3.778214,4.494334,5.2122674,6.43783,7.66158,8.887142,10.112705,11.338268,11.160598,10.982927,10.805257,10.627586,10.449916,8.950596,7.4494634,5.9501433,4.4508233,2.94969,2.572594,2.1954978,1.8165885,1.4394923,1.062396,0.97718686,0.8919776,0.80676836,0.72337204,0.63816285,0.6417888,0.64722764,0.6526665,0.65810543,0.66173136,0.58921283,0.5166943,0.44417584,0.37165734,0.2991388,0.29732585,0.2955129,0.291887,0.29007402,0.28826106,0.46774435,0.64722764,0.82671094,1.0080072,1.1874905,2.8717327,4.557788,6.24203,7.9280853,9.612328,10.767185,11.922042,13.0769,14.231756,15.386614,14.355038,13.321649,12.290073,11.256684,10.225109,10.384649,10.54419,10.705544,10.865085,11.024626,10.7273,10.429974,10.1326475,9.835322,9.537996,8.01692,6.497658,4.976582,3.4573197,1.938057,3.1382382,4.3366065,5.5367875,6.736969,7.93715,7.8247466,7.7123427,7.5999393,7.4875355,7.3751316,6.981719,6.590119,6.1967063,5.805106,5.411693,7.0959353,8.778365,10.460794,12.143224,13.825653,12.618219,11.408974,10.203354,8.99592,7.7866745,9.458226,11.127964,12.797703,14.467442,16.13718,16.691946,17.246714,17.803293,18.358059,18.912827,18.847559,18.782291,18.717026,18.651758,18.588305,17.68545,16.782595,15.879739,14.976884,14.075842,13.180238,12.284635,11.390844,10.49524,9.599637,9.066626,8.535428,8.002417,7.4694057,6.9382076,5.8431783,4.748149,3.6531196,2.5580902,1.4630609,1.3270886,1.1929294,1.0569572,0.922798,0.7868258,0.69255173,0.5982776,0.50219065,0.40791658,0.31182957,8.636953,8.571687,8.508233,8.442966,8.3777,8.312433,7.5455503,6.776854,6.009971,5.243088,4.4743915,4.3347936,4.195195,4.0555973,3.9141862,3.774588,3.6857529,3.5951047,3.5044568,3.4156215,3.3249733,2.7847104,2.2444477,1.7041848,1.1657349,0.62547207,0.80495536,0.98443866,1.1657349,1.3452182,1.5247015,1.3633479,1.2001812,1.0370146,0.87566096,0.7124943,0.99531645,1.2781386,1.5591478,1.84197,2.124792,1.8147756,1.504759,1.1947423,0.88472575,0.5747091,0.5275721,0.48043507,0.43329805,0.38434806,0.33721104,0.3245203,0.31182957,0.2991388,0.28826106,0.2755703,0.23568514,0.19579996,0.15410182,0.11421664,0.07433146,0.06707962,0.059827764,0.052575916,0.045324065,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.07795739,0.15410182,0.23205921,0.3100166,0.387974,0.34083697,0.291887,0.24474995,0.19761293,0.15047589,0.21936847,0.29007402,0.36077955,0.42967212,0.50037766,0.51306844,0.52575916,0.53663695,0.5493277,0.5620184,2.2353828,3.9069343,5.580299,7.25185,8.925215,8.009668,7.0959353,6.1803894,5.2648435,4.349297,3.5044568,2.659616,1.8147756,0.969935,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.52575916,1.0497054,1.5754645,2.0994108,2.6251698,2.1193533,1.6153497,1.1095331,0.6055295,0.099712946,0.15954071,0.21936847,0.27919623,0.34083697,0.40066472,0.39522585,0.38978696,0.38434806,0.38072214,0.37528324,0.50219065,0.629098,0.75781834,0.88472575,1.0116332,0.9300498,0.8466535,0.7650702,0.68167394,0.6000906,0.6744221,0.7505665,0.824898,0.89922947,0.97537386,0.7850128,0.5946517,0.40429065,0.21574254,0.025381476,0.0870222,0.15047589,0.21211663,0.2755703,0.33721104,1.5682126,2.7974012,4.028403,5.2575917,6.48678,5.542227,4.597673,3.6531196,2.7067533,1.7621996,1.4467441,1.1331016,0.81764615,0.50219065,0.18673515,0.25925365,0.33177215,0.40429065,0.47680917,0.5493277,0.73424983,0.91917205,1.1059072,1.2908293,1.4757515,1.2255627,0.97537386,0.72518504,0.4749962,0.22480737,0.2030518,0.1794833,0.15772775,0.13415924,0.11240368,0.1794833,0.24837588,0.3154555,0.3825351,0.44961473,0.45686656,0.46411842,0.47318324,0.48043507,0.48768693,0.43511102,0.3825351,0.32995918,0.27738327,0.22480737,0.27013144,0.3154555,0.36077955,0.40429065,0.44961473,0.36077955,0.27013144,0.1794833,0.09064813,0.0,0.0,0.0,0.0,0.0,0.0,0.25018883,0.50037766,0.7505665,1.0007553,1.2491312,1.2545701,1.260009,1.2654479,1.2708868,1.2745126,1.020698,0.7650702,0.5094425,0.25562772,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.11240368,0.17585737,0.2374981,0.2991388,0.36259252,0.29007402,0.21755551,0.14503701,0.072518505,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.19579996,0.38978696,0.5855869,0.7795739,0.97537386,1.260009,1.5446441,1.8292793,2.1157274,2.4003625,2.0105755,1.6207886,1.2291887,0.83940166,0.44961473,0.44236287,0.43511102,0.42785916,0.42060733,0.41335547,0.40791658,0.40247768,0.39703882,0.39159992,0.387974,0.3825351,0.3770962,0.37165734,0.3680314,0.36259252,0.34264994,0.32270733,0.30276474,0.28282216,0.26287958,0.27013144,0.27738327,0.28463513,0.291887,0.2991388,0.23931105,0.1794833,0.11965553,0.059827764,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.43329805,0.86478317,1.2980812,1.7295663,2.1628644,1.7966459,1.4322405,1.067835,0.7016165,0.33721104,0.27738327,0.21755551,0.15772775,0.09789998,0.038072214,0.21030366,0.3825351,0.55476654,0.726998,0.89922947,1.357909,1.8147756,2.2716422,2.7303216,3.1871881,2.5907235,1.9924458,1.3941683,0.79770356,0.19942589,0.15954071,0.11965553,0.07977036,0.03988518,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.6526665,1.305333,1.9579996,2.610666,3.2633326,3.8597972,4.458075,5.0545397,5.6528172,6.249282,6.300045,6.350808,6.399758,6.450521,6.4994707,5.710832,4.9203806,4.1299286,3.339477,2.5508385,2.619731,2.6904364,2.759329,2.8300345,2.9007401,2.4891977,2.079468,1.6697385,1.260009,0.85027945,0.81583315,0.7795739,0.7451276,0.7106813,0.6744221,0.7106813,0.7451276,0.7795739,0.81583315,0.85027945,0.81583315,0.7795739,0.7451276,0.7106813,0.6744221,0.9644961,1.2545701,1.5446441,1.8347181,2.124792,2.5073273,2.8898623,3.2723975,3.6549325,4.0374675,5.57486,7.112252,8.649645,10.1870365,11.724429,11.352772,10.979301,10.607644,10.234174,9.862516,8.488291,7.112252,5.7380266,4.361988,2.9877625,2.6269827,2.268016,1.9072367,1.54827,1.1874905,1.1349145,1.0823387,1.0297627,0.97718686,0.9246109,0.90829426,0.8901646,0.872035,0.8557183,0.8375887,0.7469406,0.65810543,0.56745726,0.47680917,0.387974,0.35171473,0.31726846,0.28282216,0.24837588,0.21211663,0.48224804,0.7523795,1.0225109,1.2926424,1.5627737,3.101979,4.6429973,6.1822023,7.723221,9.262425,10.306692,11.352772,12.397038,13.443117,14.487384,13.932617,13.377851,12.823084,12.268318,11.711739,12.377095,13.042453,13.70781,14.373167,15.036712,14.810091,14.581658,14.355038,14.126604,13.899984,11.606586,9.3150015,7.021604,4.7300196,2.4366217,3.1128569,3.787279,4.461701,5.137936,5.812358,6.350808,6.887445,7.4258947,7.9625316,8.499168,7.993352,7.4857225,6.978093,6.4704633,5.962834,7.605378,9.247922,10.890467,12.5330105,14.175554,12.995316,11.815077,10.634838,9.4546,8.274362,9.980359,11.684544,13.390542,15.094727,16.800724,17.194138,17.589363,17.984589,18.379814,18.77504,18.628191,18.479528,18.332678,18.185827,18.037165,17.252151,16.467138,15.682126,14.897114,14.112101,13.470312,12.826711,12.184921,11.543133,10.899531,10.694666,10.489801,10.284937,10.080072,9.875207,8.270736,6.6644506,5.0599785,3.4555066,1.8492218,1.647983,1.4449311,1.2418793,1.0406405,0.8375887,0.7324369,0.62728506,0.52213323,0.4169814,0.31182957,9.287807,9.518054,9.7483,9.976733,10.20698,10.437225,9.197159,7.957093,6.717026,5.47696,4.2368937,4.004834,3.7727752,3.540716,3.3068438,3.0747845,3.0675328,3.0602808,3.053029,3.045777,3.0367124,2.5544643,2.0722163,1.5899682,1.1077201,0.62547207,0.7016165,0.7795739,0.8575313,0.9354887,1.0116332,0.97537386,0.93730164,0.89922947,0.8629702,0.824898,1.1983683,1.5700256,1.9416829,2.3151531,2.6868105,2.2444477,1.8020848,1.3597219,0.91735905,0.4749962,0.42060733,0.36440548,0.3100166,0.25562772,0.19942589,0.21211663,0.22480737,0.2374981,0.25018883,0.26287958,0.23024625,0.19761293,0.16497959,0.13234627,0.099712946,0.09064813,0.07977036,0.07070554,0.059827764,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.08339628,0.16497959,0.24837588,0.32995918,0.41335547,0.36984438,0.32814622,0.28463513,0.24293698,0.19942589,0.28463513,0.36984438,0.4550536,0.5402629,0.62547207,0.6000906,0.5747091,0.5493277,0.52575916,0.50037766,1.2926424,2.084907,2.8771715,3.6694362,4.461701,4.004834,3.5479677,3.0892882,2.6324217,2.175555,1.7531348,1.3307146,0.90829426,0.48587397,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.69980353,1.3996071,2.0994108,2.7992141,3.5008307,2.8227828,2.1447346,1.4666867,0.7904517,0.11240368,0.13053331,0.14684997,0.16497959,0.18310922,0.19942589,0.25925365,0.3208944,0.38072214,0.4405499,0.50037766,0.67079616,0.83940166,1.0098201,1.1802386,1.3506571,1.2400664,1.1294757,1.020698,0.9101072,0.7995165,0.89922947,1.0007553,1.1004683,1.2001812,1.2998942,1.0424535,0.7850128,0.5275721,0.27013144,0.012690738,0.0870222,0.16316663,0.2374981,0.31182957,0.387974,1.9906329,3.5932918,5.195951,6.796797,8.399456,6.9019485,5.4044414,3.9069343,2.4094272,0.9119202,0.7541924,0.5982776,0.4405499,0.28282216,0.12509441,0.1794833,0.23568514,0.29007402,0.3444629,0.40066472,0.70524246,1.0098201,1.3143979,1.6207886,1.9253663,1.6008459,1.2745126,0.9499924,0.62547207,0.2991388,0.27013144,0.23931105,0.21030366,0.1794833,0.15047589,0.23931105,0.32995918,0.42060733,0.5094425,0.6000906,0.6091554,0.6200332,0.629098,0.6399758,0.6508536,0.58014804,0.5094425,0.4405499,0.36984438,0.2991388,0.36077955,0.42060733,0.48043507,0.5402629,0.6000906,0.48043507,0.36077955,0.23931105,0.11965553,0.0,0.0,0.0,0.0,0.0,0.0,0.12509441,0.25018883,0.37528324,0.50037766,0.62547207,0.62728506,0.629098,0.6327239,0.6345369,0.63816285,0.5094425,0.3825351,0.25562772,0.12690738,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.099712946,0.17585737,0.25018883,0.3245203,0.40066472,0.3208944,0.23931105,0.15954071,0.07977036,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.25925365,0.52032024,0.7795739,1.0406405,1.2998942,1.6298534,1.9598125,2.2897718,2.619731,2.94969,2.4547513,1.9598125,1.4648738,0.969935,0.4749962,0.45324063,0.42967212,0.40791658,0.38434806,0.36259252,0.3480888,0.33177215,0.31726846,0.30276474,0.28826106,0.32270733,0.35715362,0.39159992,0.42785916,0.46230546,0.42785916,0.39159992,0.35715362,0.32270733,0.28826106,0.3100166,0.33177215,0.35534066,0.3770962,0.40066472,0.3208944,0.23931105,0.15954071,0.07977036,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.5475147,1.0950294,1.6425442,2.1900587,2.7375734,2.2553256,1.7730774,1.2908293,0.80676836,0.3245203,0.27013144,0.21574254,0.15954071,0.10515183,0.05076295,0.23024625,0.40972954,0.58921283,0.7705091,0.9499924,1.3597219,1.7694515,2.179181,2.5907235,3.000453,2.420305,1.840157,1.260009,0.67986095,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.4949388,0.9898776,1.4848163,1.9797552,2.474694,3.2306993,3.9848917,4.740897,5.4950895,6.249282,6.5121617,6.775041,7.037921,7.3008003,7.5618668,6.454147,5.3482394,4.2405195,3.1327994,2.0250793,1.9217403,1.8202144,1.7168756,1.6153497,1.5120108,1.4068589,1.3017071,1.1983683,1.0932164,0.9880646,0.969935,0.95180535,0.9354887,0.91735905,0.89922947,0.91735905,0.9354887,0.95180535,0.969935,0.9880646,0.8575313,0.726998,0.5982776,0.46774435,0.33721104,0.79589057,1.2527572,1.7096237,2.1683033,2.6251698,2.6723068,2.7194438,2.7683938,2.8155308,2.8626678,4.7118897,6.5629244,8.412147,10.263181,12.112403,11.544946,10.9774885,10.410031,9.842574,9.275117,8.024173,6.775041,5.524097,4.274966,3.0258346,2.6831846,2.3405347,1.9978848,1.6552348,1.3125849,1.2926424,1.2726997,1.2527572,1.2328146,1.2128719,1.1729867,1.1331016,1.0932164,1.0533313,1.0116332,0.90466833,0.79770356,0.69073874,0.581961,0.4749962,0.40791658,0.34083697,0.27194437,0.20486477,0.13778515,0.49675176,0.8575313,1.2183108,1.5772774,1.938057,3.3322253,4.7282066,6.1223745,7.516543,8.912524,9.848013,10.781689,11.717177,12.652666,13.588155,13.510198,13.43224,13.354282,13.278138,13.200181,14.369541,15.540715,16.710075,17.879436,19.050611,18.892883,18.735155,18.577427,18.4197,18.261972,15.198066,12.132345,9.066626,6.002719,2.9369993,3.0874753,3.2379513,3.386614,3.53709,3.6875658,4.8750563,6.0625467,7.250037,8.437528,9.625018,9.003172,8.379513,7.757667,7.135821,6.5121617,8.1148205,9.71748,11.320138,12.922797,14.525456,13.372412,12.219368,11.068136,9.915092,8.762048,10.502492,12.242936,13.98338,15.722012,17.462456,17.698141,17.932013,18.167698,18.403383,18.637255,18.40701,18.176764,17.94833,17.718082,17.487837,16.820667,16.151684,15.484513,14.817343,14.150173,13.760386,13.370599,12.980812,12.589212,12.199425,12.322706,12.444175,12.567456,12.690738,12.812206,10.698292,8.582565,6.4668374,4.3529234,2.2371957,1.9670644,1.696933,1.4268016,1.1566701,0.8883517,0.77232206,0.65810543,0.5420758,0.42785916,0.31182957,9.936848,10.462607,10.988366,11.512312,12.038072,12.562017,10.850581,9.137331,7.424082,5.712645,3.9993954,3.6748753,3.350355,3.0258346,2.6995013,2.374981,2.4493124,2.525457,2.5997884,2.6741197,2.7502642,2.324218,1.8999848,1.4757515,1.0497054,0.62547207,0.6000906,0.5747091,0.5493277,0.52575916,0.50037766,0.5873999,0.6744221,0.76325727,0.85027945,0.93730164,1.3996071,1.8619126,2.324218,2.7883365,3.2506418,2.6741197,2.0994108,1.5247015,0.9499924,0.37528324,0.31182957,0.25018883,0.18673515,0.12509441,0.06164073,0.099712946,0.13778515,0.17585737,0.21211663,0.25018883,0.22480737,0.19942589,0.17585737,0.15047589,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0870222,0.17585737,0.26287958,0.34990177,0.43692398,0.40066472,0.36259252,0.3245203,0.28826106,0.25018883,0.34990177,0.44961473,0.5493277,0.6508536,0.7505665,0.6871128,0.62547207,0.5620184,0.50037766,0.43692398,0.34990177,0.26287958,0.17585737,0.0870222,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.87566096,1.7495089,2.6251698,3.5008307,4.3746786,3.5243993,2.6741197,1.8256533,0.97537386,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.12509441,0.25018883,0.37528324,0.50037766,0.62547207,0.8375887,1.0497054,1.261822,1.4757515,1.6878681,1.550083,1.4122978,1.2745126,1.1367276,1.0007553,1.1258497,1.2491312,1.3742256,1.49932,1.6244144,1.2998942,0.97537386,0.6508536,0.3245203,0.0,0.0870222,0.17585737,0.26287958,0.34990177,0.43692398,2.4130533,4.3873696,6.3616858,8.337815,10.312131,8.26167,6.2130227,4.162562,2.1121013,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.099712946,0.13778515,0.17585737,0.21211663,0.25018883,0.6744221,1.1004683,1.5247015,1.9507477,2.374981,1.9743162,1.5754645,1.1747998,0.774135,0.37528324,0.33721104,0.2991388,0.26287958,0.22480737,0.18673515,0.2991388,0.41335547,0.52575916,0.63816285,0.7505665,0.76325727,0.774135,0.7868258,0.7995165,0.8122072,0.72518504,0.63816285,0.5493277,0.46230546,0.37528324,0.44961473,0.52575916,0.6000906,0.6744221,0.7505665,0.6000906,0.44961473,0.2991388,0.15047589,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0870222,0.17585737,0.26287958,0.34990177,0.43692398,0.34990177,0.26287958,0.17585737,0.0870222,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.3245203,0.6508536,0.97537386,1.2998942,1.6244144,1.9996977,2.374981,2.7502642,3.1255474,3.5008307,2.9007401,2.3006494,1.7005589,1.1004683,0.50037766,0.46230546,0.42423326,0.387974,0.34990177,0.31182957,0.28826106,0.26287958,0.2374981,0.21211663,0.18673515,0.26287958,0.33721104,0.41335547,0.48768693,0.5620184,0.51306844,0.46230546,0.41335547,0.36259252,0.31182957,0.34990177,0.387974,0.42423326,0.46230546,0.50037766,0.40066472,0.2991388,0.19942589,0.099712946,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.66173136,1.3252757,1.987007,2.6505513,3.3122826,2.712192,2.1121013,1.5120108,0.9119202,0.31182957,0.26287958,0.21211663,0.16316663,0.11240368,0.06164073,0.25018883,0.43692398,0.62547207,0.8122072,1.0007553,1.3633479,1.7241274,2.08672,2.4493124,2.811905,2.2498865,1.6878681,1.1258497,0.5620184,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.33721104,0.6744221,1.0116332,1.3506571,1.6878681,2.5997884,3.5117085,4.4254417,5.337362,6.249282,6.7242785,7.1992745,7.6742706,8.149267,8.624263,7.1992745,5.774286,4.349297,2.9243085,1.49932,1.2255627,0.9499924,0.6744221,0.40066472,0.12509441,0.3245203,0.52575916,0.72518504,0.9246109,1.1258497,1.1258497,1.1258497,1.1258497,1.1258497,1.1258497,1.1258497,1.1258497,1.1258497,1.1258497,1.1258497,0.89922947,0.6744221,0.44961473,0.22480737,0.0,0.62547207,1.2491312,1.8746033,2.5000753,3.1255474,2.8372865,2.5508385,2.2625773,1.9743162,1.6878681,3.8507326,6.011784,8.174648,10.337513,12.500377,11.73712,10.975676,10.212419,9.449161,8.6877165,7.5618668,6.43783,5.3119802,4.1879435,3.0620937,2.7375734,2.4130533,2.08672,1.7621996,1.4376793,1.4503701,1.4630609,1.4757515,1.4866294,1.49932,1.4376793,1.3742256,1.3125849,1.2491312,1.1874905,1.062396,0.93730164,0.8122072,0.6871128,0.5620184,0.46230546,0.36259252,0.26287958,0.16316663,0.06164073,0.51306844,0.96268314,1.4122978,1.8619126,2.3133402,3.5624714,4.8116026,6.0625467,7.311678,8.562622,9.38752,10.212419,11.037316,11.862214,12.687112,13.087777,13.486629,13.887294,14.287958,14.68681,16.361988,18.037165,19.712341,21.38752,23.062696,22.975676,22.886839,22.799818,22.712795,22.625772,18.787731,14.94969,11.111648,7.2754188,3.437377,3.0620937,2.6868105,2.3133402,1.938057,1.5627737,3.3993049,5.237649,7.07418,8.912524,10.750868,10.012992,9.275117,8.537241,7.799365,7.063302,8.624263,10.1870365,11.74981,13.312584,14.875358,13.749508,12.625471,11.499621,10.375585,9.249735,11.024626,12.799516,14.574407,16.349297,18.124187,18.20033,18.274662,18.350807,18.425138,18.49947,18.187641,17.87581,17.562168,17.25034,16.936697,16.38737,15.838041,15.2869005,14.737573,14.188245,14.05046,13.912675,13.77489,13.637105,13.499319,13.9507475,14.400362,14.849977,15.299591,15.749206,13.124036,10.498866,7.8755093,5.2503395,2.6251698,2.2879589,1.9507477,1.6117238,1.2745126,0.93730164,0.8122072,0.6871128,0.5620184,0.43692398,0.31182957,9.438283,9.904215,10.371959,10.839704,11.307447,11.775192,10.672911,9.570629,8.4683485,7.364254,6.261973,5.9827766,5.7017674,5.422571,5.143375,4.8623657,4.7318325,4.603112,4.4725785,4.3420453,4.213325,3.7401419,3.2669585,2.7955883,2.322405,1.8492218,1.6298534,1.4104849,1.1893034,0.969935,0.7505665,0.774135,0.7995165,0.824898,0.85027945,0.87566096,1.2908293,1.7041848,2.1193533,2.5345216,2.94969,2.469255,1.9906329,1.5101979,1.0297627,0.5493277,0.533011,0.5148814,0.49675176,0.48043507,0.46230546,0.43692398,0.41335547,0.387974,0.36259252,0.33721104,0.291887,0.24837588,0.2030518,0.15772775,0.11240368,0.14503701,0.17767033,0.21030366,0.24293698,0.2755703,0.2991388,0.3245203,0.34990177,0.37528324,0.40066472,0.3245203,0.25018883,0.17585737,0.099712946,0.025381476,0.03988518,0.054388877,0.07070554,0.08520924,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.030820364,0.034446288,0.03988518,0.045324065,0.05076295,0.15410182,0.25925365,0.36440548,0.46955732,0.5747091,0.4604925,0.3444629,0.23024625,0.11421664,0.0,0.11421664,0.23024625,0.3444629,0.4604925,0.5747091,0.7995165,1.0243238,1.2491312,1.4757515,1.7005589,1.4902552,1.2799516,1.0696479,0.85934424,0.6508536,0.58921283,0.5293851,0.46955732,0.40972954,0.34990177,0.27919623,0.21030366,0.13959812,0.07070554,0.0,0.0,0.0,0.0,0.0,0.0,0.18492219,0.36984438,0.55476654,0.73968875,0.9246109,0.7451276,0.5656443,0.38434806,0.20486477,0.025381476,0.72337204,1.4195497,2.1175404,2.8155308,3.5117085,2.902553,2.2933977,1.6824293,1.0732739,0.46230546,0.43692398,0.41335547,0.387974,0.36259252,0.33721104,0.38434806,0.43329805,0.48043507,0.5275721,0.5747091,0.7324369,0.8901646,1.0478923,1.2056202,1.3633479,1.3470312,1.3325275,1.3180238,1.3017071,1.2872034,1.3125849,1.3379664,1.3633479,1.3869164,1.4122978,1.2019942,0.9916905,0.78319985,0.5728962,0.36259252,0.48224804,0.60190356,0.72337204,0.8430276,0.96268314,2.520018,4.077353,5.634688,7.192023,8.749357,7.0469856,5.3446136,3.6422417,1.93987,0.2374981,0.27013144,0.30276474,0.33539808,0.3680314,0.40066472,0.39522585,0.38978696,0.38434806,0.38072214,0.37528324,0.67986095,0.98443866,1.2908293,1.5954071,1.8999848,1.5881553,1.2745126,0.96268314,0.6508536,0.33721104,0.2991388,0.26287958,0.22480737,0.18673515,0.15047589,0.23931105,0.32995918,0.42060733,0.5094425,0.6000906,0.6091554,0.6200332,0.629098,0.6399758,0.6508536,0.59283876,0.53482395,0.47680917,0.42060733,0.36259252,0.40972954,0.45686656,0.5058166,0.5529536,0.6000906,0.48043507,0.36077955,0.23931105,0.11965553,0.0,0.027194439,0.054388877,0.08339628,0.11059072,0.13778515,0.22662032,0.31726846,0.40791658,0.49675176,0.5873999,0.52213323,0.45686656,0.3934129,0.32814622,0.26287958,0.21755551,0.17223145,0.12690738,0.08339628,0.038072214,0.11421664,0.19217403,0.27013144,0.3480888,0.42423326,0.5076295,0.58921283,0.6726091,0.7541924,0.8375887,0.8684091,0.8974165,0.92823684,0.9572442,0.9880646,0.97537386,0.96268314,0.9499924,0.93730164,0.9246109,0.7541924,0.5855869,0.41516843,0.24474995,0.07433146,0.09427405,0.11421664,0.13415924,0.15410182,0.17585737,0.15772775,0.13959812,0.12328146,0.10515183,0.0870222,0.19036107,0.291887,0.39522585,0.49675176,0.6000906,0.5855869,0.56927025,0.55476654,0.5402629,0.52575916,0.50219065,0.48043507,0.45686656,0.43511102,0.41335547,0.45686656,0.50219065,0.5475147,0.59283876,0.63816285,0.9826257,1.3270886,1.6733645,2.0178273,2.3622901,2.467442,2.572594,2.6777458,2.7828975,2.8880494,2.4021754,1.9181144,1.4322405,0.9481794,0.46230546,0.533011,0.60190356,0.6726091,0.7433147,0.8122072,0.73424983,0.65810543,0.58014804,0.50219065,0.42423326,0.4405499,0.4550536,0.46955732,0.48587397,0.50037766,0.4550536,0.40972954,0.36440548,0.3208944,0.2755703,0.31182957,0.34990177,0.387974,0.42423326,0.46230546,0.36984438,0.27738327,0.18492219,0.092461094,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.533011,1.064209,1.5972201,2.1302311,2.663242,2.1991236,1.7368182,1.2745126,0.8122072,0.34990177,0.29007402,0.23024625,0.17041849,0.11059072,0.05076295,0.21574254,0.38072214,0.54570174,0.7106813,0.87566096,1.2128719,1.550083,1.887294,2.2245052,2.561716,2.0504606,1.5373923,1.0243238,0.51306844,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.32995918,0.65991837,0.9898776,1.3198367,1.649796,2.373168,3.094727,3.8180993,4.539658,5.2630305,5.6854506,6.107871,6.530291,6.9527116,7.3751316,6.3852544,5.3953767,4.405499,3.4156215,2.4257438,1.9670644,1.5101979,1.0533313,0.5946517,0.13778515,0.3825351,0.62728506,0.872035,1.1167849,1.3633479,1.3017071,1.2418793,1.1820517,1.1222239,1.062396,1.0895905,1.1167849,1.1457924,1.1729867,1.2001812,0.96087015,0.7197462,0.48043507,0.23931105,0.0,0.5148814,1.0297627,1.5446441,2.0595255,2.5744069,2.4801328,2.3858588,2.2897718,2.1954978,2.0994108,4.0501585,5.999093,7.949841,9.900589,11.849524,11.095331,10.339326,9.585134,8.829127,8.074935,7.0342946,5.995467,4.954827,3.9141862,2.8753586,2.5290828,2.18462,1.840157,1.4956942,1.1494182,1.1602961,1.1693609,1.1802386,1.1893034,1.2001812,1.1494182,1.1004683,1.0497054,1.0007553,0.9499924,0.85027945,0.7505665,0.6508536,0.5493277,0.44961473,0.37165734,0.2955129,0.21755551,0.13959812,0.06164073,0.42060733,0.7777609,1.1349145,1.4920682,1.8492218,2.913431,3.975827,5.038223,6.1006193,7.1630154,7.8120556,8.46291,9.11195,9.762803,10.411844,11.122525,11.833207,12.542075,13.252756,13.961625,15.292339,16.623055,17.951956,19.282671,20.611572,20.491917,20.372261,20.252605,20.13295,20.013294,17.230396,14.447499,11.664601,8.883516,6.1006193,5.331923,4.5650396,3.7981565,3.0294604,2.2625773,3.5679104,4.8732433,6.1767635,7.4820967,8.78743,8.21816,7.647076,7.077806,6.506723,5.9374523,7.7776093,9.617766,11.457924,13.29808,15.138238,13.985193,12.8321495,11.679105,10.527874,9.374829,10.725487,12.07433,13.424988,14.775645,16.124489,16.294909,16.465326,16.635744,16.80435,16.97477,17.27572,17.57486,17.87581,18.17495,18.475903,17.629248,16.784407,15.939567,15.094727,14.249886,14.170115,14.090345,14.010575,13.930804,13.849221,13.852847,13.85466,13.858286,13.860099,13.861912,11.544946,9.22798,6.9092,4.592234,2.275268,1.9942589,1.7150626,1.4358664,1.1548572,0.87566096,0.7650702,0.6544795,0.54570174,0.43511102,0.3245203,8.937905,9.347635,9.757364,10.167094,10.576823,10.988366,10.49524,10.002114,9.510801,9.017676,8.52455,8.290678,8.054993,7.819308,7.5854354,7.3497505,7.0143523,6.680767,6.345369,6.009971,5.674573,5.1542525,4.6357455,4.115425,3.5951047,3.0747845,2.659616,2.2444477,1.8292793,1.4141108,1.0007553,0.96268314,0.9246109,0.8883517,0.85027945,0.8122072,1.1802386,1.54827,1.9144884,2.2825198,2.6505513,2.2643902,1.8800422,1.4956942,1.1095331,0.72518504,0.7523795,0.7795739,0.80676836,0.83577573,0.8629702,0.774135,0.6871128,0.6000906,0.51306844,0.42423326,0.36077955,0.2955129,0.23024625,0.16497959,0.099712946,0.17767033,0.25562772,0.33177215,0.40972954,0.48768693,0.5493277,0.61278135,0.6744221,0.73787576,0.7995165,0.6508536,0.50037766,0.34990177,0.19942589,0.05076295,0.07977036,0.11059072,0.13959812,0.17041849,0.19942589,0.15954071,0.11965553,0.07977036,0.03988518,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.047137026,0.045324065,0.04169814,0.03988518,0.038072214,0.25925365,0.48224804,0.70524246,0.92823684,1.1494182,0.91917205,0.69073874,0.4604925,0.23024625,0.0,0.14322405,0.28463513,0.42785916,0.56927025,0.7124943,1.2001812,1.6878681,2.175555,2.663242,3.149116,2.6306088,2.1102884,1.5899682,1.0696479,0.5493277,0.49312583,0.43511102,0.3770962,0.3208944,0.26287958,0.21030366,0.15772775,0.10515183,0.052575916,0.0,0.0,0.0,0.0,0.0,0.0,0.36984438,0.73968875,1.1095331,1.4793775,1.8492218,1.4902552,1.1294757,0.7705091,0.40972954,0.05076295,0.56927025,1.0895905,1.6099107,2.1302311,2.6505513,2.280707,1.9108626,1.5392052,1.1693609,0.7995165,0.774135,0.7505665,0.72518504,0.69980353,0.6744221,0.64541465,0.61459434,0.5855869,0.55476654,0.52575916,0.62728506,0.7306239,0.8321498,0.9354887,1.0370146,1.1457924,1.2527572,1.3597219,1.4666867,1.5754645,1.49932,1.4249886,1.3506571,1.2745126,1.2001812,1.1059072,1.0098201,0.9155461,0.8194591,0.72518504,0.8774739,1.0297627,1.1820517,1.3343405,1.4866294,2.6269827,3.7673361,4.9076896,6.0480433,7.1865835,5.8323007,4.478018,3.1219215,1.7676386,0.41335547,0.47680917,0.5420758,0.6073425,0.6726091,0.73787576,0.69073874,0.6417888,0.5946517,0.5475147,0.50037766,0.6852999,0.87022203,1.0551442,1.2400664,1.4249886,1.2001812,0.97537386,0.7505665,0.52575916,0.2991388,0.26287958,0.22480737,0.18673515,0.15047589,0.11240368,0.1794833,0.24837588,0.3154555,0.3825351,0.44961473,0.45686656,0.46411842,0.47318324,0.48043507,0.48768693,0.4604925,0.43329805,0.40429065,0.3770962,0.34990177,0.36984438,0.38978696,0.40972954,0.42967212,0.44961473,0.36077955,0.27013144,0.1794833,0.09064813,0.0,0.054388877,0.11059072,0.16497959,0.21936847,0.2755703,0.4550536,0.6345369,0.81583315,0.99531645,1.1747998,1.0442665,0.9155461,0.7850128,0.6544795,0.52575916,0.43511102,0.3444629,0.25562772,0.16497959,0.07433146,0.23024625,0.38434806,0.5402629,0.69436467,0.85027945,0.92823684,1.0043813,1.0823387,1.1602961,1.2382535,1.3851035,1.5319533,1.6806163,1.8274662,1.9743162,1.9507477,1.9253663,1.8999848,1.8746033,1.8492218,1.5101979,1.1693609,0.83033687,0.4894999,0.15047589,0.19036107,0.23024625,0.27013144,0.3100166,0.34990177,0.3154555,0.27919623,0.24474995,0.21030366,0.17585737,0.38072214,0.5855869,0.7904517,0.99531645,1.2001812,1.1693609,1.1403534,1.1095331,1.0805258,1.0497054,1.0043813,0.96087015,0.9155461,0.87022203,0.824898,0.9155461,1.0043813,1.0950294,1.1856775,1.2745126,1.6407311,2.0051367,2.3695421,2.7357605,3.100166,2.9351864,2.770207,2.6052272,2.4402475,2.275268,1.9054236,1.5355793,1.1657349,0.79589057,0.42423326,0.60190356,0.7795739,0.9572442,1.1349145,1.3125849,1.1820517,1.0533313,0.922798,0.79226464,0.66173136,0.61822027,0.5728962,0.5275721,0.48224804,0.43692398,0.39703882,0.35715362,0.31726846,0.27738327,0.2374981,0.2755703,0.31182957,0.34990177,0.387974,0.42423326,0.34083697,0.25562772,0.17041849,0.08520924,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.40247768,0.80495536,1.2074331,1.6099107,2.0123885,1.6878681,1.3633479,1.0370146,0.7124943,0.387974,0.31726846,0.24837588,0.17767033,0.10696479,0.038072214,0.1794833,0.32270733,0.46411842,0.6073425,0.7505665,1.062396,1.3742256,1.6878681,1.9996977,2.3133402,1.8492218,1.3869164,0.9246109,0.46230546,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.32270733,0.64541465,0.968122,1.2908293,1.6117238,2.1447346,2.6777458,3.2107568,3.7419548,4.274966,4.64481,5.0146546,5.384499,5.754343,6.1241875,5.569421,5.0146546,4.459888,3.9051213,3.350355,2.7103791,2.0704033,1.4304274,0.7904517,0.15047589,0.4405499,0.7306239,1.020698,1.310772,1.6008459,1.4793775,1.3597219,1.2400664,1.1204109,1.0007553,1.0551442,1.1095331,1.1657349,1.2201238,1.2745126,1.020698,0.7650702,0.5094425,0.25562772,0.0,0.40429065,0.8103943,1.214685,1.6207886,2.0250793,2.1229792,2.220879,2.3169663,2.4148662,2.5127661,4.249584,5.9882154,7.7250338,9.461852,11.200482,10.451729,9.704789,8.957849,8.209095,7.462154,6.506723,5.5531044,4.597673,3.6422417,2.6868105,2.322405,1.9579996,1.5917811,1.2273756,0.8629702,0.87022203,0.8774739,0.88472575,0.8919776,0.89922947,0.8629702,0.824898,0.7868258,0.7505665,0.7124943,0.63816285,0.5620184,0.48768693,0.41335547,0.33721104,0.28282216,0.22662032,0.17223145,0.11784257,0.06164073,0.32814622,0.59283876,0.8575313,1.1222239,1.3869164,2.2625773,3.1382382,4.0120864,4.8877473,5.7615952,6.2384043,6.7115874,7.1883965,7.66158,8.138389,9.157274,10.177972,11.1968565,12.217555,13.238253,14.222692,15.20713,16.193382,17.17782,18.16226,18.00997,17.857681,17.705393,17.553104,17.400814,15.673061,13.945308,12.217555,10.489801,8.762048,7.6017523,6.4432693,5.282973,4.122677,2.962381,3.7347028,4.507025,5.279347,6.051669,6.825804,6.4233265,6.019036,5.618371,5.2158933,4.8116026,6.930956,9.048496,11.164224,13.281764,15.399304,14.219066,13.04064,11.860401,10.680162,9.499924,10.424535,11.350959,12.27557,13.200181,14.124791,14.389484,14.654177,14.920682,15.185374,15.4500675,16.361988,17.27572,18.187641,19.099562,20.013294,18.87294,17.732588,16.592234,15.45188,14.313339,14.289771,14.268016,14.244447,14.222692,14.199123,13.754947,13.310771,12.864782,12.420607,11.974618,9.964043,7.95528,5.9447045,3.9359417,1.9253663,1.7023718,1.4793775,1.258196,1.0352017,0.8122072,0.7179332,0.62184614,0.5275721,0.43329805,0.33721104,8.437528,8.789243,9.142771,9.494485,9.848013,10.199727,10.31757,10.435412,10.553255,10.669285,10.7871275,10.596766,10.408218,10.217857,10.027496,9.837135,9.296872,8.756609,8.21816,7.6778965,7.137634,6.5701766,6.002719,5.4352617,4.8678045,4.3003473,3.6893787,3.0802233,2.469255,1.8600996,1.2491312,1.1494182,1.0497054,0.9499924,0.85027945,0.7505665,1.0696479,1.3905423,1.7096237,2.030518,2.3495996,2.0595255,1.7694515,1.4793775,1.1893034,0.89922947,0.97174793,1.0442665,1.1167849,1.1893034,1.261822,1.1131591,0.96268314,0.8122072,0.66173136,0.51306844,0.42785916,0.34264994,0.2574407,0.17223145,0.0870222,0.21030366,0.33177215,0.4550536,0.57833505,0.69980353,0.7995165,0.89922947,1.0007553,1.1004683,1.2001812,0.97537386,0.7505665,0.52575916,0.2991388,0.07433146,0.11965553,0.16497959,0.21030366,0.25562772,0.2991388,0.23931105,0.1794833,0.11965553,0.059827764,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.065266654,0.054388877,0.045324065,0.034446288,0.025381476,0.36440548,0.70524246,1.0442665,1.3851035,1.7241274,1.3796645,1.0352017,0.69073874,0.3444629,0.0,0.17041849,0.34083697,0.5094425,0.67986095,0.85027945,1.6008459,2.3495996,3.100166,3.8507326,4.599486,3.7691493,2.9406252,2.1102884,1.2799516,0.44961473,0.39522585,0.34083697,0.28463513,0.23024625,0.17585737,0.13959812,0.10515183,0.07070554,0.034446288,0.0,0.0,0.0,0.0,0.0,0.0,0.55476654,1.1095331,1.6642996,2.220879,2.7756457,2.2353828,1.69512,1.1548572,0.61459434,0.07433146,0.4169814,0.75963134,1.1022812,1.4449311,1.7875811,1.6570477,1.5283275,1.3977941,1.2672608,1.1367276,1.1131591,1.0877775,1.062396,1.0370146,1.0116332,0.90466833,0.79770356,0.69073874,0.581961,0.4749962,0.52213323,0.56927025,0.61822027,0.6653573,0.7124943,0.94274056,1.1729867,1.403233,1.6316663,1.8619126,1.6878681,1.5120108,1.3379664,1.162109,0.9880646,1.0080072,1.0279498,1.0478923,1.067835,1.0877775,1.2726997,1.4576219,1.6425442,1.8274662,2.0123885,2.7357605,3.4573197,4.1806917,4.902251,5.6256227,4.6176157,3.6096084,2.6016014,1.5954071,0.5873999,0.6852999,0.78319985,0.8792868,0.97718686,1.0750868,0.98443866,0.89560354,0.80495536,0.71430725,0.62547207,0.69073874,0.7541924,0.8194591,0.88472575,0.9499924,0.8122072,0.6744221,0.53663695,0.40066472,0.26287958,0.22480737,0.18673515,0.15047589,0.11240368,0.07433146,0.11965553,0.16497959,0.21030366,0.25562772,0.2991388,0.3045777,0.3100166,0.3154555,0.3208944,0.3245203,0.32814622,0.32995918,0.33177215,0.33539808,0.33721104,0.32995918,0.32270733,0.3154555,0.30820364,0.2991388,0.23931105,0.1794833,0.11965553,0.059827764,0.0,0.08339628,0.16497959,0.24837588,0.32995918,0.41335547,0.68167394,0.95180535,1.2219368,1.4920682,1.7621996,1.5682126,1.3724127,1.1766127,0.9826257,0.7868258,0.6526665,0.5166943,0.3825351,0.24837588,0.11240368,0.3444629,0.57833505,0.8103943,1.0424535,1.2745126,1.3470312,1.4195497,1.4920682,1.5645868,1.6371052,1.9017978,2.1683033,2.4329958,2.6976883,2.962381,2.9243085,2.8880494,2.8499773,2.811905,2.7756457,2.2643902,1.7549478,1.2455053,0.73424983,0.22480737,0.28463513,0.3444629,0.40429065,0.46411842,0.52575916,0.47318324,0.42060733,0.3680314,0.3154555,0.26287958,0.56927025,0.8774739,1.1856775,1.4920682,1.8002719,1.7549478,1.7096237,1.6642996,1.6207886,1.5754645,1.5083848,1.4394923,1.3724127,1.305333,1.2382535,1.3724127,1.5083848,1.6425442,1.7767034,1.9126755,2.2970235,2.6831846,3.0675328,3.4518807,3.8380418,3.4029307,2.9678197,2.5327086,2.0975976,1.6624867,1.4068589,1.1530442,0.8974165,0.6417888,0.387974,0.6726091,0.9572442,1.2418793,1.5283275,1.8129625,1.6298534,1.4467441,1.2654479,1.0823387,0.89922947,0.79589057,0.69073874,0.5855869,0.48043507,0.37528324,0.34083697,0.3045777,0.27013144,0.23568514,0.19942589,0.2374981,0.2755703,0.31182957,0.34990177,0.387974,0.3100166,0.23205921,0.15410182,0.07795739,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.27194437,0.54570174,0.81764615,1.0895905,1.3633479,1.1747998,0.9880646,0.7995165,0.61278135,0.42423326,0.3444629,0.26469254,0.18492219,0.10515183,0.025381476,0.14503701,0.26469254,0.38434806,0.5058166,0.62547207,0.9119202,1.2001812,1.4866294,1.7748904,2.0631514,1.649796,1.2382535,0.824898,0.41335547,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.3154555,0.629098,0.9445535,1.260009,1.5754645,1.9181144,2.2607644,2.6034143,2.9442513,3.2869012,3.6041696,3.923251,4.2405195,4.557788,4.8750563,4.7554007,4.6357455,4.514277,4.3946214,4.274966,3.4518807,2.6306088,1.8075237,0.98443866,0.16316663,0.49675176,0.8321498,1.167548,1.502946,1.8383441,1.6570477,1.4775645,1.2980812,1.1167849,0.93730164,1.020698,1.1022812,1.1856775,1.2672608,1.3506571,1.0805258,0.8103943,0.5402629,0.27013144,0.0,0.2955129,0.58921283,0.88472575,1.1802386,1.4757515,1.7658255,2.0540867,2.3441606,2.6342347,2.9243085,4.4508233,5.975525,7.500226,9.024928,10.549629,9.80994,9.070251,8.330563,7.590874,6.849373,5.979151,5.1107416,4.2405195,3.3702974,2.5000753,2.1157274,1.7295663,1.3452182,0.96087015,0.5747091,0.58014804,0.5855869,0.58921283,0.5946517,0.6000906,0.5747091,0.5493277,0.52575916,0.50037766,0.4749962,0.42423326,0.37528324,0.3245203,0.2755703,0.22480737,0.19217403,0.15954071,0.12690738,0.09427405,0.06164073,0.23568514,0.40791658,0.58014804,0.7523795,0.9246109,1.6117238,2.3006494,2.9877625,3.6748753,4.361988,4.6629395,4.9620786,5.2630305,5.562169,5.863121,7.192023,8.5227375,9.853452,11.182353,12.513068,13.153044,13.793019,14.432995,15.072971,15.712947,15.528025,15.343102,15.15818,14.973258,14.788336,14.115726,13.443117,12.770509,12.097899,11.42529,9.871581,8.319685,6.7677894,5.2158933,3.6621845,3.9033084,4.1426196,4.3819304,4.6230545,4.8623657,4.6266804,4.3928084,4.157123,3.923251,3.6875658,6.0824895,8.477413,10.872336,13.267261,15.662184,14.454751,13.247317,12.039885,10.832452,9.625018,10.125396,10.625773,11.124338,11.624716,12.125093,12.485873,12.84484,13.20562,13.564586,13.925365,15.4500675,16.97477,18.49947,20.024172,21.550686,20.11482,18.678953,17.2449,15.810846,14.37498,14.409427,14.445685,14.480132,14.514579,14.5508375,13.657047,12.76507,11.873092,10.979301,10.087324,8.384952,6.68258,4.9802084,3.2778363,1.5754645,1.4104849,1.2455053,1.0805258,0.9155461,0.7505665,0.67079616,0.58921283,0.5094425,0.42967212,0.34990177,7.93715,8.232663,8.528176,8.821876,9.117389,9.412902,10.139899,10.866898,11.595709,12.322706,13.049705,12.904668,12.75963,12.6145935,12.469557,12.32452,11.579392,10.834265,10.089137,9.345822,8.600695,7.9842873,7.369693,6.755099,6.1405044,5.52591,4.7191415,3.9141862,3.1092308,2.3042755,1.49932,1.3379664,1.1747998,1.0116332,0.85027945,0.6871128,0.96087015,1.2328146,1.504759,1.7767034,2.0504606,1.8546607,1.6606737,1.4648738,1.2708868,1.0750868,1.1929294,1.310772,1.4268016,1.5446441,1.6624867,1.4503701,1.2382535,1.0243238,0.8122072,0.6000906,0.4949388,0.38978696,0.28463513,0.1794833,0.07433146,0.24293698,0.40972954,0.57833505,0.7451276,0.9119202,1.0497054,1.1874905,1.3252757,1.4630609,1.6008459,1.2998942,1.0007553,0.69980353,0.40066472,0.099712946,0.15954071,0.21936847,0.27919623,0.34083697,0.40066472,0.3208944,0.23931105,0.15954071,0.07977036,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.08339628,0.065266654,0.047137026,0.030820364,0.012690738,0.46955732,0.92823684,1.3851035,1.84197,2.3006494,1.840157,1.3796645,0.91917205,0.4604925,0.0,0.19761293,0.39522585,0.59283876,0.7904517,0.9880646,1.9996977,3.0131438,4.024777,5.038223,6.049856,4.9095025,3.7691493,2.6306088,1.4902552,0.34990177,0.29732585,0.24474995,0.19217403,0.13959812,0.0870222,0.07070554,0.052575916,0.034446288,0.018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.73968875,1.4793775,2.220879,2.960568,3.7002566,2.9805105,2.2607644,1.5392052,0.8194591,0.099712946,0.26469254,0.42967212,0.5946517,0.75963134,0.9246109,1.0352017,1.1457924,1.2545701,1.3651608,1.4757515,1.4503701,1.4249886,1.3996071,1.3742256,1.3506571,1.1657349,0.9808127,0.79589057,0.6091554,0.42423326,0.4169814,0.40972954,0.40247768,0.39522585,0.387974,0.73968875,1.0932164,1.4449311,1.7966459,2.1501737,1.8746033,1.6008459,1.3252757,1.0497054,0.774135,0.9101072,1.0442665,1.1802386,1.3143979,1.4503701,1.6679256,1.8854811,2.1030366,2.3205922,2.5381477,2.8427253,3.147303,3.4518807,3.7582715,4.062849,3.4029307,2.7430124,2.0830941,1.4231756,0.76325727,0.8919776,1.0225109,1.1530442,1.2817645,1.4122978,1.2799516,1.1476053,1.015259,0.88291276,0.7505665,0.69436467,0.6399758,0.5855869,0.5293851,0.4749962,0.42423326,0.37528324,0.3245203,0.2755703,0.22480737,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.059827764,0.08339628,0.10515183,0.12690738,0.15047589,0.15228885,0.15410182,0.15772775,0.15954071,0.16316663,0.19579996,0.22662032,0.25925365,0.291887,0.3245203,0.29007402,0.25562772,0.21936847,0.18492219,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.11059072,0.21936847,0.32995918,0.4405499,0.5493277,0.9101072,1.2708868,1.6298534,1.9906329,2.3495996,2.0903459,1.8292793,1.5700256,1.310772,1.0497054,0.87022203,0.69073874,0.5094425,0.32995918,0.15047589,0.4604925,0.7705091,1.0805258,1.3905423,1.7005589,1.7676386,1.8347181,1.9017978,1.9706904,2.03777,2.420305,2.8028402,3.1853752,3.5679104,3.9504454,3.8996825,3.8507326,3.7999697,3.7492065,3.7002566,3.0203958,2.3405347,1.6606737,0.9808127,0.2991388,0.38072214,0.4604925,0.5402629,0.6200332,0.69980353,0.629098,0.56020546,0.4894999,0.42060733,0.34990177,0.75963134,1.1693609,1.5809034,1.9906329,2.4003625,2.3405347,2.280707,2.220879,2.1592383,2.0994108,2.0105755,1.9199274,1.8292793,1.7404441,1.649796,1.8292793,2.0105755,2.1900587,2.3695421,2.5508385,2.955129,3.3594196,3.7655232,4.169814,4.5759177,3.870675,3.1654327,2.4601903,1.7549478,1.0497054,0.9101072,0.7705091,0.629098,0.4894999,0.34990177,0.7433147,1.1349145,1.5283275,1.9199274,2.3133402,2.077655,1.84197,1.6080978,1.3724127,1.1367276,0.97174793,0.80676836,0.6417888,0.47680917,0.31182957,0.28282216,0.2520018,0.2229944,0.19217403,0.16316663,0.19942589,0.2374981,0.2755703,0.31182957,0.34990177,0.27919623,0.21030366,0.13959812,0.07070554,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14322405,0.28463513,0.42785916,0.56927025,0.7124943,0.66173136,0.61278135,0.5620184,0.51306844,0.46230546,0.37165734,0.28282216,0.19217403,0.10333887,0.012690738,0.11059072,0.20667773,0.3045777,0.40247768,0.50037766,0.76325727,1.0243238,1.2872034,1.550083,1.8129625,1.4503701,1.0877775,0.72518504,0.36259252,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.30820364,0.61459434,0.922798,1.2291887,1.5373923,1.6896812,1.84197,1.9942589,2.1483607,2.3006494,2.565342,2.8300345,3.094727,3.3594196,3.6241121,3.9395678,4.255023,4.5704784,4.8841214,5.199577,4.195195,3.1908143,2.18462,1.1802386,0.17585737,0.55476654,0.9354887,1.3143979,1.69512,2.0758421,1.8347181,1.5954071,1.3542831,1.114972,0.87566096,0.98443866,1.0950294,1.2056202,1.3143979,1.4249886,1.1403534,0.8557183,0.56927025,0.28463513,0.0,0.18492219,0.36984438,0.55476654,0.73968875,0.9246109,1.4068589,1.889107,2.373168,2.855416,3.3376641,4.650249,5.962834,7.2754188,8.588004,9.900589,9.168152,8.435715,7.703278,6.970841,6.2365913,5.4515786,4.668379,3.8833659,3.0983531,2.3133402,1.9072367,1.502946,1.0968424,0.69255173,0.28826106,0.29007402,0.291887,0.2955129,0.29732585,0.2991388,0.28826106,0.2755703,0.26287958,0.25018883,0.2374981,0.21211663,0.18673515,0.16316663,0.13778515,0.11240368,0.10333887,0.092461094,0.08339628,0.072518505,0.06164073,0.14322405,0.2229944,0.30276474,0.3825351,0.46230546,0.96268314,1.4630609,1.9616255,2.4620032,2.962381,3.0874753,3.2125697,3.3376641,3.4627585,3.587853,5.2267714,6.867502,8.508233,10.147152,11.787883,12.083396,12.377095,12.672608,12.968122,13.261822,13.044266,12.826711,12.609155,12.3916,12.175857,12.558392,12.939114,13.321649,13.704185,14.0867195,12.143224,10.197914,8.252605,6.3072968,4.361988,4.070101,3.778214,3.484514,3.1926272,2.9007401,2.8318477,2.764768,2.6976883,2.6306088,2.561716,5.235836,7.9081426,10.58045,13.252756,15.925063,14.690435,13.453996,12.219368,10.98474,9.750113,9.824444,9.900589,9.97492,10.049252,10.125396,10.58045,11.035503,11.490557,11.94561,12.400664,14.538147,16.67563,18.813112,20.950596,23.088078,21.356699,19.627132,17.897566,16.168001,14.436621,14.530895,14.623356,14.715817,14.808278,14.90074,13.559147,12.219368,10.879588,9.539809,8.200029,6.8040485,5.40988,4.0157123,2.619731,1.2255627,1.1167849,1.0098201,0.90285534,0.79589057,0.6871128,0.62184614,0.55839247,0.49312583,0.42785916,0.36259252,7.4367723,7.6742706,7.911769,8.149267,8.386765,8.624263,9.96223,11.300196,12.638163,13.974316,15.312282,15.212569,15.112856,15.013144,14.911617,14.811904,13.861912,12.91192,11.961927,11.011934,10.061942,9.400211,8.736667,8.074935,7.413204,6.7496595,5.750717,4.749962,3.7492065,2.7502642,1.7495089,1.5247015,1.2998942,1.0750868,0.85027945,0.62547207,0.85027945,1.0750868,1.2998942,1.5247015,1.7495089,1.649796,1.550083,1.4503701,1.3506571,1.2491312,1.4122978,1.5754645,1.7368182,1.8999848,2.0631514,1.7875811,1.5120108,1.2382535,0.96268314,0.6871128,0.5620184,0.43692398,0.31182957,0.18673515,0.06164073,0.2755703,0.48768693,0.69980353,0.9119202,1.1258497,1.2998942,1.4757515,1.649796,1.8256533,1.9996977,1.6244144,1.2491312,0.87566096,0.50037766,0.12509441,0.19942589,0.2755703,0.34990177,0.42423326,0.50037766,0.40066472,0.2991388,0.19942589,0.099712946,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.5747091,1.1494182,1.7241274,2.3006494,2.8753586,2.3006494,1.7241274,1.1494182,0.5747091,0.0,0.22480737,0.44961473,0.6744221,0.89922947,1.1258497,2.4003625,3.6748753,4.949388,6.2257137,7.500226,6.049856,4.599486,3.149116,1.7005589,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.9246109,1.8492218,2.7756457,3.7002566,4.6248674,3.7256382,2.8245957,1.9253663,1.0243238,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.41335547,0.76325727,1.1131591,1.4630609,1.8129625,1.7875811,1.7621996,1.7368182,1.7132497,1.6878681,1.4249886,1.162109,0.89922947,0.63816285,0.37528324,0.31182957,0.25018883,0.18673515,0.12509441,0.06164073,0.53663695,1.0116332,1.4866294,1.9616255,2.4366217,2.0631514,1.6878681,1.3125849,0.93730164,0.5620184,0.8122072,1.062396,1.3125849,1.5627737,1.8129625,2.0631514,2.3133402,2.561716,2.811905,3.0620937,2.94969,2.8372865,2.7248828,2.612479,2.5000753,2.1882458,1.8746033,1.5627737,1.2491312,0.93730164,1.1004683,1.261822,1.4249886,1.5881553,1.7495089,1.5754645,1.3996071,1.2255627,1.0497054,0.87566096,0.69980353,0.52575916,0.34990177,0.17585737,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06164073,0.12509441,0.18673515,0.25018883,0.31182957,0.25018883,0.18673515,0.12509441,0.06164073,0.0,0.0,0.0,0.0,0.0,0.0,0.13778515,0.2755703,0.41335547,0.5493277,0.6871128,1.1367276,1.5881553,2.03777,2.4873846,2.9369993,2.612479,2.2879589,1.9616255,1.6371052,1.3125849,1.0877775,0.8629702,0.63816285,0.41335547,0.18673515,0.5747091,0.96268314,1.3506571,1.7368182,2.124792,2.1882458,2.2498865,2.3133402,2.374981,2.4366217,2.9369993,3.437377,3.9377546,4.4381323,4.936697,4.8750563,4.8116026,4.749962,4.688321,4.6248674,3.774588,2.9243085,2.0758421,1.2255627,0.37528324,0.4749962,0.5747091,0.6744221,0.774135,0.87566096,0.7868258,0.69980353,0.61278135,0.52575916,0.43692398,0.9499924,1.4630609,1.9743162,2.4873846,3.000453,2.9243085,2.8499773,2.7756457,2.6995013,2.6251698,2.5127661,2.4003625,2.2879589,2.175555,2.0631514,2.2879589,2.5127661,2.7375734,2.962381,3.1871881,3.6132345,4.0374675,4.461701,4.8877473,5.3119802,4.3366065,3.3630457,2.3876717,1.4122978,0.43692398,0.41335547,0.387974,0.36259252,0.33721104,0.31182957,0.8122072,1.3125849,1.8129625,2.3133402,2.811905,2.525457,2.2371957,1.9507477,1.6624867,1.3742256,1.1494182,0.9246109,0.69980353,0.4749962,0.25018883,0.22480737,0.19942589,0.17585737,0.15047589,0.12509441,0.16316663,0.19942589,0.2374981,0.2755703,0.31182957,0.25018883,0.18673515,0.12509441,0.06164073,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.15047589,0.2374981,0.3245203,0.41335547,0.50037766,0.40066472,0.2991388,0.19942589,0.099712946,0.0,0.07433146,0.15047589,0.22480737,0.2991388,0.37528324,0.61278135,0.85027945,1.0877775,1.3252757,1.5627737,1.2491312,0.93730164,0.62547207,0.31182957,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.2991388,0.6000906,0.89922947,1.2001812,1.49932,1.4630609,1.4249886,1.3869164,1.3506571,1.3125849,1.5247015,1.7368182,1.9507477,2.1628644,2.374981,3.1255474,3.874301,4.6248674,5.375434,6.1241875,4.936697,3.7492065,2.561716,1.3742256,0.18673515,0.61278135,1.0370146,1.4630609,1.887294,2.3133402,2.0123885,1.7132497,1.4122978,1.1131591,0.8122072,0.9499924,1.0877775,1.2255627,1.3633479,1.49932,1.2001812,0.89922947,0.6000906,0.2991388,0.0,0.07433146,0.15047589,0.22480737,0.2991388,0.37528324,1.0497054,1.7241274,2.4003625,3.0747845,3.7492065,4.8496747,5.9501433,7.0506115,8.149267,9.249735,8.52455,7.799365,7.07418,6.350808,5.6256227,4.9258194,4.2242026,3.5243993,2.8245957,2.124792,1.7005589,1.2745126,0.85027945,0.42423326,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.31182957,0.62547207,0.93730164,1.2491312,1.5627737,1.5120108,1.4630609,1.4122978,1.3633479,1.3125849,3.2633326,5.2122674,7.1630154,9.11195,11.062697,11.011934,10.962985,10.912222,10.863272,10.812509,10.56232,10.312131,10.061942,9.811753,9.563377,10.999244,12.436923,13.874602,15.312282,16.749962,14.413053,12.07433,9.737422,7.400513,5.0617914,4.2368937,3.4119956,2.5870976,1.7621996,0.93730164,1.0370146,1.1367276,1.2382535,1.3379664,1.4376793,4.3873696,7.3370595,10.28675,13.23644,16.187943,14.924308,13.662486,12.400664,11.137029,9.875207,9.525306,9.175404,8.825501,8.4756,8.125698,8.675026,9.224354,9.775495,10.324821,10.874149,13.6244135,16.374678,19.124943,21.875206,24.625471,22.600391,20.575312,18.550234,16.525154,14.500074,14.650551,14.799213,14.94969,15.100165,15.250641,13.46306,11.675479,9.8878975,8.100317,6.3127356,5.224958,4.137181,3.049403,1.9634385,0.87566096,0.824898,0.774135,0.72518504,0.6744221,0.62547207,0.5747091,0.52575916,0.4749962,0.42423326,0.37528324,8.649645,8.792869,8.934279,9.077503,9.220728,9.362139,10.279498,11.1968565,12.114216,13.033388,13.9507475,13.765825,13.57909,13.394168,13.209246,13.024323,12.402477,11.780631,11.156972,10.535126,9.91328,9.612328,9.313189,9.012237,8.713099,8.412147,7.752228,7.0923095,6.432391,5.772473,5.1125546,4.267714,3.4228733,2.5780327,1.7331922,0.8883517,1.0732739,1.258196,1.4431182,1.6280404,1.8129625,1.6751775,1.5373923,1.3996071,1.261822,1.1258497,1.3397794,1.5555218,1.7694515,1.9851941,2.1991236,1.9416829,1.6842422,1.4268016,1.1693609,0.9119202,0.7850128,0.65810543,0.5293851,0.40247768,0.2755703,0.43511102,0.5946517,0.7541924,0.9155461,1.0750868,1.209246,1.3452182,1.4793775,1.6153497,1.7495089,1.5392052,1.3307146,1.1204109,0.9101072,0.69980353,0.85934424,1.020698,1.1802386,1.3397794,1.49932,1.2219368,0.9445535,0.6671702,0.38978696,0.11240368,0.12328146,0.13234627,0.14322405,0.15228885,0.16316663,0.13415924,0.10696479,0.07977036,0.052575916,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.03988518,0.054388877,0.07070554,0.08520924,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.48043507,0.96087015,1.4394923,1.9199274,2.4003625,1.9942589,1.5899682,1.1856775,0.7795739,0.37528324,0.48224804,0.58921283,0.6979906,0.80495536,0.9119202,1.9525607,2.9932013,4.0320287,5.0726695,6.11331,4.9294453,3.7473936,2.565342,1.3832904,0.19942589,0.15954071,0.11965553,0.07977036,0.03988518,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,1.2074331,2.3894846,3.5733492,4.7554007,5.9374523,4.835171,3.73289,2.6306088,1.5283275,0.42423326,0.58921283,0.7541924,0.91917205,1.0841516,1.2491312,1.7205015,2.1900587,2.659616,3.1291735,3.6005437,3.4228733,3.245203,3.0675328,2.8898623,2.712192,2.5327086,2.3532255,2.1719291,1.9924458,1.8129625,1.6443571,1.4775645,1.310772,1.1421664,0.97537386,1.1947423,1.4141108,1.6352923,1.8546607,2.0758421,2.2118144,2.3495996,2.4873846,2.6251698,2.762955,3.395679,4.028403,4.6593137,5.292038,5.924762,6.1169357,6.3109226,6.5030966,6.695271,6.887445,5.964647,5.041849,4.120864,3.198066,2.275268,2.084907,1.8945459,1.7041848,1.5156367,1.3252757,1.3669738,1.4104849,1.452183,1.4956942,1.5373923,1.3705997,1.2019942,1.0352017,0.8665961,0.69980353,0.56020546,0.42060733,0.27919623,0.13959812,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13415924,0.27013144,0.40429065,0.5402629,0.6744221,0.8430276,1.0098201,1.1784257,1.3452182,1.5120108,1.5827163,1.6534219,1.7223145,1.79302,1.8619126,2.0722163,2.2825198,2.4928236,2.7031271,2.913431,3.3231604,3.73289,4.1426196,4.552349,4.9620786,4.610364,4.256836,3.9051213,3.5534067,3.199879,2.6904364,2.179181,1.6697385,1.1602961,0.6508536,1.020698,1.3905423,1.7603867,2.1302311,2.5000753,2.6777458,2.855416,3.0330863,3.2107568,3.388427,3.5733492,3.7582715,3.9431937,4.1281157,4.313038,4.1933823,4.071914,3.9522583,3.832603,3.7129474,3.0403383,2.3677292,1.69512,1.0225109,0.34990177,0.49312583,0.6345369,0.7777609,0.91917205,1.062396,0.93911463,0.81764615,0.69436467,0.5728962,0.44961473,0.83940166,1.2291887,1.6207886,2.0105755,2.4003625,2.5544643,2.7103791,2.864481,3.0203958,3.1744974,3.002266,2.8300345,2.657803,2.4855716,2.3133402,2.3949237,2.47832,2.5599031,2.6432993,2.7248828,3.0729716,3.4192474,3.7673361,4.115425,4.461701,3.6476808,2.8318477,2.0178273,1.2019942,0.387974,0.36077955,0.33177215,0.3045777,0.27738327,0.25018883,0.6544795,1.0605831,1.4648738,1.8691645,2.275268,2.0468347,1.8202144,1.5917811,1.3651608,1.1367276,0.9826257,0.82671094,0.6726091,0.5166943,0.36259252,0.33721104,0.31182957,0.28826106,0.26287958,0.2374981,0.24474995,0.2520018,0.25925365,0.26831847,0.2755703,0.21936847,0.16497959,0.11059072,0.054388877,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.032633327,0.065266654,0.09789998,0.13053331,0.16316663,0.21030366,0.2574407,0.3045777,0.35171473,0.40066472,0.3208944,0.23931105,0.15954071,0.07977036,0.0,0.06164073,0.12509441,0.18673515,0.25018883,0.31182957,0.59283876,0.872035,1.1530442,1.4322405,1.7132497,1.3778516,1.0424535,0.7070554,0.37165734,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.23568514,0.45686656,0.67986095,0.90285534,1.1258497,1.1856775,1.2455053,1.305333,1.3651608,1.4249886,1.357909,1.2908293,1.2219368,1.1548572,1.0877775,1.6280404,2.1683033,2.7067533,3.247016,3.787279,4.942136,6.096993,7.25185,8.406708,9.563377,7.71053,5.857682,4.004834,2.1519866,0.2991388,0.6327239,0.9644961,1.2980812,1.6298534,1.9616255,1.7005589,1.4376793,1.1747998,0.9119202,0.6508536,0.7777609,0.90466833,1.0333886,1.1602961,1.2872034,1.0297627,0.77232206,0.5148814,0.2574407,0.0,0.059827764,0.11965553,0.1794833,0.23931105,0.2991388,0.85934424,1.4195497,1.9797552,2.5399606,3.100166,4.079166,5.0599785,6.0407915,7.019791,8.000604,7.36788,6.735156,6.1024323,5.469708,4.836984,4.209699,3.5824142,2.955129,2.327844,1.7005589,1.3597219,1.020698,0.67986095,0.34083697,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.25018883,0.50037766,0.7505665,1.0007553,1.2491312,1.2291887,1.209246,1.1893034,1.1693609,1.1494182,3.0222087,4.894999,6.7677894,8.640579,10.51337,10.51337,10.51337,10.51337,10.51337,10.51337,10.536939,10.56232,10.587702,10.613083,10.636651,11.731681,12.826711,13.92174,15.016769,16.1118,14.320591,12.527572,10.734551,8.943344,7.1503243,6.5556726,5.959208,5.3645563,4.7699046,4.175253,4.749962,5.3246713,5.89938,6.4759026,7.0506115,8.733041,10.41547,12.097899,13.780329,15.462758,14.19731,12.931862,11.668227,10.40278,9.137331,8.977791,8.81825,8.656897,8.497355,8.337815,8.689529,9.043057,9.394773,9.7483,10.100015,12.250188,14.400362,16.550535,18.698896,20.84907,19.572744,18.294605,17.01828,15.740141,14.462003,14.554463,14.646925,14.739386,14.831847,14.924308,13.252756,11.579392,9.907841,8.234476,6.5629244,5.582112,4.603112,3.6222992,2.6432993,1.6624867,1.4648738,1.2672608,1.0696479,0.872035,0.6744221,0.6091554,0.54570174,0.48043507,0.41516843,0.34990177,9.862516,9.909654,9.956791,10.00574,10.052877,10.100015,10.596766,11.095331,11.592083,12.090648,12.5873995,12.317267,12.047136,11.777005,11.506873,11.236742,10.943042,10.64753,10.352016,10.058316,9.762803,9.824444,9.8878975,9.949538,10.012992,10.074633,9.755551,9.434657,9.115576,8.794682,8.4756,7.0107265,5.5458527,4.079166,2.6142921,1.1494182,1.2944553,1.4394923,1.5845293,1.7295663,1.8746033,1.7005589,1.5247015,1.3506571,1.1747998,1.0007553,1.2672608,1.5355793,1.8020848,2.0704033,2.3369088,2.0975976,1.8582866,1.6171626,1.3778516,1.1367276,1.0080072,0.8774739,0.7469406,0.61822027,0.48768693,0.5946517,0.7016165,0.8103943,0.91735905,1.0243238,1.1204109,1.214685,1.310772,1.405046,1.49932,1.455809,1.4104849,1.3651608,1.3198367,1.2745126,1.5192627,1.7658255,2.0105755,2.2553256,2.5000753,2.0450218,1.5899682,1.1349145,0.67986095,0.22480737,0.24474995,0.26469254,0.28463513,0.3045777,0.3245203,0.27013144,0.21574254,0.15954071,0.10515183,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.054388877,0.059827764,0.065266654,0.07070554,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.38434806,0.7705091,1.1548572,1.5392052,1.9253663,1.6896812,1.455809,1.2201238,0.98443866,0.7505665,0.73968875,0.7306239,0.7197462,0.7106813,0.69980353,1.504759,2.3097143,3.1146698,3.919625,4.7245803,3.8108473,2.8953013,1.9797552,1.064209,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,1.4902552,2.9297476,4.36924,5.810545,7.250037,5.9447045,4.6393714,3.3358512,2.030518,0.72518504,1.067835,1.4104849,1.7531348,2.0957847,2.4366217,3.0276475,3.6168604,4.207886,4.797099,5.388125,5.0581656,4.7282066,4.3982472,4.068288,3.738329,3.6404288,3.5425289,3.444629,3.346729,3.2506418,2.9768846,2.70494,2.4329958,2.1592383,1.887294,1.8528478,1.8184015,1.7821422,1.7476959,1.7132497,2.3622901,3.0131438,3.6621845,4.313038,4.9620786,5.977338,6.9925966,8.007855,9.023115,10.038374,10.172533,10.306692,10.442664,10.576823,10.712796,8.979604,7.2482243,5.5150323,3.7818398,2.0504606,1.983381,1.9144884,1.8474089,1.7803292,1.7132497,1.6352923,1.5573349,1.4793775,1.403233,1.3252757,1.1657349,1.0043813,0.8448406,0.6852999,0.52575916,0.42060733,0.3154555,0.21030366,0.10515183,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.09064813,0.06707962,0.045324065,0.02175555,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.20667773,0.41516843,0.62184614,0.83033687,1.0370146,1.4358664,1.8329052,2.229944,2.6269827,3.0258346,3.1654327,3.3050308,3.444629,3.584227,3.7256382,4.006647,4.2894692,4.572292,4.855114,5.137936,5.5077806,5.8776245,6.247469,6.6173134,6.987158,6.6082487,6.2275267,5.846804,5.467895,5.087173,4.2930956,3.4972048,2.7031271,1.9072367,1.1131591,1.4648738,1.8165885,2.1701162,2.521831,2.8753586,3.1672456,3.4591327,3.7528327,4.0447197,4.3366065,4.207886,4.077353,3.9468195,3.8180993,3.6875658,3.5098956,3.3322253,3.1545548,2.9768846,2.7992141,2.3042755,1.8093367,1.3143979,0.8194591,0.3245203,0.5094425,0.69436467,0.8792868,1.064209,1.2491312,1.0932164,0.9354887,0.7777609,0.6200332,0.46230546,0.7306239,0.99712944,1.2654479,1.5319533,1.8002719,2.18462,2.570781,2.955129,3.339477,3.7256382,3.491766,3.2597067,3.0276475,2.7955883,2.561716,2.5018883,2.4420607,2.382233,2.322405,2.2625773,2.5327086,2.8028402,3.0729716,3.343103,3.6132345,2.956942,2.3024626,1.647983,0.9916905,0.33721104,0.30820364,0.27738327,0.24837588,0.21755551,0.18673515,0.49675176,0.80676836,1.1167849,1.4268016,1.7368182,1.5700256,1.403233,1.2346275,1.067835,0.89922947,0.81583315,0.7306239,0.64541465,0.56020546,0.4749962,0.44961473,0.42423326,0.40066472,0.37528324,0.34990177,0.32814622,0.3045777,0.28282216,0.25925365,0.2374981,0.19036107,0.14322405,0.09427405,0.047137026,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.052575916,0.10515183,0.15772775,0.21030366,0.26287958,0.27013144,0.27738327,0.28463513,0.291887,0.2991388,0.23931105,0.1794833,0.11965553,0.059827764,0.0,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,0.5728962,0.89560354,1.2183108,1.5392052,1.8619126,1.504759,1.1476053,0.7904517,0.43329805,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.46955732,0.9155461,1.3597219,1.8057107,2.2498865,2.0704033,1.889107,1.7096237,1.5301404,1.3506571,1.2527572,1.1548572,1.0569572,0.96087015,0.8629702,1.7295663,2.5979755,3.4645715,4.3329806,5.199577,6.7605376,8.319685,9.880646,11.439794,13.000754,10.48255,7.9643445,5.4479527,2.9297476,0.41335547,0.6526665,0.8919776,1.1331016,1.3724127,1.6117238,1.3869164,1.162109,0.93730164,0.7124943,0.48768693,0.6055295,0.72337204,0.83940166,0.9572442,1.0750868,0.85934424,0.64541465,0.42967212,0.21574254,0.0,0.045324065,0.09064813,0.13415924,0.1794833,0.22480737,0.67079616,1.114972,1.5591478,2.0051367,2.4493124,3.3104696,4.169814,5.029158,5.8903155,6.7496595,6.209397,5.669134,5.130684,4.590421,4.0501585,3.4953918,2.9406252,2.3858588,1.8292793,1.2745126,1.020698,0.7650702,0.5094425,0.25562772,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.18673515,0.37528324,0.5620184,0.7505665,0.93730164,0.9481794,0.9572442,0.968122,0.97718686,0.9880646,2.7828975,4.5777307,6.3725634,8.167397,9.96223,10.012992,10.061942,10.112705,10.161655,10.212419,10.51337,10.812509,11.111648,11.4126,11.711739,12.465931,13.21831,13.97069,14.723069,15.475449,14.22813,12.980812,11.731681,10.484363,9.237044,8.872639,8.508233,8.1420145,7.7776093,7.413204,8.46291,9.512614,10.56232,11.612025,12.661731,13.0769,13.492067,13.907236,14.322405,14.737573,13.470312,12.203052,10.93579,9.666717,8.399456,8.430276,8.459284,8.490104,8.519112,8.549932,8.705847,8.859948,9.015862,9.169965,9.325879,10.875962,12.426045,13.974316,15.524399,17.074482,16.545097,16.01571,15.484513,14.955129,14.425743,14.46019,14.494636,14.530895,14.565341,14.599788,13.042453,11.485118,9.927783,8.370448,6.813113,5.9392653,5.06723,4.195195,3.3231604,2.4493124,2.1048496,1.7603867,1.4141108,1.0696479,0.72518504,0.64541465,0.5656443,0.48587397,0.40429065,0.3245203,11.075388,11.028252,10.979301,10.932164,10.885027,10.837891,10.915848,10.991992,11.069949,11.147907,11.225864,10.870523,10.515183,10.1598425,9.804502,9.449161,9.481794,9.514427,9.547061,9.579695,9.612328,10.038374,10.462607,10.88684,11.312886,11.73712,11.757062,11.777005,11.7969475,11.81689,11.836833,9.751925,7.667019,5.582112,3.4972048,1.4122978,1.5174497,1.6226015,1.7277533,1.8329052,1.938057,1.7241274,1.5120108,1.2998942,1.0877775,0.87566096,1.1947423,1.5156367,1.8347181,2.1556125,2.474694,2.2516994,2.030518,1.8075237,1.5845293,1.3633479,1.2291887,1.0968424,0.9644961,0.8321498,0.69980353,0.7541924,0.8103943,0.86478317,0.91917205,0.97537386,1.0297627,1.0841516,1.1403534,1.1947423,1.2491312,1.3705997,1.4902552,1.6099107,1.7295663,1.8492218,2.179181,2.5091403,2.8390994,3.1708715,3.5008307,2.8681068,2.2353828,1.6026589,0.969935,0.33721104,0.3680314,0.39703882,0.42785916,0.45686656,0.48768693,0.40429065,0.32270733,0.23931105,0.15772775,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.07070554,0.065266654,0.059827764,0.054388877,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.29007402,0.58014804,0.87022203,1.1602961,1.4503701,1.3851035,1.3198367,1.2545701,1.1893034,1.1258497,0.99712944,0.87022203,0.7433147,0.61459434,0.48768693,1.0569572,1.6280404,2.1973107,2.7683938,3.3376641,2.6904364,2.0432088,1.3941683,0.7469406,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,1.7730774,3.4700103,5.1669436,6.8656893,8.562622,7.0542374,5.5476656,4.0392804,2.5327086,1.0243238,1.5446441,2.0649643,2.5852847,3.105605,3.6241121,4.3347936,5.045475,5.754343,6.4650245,7.175706,6.6916447,6.209397,5.727149,5.2449007,4.762653,4.748149,4.7318325,4.7173285,4.702825,4.688321,4.309412,3.9323158,3.5552197,3.1781235,2.7992141,2.5091403,2.220879,1.9308052,1.6407311,1.3506571,2.5127661,3.6748753,4.836984,6.000906,7.1630154,8.560809,9.956791,11.354585,12.752378,14.150173,14.22813,14.304275,14.382232,14.46019,14.538147,11.99456,9.452786,6.9092,4.367427,1.8256533,1.8800422,1.9344311,1.9906329,2.0450218,2.0994108,1.9017978,1.7041848,1.5083848,1.310772,1.1131591,0.96087015,0.80676836,0.6544795,0.50219065,0.34990177,0.27919623,0.21030366,0.13959812,0.07070554,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.27919623,0.56020546,0.83940166,1.1204109,1.3996071,2.0268922,2.6541772,3.2832751,3.9105604,4.537845,4.748149,4.95664,5.1669436,5.377247,5.5875506,5.942891,6.298232,6.6517596,7.0071006,7.362441,7.6924005,8.02236,8.352319,8.682278,9.012237,8.604321,8.198216,7.7903004,7.382384,6.9744673,5.8957543,4.8152285,3.7347028,2.6541772,1.5754645,1.9108626,2.2444477,2.5798457,2.9152439,3.2506418,3.6567454,4.064662,4.4725785,4.880495,5.2865987,4.842423,4.3982472,3.9522583,3.5080826,3.0620937,2.8282216,2.5925364,2.3568513,2.1229792,1.887294,1.5700256,1.2527572,0.9354887,0.61822027,0.2991388,0.5275721,0.7541924,0.9826257,1.209246,1.4376793,1.2455053,1.0533313,0.85934424,0.6671702,0.4749962,0.6200332,0.7650702,0.9101072,1.0551442,1.2001812,1.8147756,2.42937,3.045777,3.6603715,4.274966,3.9830787,3.6893787,3.397492,3.105605,2.811905,2.610666,2.4076142,2.2045624,2.0033236,1.8002719,1.9924458,2.18462,2.3767939,2.570781,2.762955,2.268016,1.7730774,1.2781386,0.78319985,0.28826106,0.25562772,0.2229944,0.19036107,0.15772775,0.12509441,0.34083697,0.55476654,0.7705091,0.98443866,1.2001812,1.0932164,0.98443866,0.8774739,0.7705091,0.66173136,0.64722764,0.6327239,0.61822027,0.60190356,0.5873999,0.5620184,0.53663695,0.51306844,0.48768693,0.46230546,0.40972954,0.35715362,0.3045777,0.2520018,0.19942589,0.15954071,0.11965553,0.07977036,0.03988518,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.072518505,0.14503701,0.21755551,0.29007402,0.36259252,0.32995918,0.29732585,0.26469254,0.23205921,0.19942589,0.15954071,0.11965553,0.07977036,0.03988518,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.5529536,0.91735905,1.2817645,1.647983,2.0123885,1.6316663,1.2527572,0.872035,0.49312583,0.11240368,0.09064813,0.06707962,0.045324065,0.02175555,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.70524246,1.3724127,2.039583,2.7067533,3.3757362,2.955129,2.5345216,2.1157274,1.69512,1.2745126,1.1476053,1.020698,0.8919776,0.7650702,0.63816285,1.8329052,3.0276475,4.2223897,5.4171324,6.6118746,8.577126,10.542377,12.507628,14.47288,16.438131,13.254569,10.07282,6.889258,3.7075086,0.52575916,0.6726091,0.8194591,0.968122,1.114972,1.261822,1.0750868,0.8883517,0.69980353,0.51306844,0.3245203,0.43329805,0.5402629,0.64722764,0.7541924,0.8629702,0.69073874,0.5166943,0.3444629,0.17223145,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.48043507,0.8103943,1.1403534,1.4703126,1.8002719,2.5399606,3.2796493,4.019338,4.76084,5.5005283,5.0527267,4.604925,4.157123,3.7093215,3.2633326,2.7792716,2.2970235,1.8147756,1.3325275,0.85027945,0.67986095,0.5094425,0.34083697,0.17041849,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.12509441,0.25018883,0.37528324,0.50037766,0.62547207,0.6653573,0.70524246,0.7451276,0.7850128,0.824898,2.5417736,4.2604623,5.977338,7.6942134,9.412902,9.512614,9.612328,9.712041,9.811753,9.91328,10.487988,11.062697,11.637406,12.212116,12.786825,13.198368,13.608097,14.017827,14.427556,14.837286,14.13567,13.43224,12.730623,12.027194,11.325577,11.189605,11.055446,10.919474,10.785315,10.649343,12.175857,13.700559,15.22526,16.749962,18.274662,17.422571,16.570478,15.716573,14.86448,14.012388,12.743314,11.472427,10.203354,8.9324665,7.663393,7.8827615,8.10213,8.323311,8.54268,8.762048,8.72035,8.676839,8.63514,8.59163,8.549932,9.499924,10.449916,11.399909,12.349901,13.299893,13.517449,13.735004,13.95256,14.170115,14.387671,14.364102,14.342347,14.320591,14.297023,14.275268,12.8321495,11.389031,9.947725,8.504607,7.063302,6.298232,5.5331616,4.7680917,4.0030212,3.2379513,2.7448254,2.2516994,1.7603867,1.2672608,0.774135,0.67986095,0.5855869,0.4894999,0.39522585,0.2991388,12.28826,12.145037,12.001812,11.860401,11.717177,11.575767,11.233116,10.890467,10.547816,10.205167,9.862516,9.421967,8.98323,8.54268,8.10213,7.66158,8.02236,8.383139,8.7421055,9.102885,9.461852,10.25049,11.037316,11.8241415,12.612781,13.399607,13.760386,14.119352,14.480132,14.840912,15.199879,12.494938,9.789998,7.0850577,4.3801174,1.6751775,1.7404441,1.8057107,1.8691645,1.9344311,1.9996977,1.7495089,1.49932,1.2491312,1.0007553,0.7505665,1.1222239,1.4956942,1.8673514,2.2408218,2.612479,2.4076142,2.2027495,1.9978848,1.79302,1.5881553,1.452183,1.3180238,1.1820517,1.0478923,0.9119202,0.9155461,0.91735905,0.91917205,0.922798,0.9246109,0.93911463,0.9554313,0.969935,0.98443866,1.0007553,1.2853905,1.5700256,1.8546607,2.1392958,2.4257438,2.8390994,3.254268,3.6694362,4.0846047,4.499773,3.6893787,2.8807976,2.0704033,1.260009,0.44961473,0.4894999,0.5293851,0.56927025,0.6091554,0.6508536,0.5402629,0.42967212,0.3208944,0.21030366,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.08520924,0.07070554,0.054388877,0.03988518,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.19579996,0.38978696,0.5855869,0.7795739,0.97537386,1.0805258,1.1856775,1.2908293,1.3941683,1.49932,1.2545701,1.0098201,0.7650702,0.52032024,0.2755703,0.6091554,0.9445535,1.2799516,1.6153497,1.9507477,1.5700256,1.1893034,0.8103943,0.42967212,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,2.0540867,4.0102735,5.964647,7.9208336,9.875207,8.165584,6.45596,4.744523,3.0348995,1.3252757,2.0232663,2.7194438,3.4174345,4.115425,4.8134155,5.6419396,6.472276,7.3026133,8.13295,8.963287,8.326937,7.6924005,7.057863,6.4233265,5.7869763,5.8558693,5.922949,5.9900284,6.057108,6.1241875,5.6419396,5.1596913,4.6774435,4.195195,3.7129474,3.1672456,2.6233568,2.077655,1.5319533,0.9880646,2.663242,4.3366065,6.011784,7.686961,9.362139,11.142468,12.922797,14.703127,16.483456,18.261972,18.281914,18.301857,18.3218,18.341742,18.361685,15.009518,11.65735,8.3051815,4.953014,1.6008459,1.7767034,1.9543737,2.132044,2.3097143,2.4873846,2.1701162,1.8528478,1.5355793,1.2183108,0.89922947,0.7541924,0.6091554,0.46411842,0.3208944,0.17585737,0.13959812,0.10515183,0.07070554,0.034446288,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.35171473,0.70524246,1.0569572,1.4104849,1.7621996,2.619731,3.4772623,4.3347936,5.1923246,6.049856,6.3308654,6.6100616,6.889258,7.170267,7.4494634,7.877322,8.3051815,8.733041,9.1609,9.5869465,9.87702,10.167094,10.457169,10.747242,11.037316,10.602205,10.167094,9.731983,9.296872,8.861761,7.498413,6.1332526,4.7680917,3.4029307,2.03777,2.3550384,2.6723068,2.9895754,3.3068438,3.6241121,4.1480584,4.670192,5.1923246,5.714458,6.2384043,5.47696,4.7173285,3.9576974,3.198066,2.4366217,2.1447346,1.8528478,1.5591478,1.2672608,0.97537386,0.83577573,0.69436467,0.55476654,0.41516843,0.2755703,0.54570174,0.81583315,1.0841516,1.3542831,1.6244144,1.3977941,1.1693609,0.94274056,0.71430725,0.48768693,0.5094425,0.533011,0.55476654,0.57833505,0.6000906,1.4449311,2.2897718,3.1346123,3.9794528,4.8242936,4.4725785,4.120864,3.7673361,3.4156215,3.0620937,2.7176309,2.373168,2.0268922,1.6824293,1.3379664,1.452183,1.5682126,1.6824293,1.7966459,1.9126755,1.5772774,1.2418793,0.90829426,0.5728962,0.2374981,0.2030518,0.16679256,0.13234627,0.09789998,0.06164073,0.18310922,0.30276474,0.4224203,0.5420758,0.66173136,0.61459434,0.56745726,0.52032024,0.47318324,0.42423326,0.48043507,0.53482395,0.58921283,0.64541465,0.69980353,0.6744221,0.6508536,0.62547207,0.6000906,0.5747091,0.49312583,0.40972954,0.32814622,0.24474995,0.16316663,0.13053331,0.09789998,0.065266654,0.032633327,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.092461094,0.18492219,0.27738327,0.36984438,0.46230546,0.38978696,0.31726846,0.24474995,0.17223145,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.533011,0.93911463,1.3470312,1.7549478,2.1628644,1.7603867,1.357909,0.9554313,0.5529536,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.94092757,1.8292793,2.7194438,3.6096084,4.499773,3.8398547,3.1799364,2.520018,1.8600996,1.2001812,1.0424535,0.88472575,0.726998,0.56927025,0.41335547,1.9344311,3.4573197,4.9802084,6.5030966,8.024173,10.395528,12.76507,15.134612,17.505966,19.87551,16.026588,12.179482,8.3323765,4.4852695,0.63816285,0.69255173,0.7469406,0.8031424,0.8575313,0.9119202,0.76325727,0.61278135,0.46230546,0.31182957,0.16316663,0.25925365,0.35715362,0.4550536,0.5529536,0.6508536,0.52032024,0.38978696,0.25925365,0.13053331,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.29007402,0.5058166,0.7197462,0.9354887,1.1494182,1.7694515,2.3894846,3.009518,3.6295512,4.249584,3.8942437,3.540716,3.1853752,2.8300345,2.474694,2.0649643,1.6552348,1.2455053,0.83577573,0.42423326,0.34083697,0.25562772,0.17041849,0.08520924,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.06164073,0.12509441,0.18673515,0.25018883,0.31182957,0.3825351,0.45324063,0.52213323,0.59283876,0.66173136,2.3024626,3.9431937,5.582112,7.2228427,8.861761,9.012237,9.162713,9.313189,9.461852,9.612328,10.462607,11.312886,12.163166,13.011633,13.861912,13.930804,13.997884,14.064963,14.132043,14.199123,14.043208,13.885481,13.727753,13.5700245,13.412297,13.508384,13.602658,13.696932,13.793019,13.887294,15.8869915,17.888502,19.888199,21.887897,23.887594,21.768242,19.647076,17.527721,15.408369,13.287203,12.0145035,10.741803,9.469104,8.198216,6.925517,7.3352466,7.744976,8.154706,8.564435,8.974165,8.734854,8.495543,8.254418,8.015107,7.7757964,8.125698,8.4756,8.825501,9.175404,9.525306,10.489801,11.454298,12.420607,13.385102,14.349599,14.269829,14.190058,14.110288,14.030518,13.9507475,12.621845,11.294757,9.967669,8.640579,7.311678,6.6553855,5.99728,5.3391747,4.6828823,4.024777,3.3848011,2.7448254,2.1048496,1.4648738,0.824898,0.71430725,0.6055295,0.4949388,0.38434806,0.2755703,13.499319,13.261822,13.024323,12.786825,12.549327,12.311829,11.5503845,10.7871275,10.025683,9.262425,8.499168,7.9752226,7.4494634,6.925517,6.399758,5.8758116,6.5629244,7.250037,7.93715,8.624263,9.313189,10.462607,11.612025,12.763257,13.912675,15.062093,15.761897,16.4617,17.163317,17.863121,18.562923,15.23795,11.912977,8.588004,5.2630305,1.938057,1.9616255,1.987007,2.0123885,2.03777,2.0631514,1.7748904,1.4866294,1.2001812,0.9119202,0.62547207,1.0497054,1.4757515,1.8999848,2.324218,2.7502642,2.561716,2.374981,2.1882458,1.9996977,1.8129625,1.6751775,1.5373923,1.3996071,1.261822,1.1258497,1.0750868,1.0243238,0.97537386,0.9246109,0.87566096,0.85027945,0.824898,0.7995165,0.774135,0.7505665,1.2001812,1.649796,2.0994108,2.5508385,3.000453,3.5008307,3.9993954,4.499773,5.0001507,5.5005283,4.512464,3.5243993,2.5381477,1.550083,0.5620184,0.61278135,0.66173136,0.7124943,0.76325727,0.8122072,0.6744221,0.53663695,0.40066472,0.26287958,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.099712946,0.19942589,0.2991388,0.40066472,0.50037766,0.774135,1.0497054,1.3252757,1.6008459,1.8746033,1.5120108,1.1494182,0.7868258,0.42423326,0.06164073,0.16316663,0.26287958,0.36259252,0.46230546,0.5620184,0.44961473,0.33721104,0.22480737,0.11240368,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,2.3369088,4.550536,6.7623506,8.974165,11.187792,9.275117,7.362441,5.4497657,3.53709,1.6244144,2.5000753,3.3757362,4.249584,5.125245,6.000906,6.9490857,7.899078,8.8508835,9.800876,10.750868,9.96223,9.175404,8.386765,7.5999393,6.813113,6.9617763,7.112252,7.262728,7.413204,7.5618668,6.9744673,6.3870673,5.7996674,5.2122674,4.6248674,3.825351,3.0258346,2.2245052,1.4249886,0.62547207,2.811905,5.0001507,7.1883965,9.374829,11.563075,13.724127,15.8869915,18.049856,20.212719,22.375584,22.337511,22.29944,22.26318,22.22511,22.187037,18.024473,13.861912,9.699349,5.5367875,1.3742256,1.6751775,1.9743162,2.275268,2.5744069,2.8753586,2.4366217,1.9996977,1.5627737,1.1258497,0.6871128,0.5493277,0.41335547,0.2755703,0.13778515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.42423326,0.85027945,1.2745126,1.7005589,2.124792,3.2125697,4.3003473,5.388125,6.4759026,7.5618668,7.911769,8.26167,8.613385,8.963287,9.313189,9.811753,10.312131,10.812509,11.312886,11.813264,12.06164,12.311829,12.562017,12.812206,13.062395,12.60009,12.137785,11.675479,11.213174,10.750868,9.099259,7.4494634,5.7996674,4.1498713,2.5000753,2.7992141,3.100166,3.3993049,3.7002566,3.9993954,4.6375585,5.275721,5.9120708,6.550234,7.1883965,6.11331,5.038223,3.9631362,2.8880494,1.8129625,1.4630609,1.1131591,0.76325727,0.41335547,0.06164073,0.099712946,0.13778515,0.17585737,0.21211663,0.25018883,0.5620184,0.87566096,1.1874905,1.49932,1.8129625,1.550083,1.2872034,1.0243238,0.76325727,0.50037766,0.40066472,0.2991388,0.19942589,0.099712946,0.0,1.0750868,2.1501737,3.2252605,4.3003473,5.375434,4.9620786,4.550536,4.137181,3.7256382,3.3122826,2.8245957,2.3369088,1.8492218,1.3633479,0.87566096,0.9119202,0.9499924,0.9880646,1.0243238,1.062396,0.8883517,0.7124943,0.53663695,0.36259252,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.13778515,0.15047589,0.16316663,0.17585737,0.18673515,0.31182957,0.43692398,0.5620184,0.6871128,0.8122072,0.7868258,0.76325727,0.73787576,0.7124943,0.6871128,0.5747091,0.46230546,0.34990177,0.2374981,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.11240368,0.22480737,0.33721104,0.44961473,0.5620184,0.44961473,0.33721104,0.22480737,0.11240368,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.51306844,0.96268314,1.4122978,1.8619126,2.3133402,1.887294,1.4630609,1.0370146,0.61278135,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,1.1747998,2.2879589,3.3993049,4.512464,5.6256227,4.7245803,3.825351,2.9243085,2.0250793,1.1258497,0.93730164,0.7505665,0.5620184,0.37528324,0.18673515,2.03777,3.8869917,5.7380266,7.5872483,9.438283,12.212116,14.9877615,17.763407,20.537241,23.312885,18.800423,14.287958,9.775495,5.2630305,0.7505665,0.7124943,0.6744221,0.63816285,0.6000906,0.5620184,0.44961473,0.33721104,0.22480737,0.11240368,0.0,0.0870222,0.17585737,0.26287958,0.34990177,0.43692398,0.34990177,0.26287958,0.17585737,0.0870222,0.0,0.0,0.0,0.0,0.0,0.0,0.099712946,0.19942589,0.2991388,0.40066472,0.50037766,1.0007553,1.49932,1.9996977,2.5000753,3.000453,2.7375734,2.474694,2.2118144,1.9507477,1.6878681,1.3506571,1.0116332,0.6744221,0.33721104,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.099712946,0.19942589,0.2991388,0.40066472,0.50037766,2.0631514,3.6241121,5.186886,6.7496595,8.312433,8.511859,8.713099,8.912524,9.11195,9.313189,10.437225,11.563075,12.687112,13.812962,14.936998,14.663241,14.387671,14.112101,13.838344,13.562773,13.9507475,14.336908,14.724882,15.112856,15.50083,15.825351,16.14987,16.474392,16.800724,17.125244,19.59994,22.074633,24.549326,27.024021,29.500526,26.1121,22.725487,19.337059,15.950445,12.562017,11.287505,10.012992,8.736667,7.462154,6.187641,6.787732,7.3878226,7.987913,8.588004,9.188094,8.749357,8.312433,7.8755093,7.4367723,6.9998484,6.7496595,6.4994707,6.249282,6.000906,5.750717,7.462154,9.175404,10.88684,12.60009,14.313339,14.175554,14.037769,13.899984,13.762199,13.6244135,12.411542,11.200482,9.987611,8.774739,7.5618668,7.0125394,6.4632115,5.9120708,5.3627434,4.8116026,4.024777,3.2379513,2.4493124,1.6624867,0.87566096,0.7505665,0.62547207,0.50037766,0.37528324,0.25018883,13.874602,13.6244135,13.374225,13.125849,12.87566,12.625471,11.949236,11.274815,10.600392,9.924157,9.249735,8.584378,7.9208336,7.2554765,6.590119,5.924762,6.2927933,6.6608243,7.027043,7.3950744,7.763106,8.682278,9.603263,10.522435,11.4416065,12.362592,13.325275,14.287958,15.250641,16.213324,17.174194,14.282519,11.390844,8.497355,5.6056805,2.712192,2.514579,2.3169663,2.1193533,1.9217403,1.7241274,1.4902552,1.2545701,1.020698,0.7850128,0.5493277,0.95180535,1.3542831,1.7567607,2.1592383,2.561716,2.3767939,2.1918716,2.0069497,1.8220274,1.6371052,1.5319533,1.4268016,1.3216497,1.2183108,1.1131591,1.0406405,0.968122,0.89560354,0.823085,0.7505665,0.7433147,0.73424983,0.726998,0.7197462,0.7124943,1.0569572,1.403233,1.7476959,2.0921588,2.4366217,2.907992,3.3775494,3.8471067,4.3166637,4.788034,3.9377546,3.0874753,2.2371957,1.3869164,0.53663695,0.62728506,0.7179332,0.80676836,0.8974165,0.9880646,0.8575313,0.726998,0.5982776,0.46774435,0.33721104,0.27194437,0.20667773,0.14322405,0.07795739,0.012690738,0.05076295,0.0870222,0.12509441,0.16316663,0.19942589,0.19579996,0.19036107,0.18492219,0.1794833,0.17585737,0.13959812,0.10515183,0.07070554,0.034446288,0.0,0.07977036,0.15954071,0.23931105,0.3208944,0.40066472,0.6200332,0.83940166,1.0605831,1.2799516,1.49932,1.3270886,1.1548572,0.9826257,0.8103943,0.63816285,1.2291887,1.8220274,2.4148662,3.007705,3.6005437,2.955129,2.3097143,1.6642996,1.020698,0.37528324,0.33721104,0.2991388,0.26287958,0.22480737,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.027194439,0.054388877,0.08339628,0.11059072,0.13778515,1.9253663,3.7129474,5.5005283,7.28811,9.07569,7.520169,5.964647,4.409125,2.855416,1.2998942,1.9996977,2.6995013,3.3993049,4.099108,4.800725,6.1296263,7.460341,8.789243,10.119957,11.450671,10.460794,9.470917,8.479226,7.4893484,6.4994707,7.400513,8.299743,9.200785,10.100015,10.999244,9.817192,8.63514,7.453089,6.2692246,5.087173,5.185073,5.282973,5.3808727,5.47696,5.57486,6.3109226,7.0451727,7.7794223,8.515485,9.249735,11.022813,12.794077,14.567154,16.34023,18.11331,18.280102,18.446894,18.6155,18.782291,18.949085,15.5606575,12.170418,8.780178,5.389938,1.9996977,2.2408218,2.4801328,2.7194438,2.960568,3.199879,3.1182957,3.0348995,2.953316,2.8699198,2.7883365,2.2625773,1.7368182,1.2128719,0.6871128,0.16316663,0.15410182,0.14684997,0.13959812,0.13234627,0.12509441,0.12328146,0.11965553,0.11784257,0.11421664,0.11240368,0.10696479,0.10333887,0.09789998,0.092461094,0.0870222,0.07070554,0.052575916,0.034446288,0.018129626,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.4405499,0.8665961,1.2944553,1.7223145,2.1501737,2.9297476,3.7093215,4.4907084,5.2702823,6.049856,6.338117,6.624565,6.9128265,7.1992745,7.4875355,7.995165,8.502794,9.010424,9.518054,10.025683,10.130835,10.234174,10.339326,10.444477,10.549629,10.230548,9.909654,9.590572,9.269678,8.950596,7.6380115,6.3254266,5.0128417,3.7002566,2.3876717,2.5508385,2.712192,2.8753586,3.0367124,3.199879,3.7093215,4.220577,4.7300196,5.239462,5.750717,4.88956,4.0302157,3.1690586,2.3097143,1.4503701,1.1766127,0.90466833,0.6327239,0.36077955,0.0870222,0.11059072,0.13234627,0.15410182,0.17767033,0.19942589,0.47680917,0.7541924,1.0333886,1.310772,1.5881553,1.3977941,1.2074331,1.017072,0.82671094,0.63816285,0.67986095,0.72337204,0.7650702,0.80676836,0.85027945,1.9453088,3.0403383,4.135368,5.230397,6.3254266,5.77066,5.2158933,4.6593137,4.1045475,3.5497808,3.0167696,2.4855716,1.9525607,1.4195497,0.8883517,0.89560354,0.90285534,0.9101072,0.91735905,0.9246109,0.79226464,0.65991837,0.5275721,0.39522585,0.26287958,0.21574254,0.16679256,0.11965553,0.072518505,0.025381476,0.03988518,0.054388877,0.07070554,0.08520924,0.099712946,0.11421664,0.13053331,0.14503701,0.15954071,0.17585737,0.27194437,0.36984438,0.46774435,0.5656443,0.66173136,0.6544795,0.64722764,0.6399758,0.6327239,0.62547207,0.5493277,0.4749962,0.40066472,0.3245203,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.11965553,0.2030518,0.28463513,0.3680314,0.44961473,0.36077955,0.27013144,0.1794833,0.09064813,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.40972954,0.7705091,1.1294757,1.4902552,1.8492218,1.5101979,1.1693609,0.83033687,0.4894999,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.018129626,0.034446288,0.052575916,0.07070554,0.0870222,1.1893034,2.2915847,3.395679,4.49796,5.600241,4.710077,3.8199122,2.9297476,2.039583,1.1494182,1.1693609,1.1893034,1.209246,1.2291887,1.2491312,3.4518807,5.65463,7.85738,10.060129,12.262879,14.447499,16.632118,18.816738,21.003172,23.187792,18.809486,14.432995,10.05469,5.678199,1.2998942,1.1294757,0.96087015,0.7904517,0.6200332,0.44961473,0.36077955,0.27013144,0.1794833,0.09064813,0.0,0.072518505,0.14503701,0.21755551,0.29007402,0.36259252,0.2955129,0.22662032,0.15954071,0.092461094,0.025381476,0.02175555,0.01994259,0.018129626,0.014503701,0.012690738,0.09064813,0.16679256,0.24474995,0.32270733,0.40066472,0.7995165,1.2001812,1.6008459,1.9996977,2.4003625,2.1991236,1.9996977,1.8002719,1.6008459,1.3996071,1.1204109,0.83940166,0.56020546,0.27919623,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.11421664,0.23024625,0.3444629,0.4604925,0.5747091,1.887294,3.199879,4.512464,5.825049,7.137634,7.817495,8.497355,9.177217,9.857078,10.536939,11.439794,12.342649,13.245504,14.146547,15.049402,14.973258,14.895301,14.817343,14.739386,14.663241,15.31772,15.9722,16.62668,17.282972,17.937452,17.7344,17.533161,17.330109,17.127058,16.92582,18.265598,19.605377,20.945156,22.284937,23.624716,21.347635,19.06874,16.79166,14.514579,12.237497,11.780631,11.321951,10.865085,10.408218,9.949538,9.452786,8.954222,8.457471,7.9607186,7.462154,7.322556,7.1829576,7.0433598,6.9019485,6.7623506,6.5230393,6.281915,6.0426044,5.803293,5.562169,7.1430726,8.722163,10.303066,11.882156,13.46306,13.113158,12.763257,12.413355,12.06164,11.711739,10.680162,9.646774,8.615198,7.5818095,6.550234,7.518356,8.484665,9.452786,10.420909,11.3872175,10.065568,8.7421055,7.420456,6.096993,4.7753434,4.4508233,4.12449,3.7999697,3.4754493,3.150929,14.249886,13.987006,13.724127,13.46306,13.200181,12.937301,12.349901,11.762501,11.175101,10.587702,10.000301,9.195346,8.39039,7.5854354,6.78048,5.975525,6.0226617,6.069799,6.1169357,6.165886,6.2130227,6.9019485,7.592687,8.281613,8.972352,9.663091,10.88684,12.112403,13.337966,14.561715,15.787278,13.327088,10.866898,8.406708,5.9483304,3.48814,3.0675328,2.6469254,2.228131,1.8075237,1.3869164,1.2056202,1.0225109,0.83940166,0.65810543,0.4749962,0.8557183,1.2346275,1.6153497,1.9942589,2.374981,2.1918716,2.0105755,1.8274662,1.6443571,1.4630609,1.3905423,1.3180238,1.2455053,1.1729867,1.1004683,1.0043813,0.9101072,0.81583315,0.7197462,0.62547207,0.6345369,0.64541465,0.6544795,0.6653573,0.6744221,0.9155461,1.1548572,1.3941683,1.6352923,1.8746033,2.3151531,2.7557032,3.1944401,3.63499,4.07554,3.3630457,2.6505513,1.938057,1.2255627,0.51306844,0.6417888,0.77232206,0.90285534,1.0333886,1.162109,1.0406405,0.91735905,0.79589057,0.6726091,0.5493277,0.44417584,0.34083697,0.23568514,0.13053331,0.025381476,0.07433146,0.12509441,0.17585737,0.22480737,0.2755703,0.29007402,0.3045777,0.3208944,0.33539808,0.34990177,0.27919623,0.21030366,0.13959812,0.07070554,0.0,0.059827764,0.11965553,0.1794833,0.23931105,0.2991388,0.46411842,0.629098,0.79589057,0.96087015,1.1258497,1.1421664,1.1602961,1.1766127,1.1947423,1.2128719,2.2970235,3.3829882,4.4671397,5.5531044,6.637256,5.4606433,4.2822175,3.105605,1.9271792,0.7505665,0.6744221,0.6000906,0.52575916,0.44961473,0.37528324,0.2991388,0.22480737,0.15047589,0.07433146,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,1.5120108,2.8753586,4.2368937,5.600241,6.9617763,5.765221,4.5668526,3.3702974,2.1719291,0.97537386,1.49932,2.0250793,2.5508385,3.0747845,3.6005437,5.3101673,7.019791,8.729415,10.440851,12.1504755,10.957546,9.764616,8.571687,7.380571,6.187641,7.837437,9.487233,11.137029,12.786825,14.436621,12.659918,10.883214,9.104698,7.327995,5.5494785,6.544795,7.5401115,8.535428,9.530745,10.524248,9.808127,9.090195,8.372261,7.654328,6.9382076,8.319685,9.702975,11.084454,12.467744,13.849221,14.222692,14.594349,14.967819,15.339477,15.712947,13.095029,10.477111,7.859193,5.243088,2.6251698,2.8046532,2.9841363,3.1654327,3.3449159,3.5243993,3.7981565,4.070101,4.3420453,4.615803,4.8877473,3.975827,3.0620937,2.1501737,1.2382535,0.3245203,0.3100166,0.2955129,0.27919623,0.26469254,0.25018883,0.24474995,0.23931105,0.23568514,0.23024625,0.22480737,0.21574254,0.20486477,0.19579996,0.18492219,0.17585737,0.13959812,0.10515183,0.07070554,0.034446288,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.4550536,0.88472575,1.3143979,1.745883,2.175555,2.6469254,3.1201086,3.5932918,4.064662,4.537845,4.762653,4.98746,5.2122674,5.4370747,5.661882,6.1767635,6.6916447,7.208339,7.723221,8.238102,8.198216,8.158332,8.116633,8.076748,8.036863,7.859193,7.6833353,7.5056653,7.327995,7.1503243,6.1749506,5.199577,4.2242026,3.2506418,2.275268,2.3006494,2.324218,2.3495996,2.374981,2.4003625,2.7828975,3.1654327,3.5479677,3.930503,4.313038,3.6676233,3.0222087,2.3767939,1.7331922,1.0877775,0.8919776,0.6979906,0.50219065,0.30820364,0.11240368,0.11965553,0.12690738,0.13415924,0.14322405,0.15047589,0.39159992,0.6345369,0.8774739,1.1204109,1.3633479,1.2455053,1.1276628,1.0098201,0.8919776,0.774135,0.96087015,1.1457924,1.3307146,1.5156367,1.7005589,2.8155308,3.930503,5.045475,6.1604466,7.2754188,6.5774283,5.8794374,5.18326,4.4852695,3.787279,3.2107568,2.6324217,2.0540867,1.4775645,0.89922947,0.8774739,0.8557183,0.8321498,0.8103943,0.7868258,0.6979906,0.6073425,0.5166943,0.42785916,0.33721104,0.27919623,0.2229944,0.16497959,0.10696479,0.05076295,0.054388877,0.059827764,0.065266654,0.07070554,0.07433146,0.092461094,0.11059072,0.12690738,0.14503701,0.16316663,0.23205921,0.30276474,0.37165734,0.44236287,0.51306844,0.52213323,0.533011,0.5420758,0.5529536,0.5620184,0.52575916,0.48768693,0.44961473,0.41335547,0.37528324,0.2991388,0.22480737,0.15047589,0.07433146,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.12690738,0.1794833,0.23205921,0.28463513,0.33721104,0.27013144,0.2030518,0.13415924,0.06707962,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.30820364,0.57833505,0.8466535,1.1167849,1.3869164,1.1331016,0.8774739,0.62184614,0.3680314,0.11240368,0.09064813,0.06707962,0.045324065,0.02175555,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,1.2056202,2.2970235,3.39024,4.4816437,5.57486,4.695573,3.8144734,2.9351864,2.0540867,1.1747998,1.403233,1.6298534,1.8582866,2.084907,2.3133402,4.8678045,7.422269,9.976733,12.5330105,15.087475,16.682882,18.278288,19.871883,21.46729,23.062696,18.820364,14.5780325,10.3357,6.091554,1.8492218,1.54827,1.2455053,0.94274056,0.6399758,0.33721104,0.27013144,0.2030518,0.13415924,0.06707962,0.0,0.058014803,0.11421664,0.17223145,0.23024625,0.28826106,0.23931105,0.19217403,0.14503701,0.09789998,0.05076295,0.045324065,0.03988518,0.034446288,0.030820364,0.025381476,0.07977036,0.13415924,0.19036107,0.24474995,0.2991388,0.6000906,0.89922947,1.2001812,1.49932,1.8002719,1.6624867,1.5247015,1.3869164,1.2491312,1.1131591,0.8901646,0.6671702,0.44417584,0.2229944,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13053331,0.25925365,0.38978696,0.52032024,0.6508536,1.7132497,2.7756457,3.8380418,4.900438,5.962834,7.12313,8.281613,9.441909,10.602205,11.762501,12.442362,13.122223,13.802084,14.481945,15.161806,15.283275,15.40293,15.522586,15.6422415,15.761897,16.684694,17.607492,18.53029,19.453089,20.375887,19.645262,18.914639,18.185827,17.455204,16.72458,16.929445,17.13431,17.339174,17.545853,17.750717,16.583168,15.415621,14.248073,13.080525,11.912977,12.271944,12.632723,12.99169,13.352469,13.713249,12.117842,10.522435,8.927028,7.3334336,5.7380266,5.8957543,6.051669,6.209397,6.3671246,6.5248523,6.294606,6.0643597,5.8341136,5.6056805,5.375434,6.8221784,8.270736,9.71748,11.164224,12.612781,12.050762,11.486931,10.924912,10.362894,9.800876,8.94697,8.094878,7.2427855,6.390693,5.5367875,8.02236,10.507931,12.993503,15.477262,17.962833,16.104548,14.248073,12.389787,10.533313,8.675026,8.149267,7.6253204,7.0995617,6.5756154,6.049856,14.625169,14.349599,14.075842,13.800271,13.524701,13.24913,12.750566,12.250188,11.74981,11.249433,10.750868,9.804502,8.859948,7.915395,6.970841,6.0244746,5.75253,5.480586,5.2068286,4.934884,4.6629395,5.121619,5.582112,6.0426044,6.5030966,6.9617763,8.450218,9.936848,11.42529,12.91192,14.400362,12.371656,10.344765,8.317872,6.2891674,4.262275,3.6204863,2.9768846,2.335096,1.693307,1.0497054,0.91917205,0.7904517,0.65991837,0.5293851,0.40066472,0.75781834,1.114972,1.4721256,1.8292793,2.1882458,2.0069497,1.8274662,1.647983,1.4666867,1.2872034,1.2473183,1.2074331,1.167548,1.1276628,1.0877775,0.969935,0.8520924,0.73424983,0.61822027,0.50037766,0.5275721,0.55476654,0.581961,0.6091554,0.63816285,0.77232206,0.90829426,1.0424535,1.1766127,1.3125849,1.7223145,2.132044,2.5417736,2.953316,3.3630457,2.7883365,2.2118144,1.6371052,1.062396,0.48768693,0.65810543,0.82671094,0.99712944,1.167548,1.3379664,1.2219368,1.1077201,0.9916905,0.8774739,0.76325727,0.61822027,0.47318324,0.32814622,0.18310922,0.038072214,0.099712946,0.16316663,0.22480737,0.28826106,0.34990177,0.38434806,0.42060733,0.4550536,0.4894999,0.52575916,0.42060733,0.3154555,0.21030366,0.10515183,0.0,0.03988518,0.07977036,0.11965553,0.15954071,0.19942589,0.3100166,0.42060733,0.5293851,0.6399758,0.7505665,0.9572442,1.1657349,1.3724127,1.5809034,1.7875811,3.3648586,4.942136,6.5194135,8.096691,9.675781,7.9643445,6.2547207,4.5450974,2.8354735,1.1258497,1.0116332,0.89922947,0.7868258,0.6744221,0.5620184,0.44961473,0.33721104,0.22480737,0.11240368,0.0,0.032633327,0.065266654,0.09789998,0.13053331,0.16316663,1.1004683,2.03777,2.9750717,3.9123733,4.8496747,4.0102735,3.1708715,2.3296568,1.4902552,0.6508536,1.0007553,1.3506571,1.7005589,2.0504606,2.4003625,4.4907084,6.5792413,8.669587,10.7599325,12.850279,11.454298,10.060129,8.664148,7.26998,5.8758116,8.274362,10.674724,13.075087,15.475449,17.87581,15.502643,13.129475,10.75812,8.384952,6.011784,7.9045167,9.79725,11.689982,13.582716,15.475449,13.305332,11.135216,8.9651,6.794984,4.6248674,5.618371,6.6100616,7.6017523,8.595256,9.5869465,10.165281,10.741803,11.320138,11.896661,12.474996,10.629399,8.785617,6.9400206,5.0944247,3.2506418,3.3702974,3.489953,3.6096084,3.729264,3.8507326,4.478018,5.105303,5.732588,6.359873,6.987158,5.6872635,4.3873696,3.0874753,1.7875811,0.48768693,0.46411842,0.44236287,0.42060733,0.39703882,0.37528324,0.3680314,0.36077955,0.35171473,0.3444629,0.33721104,0.32270733,0.30820364,0.291887,0.27738327,0.26287958,0.21030366,0.15772775,0.10515183,0.052575916,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.46955732,0.90285534,1.3343405,1.7676386,2.1991236,2.3641033,2.5308957,2.6958754,2.8608549,3.0258346,3.1871881,3.350355,3.5117085,3.6748753,3.8380418,4.360175,4.882308,5.4044414,5.9283876,6.450521,6.265599,6.0806766,5.8957543,5.710832,5.52591,5.4896507,5.4552045,5.4207582,5.384499,5.3500524,4.7118897,4.07554,3.437377,2.7992141,2.1628644,2.0504606,1.938057,1.8256533,1.7132497,1.6008459,1.8546607,2.1102884,2.3659163,2.619731,2.8753586,2.4456866,2.0142014,1.5845293,1.1548572,0.72518504,0.6073425,0.4894999,0.37165734,0.25562772,0.13778515,0.13053331,0.12328146,0.11421664,0.10696479,0.099712946,0.30820364,0.5148814,0.72337204,0.9300498,1.1367276,1.0932164,1.0478923,1.0025684,0.9572442,0.9119202,1.2400664,1.5682126,1.8945459,2.222692,2.5508385,3.6857529,4.8206677,5.955582,7.0904965,8.225411,7.3841968,6.544795,5.7053933,4.8641787,4.024777,3.4029307,2.7792716,2.1574254,1.5355793,0.9119202,0.85934424,0.80676836,0.7541924,0.7016165,0.6508536,0.60190356,0.55476654,0.5076295,0.4604925,0.41335547,0.3444629,0.27738327,0.21030366,0.14322405,0.07433146,0.07070554,0.065266654,0.059827764,0.054388877,0.05076295,0.07070554,0.09064813,0.11059072,0.13053331,0.15047589,0.19217403,0.23568514,0.27738327,0.3208944,0.36259252,0.38978696,0.4169814,0.44417584,0.47318324,0.50037766,0.50037766,0.50037766,0.50037766,0.50037766,0.50037766,0.40066472,0.2991388,0.19942589,0.099712946,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.13415924,0.15772775,0.1794833,0.2030518,0.22480737,0.1794833,0.13415924,0.09064813,0.045324065,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.20486477,0.38434806,0.5656443,0.7451276,0.9246109,0.7541924,0.5855869,0.41516843,0.24474995,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.027194439,0.054388877,0.08339628,0.11059072,0.13778515,1.2201238,2.3024626,3.3848011,4.4671397,5.5494785,4.6792564,3.8108473,2.9406252,2.0704033,1.2001812,1.6352923,2.0704033,2.5055144,2.9406252,3.3757362,6.281915,9.189907,12.097899,15.005891,17.912071,18.918264,19.922646,20.927027,21.933222,22.937603,18.82943,14.723069,10.614896,6.506723,2.4003625,1.9652514,1.5301404,1.0950294,0.65991837,0.22480737,0.1794833,0.13415924,0.09064813,0.045324065,0.0,0.04169814,0.08520924,0.12690738,0.17041849,0.21211663,0.18492219,0.15772775,0.13053331,0.10333887,0.07433146,0.06707962,0.059827764,0.052575916,0.045324065,0.038072214,0.07070554,0.10333887,0.13415924,0.16679256,0.19942589,0.40066472,0.6000906,0.7995165,1.0007553,1.2001812,1.1258497,1.0497054,0.97537386,0.89922947,0.824898,0.65991837,0.4949388,0.32995918,0.16497959,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14503701,0.29007402,0.43511102,0.58014804,0.72518504,1.5373923,2.3495996,3.1618068,3.975827,4.788034,6.4269524,8.067683,9.708415,11.347333,12.988064,13.44493,13.901797,14.3604765,14.817343,15.27421,15.593291,15.91056,16.227829,16.545097,16.862366,18.051668,19.242785,20.432089,21.623205,22.812508,21.554312,20.29793,19.039734,17.78335,16.525154,15.595104,14.665054,13.735004,12.804955,11.874905,11.81689,11.760688,11.702674,11.644659,11.586644,12.76507,13.943495,15.120108,16.29672,17.475147,14.782897,12.088835,9.396585,6.7043357,4.0120864,4.4671397,4.9221935,5.377247,5.8323007,6.2873545,6.0679855,5.846804,5.6274357,5.408067,5.186886,6.5030966,7.817495,9.131892,10.448103,11.762501,10.988366,10.212419,9.438283,8.662335,7.8882003,7.215591,6.542982,5.870373,5.197764,4.5251546,8.528176,12.531198,16.532406,20.535427,24.536636,22.145338,19.752228,17.359118,14.967819,12.574709,11.849524,11.124338,10.399154,9.675781,8.950596,15.000452,14.712192,14.425743,14.137483,13.849221,13.562773,13.149418,12.737875,12.32452,11.912977,11.499621,10.41547,9.329506,8.245354,7.159389,6.0752378,5.482399,4.88956,4.2967215,3.7056956,3.1128569,3.343103,3.5733492,3.8017826,4.0320287,4.262275,6.011784,7.763106,9.512614,11.262123,13.011633,11.418038,9.822631,8.227224,6.6318173,5.038223,4.171627,3.3068438,2.4420607,1.5772774,0.7124943,0.6345369,0.55839247,0.48043507,0.40247768,0.3245203,0.65991837,0.99531645,1.3307146,1.6642996,1.9996977,1.8220274,1.6443571,1.4666867,1.2908293,1.1131591,1.1040943,1.0968424,1.0895905,1.0823387,1.0750868,0.9354887,0.79589057,0.6544795,0.5148814,0.37528324,0.42060733,0.46411842,0.5094425,0.55476654,0.6000906,0.629098,0.65991837,0.69073874,0.7197462,0.7505665,1.1294757,1.5101979,1.889107,2.269829,2.6505513,2.2118144,1.7748904,1.3379664,0.89922947,0.46230546,0.6726091,0.88291276,1.0932164,1.3017071,1.5120108,1.405046,1.2980812,1.1893034,1.0823387,0.97537386,0.7904517,0.6055295,0.42060733,0.23568514,0.05076295,0.12509441,0.19942589,0.2755703,0.34990177,0.42423326,0.48043507,0.53482395,0.58921283,0.64541465,0.69980353,0.56020546,0.42060733,0.27919623,0.13959812,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.15410182,0.21030366,0.26469254,0.3208944,0.37528324,0.77232206,1.1693609,1.5682126,1.9652514,2.3622901,4.4326935,6.5030966,8.5735,10.642091,12.712494,10.469859,8.227224,5.9845896,3.7419548,1.49932,1.3506571,1.2001812,1.0497054,0.89922947,0.7505665,0.6000906,0.44961473,0.2991388,0.15047589,0.0,0.034446288,0.07070554,0.10515183,0.13959812,0.17585737,0.6871128,1.2001812,1.7132497,2.2245052,2.7375734,2.2553256,1.7730774,1.2908293,0.80676836,0.3245203,0.50037766,0.6744221,0.85027945,1.0243238,1.2001812,3.6694362,6.1405044,8.609759,11.080828,13.550082,11.952863,10.355642,8.756609,7.159389,5.562169,8.713099,11.862214,15.013144,18.16226,21.313189,18.345367,15.377548,12.409729,9.441909,6.4759026,9.264238,12.054388,14.844538,17.634687,20.424837,16.802538,13.180238,9.557939,5.9356394,2.3133402,2.9152439,3.5171473,4.120864,4.7227674,5.3246713,6.107871,6.889258,7.6724577,8.455658,9.237044,8.165584,7.0923095,6.0208488,4.947575,3.874301,3.9341288,3.9957695,4.0555973,4.115425,4.175253,5.1578784,6.1405044,7.12313,8.105756,9.088382,7.400513,5.712645,4.024777,2.3369088,0.6508536,0.6200332,0.58921283,0.56020546,0.5293851,0.50037766,0.4894999,0.48043507,0.46955732,0.4604925,0.44961473,0.42967212,0.40972954,0.38978696,0.36984438,0.34990177,0.27919623,0.21030366,0.13959812,0.07070554,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.48587397,0.91917205,1.3542831,1.789394,2.2245052,2.0830941,1.93987,1.7966459,1.6552348,1.5120108,1.6117238,1.7132497,1.8129625,1.9126755,2.0123885,2.5417736,3.0729716,3.6023567,4.1317415,4.6629395,4.3329806,4.0030212,3.673062,3.343103,3.0131438,3.1201086,3.2270734,3.3358512,3.442816,3.5497808,3.2506418,2.94969,2.6505513,2.3495996,2.0504606,1.8002719,1.550083,1.2998942,1.0497054,0.7995165,0.92823684,1.0551442,1.1820517,1.310772,1.4376793,1.2219368,1.0080072,0.79226464,0.57833505,0.36259252,0.32270733,0.28282216,0.24293698,0.2030518,0.16316663,0.13959812,0.11784257,0.09427405,0.072518505,0.05076295,0.2229944,0.39522585,0.56745726,0.73968875,0.9119202,0.93911463,0.968122,0.99531645,1.0225109,1.0497054,1.5192627,1.9906329,2.4601903,2.9297476,3.3993049,4.555975,5.710832,6.8656893,8.020547,9.175404,8.192778,7.210152,6.2275267,5.2449007,4.262275,3.5951047,2.9279346,2.2607644,1.5917811,0.9246109,0.8430276,0.75963134,0.678048,0.5946517,0.51306844,0.5076295,0.50219065,0.49675176,0.49312583,0.48768693,0.40972954,0.33177215,0.25562772,0.17767033,0.099712946,0.08520924,0.07070554,0.054388877,0.03988518,0.025381476,0.047137026,0.07070554,0.092461094,0.11421664,0.13778515,0.15228885,0.16679256,0.18310922,0.19761293,0.21211663,0.2574407,0.30276474,0.3480888,0.39159992,0.43692398,0.4749962,0.51306844,0.5493277,0.5873999,0.62547207,0.50037766,0.37528324,0.25018883,0.12509441,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.14322405,0.13415924,0.12690738,0.11965553,0.11240368,0.09064813,0.06707962,0.045324065,0.02175555,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.10333887,0.19217403,0.28282216,0.37165734,0.46230546,0.3770962,0.291887,0.20667773,0.12328146,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.032633327,0.065266654,0.09789998,0.13053331,0.16316663,1.2346275,2.3079014,3.3793623,4.4526362,5.524097,4.664753,3.8054085,2.9442513,2.084907,1.2255627,1.8673514,2.5091403,3.152742,3.7945306,4.4381323,7.6978393,10.957546,14.217253,17.47696,20.736666,21.151834,21.567003,21.982172,22.397339,22.812508,18.840307,14.868106,10.894093,6.921891,2.94969,2.382233,1.8147756,1.2473183,0.67986095,0.11240368,0.09064813,0.06707962,0.045324065,0.02175555,0.0,0.027194439,0.054388877,0.08339628,0.11059072,0.13778515,0.13053331,0.12328146,0.11421664,0.10696479,0.099712946,0.09064813,0.07977036,0.07070554,0.059827764,0.05076295,0.059827764,0.07070554,0.07977036,0.09064813,0.099712946,0.19942589,0.2991388,0.40066472,0.50037766,0.6000906,0.5873999,0.5747091,0.5620184,0.5493277,0.53663695,0.42967212,0.32270733,0.21574254,0.10696479,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.15954071,0.3208944,0.48043507,0.6399758,0.7995165,1.3633479,1.9253663,2.4873846,3.049403,3.6132345,5.732588,7.851941,9.973107,12.092461,14.211814,14.447499,14.683184,14.917056,15.152741,15.386614,15.903308,16.41819,16.933071,17.447952,17.962833,19.420456,20.878077,22.3357,23.793322,25.250942,23.465176,21.679407,19.89545,18.109684,16.325727,14.25895,12.193986,10.129022,8.06587,5.999093,7.0524244,8.105756,9.157274,10.210606,11.262123,13.258195,15.252454,17.246714,19.242785,21.237043,17.447952,13.657047,9.867955,6.0770507,2.2879589,3.0403383,3.7927177,4.5450974,5.297477,6.049856,5.8395524,5.6292486,5.4207582,5.2104545,5.0001507,6.1822023,7.364254,8.548119,9.73017,10.912222,9.924157,8.937905,7.949841,6.9617763,5.975525,5.482399,4.989273,4.49796,4.004834,3.5117085,9.03218,14.55265,20.073122,25.59178,31.112251,28.184317,25.256382,22.33026,19.402325,16.474392,15.54978,14.625169,13.700559,12.775948,11.849524,15.375735,15.074784,14.775645,14.474693,14.175554,13.874602,13.550082,13.225562,12.899229,12.574709,12.250188,11.024626,9.800876,8.575313,7.3497505,6.1241875,5.2122674,4.3003473,3.386614,2.474694,1.5627737,1.5627737,1.5627737,1.5627737,1.5627737,1.5627737,3.5751622,5.5875506,7.5999393,9.612328,11.624716,10.462607,9.300498,8.136576,6.9744673,5.812358,4.7245803,3.636803,2.5508385,1.4630609,0.37528324,0.34990177,0.3245203,0.2991388,0.2755703,0.25018883,0.5620184,0.87566096,1.1874905,1.49932,1.8129625,1.6371052,1.4630609,1.2872034,1.1131591,0.93730164,0.96268314,0.9880646,1.0116332,1.0370146,1.062396,0.89922947,0.73787576,0.5747091,0.41335547,0.25018883,0.31182957,0.37528324,0.43692398,0.50037766,0.5620184,0.48768693,0.41335547,0.33721104,0.26287958,0.18673515,0.53663695,0.8883517,1.2382535,1.5881553,1.938057,1.6371052,1.3379664,1.0370146,0.73787576,0.43692398,0.6871128,0.93730164,1.1874905,1.4376793,1.6878681,1.5881553,1.4866294,1.3869164,1.2872034,1.1874905,0.96268314,0.73787576,0.51306844,0.28826106,0.06164073,0.15047589,0.2374981,0.3245203,0.41335547,0.50037766,0.5747091,0.6508536,0.72518504,0.7995165,0.87566096,0.69980353,0.52575916,0.34990177,0.17585737,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.5873999,1.1747998,1.7621996,2.3495996,2.9369993,5.5005283,8.062244,10.625773,13.1874895,15.749206,12.975373,10.199727,7.424082,4.650249,1.8746033,1.6878681,1.49932,1.3125849,1.1258497,0.93730164,0.7505665,0.5620184,0.37528324,0.18673515,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.2755703,0.36259252,0.44961473,0.53663695,0.62547207,0.50037766,0.37528324,0.25018883,0.12509441,0.0,0.0,0.0,0.0,0.0,0.0,2.8499773,5.6999545,8.549932,11.399909,14.249886,12.449615,10.649343,8.849071,7.0506115,5.2503395,9.1500225,13.049705,16.949387,20.850883,24.750565,21.188093,17.625622,14.06315,10.500679,6.9382076,10.625773,14.311526,18.000906,21.686659,25.374224,20.299742,15.22526,10.148965,5.0744824,0.0,0.21211663,0.42423326,0.63816285,0.85027945,1.062396,2.0504606,3.0367124,4.024777,5.0128417,6.000906,5.6999545,5.4008155,5.0998635,4.800725,4.499773,4.499773,4.499773,4.499773,4.499773,4.499773,5.8377395,7.175706,8.511859,9.849826,11.187792,9.11195,7.037921,4.9620786,2.8880494,0.8122072,0.774135,0.73787576,0.69980353,0.66173136,0.62547207,0.61278135,0.6000906,0.5873999,0.5747091,0.5620184,0.53663695,0.51306844,0.48768693,0.46230546,0.43692398,0.34990177,0.26287958,0.17585737,0.0870222,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.50037766,0.93730164,1.3742256,1.8129625,2.2498865,1.8002719,1.3506571,0.89922947,0.44961473,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.72518504,1.261822,1.8002719,2.3369088,2.8753586,2.4003625,1.9253663,1.4503701,0.97537386,0.50037766,0.7505665,1.0007553,1.2491312,1.49932,1.7495089,1.7875811,1.8256533,1.8619126,1.8999848,1.938057,1.550083,1.162109,0.774135,0.387974,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.13778515,0.2755703,0.41335547,0.5493277,0.6871128,0.7868258,0.8883517,0.9880646,1.0877775,1.1874905,1.8002719,2.4130533,3.0258346,3.636803,4.249584,5.424384,6.599184,7.7757964,8.950596,10.125396,8.999546,7.8755093,6.7496595,5.6256227,4.499773,3.787279,3.0747845,2.3622901,1.649796,0.93730164,0.824898,0.7124943,0.6000906,0.48768693,0.37528324,0.41335547,0.44961473,0.48768693,0.52575916,0.5620184,0.4749962,0.387974,0.2991388,0.21211663,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.12509441,0.18673515,0.25018883,0.31182957,0.37528324,0.44961473,0.52575916,0.6000906,0.6744221,0.7505665,0.6000906,0.44961473,0.2991388,0.15047589,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,1.2509441,2.3133402,3.3757362,4.4381323,5.5005283,4.650249,3.7999697,2.94969,2.0994108,1.2491312,2.0994108,2.94969,3.7999697,4.650249,5.5005283,9.11195,12.725184,16.338419,19.94984,23.563074,23.387217,23.213173,23.037315,22.863272,22.687414,18.849373,15.013144,11.175101,7.3370595,3.5008307,2.7992141,2.0994108,1.3996071,0.69980353,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.17585737,0.34990177,0.52575916,0.69980353,0.87566096,1.1874905,1.49932,1.8129625,2.124792,2.4366217,5.038223,7.6380115,10.2378,12.837588,15.437376,15.4500675,15.462758,15.475449,15.488139,15.50083,16.213324,16.92582,17.638313,18.350807,19.063301,20.78743,22.511557,24.237497,25.961624,27.687565,25.374224,23.062696,20.749357,18.43783,16.124489,12.92461,9.724731,6.5248523,3.3249733,0.12509441,2.2879589,4.4508233,6.6118746,8.774739,10.937603,13.749508,16.563227,19.375132,22.187037,25.000753,20.113007,15.22526,10.337513,5.4497657,0.5620184,1.6117238,2.663242,3.7129474,4.762653,5.812358,5.612932,5.411693,5.2122674,5.0128417,4.8116026,5.863121,6.9128265,7.9625316,9.012237,10.061942,8.861761,7.66158,6.4632115,5.2630305,4.062849,3.7492065,3.437377,3.1255474,2.811905,2.5000753,9.537996,16.575916,23.612024,30.649946,37.687866,34.22511,30.762348,27.299591,23.836832,20.375887,19.250036,18.124187,17.00015,15.8743,14.750263,16.187943,15.71476,15.243389,14.770206,14.297023,13.825653,13.657047,13.490254,13.321649,13.154857,12.988064,12.019942,11.05182,10.085511,9.117389,8.149267,6.9907837,5.8304877,4.670192,3.5098956,2.3495996,2.2118144,2.0758421,1.938057,1.8002719,1.6624867,3.2597067,4.856927,6.454147,8.05318,9.6504,8.821876,7.995165,7.166641,6.33993,5.5132194,4.5632267,3.6132345,2.663242,1.7132497,0.76325727,0.7124943,0.66173136,0.61278135,0.5620184,0.51306844,0.72337204,0.9318628,1.1421664,1.35247,1.5627737,1.5101979,1.4576219,1.405046,1.35247,1.2998942,1.2128719,1.1258497,1.0370146,0.9499924,0.8629702,0.7650702,0.6671702,0.56927025,0.47318324,0.37528324,0.40972954,0.44417584,0.48043507,0.5148814,0.5493277,0.46955732,0.38978696,0.3100166,0.23024625,0.15047589,0.43329805,0.71430725,0.99712944,1.2799516,1.5627737,1.4376793,1.3125849,1.1874905,1.062396,0.93730164,1.1258497,1.3125849,1.49932,1.6878681,1.8746033,1.7295663,1.5845293,1.4394923,1.2944553,1.1494182,0.94274056,0.73424983,0.5275721,0.3208944,0.11240368,0.23568514,0.35715362,0.48043507,0.60190356,0.72518504,0.73968875,0.7541924,0.7705091,0.7850128,0.7995165,0.6399758,0.48043507,0.3208944,0.15954071,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.6852999,1.3705997,2.0558996,2.7393866,3.4246864,5.282973,7.1394467,8.997733,10.854207,12.712494,10.924912,9.137331,7.3497505,5.562169,3.774588,3.6531196,3.529838,3.4083695,3.2850883,3.1618068,3.2597067,3.3576066,3.4555066,3.5534067,3.6494937,3.4500678,3.2506418,3.049403,2.8499773,2.6505513,2.2408218,1.8292793,1.4195497,1.0098201,0.6000906,3.7727752,6.94546,10.118144,13.290829,16.463512,13.172986,9.882459,6.591932,3.303218,0.012690738,2.5798457,5.147001,7.7141557,10.283124,12.850279,11.483305,10.114518,8.747544,7.380571,6.011784,8.898021,11.782444,14.666867,17.553104,20.437527,18.093367,15.747393,13.403233,11.057259,8.713099,11.648285,14.581658,17.516844,20.45203,23.387217,19.4549,15.522586,11.59027,7.6579537,3.7256382,3.3104696,2.8953013,2.4801328,2.0649643,1.649796,2.764768,3.87974,4.994712,6.109684,7.224656,6.506723,5.7906027,5.0726695,4.3547363,3.636803,3.9957695,4.3529234,4.710077,5.06723,5.424384,6.1296263,6.834869,7.5401115,8.245354,8.950596,7.2899227,5.6292486,3.9703882,2.3097143,0.6508536,0.6200332,0.58921283,0.56020546,0.5293851,0.50037766,0.4894999,0.48043507,0.46955732,0.4604925,0.44961473,0.42967212,0.40972954,0.38978696,0.36984438,0.34990177,0.27919623,0.21030366,0.13959812,0.07070554,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.40066472,0.7505665,1.1004683,1.4503701,1.8002719,1.4394923,1.0805258,0.7197462,0.36077955,0.0,0.15954071,0.3208944,0.48043507,0.6399758,0.7995165,1.2273756,1.6552348,2.0830941,2.5091403,2.9369993,2.4420607,1.9471219,1.452183,0.9572442,0.46230546,0.6852999,0.90829426,1.1294757,1.35247,1.5754645,1.5754645,1.5754645,1.5754645,1.5754645,1.5754645,1.260009,0.9445535,0.629098,0.3154555,0.0,0.26469254,0.5293851,0.79589057,1.0605831,1.3252757,1.209246,1.0950294,0.9808127,0.86478317,0.7505665,0.8629702,0.97537386,1.0877775,1.2001812,1.3125849,1.2328146,1.1530442,1.0732739,0.9916905,0.9119202,1.0333886,1.1530442,1.2726997,1.3923552,1.5120108,1.5573349,1.6026589,1.647983,1.693307,1.7368182,2.179181,2.6233568,3.0657198,3.5080826,3.9504454,4.936697,5.924762,6.9128265,7.900891,8.887142,7.897265,6.9073873,5.91751,4.9276323,3.9377546,3.299592,2.663242,2.0250793,1.3869164,0.7505665,0.65991837,0.56927025,0.48043507,0.38978696,0.2991388,0.32995918,0.36077955,0.38978696,0.42060733,0.44961473,0.38072214,0.3100166,0.23931105,0.17041849,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.09064813,0.07977036,0.07070554,0.059827764,0.05076295,0.15047589,0.25018883,0.34990177,0.44961473,0.5493277,0.56020546,0.56927025,0.58014804,0.58921283,0.6000906,0.48043507,0.36077955,0.23931105,0.11965553,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.027194439,0.054388877,0.08339628,0.11059072,0.13778515,0.13959812,0.14322405,0.14503701,0.14684997,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,1.0007553,1.8492218,2.6995013,3.5497808,4.40006,3.7655232,3.1291735,2.4946365,1.8600996,1.2255627,1.9271792,2.6306088,3.3322253,4.0356545,4.7372713,7.706904,10.676537,13.647983,16.617615,19.587248,19.505665,19.422268,19.340685,19.257288,19.175705,15.912373,12.650853,9.38752,6.1241875,2.8626678,2.2897718,1.7168756,1.1457924,0.5728962,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.065266654,0.07977036,0.09427405,0.11059072,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.19942589,0.2755703,0.34990177,0.42423326,0.50037766,0.40066472,0.2991388,0.19942589,0.099712946,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.07070554,0.12690738,0.18492219,0.24293698,0.2991388,0.23931105,0.1794833,0.11965553,0.059827764,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13959812,0.27919623,0.42060733,0.56020546,0.69980353,0.99531645,1.2908293,1.5845293,1.8800422,2.175555,4.550536,6.925517,9.300498,11.675479,14.05046,13.9779415,13.905423,13.832905,13.760386,13.687867,14.327844,14.967819,15.607795,16.24777,16.887747,18.425138,19.96253,21.499924,23.037315,24.574707,22.359268,20.14564,17.9302,15.71476,13.499319,12.473183,11.445232,10.417283,9.389333,8.363196,8.937905,9.512614,10.087324,10.662033,11.236742,13.174799,15.112856,17.0491,18.987158,20.925215,16.962078,12.998941,9.037619,5.0744824,1.1131591,1.987007,2.8626678,3.738329,4.612177,5.487838,5.5531044,5.618371,5.6818247,5.7470913,5.812358,6.644508,7.478471,8.31062,9.142771,9.97492,10.277685,10.58045,10.883214,11.185979,11.486931,10.145339,8.801933,7.460341,6.1169357,4.7753434,9.953164,15.130985,20.306993,25.484816,30.662636,27.848919,25.037014,22.22511,19.413204,16.599485,15.8326025,15.065719,14.297023,13.53014,12.763257,17.00015,16.354736,15.709321,15.065719,14.420304,13.77489,13.765825,13.754947,13.745882,13.735004,13.724127,13.015259,12.304577,11.595709,10.885027,10.174346,8.767487,7.360628,5.9519563,4.5450974,3.1382382,2.8626678,2.5870976,2.3133402,2.03777,1.7621996,2.9442513,4.1281157,5.3101673,6.492219,7.6742706,7.1829576,6.6898317,6.1967063,5.7053933,5.2122674,4.40006,3.587853,2.7756457,1.9616255,1.1494182,1.0750868,1.0007553,0.9246109,0.85027945,0.774135,0.88291276,0.9898776,1.0968424,1.2056202,1.3125849,1.3832904,1.452183,1.5228885,1.5917811,1.6624867,1.4630609,1.261822,1.062396,0.8629702,0.66173136,0.629098,0.5982776,0.5656443,0.533011,0.50037766,0.5076295,0.5148814,0.52213323,0.5293851,0.53663695,0.45324063,0.3680314,0.28282216,0.19761293,0.11240368,0.32814622,0.5420758,0.75781834,0.97174793,1.1874905,1.2382535,1.2872034,1.3379664,1.3869164,1.4376793,1.5627737,1.6878681,1.8129625,1.938057,2.0631514,1.8727903,1.6824293,1.4920682,1.3017071,1.1131591,0.922798,0.7324369,0.5420758,0.35171473,0.16316663,0.3208944,0.47680917,0.6345369,0.79226464,0.9499924,0.90466833,0.85934424,0.81583315,0.7705091,0.72518504,0.58014804,0.43511102,0.29007402,0.14503701,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.78319985,1.5645868,2.3477864,3.1291735,3.9123733,5.0654173,6.2166486,7.369693,8.5227375,9.675781,8.874452,8.074935,7.2754188,6.474089,5.674573,5.618371,5.560356,5.5023413,5.4443264,5.388125,5.77066,6.153195,6.53573,6.9182653,7.3008003,6.8620634,6.4251394,5.9882154,5.5494785,5.1125546,4.2042603,3.2977788,2.3894846,1.4830034,0.5747091,7.0451727,13.515636,19.9861,26.45475,32.925213,26.345972,19.764917,13.185677,6.604623,0.025381476,2.3097143,4.594047,6.880193,9.164526,11.450671,10.515183,9.579695,8.644206,7.71053,6.775041,8.644206,10.515183,12.384347,14.255324,16.124489,14.996826,13.8691635,12.743314,11.615651,10.487988,12.670795,14.851789,17.034595,19.217403,21.40021,18.610062,15.819912,13.029762,10.239613,7.4494634,6.4070096,5.3645563,4.322103,3.2796493,2.2371957,3.4808881,4.7227674,5.964647,7.208339,8.450218,7.315304,6.1803894,5.045475,3.9105604,2.7756457,3.489953,4.2042603,4.9203806,5.634688,6.350808,6.4233265,6.495845,6.5683637,6.640882,6.7115874,5.467895,4.2223897,2.9768846,1.7331922,0.48768693,0.46411842,0.44236287,0.42060733,0.39703882,0.37528324,0.3680314,0.36077955,0.35171473,0.3444629,0.33721104,0.32270733,0.30820364,0.291887,0.27738327,0.26287958,0.21030366,0.15772775,0.10515183,0.052575916,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.2991388,0.5620184,0.824898,1.0877775,1.3506571,1.0805258,0.8103943,0.5402629,0.27013144,0.0,0.28282216,0.5656443,0.8466535,1.1294757,1.4122978,1.7295663,2.0468347,2.3659163,2.6831846,3.000453,2.4855716,1.9706904,1.455809,0.93911463,0.42423326,0.6200332,0.81583315,1.0098201,1.2056202,1.3996071,1.3633479,1.3252757,1.2872034,1.2491312,1.2128719,0.969935,0.726998,0.48587397,0.24293698,0.0,0.5293851,1.0605831,1.5899682,2.1193533,2.6505513,2.420305,2.1900587,1.9598125,1.7295663,1.49932,1.6878681,1.8746033,2.0631514,2.2498865,2.4366217,2.3151531,2.1918716,2.0704033,1.9471219,1.8256533,1.9271792,2.030518,2.132044,2.2353828,2.3369088,2.327844,2.3169663,2.3079014,2.2970235,2.2879589,2.5599031,2.8318477,3.105605,3.3775494,3.6494937,4.4508233,5.2503395,6.049856,6.849373,7.650702,6.794984,5.9392653,5.08536,4.229642,3.3757362,2.811905,2.2498865,1.6878681,1.1258497,0.5620184,0.4949388,0.42785916,0.36077955,0.291887,0.22480737,0.24837588,0.27013144,0.291887,0.3154555,0.33721104,0.28463513,0.23205921,0.1794833,0.12690738,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.06707962,0.059827764,0.052575916,0.045324065,0.038072214,0.17585737,0.31182957,0.44961473,0.5873999,0.72518504,0.67079616,0.61459434,0.56020546,0.5058166,0.44961473,0.36077955,0.27013144,0.1794833,0.09064813,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.054388877,0.11059072,0.16497959,0.21936847,0.2755703,0.24293698,0.21030366,0.17767033,0.14503701,0.11240368,0.09064813,0.06707962,0.045324065,0.02175555,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.7505665,1.3869164,2.0250793,2.663242,3.299592,2.8807976,2.4601903,2.039583,1.6207886,1.2001812,1.7549478,2.3097143,2.864481,3.4192474,3.975827,6.301858,8.629702,10.957546,13.28539,15.613234,15.622298,15.633177,15.6422415,15.653119,15.662184,12.975373,10.28675,7.5999393,4.9131284,2.2245052,1.7803292,1.3343405,0.8901646,0.44417584,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.11784257,0.13415924,0.15228885,0.17041849,0.18673515,0.17585737,0.16316663,0.15047589,0.13778515,0.12509441,0.28826106,0.44961473,0.61278135,0.774135,0.93730164,0.7505665,0.5620184,0.37528324,0.18673515,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.09064813,0.15410182,0.21936847,0.28463513,0.34990177,0.27919623,0.21030366,0.13959812,0.07070554,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.10515183,0.21030366,0.3154555,0.42060733,0.52575916,0.8031424,1.0805258,1.357909,1.6352923,1.9126755,4.062849,6.2130227,8.363196,10.511557,12.661731,12.5058155,12.348088,12.19036,12.032633,11.874905,12.442362,13.009819,13.577277,14.144734,14.712192,16.062849,17.411694,18.76235,20.113007,21.461851,19.34431,17.22677,15.10923,12.993503,10.874149,12.019942,13.165734,14.309713,15.455506,16.599485,15.5878525,14.574407,13.562773,12.549327,11.537694,12.60009,13.662486,14.724882,15.787278,16.849674,13.812962,10.774437,7.7377243,4.701012,1.6624867,2.3622901,3.0620937,3.7618973,4.461701,5.163317,5.4932766,5.823236,6.153195,6.4831543,6.813113,7.4277077,8.042302,8.656897,9.273304,9.8878975,11.691795,13.497506,15.303217,17.107115,18.912827,16.539658,14.16649,11.795135,9.421967,7.0506115,10.368333,13.686054,17.001963,20.319685,23.637405,21.474543,19.311678,17.150625,14.9877615,12.824898,12.415168,12.005438,11.595709,11.184166,10.774437,17.812357,16.99471,16.177065,15.359419,14.541773,13.724127,13.872789,14.01964,14.168303,14.315152,14.462003,14.010575,13.557334,13.104094,12.652666,12.199425,10.54419,8.890768,7.2355337,5.580299,3.925064,3.5117085,3.100166,2.6868105,2.275268,1.8619126,2.6306088,3.397492,4.164375,4.933071,5.6999545,5.542227,5.384499,5.2267714,5.0708566,4.9131284,4.2368937,3.5624714,2.8880494,2.2118144,1.5373923,1.4376793,1.3379664,1.2382535,1.1367276,1.0370146,1.0424535,1.0478923,1.0533313,1.0569572,1.062396,1.2545701,1.4467441,1.6407311,1.8329052,2.0250793,1.7132497,1.3996071,1.0877775,0.774135,0.46230546,0.4949388,0.5275721,0.56020546,0.59283876,0.62547207,0.6055295,0.5855869,0.5656443,0.54570174,0.52575916,0.43511102,0.3444629,0.25562772,0.16497959,0.07433146,0.2229944,0.36984438,0.5166943,0.6653573,0.8122072,1.0370146,1.261822,1.4866294,1.7132497,1.938057,1.9996977,2.0631514,2.124792,2.1882458,2.2498865,2.0142014,1.7803292,1.5446441,1.310772,1.0750868,0.90285534,0.7306239,0.55839247,0.38434806,0.21211663,0.40429065,0.5982776,0.7904517,0.9826257,1.1747998,1.0696479,0.9644961,0.85934424,0.7541924,0.6508536,0.52032024,0.38978696,0.25925365,0.13053331,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.8792868,1.7603867,2.6396735,3.5207734,4.40006,4.847862,5.295664,5.7416525,6.189454,6.637256,6.825804,7.0125394,7.1992745,7.3878226,7.574558,7.5818095,7.590874,7.5981264,7.605378,7.61263,8.2798,8.94697,9.6141405,10.283124,10.950294,10.275872,9.599637,8.925215,8.2507925,7.574558,6.169512,4.764466,3.3594196,1.9543737,0.5493277,10.31757,20.084,29.852242,39.620483,49.386913,39.517147,29.647377,19.777609,9.907841,0.038072214,2.039583,4.0429068,6.0444174,8.047741,10.049252,9.547061,9.04487,8.54268,8.040489,7.5382986,8.392203,9.247922,10.101828,10.957546,11.813264,11.9021,11.992747,12.083396,12.172231,12.262879,13.693306,15.121921,16.55235,17.982777,19.413204,17.76522,16.117237,14.4692545,12.823084,11.175101,9.5053625,7.835624,6.164073,4.494334,2.8245957,4.195195,5.565795,6.9345818,8.3051815,9.675781,8.122072,6.5701766,5.0182805,3.4645715,1.9126755,2.9841363,4.0574102,5.130684,6.202145,7.2754188,6.7152133,6.155008,5.5948024,5.034597,4.4743915,3.6458678,2.8155308,1.9851941,1.1548572,0.3245203,0.3100166,0.2955129,0.27919623,0.26469254,0.25018883,0.24474995,0.23931105,0.23568514,0.23024625,0.22480737,0.21574254,0.20486477,0.19579996,0.18492219,0.17585737,0.13959812,0.10515183,0.07070554,0.034446288,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.19942589,0.37528324,0.5493277,0.72518504,0.89922947,0.7197462,0.5402629,0.36077955,0.1794833,0.0,0.40429065,0.8103943,1.214685,1.6207886,2.0250793,2.231757,2.4402475,2.6469254,2.855416,3.0620937,2.5272698,1.9924458,1.4576219,0.922798,0.387974,0.55476654,0.72337204,0.8901646,1.0569572,1.2255627,1.1494182,1.0750868,1.0007553,0.9246109,0.85027945,0.67986095,0.5094425,0.34083697,0.17041849,0.0,0.79589057,1.5899682,2.3858588,3.1799364,3.975827,3.6295512,3.2850883,2.9406252,2.5943494,2.2498865,2.5127661,2.7756457,3.0367124,3.299592,3.5624714,3.397492,3.2325122,3.0675328,2.902553,2.7375734,2.8227828,2.907992,2.9932013,3.0765975,3.1618068,3.0983531,3.0330863,2.9678197,2.902553,2.8372865,2.9406252,3.0421512,3.1454902,3.247016,3.350355,3.9631362,4.574105,5.186886,5.7996674,6.412449,5.6927023,4.972956,4.25321,3.531651,2.811905,2.324218,1.8383441,1.3506571,0.8629702,0.37528324,0.32995918,0.28463513,0.23931105,0.19579996,0.15047589,0.16497959,0.1794833,0.19579996,0.21030366,0.22480737,0.19036107,0.15410182,0.11965553,0.08520924,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.045324065,0.03988518,0.034446288,0.030820364,0.025381476,0.19942589,0.37528324,0.5493277,0.72518504,0.89922947,0.7795739,0.65991837,0.5402629,0.42060733,0.2991388,0.23931105,0.1794833,0.11965553,0.059827764,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08339628,0.16497959,0.24837588,0.32995918,0.41335547,0.3444629,0.27738327,0.21030366,0.14322405,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.50037766,0.9246109,1.3506571,1.7748904,2.1991236,1.9942589,1.789394,1.5845293,1.3796645,1.1747998,1.5827163,1.9906329,2.3967366,2.8046532,3.2125697,4.896812,6.582867,8.267109,9.953164,11.637406,11.740746,11.842272,11.94561,12.047136,12.1504755,10.036561,7.9244595,5.812358,3.7002566,1.5881553,1.2708868,0.95180535,0.6345369,0.31726846,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.17041849,0.19036107,0.21030366,0.23024625,0.25018883,0.22480737,0.19942589,0.17585737,0.15047589,0.12509441,0.37528324,0.62547207,0.87566096,1.1258497,1.3742256,1.1004683,0.824898,0.5493277,0.2755703,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.11059072,0.18310922,0.25562772,0.32814622,0.40066472,0.3208944,0.23931105,0.15954071,0.07977036,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07070554,0.13959812,0.21030366,0.27919623,0.34990177,0.6091554,0.87022203,1.1294757,1.3905423,1.649796,3.5751622,5.5005283,7.4258947,9.349448,11.274815,11.0318775,10.790753,10.547816,10.304879,10.061942,10.556881,11.05182,11.546759,12.0416975,12.536636,13.700559,14.862667,16.024776,17.186886,18.350807,16.329353,14.309713,12.290073,10.270433,8.2507925,11.568514,14.886236,18.202145,21.519865,24.837587,22.237799,19.63801,17.038223,14.438434,11.836833,12.025381,12.212116,12.400664,12.5873995,12.774135,10.662033,8.549932,6.43783,4.325729,2.2118144,2.7375734,3.2633326,3.787279,4.313038,4.836984,5.431636,6.0281005,6.622752,7.217404,7.8120556,8.210908,8.607946,9.004985,9.402024,9.800876,13.107719,16.414564,19.72322,23.030064,26.336908,22.933977,19.53286,16.129929,12.726997,9.325879,10.781689,12.23931,13.696932,15.154554,16.612177,15.100165,13.588155,12.07433,10.56232,9.050309,8.997733,8.945157,8.892582,8.840006,8.78743,18.624565,17.634687,16.64481,15.654932,14.665054,13.675177,13.979754,14.284332,14.590723,14.895301,15.199879,15.005891,14.810091,14.614291,14.420304,14.224504,12.322706,10.420909,8.517298,6.6155005,4.7118897,4.162562,3.6132345,3.0620937,2.5127661,1.9616255,2.3151531,2.666868,3.0203958,3.3721104,3.7256382,3.9033084,4.079166,4.256836,4.4345064,4.612177,4.07554,3.53709,3.000453,2.4620032,1.9253663,1.8002719,1.6751775,1.550083,1.4249886,1.2998942,1.2019942,1.1059072,1.0080072,0.9101072,0.8122072,1.1276628,1.4431182,1.7567607,2.0722163,2.3876717,1.9616255,1.5373923,1.1131591,0.6871128,0.26287958,0.36077955,0.45686656,0.55476654,0.6526665,0.7505665,0.7016165,0.6544795,0.6073425,0.56020546,0.51306844,0.4169814,0.32270733,0.22662032,0.13234627,0.038072214,0.11784257,0.19761293,0.27738327,0.35715362,0.43692398,0.8375887,1.2382535,1.6371052,2.03777,2.4366217,2.4366217,2.4366217,2.4366217,2.4366217,2.4366217,2.1574254,1.8782293,1.5972201,1.3180238,1.0370146,0.88291276,0.726998,0.5728962,0.4169814,0.26287958,0.4894999,0.7179332,0.9445535,1.1729867,1.3996071,1.2346275,1.0696479,0.90466833,0.73968875,0.5747091,0.4604925,0.3444629,0.23024625,0.11421664,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.97718686,1.9543737,2.9333735,3.9105604,4.8877473,4.6303062,4.3728657,4.115425,3.8579843,3.6005437,4.7753434,5.9501433,7.124943,8.299743,9.474543,9.547061,9.619579,9.692098,9.764616,9.837135,10.790753,11.7425585,12.694364,13.647983,14.599788,13.687867,12.775948,11.862214,10.950294,10.038374,8.134763,6.2329655,4.329355,2.427557,0.52575916,13.589968,26.654177,39.720196,52.786217,65.850426,52.690132,39.529835,26.369541,13.209246,0.05076295,1.7694515,3.489953,5.2104545,6.929143,8.649645,8.580752,8.510046,8.439341,8.370448,8.299743,8.140202,7.9806614,7.819308,7.6597667,7.500226,8.807372,10.114518,11.421664,12.730623,14.037769,14.715817,15.392053,16.0701,16.748148,17.424383,16.92038,16.414564,15.91056,15.404743,14.90074,12.601903,10.304879,8.007855,5.710832,3.4119956,4.9095025,6.4070096,7.9045167,9.402024,10.899531,8.930654,6.9599633,4.989273,3.0203958,1.0497054,2.4801328,3.9105604,5.3391747,6.7696023,8.200029,7.0071006,5.814171,4.6230545,3.4301252,2.2371957,1.8220274,1.4068589,0.9916905,0.57833505,0.16316663,0.15410182,0.14684997,0.13959812,0.13234627,0.12509441,0.12328146,0.11965553,0.11784257,0.11421664,0.11240368,0.10696479,0.10333887,0.09789998,0.092461094,0.0870222,0.07070554,0.052575916,0.034446288,0.018129626,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.099712946,0.18673515,0.2755703,0.36259252,0.44961473,0.36077955,0.27013144,0.1794833,0.09064813,0.0,0.5275721,1.0551442,1.5827163,2.1102884,2.6378605,2.7357605,2.8318477,2.9297476,3.0276475,3.1255474,2.570781,2.0142014,1.4594349,0.90466833,0.34990177,0.4894999,0.629098,0.7705091,0.9101072,1.0497054,0.93730164,0.824898,0.7124943,0.6000906,0.48768693,0.38978696,0.291887,0.19579996,0.09789998,0.0,1.0605831,2.1193533,3.1799364,4.2405195,5.2992897,4.84061,4.3801174,3.919625,3.4591327,3.000453,3.3376641,3.6748753,4.0120864,4.349297,4.688321,4.4798307,4.273153,4.064662,3.8579843,3.6494937,3.7183862,3.785466,3.8525455,3.919625,3.9867048,3.8670492,3.7473936,3.6277382,3.5080826,3.386614,3.3195345,3.2524548,3.1853752,3.1182957,3.049403,3.4754493,3.8996825,4.325729,4.749962,5.1741953,4.590421,4.004834,3.4192474,2.8354735,2.2498865,1.8383441,1.4249886,1.0116332,0.6000906,0.18673515,0.16497959,0.14322405,0.11965553,0.09789998,0.07433146,0.08339628,0.09064813,0.09789998,0.10515183,0.11240368,0.09427405,0.07795739,0.059827764,0.04169814,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.02175555,0.01994259,0.018129626,0.014503701,0.012690738,0.22480737,0.43692398,0.6508536,0.8629702,1.0750868,0.8901646,0.70524246,0.52032024,0.33539808,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.11059072,0.21936847,0.32995918,0.4405499,0.5493277,0.44780177,0.3444629,0.24293698,0.13959812,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.25018883,0.46230546,0.6744221,0.8883517,1.1004683,1.1095331,1.1204109,1.1294757,1.1403534,1.1494182,1.4104849,1.6697385,1.9308052,2.1900587,2.4493124,3.491766,4.5342193,5.576673,6.6191263,7.66158,7.85738,8.05318,8.247167,8.442966,8.636953,7.0995617,5.562169,4.024777,2.4873846,0.9499924,0.75963134,0.56927025,0.38072214,0.19036107,0.0,0.03988518,0.07977036,0.11965553,0.15954071,0.19942589,0.2229944,0.24474995,0.26831847,0.29007402,0.31182957,0.2755703,0.2374981,0.19942589,0.16316663,0.12509441,0.46230546,0.7995165,1.1367276,1.4757515,1.8129625,1.4503701,1.0877775,0.72518504,0.36259252,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.13053331,0.21030366,0.29007402,0.36984438,0.44961473,0.36077955,0.27013144,0.1794833,0.09064813,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.034446288,0.07070554,0.10515183,0.13959812,0.17585737,0.4169814,0.65991837,0.90285534,1.1457924,1.3869164,3.0874753,4.788034,6.48678,8.187339,9.8878975,9.5597515,9.231606,8.9052725,8.577126,8.2507925,8.673213,9.0956335,9.518054,9.940474,10.362894,11.338268,12.311829,13.287203,14.262577,15.23795,13.314397,11.392657,9.469104,7.5473633,5.6256227,11.115273,16.604925,22.094576,27.584227,33.07569,28.887745,24.699802,20.511858,16.325727,12.137785,11.450671,10.761745,10.074633,9.38752,8.700407,7.512917,6.3254266,5.137936,3.9504454,2.762955,3.1128569,3.4627585,3.8126602,4.162562,4.512464,5.371808,6.2329655,7.0923095,7.951654,8.812811,8.992294,9.171778,9.353074,9.5325575,9.712041,14.5236435,19.333433,24.143223,28.953012,33.762802,29.330109,24.897415,20.464722,16.032028,11.599335,11.1968565,10.794379,10.391902,9.989424,9.5869465,8.723976,7.8628187,6.9998484,6.1368785,5.275721,5.580299,5.8848767,6.189454,6.495845,6.8004227,19.436771,18.274662,17.112555,15.950445,14.788336,13.6244135,14.0867195,14.5508375,15.013144,15.475449,15.937754,15.999394,16.062849,16.124489,16.187943,16.249584,14.09941,11.949236,9.799063,7.650702,5.5005283,4.8134155,4.12449,3.437377,2.7502642,2.0631514,1.9996977,1.938057,1.8746033,1.8129625,1.7495089,2.2625773,2.7756457,3.2869012,3.7999697,4.313038,3.9123733,3.5117085,3.1128569,2.712192,2.3133402,2.1628644,2.0123885,1.8619126,1.7132497,1.5627737,1.3633479,1.162109,0.96268314,0.76325727,0.5620184,1.0007553,1.4376793,1.8746033,2.3133402,2.7502642,2.2118144,1.6751775,1.1367276,0.6000906,0.06164073,0.22480737,0.387974,0.5493277,0.7124943,0.87566096,0.7995165,0.72518504,0.6508536,0.5747091,0.50037766,0.40066472,0.2991388,0.19942589,0.099712946,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.63816285,1.2128719,1.7875811,2.3622901,2.9369993,2.8753586,2.811905,2.7502642,2.6868105,2.6251698,2.3006494,1.9743162,1.649796,1.3252757,1.0007553,0.8629702,0.72518504,0.5873999,0.44961473,0.31182957,0.5747091,0.8375887,1.1004683,1.3633479,1.6244144,1.3996071,1.1747998,0.9499924,0.72518504,0.50037766,0.40066472,0.2991388,0.19942589,0.099712946,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.0750868,2.1501737,3.2252605,4.3003473,5.375434,4.4127507,3.4500678,2.4873846,1.5247015,0.5620184,2.7248828,4.8877473,7.0506115,9.211663,11.374527,11.512312,11.650098,11.787883,11.925668,12.06164,13.299893,14.538147,15.774588,17.01284,18.24928,17.099863,15.950445,14.799213,13.649796,12.500377,10.100015,7.699652,5.2992897,2.9007401,0.50037766,16.862366,33.224354,49.588154,65.95014,82.312126,65.86312,49.412296,32.96147,16.512463,0.06164073,1.49932,2.9369993,4.3746786,5.812358,7.250037,7.61263,7.9752226,8.337815,8.700407,9.063,7.8882003,6.7134004,5.5367875,4.361988,3.1871881,5.712645,8.238102,10.761745,13.287203,15.812659,15.738328,15.662184,15.5878525,15.511708,15.437376,16.075539,16.71189,17.350052,17.988214,18.624565,15.700256,12.775948,9.849826,6.925517,3.9993954,5.6256227,7.250037,8.874452,10.500679,12.125093,9.737422,7.3497505,4.9620786,2.5744069,0.18673515,1.9743162,3.7618973,5.5494785,7.3370595,9.12464,7.3008003,5.475147,3.6494937,1.8256533,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.6508536,1.2998942,1.9507477,2.5997884,3.2506418,3.2379513,3.2252605,3.2125697,3.199879,3.1871881,2.612479,2.03777,1.4630609,0.8883517,0.31182957,0.42423326,0.53663695,0.6508536,0.76325727,0.87566096,0.72518504,0.5747091,0.42423326,0.2755703,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,1.3252757,2.6505513,3.975827,5.2992897,6.624565,6.049856,5.475147,4.900438,4.325729,3.7492065,4.162562,4.574105,4.98746,5.4008155,5.812358,5.562169,5.3119802,5.0617914,4.8116026,4.5632267,4.612177,4.6629395,4.7118897,4.762653,4.8116026,4.6375585,4.461701,4.2876563,4.1117992,3.9377546,3.7002566,3.4627585,3.2252605,2.9877625,2.7502642,2.9877625,3.2252605,3.4627585,3.7002566,3.9377546,3.48814,3.0367124,2.5870976,2.137483,1.6878681,1.3506571,1.0116332,0.6744221,0.33721104,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.25018883,0.50037766,0.7505665,1.0007553,1.2491312,1.0007553,0.7505665,0.50037766,0.25018883,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13778515,0.2755703,0.41335547,0.5493277,0.6871128,0.5493277,0.41335547,0.2755703,0.13778515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.22480737,0.44961473,0.6744221,0.89922947,1.1258497,1.2382535,1.3506571,1.4630609,1.5754645,1.6878681,2.08672,2.4873846,2.8880494,3.2869012,3.6875658,3.975827,4.262275,4.550536,4.836984,5.125245,4.162562,3.199879,2.2371957,1.2745126,0.31182957,0.25018883,0.18673515,0.12509441,0.06164073,0.0,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,0.2755703,0.2991388,0.3245203,0.34990177,0.37528324,0.3245203,0.2755703,0.22480737,0.17585737,0.12509441,0.5493277,0.97537386,1.3996071,1.8256533,2.2498865,1.8002719,1.3506571,0.89922947,0.44961473,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.15047589,0.2374981,0.3245203,0.41335547,0.50037766,0.40066472,0.2991388,0.19942589,0.099712946,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.22480737,0.44961473,0.6744221,0.89922947,1.1258497,2.5997884,4.07554,5.5494785,7.02523,8.499168,8.087626,7.6742706,7.262728,6.849373,6.43783,6.787732,7.137634,7.4875355,7.837437,8.187339,8.974165,9.762803,10.549629,11.338268,12.125093,10.29944,8.4756,6.6499467,4.8242936,3.000453,10.663846,18.325426,25.987005,33.6504,41.311977,35.537693,29.761593,23.987309,18.213022,12.436923,10.874149,9.313189,7.750415,6.187641,4.6248674,4.361988,4.099108,3.8380418,3.5751622,3.3122826,3.48814,3.6621845,3.8380418,4.0120864,4.1879435,5.3119802,6.43783,7.5618668,8.6877165,9.811753,9.775495,9.737422,9.699349,9.663091,9.625018,15.937754,22.25049,28.563225,34.87415,41.186886,35.724426,30.26197,24.799515,19.337059,13.874602,11.612025,9.349448,7.0868707,4.8242936,2.561716,2.3495996,2.137483,1.9253663,1.7132497,1.49932,2.1628644,2.8245957,3.48814,4.1498713,4.8116026,19.449463,18.577427,17.705393,16.833357,15.95951,15.087475,15.511708,15.937754,16.361988,16.788034,17.212267,17.147,17.081734,17.01828,16.953012,16.887747,14.955129,13.022511,11.089892,9.157274,7.224656,6.48678,5.750717,5.0128417,4.274966,3.53709,3.4192474,3.303218,3.1853752,3.0675328,2.94969,3.3322253,3.7147603,4.0972953,4.4798307,4.8623657,4.269527,3.6766882,3.0856624,2.4928236,1.8999848,1.887294,1.8746033,1.8619126,1.8492218,1.8383441,1.5645868,1.2926424,1.020698,0.7469406,0.4749962,0.9572442,1.4394923,1.9217403,2.4058013,2.8880494,2.3967366,1.9072367,1.4177368,0.92823684,0.43692398,0.4894999,0.5420758,0.5946517,0.64722764,0.69980353,0.7016165,0.70524246,0.7070554,0.7106813,0.7124943,0.78319985,0.8520924,0.922798,0.9916905,1.062396,0.94092757,0.81764615,0.69436467,0.5728962,0.44961473,0.9445535,1.4394923,1.9344311,2.42937,2.9243085,2.8608549,2.7955883,2.7303216,2.665055,2.5997884,2.3369088,2.0758421,1.8129625,1.550083,1.2872034,1.0877775,0.8883517,0.6871128,0.48768693,0.28826106,0.4894999,0.69255173,0.89560354,1.0968424,1.2998942,1.1204109,0.93911463,0.75963134,0.58014804,0.40066472,0.3208944,0.23931105,0.15954071,0.07977036,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.8901646,1.742257,2.5943494,3.4482548,4.3003473,3.5932918,2.8844235,2.1773682,1.4703126,0.76325727,2.5798457,4.3982472,6.2148356,8.033237,9.849826,10.444477,11.039129,11.635593,12.230246,12.824898,13.7875805,14.750263,15.712947,16.67563,17.638313,16.360174,15.082036,13.80571,12.527572,11.249433,9.169965,7.0904965,5.009216,2.9297476,0.85027945,13.994258,27.140049,40.285843,53.42982,66.5738,53.678196,40.78078,27.881552,14.984136,2.08672,2.94969,3.8126602,4.6756306,5.5367875,6.399758,6.773228,7.1448855,7.518356,7.890013,8.26167,7.454902,6.6481338,5.8395524,5.032784,4.2242026,5.995467,7.764919,9.53437,11.3056345,13.075087,12.931862,12.790451,12.647227,12.5058155,12.362592,12.870221,13.377851,13.885481,14.39311,14.90074,12.5602045,10.21967,7.8791356,5.540414,3.199879,4.646623,6.09518,7.5419245,8.990481,10.437225,8.450218,6.4632115,4.4743915,2.4873846,0.50037766,1.8600996,3.2198215,4.5795436,5.9392653,7.3008003,6.205771,5.1107416,4.0157123,2.9206827,1.8256533,1.6733645,1.5192627,1.3669738,1.214685,1.062396,0.8520924,0.6417888,0.43329805,0.2229944,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.09064813,0.1794833,0.27013144,0.36077955,0.44961473,0.46774435,0.48587397,0.50219065,0.52032024,0.53663695,0.5148814,0.49312583,0.46955732,0.44780177,0.42423326,0.968122,1.5101979,2.0522738,2.5943494,3.1382382,3.0675328,2.9968271,2.9279346,2.857229,2.7883365,2.2843328,1.7821422,1.2799516,0.7777609,0.2755703,0.40066472,0.52575916,0.6508536,0.774135,0.89922947,0.7868258,0.6744221,0.5620184,0.44961473,0.33721104,0.58014804,0.823085,1.064209,1.3071461,1.550083,2.3151531,3.0802233,3.8452935,4.610364,5.375434,4.900438,4.4254417,3.9504454,3.4754493,3.000453,3.4047437,3.8108473,4.215138,4.6194286,5.0255322,4.940323,4.855114,4.7699046,4.6846952,4.599486,4.9820213,5.3645563,5.7470913,6.1296263,6.5121617,6.1368785,5.763408,5.388125,5.0128417,4.6375585,4.3202896,4.0030212,3.6857529,3.3666716,3.049403,3.152742,3.254268,3.3576066,3.4591327,3.5624714,3.1219215,2.6831846,2.2426348,1.8020848,1.3633479,1.0895905,0.81764615,0.54570174,0.27194437,0.0,0.09064813,0.1794833,0.27013144,0.36077955,0.44961473,0.4550536,0.4604925,0.46411842,0.46955732,0.4749962,0.38434806,0.2955129,0.20486477,0.11421664,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.21755551,0.43511102,0.6526665,0.87022203,1.0877775,0.87022203,0.6526665,0.43511102,0.21755551,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.11059072,0.21936847,0.32995918,0.4405499,0.5493277,0.4405499,0.32995918,0.21936847,0.11059072,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.18492219,0.36984438,0.55476654,0.73968875,0.9246109,1.0605831,1.1947423,1.3307146,1.4648738,1.6008459,1.9725033,2.3441606,2.7176309,3.0892882,3.4627585,3.7020695,3.9431937,4.1825047,4.421816,4.6629395,4.510651,4.358362,4.2042603,4.0519714,3.8996825,3.2107568,2.520018,1.8292793,1.1403534,0.44961473,0.40066472,0.34990177,0.2991388,0.25018883,0.19942589,0.21936847,0.23931105,0.25925365,0.27919623,0.2991388,0.25925365,0.21936847,0.1794833,0.13959812,0.099712946,0.4405499,0.7795739,1.1204109,1.4594349,1.8002719,1.4431182,1.0841516,0.726998,0.36984438,0.012690738,0.065266654,0.11784257,0.17041849,0.2229944,0.2755703,0.3154555,0.35534066,0.39522585,0.43511102,0.4749962,0.3825351,0.29007402,0.19761293,0.10515183,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1794833,0.36077955,0.5402629,0.7197462,0.89922947,2.1519866,3.4047437,4.6575007,5.910258,7.1630154,6.9980354,6.833056,6.6680765,6.5030966,6.338117,7.083245,7.8283725,8.571687,9.316814,10.061942,10.58045,11.097144,11.615651,12.132345,12.650853,10.9774885,9.305937,7.6325727,5.961021,4.2876563,10.167094,16.048346,21.927782,27.80722,33.686657,30.23659,26.786522,23.338266,19.888199,16.438131,15.054841,13.671551,12.290073,10.908596,9.525306,8.890768,8.254418,7.6198816,6.985345,6.350808,6.2746634,6.200332,6.1241875,6.049856,5.975525,6.6571984,7.3406854,8.02236,8.705847,9.38752,9.253361,9.117389,8.98323,8.847258,8.713099,13.647983,18.582867,23.51775,28.452635,33.38752,29.31198,25.236439,21.162712,17.087172,13.011633,11.617464,10.221483,8.827314,7.4331465,6.037165,5.422571,4.8079767,4.1933823,3.576975,2.962381,3.29234,3.6222992,3.9522583,4.2822175,4.612177,19.462152,18.880192,18.298231,17.714457,17.132496,16.550535,16.936697,17.32467,17.712645,18.100618,18.48678,18.294605,18.102432,17.910257,17.718082,17.52591,15.810846,14.095784,12.380721,10.665659,8.950596,8.161958,7.3751316,6.588306,5.7996674,5.0128417,4.84061,4.668379,4.494334,4.322103,4.1498713,4.401873,4.655688,4.9076896,5.1596913,5.411693,4.6266804,3.8416677,3.056655,2.2716422,1.4866294,1.6117238,1.7368182,1.8619126,1.987007,2.1121013,1.7676386,1.4231756,1.0768998,0.7324369,0.387974,0.9155461,1.4431182,1.9706904,2.4982624,3.0258346,2.5816586,2.1392958,1.696933,1.2545701,0.8122072,0.7541924,0.6979906,0.6399758,0.581961,0.52575916,0.6055295,0.6852999,0.7650702,0.8448406,0.9246109,1.1657349,1.405046,1.6443571,1.8854811,2.124792,1.8673514,1.6099107,1.35247,1.0950294,0.8375887,1.2527572,1.6679256,2.0830941,2.4982624,2.911618,2.8445382,2.7774587,2.7103791,2.6432993,2.5744069,2.374981,2.175555,1.9743162,1.7748904,1.5754645,1.3125849,1.0497054,0.7868258,0.52575916,0.26287958,0.40429065,0.5475147,0.69073874,0.8321498,0.97537386,0.83940166,0.70524246,0.56927025,0.43511102,0.2991388,0.23931105,0.1794833,0.11965553,0.059827764,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.70524246,1.3343405,1.9652514,2.5943494,3.2252605,2.7720199,2.3205922,1.8673514,1.4141108,0.96268314,2.4348087,3.9069343,5.3808727,6.8529987,8.325124,9.376642,10.429974,11.483305,12.534823,13.588155,14.275268,14.96238,15.649493,16.336605,17.025532,15.620485,14.21544,12.810393,11.405348,10.000301,8.239915,6.4795284,4.7191415,2.960568,1.2001812,11.127964,21.053934,30.98353,40.9095,50.837284,41.493275,32.147453,22.80163,13.457622,4.1117992,4.40006,4.688321,4.974769,5.2630305,5.5494785,5.9320135,6.3145485,6.697084,7.079619,7.462154,7.021604,6.582867,6.1423173,5.7017674,5.2630305,6.2782893,7.2917356,8.306994,9.322253,10.337513,10.127209,9.916905,9.706602,9.498111,9.287807,9.664904,10.042,10.419096,10.798005,11.175101,9.420154,7.665206,5.910258,4.15531,2.4003625,3.6694362,4.940323,6.209397,7.4802837,8.749357,7.1630154,5.57486,3.9867048,2.4003625,0.8122072,1.745883,2.6777458,3.6096084,4.5432844,5.475147,5.1107416,4.744523,4.3801174,4.0157123,3.6494937,3.3449159,3.0403383,2.7357605,2.42937,2.124792,1.7041848,1.2853905,0.86478317,0.44417584,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.1794833,0.36077955,0.5402629,0.7197462,0.89922947,0.9354887,0.969935,1.0043813,1.0406405,1.0750868,1.0297627,0.98443866,0.93911463,0.89560354,0.85027945,1.2853905,1.7205015,2.1556125,2.5907235,3.0258346,2.8971143,2.770207,2.6432993,2.514579,2.3876717,1.9579996,1.5283275,1.0968424,0.6671702,0.2374981,0.37528324,0.51306844,0.6508536,0.7868258,0.9246109,0.85027945,0.774135,0.69980353,0.62547207,0.5493277,1.0605831,1.5700256,2.079468,2.5907235,3.100166,3.3050308,3.5098956,3.7147603,3.919625,4.12449,3.7492065,3.3757362,3.000453,2.6251698,2.2498865,2.6469254,3.045777,3.442816,3.8398547,4.2368937,4.3166637,4.3982472,4.478018,4.557788,4.6375585,5.351866,6.0679855,6.782293,7.498413,8.212721,7.6380115,7.063302,6.48678,5.9120708,5.337362,4.940323,4.5432844,4.1444325,3.7473936,3.350355,3.3177216,3.2850883,3.2524548,3.2198215,3.1871881,2.7575161,2.327844,1.8981718,1.4666867,1.0370146,0.83033687,0.62184614,0.41516843,0.20667773,0.0,0.1794833,0.36077955,0.5402629,0.7197462,0.89922947,0.9101072,0.91917205,0.9300498,0.93911463,0.9499924,0.7705091,0.58921283,0.40972954,0.23024625,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.18492219,0.36984438,0.55476654,0.73968875,0.9246109,0.73968875,0.55476654,0.36984438,0.18492219,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08339628,0.16497959,0.24837588,0.32995918,0.41335547,0.32995918,0.24837588,0.16497959,0.08339628,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14503701,0.29007402,0.43511102,0.58014804,0.72518504,0.88291276,1.0406405,1.1983683,1.3542831,1.5120108,1.8582866,2.2027495,2.5472124,2.8916752,3.2379513,3.4301252,3.6222992,3.8144734,4.006647,4.2006345,4.856927,5.5150323,6.1731377,6.82943,7.4875355,6.169512,4.853301,3.5352771,2.2172532,0.89922947,0.7505665,0.6000906,0.44961473,0.2991388,0.15047589,0.16497959,0.1794833,0.19579996,0.21030366,0.22480737,0.19579996,0.16497959,0.13415924,0.10515183,0.07433146,0.32995918,0.5855869,0.83940166,1.0950294,1.3506571,1.0841516,0.8194591,0.55476654,0.29007402,0.025381476,0.11784257,0.21030366,0.30276474,0.39522585,0.48768693,0.48043507,0.47318324,0.46411842,0.45686656,0.44961473,0.36440548,0.27919623,0.19579996,0.11059072,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13415924,0.27013144,0.40429065,0.5402629,0.6744221,1.7041848,2.7357605,3.7655232,4.795286,5.825049,5.906632,5.9900284,6.071612,6.155008,6.2384043,7.3769445,8.517298,9.657652,10.798005,11.938358,12.184921,12.433297,12.67986,12.928236,13.174799,11.655537,10.13446,8.615198,7.0959353,5.57486,9.672155,13.771264,17.866747,21.96404,26.06315,24.9373,23.811451,22.687414,21.563377,20.437527,19.235533,18.031725,16.829731,15.627737,14.425743,13.417736,12.409729,11.401722,10.395528,9.38752,9.063,8.736667,8.412147,8.087626,7.763106,8.002417,8.241728,8.482852,8.722163,8.963287,8.729415,8.497355,8.265296,8.033237,7.799365,11.358211,14.915243,18.472277,22.029308,25.588154,22.89953,20.212719,17.524096,14.837286,12.1504755,11.622903,11.095331,10.567759,10.040187,9.512614,8.495543,7.476658,6.4595857,5.4425135,4.4254417,4.421816,4.420003,4.41819,4.4145637,4.4127507,19.474844,19.182957,18.889257,10258.0,18.305483,18.011784,18.361685,18.711586,19.063301,19.413204,19.763105,19.442211,19.123129,18.802235,18.483154,18.16226,16.664753,15.167245,13.669738,12.172231,10.674724,9.837135,8.999546,8.161958,7.324369,6.48678,6.26016,6.0317264,5.805106,5.576673,5.3500524,5.473334,5.5948024,5.718084,5.8395524,5.962834,4.985647,4.006647,3.0294604,2.0522738,1.0750868,1.3379664,1.6008459,1.8619126,2.124792,2.3876717,1.9706904,1.551896,1.1349145,0.7179332,0.2991388,0.872035,1.4449311,2.0178273,2.5907235,3.1618068,2.7683938,2.373168,1.9779422,1.5827163,1.1874905,1.020698,0.8520924,0.6852999,0.5166943,0.34990177,0.5076295,0.6653573,0.823085,0.9808127,1.1367276,1.54827,1.9579996,2.3677292,2.7774587,3.1871881,2.7955883,2.4021754,2.0105755,1.6171626,1.2255627,1.5591478,1.8945459,2.229944,2.565342,2.9007401,2.8300345,2.759329,2.6904364,2.619731,2.5508385,2.4130533,2.275268,2.137483,1.9996977,1.8619126,1.5373923,1.2128719,0.8883517,0.5620184,0.2374981,0.3208944,0.40247768,0.48587397,0.56745726,0.6508536,0.56020546,0.46955732,0.38072214,0.29007402,0.19942589,0.15954071,0.11965553,0.07977036,0.03988518,0.0,0.0,0.0,0.0,0.0,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.52032024,0.92823684,1.3343405,1.742257,2.1501737,1.9525607,1.7549478,1.5573349,1.3597219,1.162109,2.2897718,3.4174345,4.5450974,5.67276,6.8004227,8.31062,9.820818,11.329204,12.839401,14.349599,14.762955,15.174497,15.5878525,15.999394,16.41275,14.880796,13.347031,11.815077,10.283124,8.749357,7.309865,5.870373,4.4290676,2.9895754,1.550083,8.259857,14.969632,21.679407,28.390993,35.10077,29.308353,23.515938,17.721708,11.929294,6.1368785,5.8504305,5.562169,5.275721,4.98746,4.699199,5.092612,5.484212,5.8776245,6.2692246,6.6626377,6.590119,6.5176005,6.445082,6.3725634,6.300045,6.5592985,6.8203654,7.079619,7.3406854,7.5999393,7.322556,7.0451727,6.7677894,6.490406,6.2130227,6.4595857,6.7079616,6.9545245,7.2029004,7.4494634,6.2801023,5.1107416,3.9395678,2.770207,1.6008459,2.6922495,3.785466,4.876869,5.9700856,7.063302,5.8758116,4.688321,3.5008307,2.3133402,1.1258497,1.6298534,2.13567,2.6396735,3.1454902,3.6494937,4.0157123,4.3801174,4.744523,5.1107416,5.475147,5.0182805,4.559601,4.102734,3.6458678,3.1871881,2.5580902,1.9271792,1.2980812,0.6671702,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.27013144,0.5402629,0.8103943,1.0805258,1.3506571,1.403233,1.455809,1.5083848,1.5591478,1.6117238,1.5446441,1.4775645,1.4104849,1.3415923,1.2745126,1.6026589,1.9308052,2.2571385,2.5852847,2.911618,2.7266958,2.5417736,2.3568513,2.1719291,1.987007,1.6298534,1.2726997,0.9155461,0.55839247,0.19942589,0.34990177,0.50037766,0.6508536,0.7995165,0.9499924,0.9119202,0.87566096,0.8375887,0.7995165,0.76325727,1.5392052,2.3169663,3.094727,3.872488,4.650249,4.2949085,3.9395678,3.584227,3.2306993,2.8753586,2.5997884,2.324218,2.0504606,1.7748904,1.49932,1.889107,2.280707,2.6704938,3.0602808,3.4500678,3.6948178,3.9395678,4.1843176,4.4308805,4.6756306,5.7217097,6.7696023,7.817495,8.865387,9.91328,9.137331,8.363196,7.5872483,6.813113,6.037165,5.560356,5.081734,4.604925,4.1281157,3.6494937,3.482701,3.3159087,3.147303,2.9805105,2.811905,2.3931105,1.9725033,1.551896,1.1331016,0.7124943,0.56927025,0.42785916,0.28463513,0.14322405,0.0,0.27013144,0.5402629,0.8103943,1.0805258,1.3506571,1.3651608,1.3796645,1.3941683,1.4104849,1.4249886,1.1548572,0.88472575,0.61459434,0.3444629,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.15228885,0.3045777,0.45686656,0.6091554,0.76325727,0.6091554,0.45686656,0.3045777,0.15228885,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.22480737,0.1794833,0.13415924,0.09064813,0.045324065,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.054388877,0.11059072,0.16497959,0.21936847,0.2755703,0.21936847,0.16497959,0.11059072,0.054388877,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.10515183,0.21030366,0.3154555,0.42060733,0.52575916,0.70524246,0.88472575,1.064209,1.2455053,1.4249886,1.742257,2.0595255,2.3767939,2.6958754,3.0131438,3.1581807,3.303218,3.4482548,3.5932918,3.738329,5.2050157,6.6717024,8.140202,9.606889,11.075388,9.130079,7.1847706,5.239462,3.294153,1.3506571,1.1004683,0.85027945,0.6000906,0.34990177,0.099712946,0.11059072,0.11965553,0.13053331,0.13959812,0.15047589,0.13053331,0.11059072,0.09064813,0.07070554,0.05076295,0.21936847,0.38978696,0.56020546,0.7306239,0.89922947,0.726998,0.55476654,0.3825351,0.21030366,0.038072214,0.17041849,0.30276474,0.43511102,0.56745726,0.69980353,0.64541465,0.58921283,0.53482395,0.48043507,0.42423326,0.3480888,0.27013144,0.19217403,0.11421664,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.09064813,0.1794833,0.27013144,0.36077955,0.44961473,1.258196,2.0649643,2.8717327,3.680314,4.4870825,4.8170414,5.147001,5.47696,5.806919,6.1368785,7.6724577,9.208037,10.741803,12.277383,13.812962,13.789393,13.767638,13.745882,13.722314,13.700559,12.331772,10.964798,9.597824,8.23085,6.8620634,9.177217,11.49237,13.807523,16.122677,18.43783,19.63801,20.838192,22.038374,23.236742,24.436922,23.414412,22.391901,21.36939,20.34688,19.324368,17.944704,16.565039,15.185374,13.80571,12.4242325,11.849524,11.274815,10.700105,10.125396,9.550687,9.347635,9.144584,8.943344,8.740293,8.537241,8.207282,7.877322,7.5473633,7.217404,6.887445,9.068439,11.24762,13.426801,15.607795,17.786976,16.487082,15.187187,13.887294,12.5873995,11.287505,11.628342,11.967366,12.308203,12.647227,12.988064,11.566701,10.147152,8.727602,7.308052,5.8866897,5.5531044,5.217706,4.882308,4.5469103,4.213325,19.487535,19.485722,19.482096,19.480284,19.476658,19.474844,19.786674,20.100317,20.412146,20.725788,21.037619,20.589815,20.142014,19.694212,19.248224,18.800423,17.52047,16.240519,14.960567,13.680615,12.400664,11.512312,10.625773,9.737422,8.8508835,7.9625316,7.6797094,7.3968873,7.115878,6.833056,6.550234,6.542982,6.53573,6.526665,6.5194135,6.5121617,5.3428006,4.17344,3.002266,1.8329052,0.66173136,1.062396,1.4630609,1.8619126,2.2625773,2.663242,2.1719291,1.6824293,1.1929294,0.7016165,0.21211663,0.83033687,1.4467441,2.0649643,2.6831846,3.299592,2.953316,2.6052272,2.2571385,1.9108626,1.5627737,1.2853905,1.0080072,0.7306239,0.45324063,0.17585737,0.40972954,0.64541465,0.8792868,1.114972,1.3506571,1.9308052,2.5091403,3.0892882,3.6694362,4.249584,3.7220123,3.1944401,2.666868,2.1392958,1.6117238,1.8673514,2.1229792,2.3767939,2.6324217,2.8880494,2.8155308,2.7430124,2.6704938,2.5979755,2.525457,2.4493124,2.374981,2.3006494,2.2245052,2.1501737,1.7621996,1.3742256,0.9880646,0.6000906,0.21211663,0.23568514,0.2574407,0.27919623,0.30276474,0.3245203,0.27919623,0.23568514,0.19036107,0.14503701,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0,0.0,0.0,0.0,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.33539808,0.52032024,0.70524246,0.8901646,1.0750868,1.1331016,1.1893034,1.2473183,1.305333,1.3633479,2.1447346,2.9279346,3.7093215,4.4925213,5.275721,7.2427855,9.20985,11.176914,13.145792,15.112856,15.250641,15.386614,15.524399,15.662184,15.799969,14.139296,12.480434,10.81976,9.159087,7.500226,6.379815,5.2594047,4.1408067,3.0203958,1.8999848,5.391751,8.885329,12.377095,15.870674,19.36244,17.121618,14.882609,12.6417885,10.40278,8.161958,7.3008003,6.43783,5.57486,4.7118897,3.8507326,4.25321,4.655688,5.0581656,5.4606433,5.863121,6.156821,6.452334,6.7478466,7.0433598,7.3370595,6.8421206,6.347182,5.8522434,5.3573046,4.8623657,4.517903,4.171627,3.827164,3.482701,3.1382382,3.254268,3.3721104,3.489953,3.6077955,3.7256382,3.1400511,2.5544643,1.9706904,1.3851035,0.7995165,1.7150626,2.6306088,3.5443418,4.459888,5.375434,4.5867953,3.7999697,3.0131438,2.2245052,1.4376793,1.5156367,1.5917811,1.6697385,1.7476959,1.8256533,2.9206827,4.0157123,5.1107416,6.205771,7.3008003,6.6898317,6.0806766,5.469708,4.860553,4.249584,3.4101827,2.570781,1.7295663,0.8901646,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.36077955,0.7197462,1.0805258,1.4394923,1.8002719,1.8691645,1.93987,2.0105755,2.079468,2.1501737,2.0595255,1.9706904,1.8800422,1.789394,1.7005589,1.9199274,2.1392958,2.3604772,2.5798457,2.7992141,2.5580902,2.3151531,2.0722163,1.8292793,1.5881553,1.3017071,1.017072,0.7324369,0.44780177,0.16316663,0.3245203,0.48768693,0.6508536,0.8122072,0.97537386,0.97537386,0.97537386,0.97537386,0.97537386,0.97537386,2.0196402,3.0657198,4.1099863,5.1542525,6.200332,5.2847857,4.36924,3.4555066,2.5399606,1.6244144,1.4503701,1.2745126,1.1004683,0.9246109,0.7505665,1.1331016,1.5156367,1.8981718,2.280707,2.663242,3.0729716,3.482701,3.8924308,4.3021603,4.7118897,6.093367,7.473032,8.852696,10.232361,11.612025,10.636651,9.663091,8.6877165,7.7123427,6.736969,6.1803894,5.621997,5.0654173,4.507025,3.9504454,3.6476808,3.3449159,3.0421512,2.7393866,2.4366217,2.0268922,1.6171626,1.2074331,0.79770356,0.387974,0.3100166,0.23205921,0.15410182,0.07795739,0.0,0.36077955,0.7197462,1.0805258,1.4394923,1.8002719,1.8202144,1.840157,1.8600996,1.8800422,1.8999848,1.5392052,1.1802386,0.8194591,0.4604925,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.03988518,0.07977036,0.11965553,0.15954071,0.19942589,0.15954071,0.11965553,0.07977036,0.03988518,0.0,0.11965553,0.23931105,0.36077955,0.48043507,0.6000906,0.48043507,0.36077955,0.23931105,0.11965553,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,0.2991388,0.23931105,0.1794833,0.11965553,0.059827764,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.027194439,0.054388877,0.08339628,0.11059072,0.13778515,0.11059072,0.08339628,0.054388877,0.027194439,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.065266654,0.13053331,0.19579996,0.25925365,0.3245203,0.5275721,0.7306239,0.9318628,1.1349145,1.3379664,1.6280404,1.9181144,2.2081885,2.4982624,2.7883365,2.8844235,2.9823234,3.0802233,3.1781235,3.2742105,5.5531044,7.8301854,10.107266,12.384347,14.663241,12.090648,9.518054,6.94546,4.3728657,1.8002719,1.4503701,1.1004683,0.7505665,0.40066472,0.05076295,0.054388877,0.059827764,0.065266654,0.07070554,0.07433146,0.065266654,0.054388877,0.045324065,0.034446288,0.025381476,0.11059072,0.19579996,0.27919623,0.36440548,0.44961473,0.36984438,0.29007402,0.21030366,0.13053331,0.05076295,0.2229944,0.39522585,0.56745726,0.73968875,0.9119202,0.8103943,0.7070554,0.6055295,0.50219065,0.40066472,0.32995918,0.25925365,0.19036107,0.11965553,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.045324065,0.09064813,0.13415924,0.1794833,0.22480737,0.8103943,1.3941683,1.9797552,2.565342,3.149116,3.727451,4.305786,4.882308,5.4606433,6.037165,7.9679704,9.896963,11.827768,13.75676,15.687565,15.3956785,15.101978,14.810091,14.518205,14.224504,13.009819,11.795135,10.58045,9.365765,8.149267,8.682278,9.215289,9.7483,10.279498,10.812509,14.336908,17.863121,21.38752,24.911919,28.438131,27.595104,26.752075,25.910862,25.067833,24.224806,22.471672,20.72035,18.967215,17.215893,15.462758,14.63786,13.812962,12.988064,12.163166,11.338268,10.692853,10.047439,9.402024,8.758422,8.113008,7.6851482,7.2572894,6.82943,6.4033837,5.975525,6.776854,7.5799966,8.383139,9.184468,9.987611,10.074633,10.161655,10.25049,10.337513,10.424535,11.631968,12.839401,14.046834,15.254267,16.4617,14.639673,12.817645,10.995618,9.171778,7.3497505,6.68258,6.01541,5.3482394,4.6792564,4.0120864,19.500225,19.786674,20.074934,20.363195,20.649643,20.937904,21.211662,21.487232,21.762802,22.038374,22.31213,21.737421,21.162712,20.588003,20.013294,19.436771,18.374376,17.31198,16.249584,15.187187,14.124791,13.1874895,12.250188,11.312886,10.375585,9.438283,9.099259,8.762048,8.424837,8.087626,7.750415,7.61263,7.474845,7.3370595,7.1992745,7.063302,5.6999545,4.3384194,2.9750717,1.6117238,0.25018883,0.7868258,1.3252757,1.8619126,2.4003625,2.9369993,2.374981,1.8129625,1.2491312,0.6871128,0.12509441,0.7868258,1.4503701,2.1121013,2.7756457,3.437377,3.1382382,2.8372865,2.5381477,2.2371957,1.938057,1.550083,1.162109,0.774135,0.387974,0.0,0.31182957,0.62547207,0.93730164,1.2491312,1.5627737,2.3133402,3.0620937,3.8126602,4.5632267,5.3119802,4.650249,3.9867048,3.3249733,2.663242,1.9996977,2.175555,2.3495996,2.525457,2.6995013,2.8753586,2.7992141,2.7248828,2.6505513,2.5744069,2.5000753,2.4873846,2.474694,2.4620032,2.4493124,2.4366217,1.987007,1.5373923,1.0877775,0.63816285,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.31182957,0.62547207,0.93730164,1.2491312,1.5627737,1.9996977,2.4366217,2.8753586,3.3122826,3.7492065,6.1749506,8.600695,11.024626,13.45037,15.8743,15.738328,15.600543,15.462758,15.324973,15.187187,13.399607,11.612025,9.824444,8.036863,6.249282,5.4497657,4.650249,3.8507326,3.049403,2.2498865,2.525457,2.7992141,3.0747845,3.350355,3.6241121,4.936697,6.249282,7.5618668,8.874452,10.1870365,8.749357,7.311678,5.8758116,4.4381323,3.000453,3.4119956,3.825351,4.2368937,4.650249,5.0617914,5.7253356,6.3870673,7.0506115,7.7123427,8.375887,7.124943,5.8758116,4.6248674,3.3757362,2.124792,1.7132497,1.2998942,0.8883517,0.4749962,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.73787576,1.4757515,2.2118144,2.94969,3.6875658,3.299592,2.911618,2.525457,2.137483,1.7495089,1.3996071,1.0497054,0.69980353,0.34990177,0.0,1.8256533,3.6494937,5.475147,7.3008003,9.12464,8.363196,7.5999393,6.836682,6.0752378,5.3119802,4.262275,3.2125697,2.1628644,1.1131591,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.44961473,0.89922947,1.3506571,1.8002719,2.2498865,2.3369088,2.4257438,2.5127661,2.5997884,2.6868105,2.5744069,2.4620032,2.3495996,2.2371957,2.124792,2.2371957,2.3495996,2.4620032,2.5744069,2.6868105,2.3876717,2.08672,1.7875811,1.4866294,1.1874905,0.97537386,0.76325727,0.5493277,0.33721104,0.12509441,0.2991388,0.4749962,0.6508536,0.824898,1.0007553,1.0370146,1.0750868,1.1131591,1.1494182,1.1874905,2.5000753,3.8126602,5.125245,6.43783,7.750415,6.2746634,4.800725,3.3249733,1.8492218,0.37528324,0.2991388,0.22480737,0.15047589,0.07433146,0.0,0.37528324,0.7505665,1.1258497,1.49932,1.8746033,2.4493124,3.0258346,3.6005437,4.175253,4.749962,6.4632115,8.174648,9.8878975,11.599335,13.312584,12.137785,10.962985,9.788185,8.613385,7.4367723,6.8004227,6.16226,5.524097,4.8877473,4.249584,3.8126602,3.3757362,2.9369993,2.5000753,2.0631514,1.6624867,1.261822,0.8629702,0.46230546,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.44961473,0.89922947,1.3506571,1.8002719,2.2498865,2.275268,2.3006494,2.324218,2.3495996,2.374981,1.9253663,1.4757515,1.0243238,0.5747091,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.0870222,0.17585737,0.26287958,0.34990177,0.43692398,0.34990177,0.26287958,0.17585737,0.0870222,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.12509441,0.18673515,0.25018883,0.31182957,0.37528324,0.2991388,0.22480737,0.15047589,0.07433146,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.34990177,0.5747091,0.7995165,1.0243238,1.2491312,1.5120108,1.7748904,2.03777,2.3006494,2.561716,2.612479,2.663242,2.712192,2.762955,2.811905,5.89938,8.9868555,12.07433,15.161806,18.24928,15.049402,11.849524,8.649645,5.4497657,2.2498865,1.8002719,1.3506571,0.89922947,0.44961473,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.2755703,0.48768693,0.69980353,0.9119202,1.1258497,0.97537386,0.824898,0.6744221,0.52575916,0.37528324,0.31182957,0.25018883,0.18673515,0.12509441,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.36259252,0.72518504,1.0877775,1.4503701,1.8129625,2.6378605,3.4627585,4.2876563,5.1125546,5.9374523,8.263483,10.587702,12.91192,15.23795,17.562168,17.00015,16.438131,15.8743,15.312282,14.750263,13.687867,12.625471,11.563075,10.500679,9.438283,8.187339,6.9382076,5.6872635,4.4381323,3.1871881,9.037619,14.888049,20.73848,26.587097,32.437527,31.775795,31.112251,30.45052,29.786976,29.125244,27.000452,24.873846,22.749054,20.624262,18.49947,17.424383,16.349297,15.27421,14.200936,13.125849,12.038072,10.950294,9.862516,8.774739,7.686961,7.1630154,6.637256,6.11331,5.5875506,5.0617914,4.4870825,3.9123733,3.3376641,2.762955,2.1882458,3.6621845,5.137936,6.6118746,8.087626,9.563377,11.637406,13.713249,15.787278,17.863121,19.93715,17.712645,15.486326,13.261822,11.037316,8.812811,7.8120556,6.813113,5.812358,4.8134155,3.8126602,17.725336,17.937452,18.149569,18.361685,18.575615,18.787731,18.635443,18.483154,18.329052,18.176764,18.024473,17.82686,17.629248,17.431635,17.235836,17.038223,16.565039,16.091856,15.620485,15.147303,14.674119,13.722314,12.770509,11.81689,10.865085,9.91328,9.498111,9.082943,8.667774,8.252605,7.837437,7.750415,7.663393,7.574558,7.4875355,7.400513,6.004532,4.610364,3.2143826,1.8202144,0.42423326,0.8194591,1.214685,1.6099107,2.0051367,2.4003625,2.0595255,1.7205015,1.3796645,1.0406405,0.69980353,1.4775645,2.2553256,3.0330863,3.8108473,4.5867953,4.135368,3.682127,3.2306993,2.7774587,2.324218,1.8655385,1.405046,0.9445535,0.48587397,0.025381476,0.3480888,0.67079616,0.9916905,1.3143979,1.6371052,2.2952106,2.953316,3.6096084,4.267714,4.9258194,4.2804046,3.63499,2.9895754,2.3441606,1.7005589,1.9217403,2.1447346,2.3677292,2.5907235,2.811905,2.7393866,2.666868,2.5943494,2.521831,2.4493124,2.4474995,2.4456866,2.4420607,2.4402475,2.4366217,1.9942589,1.551896,1.1095331,0.6671702,0.22480737,0.1794833,0.13415924,0.09064813,0.045324065,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.14503701,0.13959812,0.13415924,0.13053331,0.12509441,0.40791658,0.69073874,0.97174793,1.2545701,1.5373923,1.9507477,2.3622901,2.7756457,3.1871881,3.6005437,5.573047,7.5455503,9.518054,11.490557,13.46306,13.669738,13.878228,14.084907,14.291584,14.500074,12.823084,11.144281,9.467291,7.7903004,6.11331,5.8522434,5.5929894,5.331923,5.0726695,4.8134155,4.652062,4.4925213,4.3329806,4.171627,4.0120864,4.8623657,5.712645,6.5629244,7.413204,8.26167,7.9824743,7.703278,7.422269,7.1430726,6.8620634,6.6553855,6.446895,6.240217,6.0317264,5.825049,6.378002,6.929143,7.4820967,8.03505,8.588004,7.2899227,5.9918413,4.695573,3.397492,2.0994108,2.1048496,2.1102884,2.1157274,2.1193533,2.124792,1.7132497,1.2998942,0.8883517,0.4749962,0.06164073,0.058014803,0.052575916,0.047137026,0.04169814,0.038072214,0.99531645,1.9525607,2.909805,3.8670492,4.8242936,4.1897564,3.5552197,2.9206827,2.2843328,1.649796,1.4304274,1.209246,0.9898776,0.7705091,0.5493277,1.9054236,3.2597067,4.615803,5.9700856,7.324369,7.6597667,7.995165,8.330563,8.665961,8.999546,7.217404,5.4352617,3.6531196,1.8691645,0.0870222,0.08339628,0.07795739,0.072518505,0.06707962,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.36984438,0.73968875,1.1095331,1.4793775,1.8492218,1.9906329,2.1302311,2.269829,2.4094272,2.5508385,2.3949237,2.2408218,2.084907,1.9308052,1.7748904,1.8673514,1.9598125,2.0522738,2.1447346,2.2371957,2.132044,2.0268922,1.9217403,1.8184015,1.7132497,1.7205015,1.7277533,1.7350051,1.742257,1.7495089,1.7730774,1.794833,1.8184015,1.840157,1.8619126,1.8184015,1.7730774,1.7277533,1.6824293,1.6371052,2.5580902,3.4772623,4.3982472,5.317419,6.2365913,5.049101,3.8616104,2.6741197,1.4866294,0.2991388,0.42423326,0.5493277,0.6744221,0.7995165,0.9246109,1.6171626,2.3097143,3.002266,3.6948178,4.3873696,5.139749,5.8921285,6.644508,7.3968873,8.149267,8.972352,9.795437,10.616709,11.439794,12.262879,11.108022,9.953164,8.798307,7.6416373,6.48678,5.870373,5.2521524,4.6357455,4.017525,3.3993049,3.049403,2.6995013,2.3495996,1.9996977,1.649796,1.3307146,1.0098201,0.69073874,0.36984438,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.36077955,0.7197462,1.0805258,1.4394923,1.8002719,1.8256533,1.8492218,1.8746033,1.8999848,1.9253663,1.5772774,1.2291887,0.88291276,0.53482395,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.03988518,0.07977036,0.11965553,0.15954071,0.19942589,0.2229944,0.24474995,0.26831847,0.29007402,0.31182957,0.3208944,0.32814622,0.33539808,0.34264994,0.34990177,0.2955129,0.23931105,0.18492219,0.13053331,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.018129626,0.034446288,0.052575916,0.07070554,0.0870222,0.13053331,0.17223145,0.21574254,0.2574407,0.2991388,0.23931105,0.1794833,0.11965553,0.059827764,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.027194439,0.054388877,0.08339628,0.11059072,0.13778515,0.11059072,0.08339628,0.054388877,0.027194439,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.059827764,0.058014803,0.054388877,0.052575916,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,1.2019942,2.2933977,3.3829882,4.4725785,5.562169,5.522284,5.482399,5.4425135,5.4026284,5.3627434,5.823236,6.281915,6.742408,7.2029004,7.663393,10.034748,12.407916,14.779271,17.15244,19.525606,16.623055,13.720501,10.817947,7.915395,5.0128417,4.4798307,3.9468195,3.4156215,2.8826106,2.3495996,1.983381,1.6153497,1.2473183,0.8792868,0.51306844,0.51306844,0.51306844,0.51306844,0.51306844,0.51306844,0.48043507,0.44780177,0.41516843,0.3825351,0.34990177,0.35715362,0.36440548,0.37165734,0.38072214,0.387974,0.52213323,0.65810543,0.79226464,0.92823684,1.062396,0.95180535,0.8430276,0.7324369,0.62184614,0.51306844,0.44780177,0.3825351,0.31726846,0.2520018,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.29007402,0.58014804,0.87022203,1.1602961,1.4503701,2.3079014,3.1654327,4.022964,4.880495,5.7380266,7.5999393,9.461852,11.325577,13.1874895,15.049402,14.694061,14.340534,13.985193,13.629852,13.274512,12.692551,12.11059,11.526816,10.944855,10.362894,9.329506,8.29793,7.264541,6.2329655,5.199577,9.958604,14.715817,19.473032,24.230246,28.98746,28.070099,27.15274,26.235382,25.318022,24.400663,22.90497,21.409275,19.915394,18.4197,16.92582,16.162561,15.399304,14.63786,13.874602,13.113158,12.07977,11.048194,10.014805,8.98323,7.949841,7.83925,7.7304726,7.6198816,7.509291,7.400513,6.58468,5.77066,4.954827,4.1408067,3.3249733,4.2423325,5.1596913,6.0770507,6.9944096,7.911769,9.702975,11.49237,13.281764,15.072971,16.862366,15.189,13.517449,11.844085,10.172533,8.499168,8.00423,7.509291,7.0143523,6.5194135,6.0244746,15.950445,16.08823,16.224201,16.361988,16.499773,16.637558,16.05741,15.477262,14.897114,14.316965,13.736817,13.918114,14.097597,14.277081,14.458377,14.63786,14.755702,14.871732,14.989574,15.107417,15.22526,14.257137,13.290829,12.322706,11.354585,10.388275,9.89515,9.402024,8.910711,8.417585,7.9244595,7.8882003,7.850128,7.8120556,7.7757964,7.7377243,6.3109226,4.882308,3.4555066,2.0268922,0.6000906,0.8520924,1.1040943,1.357909,1.6099107,1.8619126,1.745883,1.6280404,1.5101979,1.3923552,1.2745126,2.1683033,3.0602808,3.9522583,4.844236,5.7380266,5.132497,4.5269675,3.923251,3.3177216,2.712192,2.179181,1.647983,1.114972,0.581961,0.05076295,0.3825351,0.71430725,1.0478923,1.3796645,1.7132497,2.277081,2.8427253,3.4083695,3.972201,4.537845,3.9105604,3.2832751,2.6541772,2.0268922,1.3996071,1.6697385,1.93987,2.2100015,2.4801328,2.7502642,2.6795588,2.610666,2.5399606,2.469255,2.4003625,2.4076142,2.4148662,2.422118,2.42937,2.4366217,2.0033236,1.5682126,1.1331016,0.6979906,0.26287958,0.21030366,0.15772775,0.10515183,0.052575916,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.13959812,0.16679256,0.19579996,0.2229944,0.25018883,0.50219065,0.7541924,1.0080072,1.260009,1.5120108,1.8999848,2.2879589,2.6741197,3.0620937,3.4500678,4.9693303,6.490406,8.009668,9.530745,11.050007,11.602961,12.154101,12.707055,13.260008,13.812962,12.244749,10.6783495,9.110137,7.5419245,5.975525,6.2547207,6.53573,6.814926,7.0941224,7.3751316,6.78048,6.185828,5.5893636,4.994712,4.40006,4.788034,5.1741953,5.562169,5.9501433,6.338117,7.215591,8.093065,8.970539,9.848013,10.725487,9.896963,9.070251,8.241728,7.415017,6.588306,7.0306687,7.473032,7.915395,8.357758,8.80012,7.454902,6.109684,4.764466,3.4192474,2.0758421,2.4982624,2.9206827,3.343103,3.7655232,4.1879435,3.3757362,2.561716,1.7495089,0.93730164,0.12509441,0.11421664,0.10515183,0.09427405,0.08520924,0.07433146,1.2527572,2.42937,3.6077955,4.784408,5.962834,5.0799212,4.1970086,3.3140955,2.4329958,1.550083,1.4594349,1.3705997,1.2799516,1.1893034,1.1004683,1.9851941,2.8699198,3.7546456,4.6393714,5.524097,6.9581504,8.39039,9.822631,11.254871,12.687112,10.172533,7.6579537,5.141562,2.6269827,0.11240368,0.10333887,0.092461094,0.08339628,0.072518505,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.29007402,0.58014804,0.87022203,1.1602961,1.4503701,1.6425442,1.8347181,2.0268922,2.220879,2.4130533,2.2154403,2.0178273,1.8202144,1.6226015,1.4249886,1.4975071,1.5700256,1.6425442,1.7150626,1.7875811,1.8782293,1.9670644,2.0577126,2.1483607,2.2371957,2.465629,2.6922495,2.9206827,3.147303,3.3757362,3.245203,3.1146698,2.9841363,2.855416,2.7248828,2.5979755,2.469255,2.3423476,2.2154403,2.08672,2.6142921,3.141864,3.6694362,4.1970086,4.7245803,3.825351,2.9243085,2.0250793,1.1258497,0.22480737,0.5493277,0.87566096,1.2001812,1.5247015,1.8492218,2.8608549,3.870675,4.880495,5.8903155,6.9001355,7.8301854,8.760235,9.690285,10.620335,11.5503845,11.483305,11.4144125,11.347333,11.280253,11.213174,10.078259,8.943344,7.806617,6.6717024,5.5367875,4.940323,4.3420453,3.7455807,3.147303,2.5508385,2.2879589,2.0250793,1.7621996,1.49932,1.2382535,0.99712944,0.75781834,0.5166943,0.27738327,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.27013144,0.5402629,0.8103943,1.0805258,1.3506571,1.3742256,1.3996071,1.4249886,1.4503701,1.4757515,1.2291887,0.98443866,0.73968875,0.4949388,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.24474995,0.34083697,0.43511102,0.5293851,0.62547207,0.5529536,0.48043507,0.40791658,0.33539808,0.26287958,0.23931105,0.21755551,0.19579996,0.17223145,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.13415924,0.15772775,0.1794833,0.2030518,0.22480737,0.1794833,0.13415924,0.09064813,0.045324065,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.054388877,0.11059072,0.16497959,0.21936847,0.2755703,0.21936847,0.16497959,0.11059072,0.054388877,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.11965553,0.11421664,0.11059072,0.10515183,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0,0.0,0.0,0.0,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,2.0558996,4.0102735,5.964647,7.9208336,9.875207,9.5325575,9.189907,8.847258,8.504607,8.161958,9.03218,9.902402,10.772624,11.642846,12.513068,14.170115,15.827164,17.484211,19.143072,20.80012,18.194893,15.589665,12.984438,10.37921,7.7757964,7.159389,6.544795,5.9302006,5.315606,4.699199,3.9649491,3.2306993,2.4946365,1.7603867,1.0243238,1.0243238,1.0243238,1.0243238,1.0243238,1.0243238,0.96087015,0.89560354,0.83033687,0.7650702,0.69980353,0.7016165,0.70524246,0.7070554,0.7106813,0.7124943,0.7705091,0.82671094,0.88472575,0.94274056,1.0007553,0.9300498,0.85934424,0.7904517,0.7197462,0.6508536,0.581961,0.5148814,0.44780177,0.38072214,0.31182957,0.25018883,0.18673515,0.12509441,0.06164073,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.21755551,0.43511102,0.6526665,0.87022203,1.0877775,1.9779422,2.8681068,3.7582715,4.646623,5.5367875,6.9382076,8.337815,9.737422,11.137029,12.536636,12.389787,12.242936,12.094274,11.947423,11.800573,11.697234,11.595709,11.49237,11.390844,11.287505,10.471672,9.657652,8.841819,8.027799,7.211965,10.877775,14.543586,18.207582,21.87158,25.537392,24.364405,23.19323,22.020243,20.847258,19.67427,18.809486,17.944704,17.07992,16.215137,15.350354,14.90074,14.449312,13.999697,13.550082,13.100468,12.123281,11.144281,10.167094,9.189907,8.212721,8.517298,8.821876,9.128266,9.432844,9.737422,8.682278,7.6271334,6.5719895,5.516845,4.461701,4.8224807,5.18326,5.542227,5.903006,6.261973,7.7667317,9.273304,10.778063,12.282822,13.7875805,12.66717,11.546759,10.428161,9.30775,8.187339,8.198216,8.207282,8.21816,8.227224,8.238102,14.175554,14.237195,14.300649,14.362289,14.425743,14.487384,13.479377,12.473183,11.465176,10.457169,9.449161,10.007553,10.564133,11.122525,11.680918,12.237497,12.944552,13.651608,14.3604765,15.067532,15.774588,14.791962,13.809336,12.826711,11.844085,10.863272,10.292189,9.7229185,9.151835,8.582565,8.013294,8.024173,8.036863,8.049554,8.062244,8.074935,6.6155005,5.1542525,3.6948178,2.2353828,0.774135,0.88472575,0.99531645,1.1059072,1.214685,1.3252757,1.4304274,1.5355793,1.6407311,1.745883,1.8492218,2.857229,3.8652363,4.8732433,5.8794374,6.887445,6.1296263,5.371808,4.615803,3.8579843,3.100166,2.4946365,1.8909199,1.2853905,0.67986095,0.07433146,0.4169814,0.75963134,1.1022812,1.4449311,1.7875811,2.2607644,2.7321346,3.2053177,3.6766882,4.1498713,3.540716,2.9297476,2.3205922,1.7096237,1.1004683,1.4177368,1.7350051,2.0522738,2.3695421,2.6868105,2.619731,2.5526514,2.4855716,2.4166791,2.3495996,2.3677292,2.3858588,2.4021754,2.420305,2.4366217,2.0105755,1.5827163,1.1548572,0.726998,0.2991388,0.23931105,0.1794833,0.11965553,0.059827764,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.13415924,0.19579996,0.25562772,0.3154555,0.37528324,0.5982776,0.8194591,1.0424535,1.2654479,1.4866294,1.8492218,2.2118144,2.5744069,2.9369993,3.299592,4.367427,5.4352617,6.5030966,7.570932,8.636953,9.53437,10.431787,11.329204,12.22662,13.125849,11.668227,10.210606,8.752983,7.2953615,5.8377395,6.6571984,7.476658,8.29793,9.117389,9.936848,8.907085,7.877322,6.8475595,5.8177967,4.788034,4.7118897,4.6375585,4.5632267,4.4870825,4.4127507,6.446895,8.482852,10.516996,12.552953,14.587097,13.140353,11.691795,10.245051,8.798307,7.3497505,7.6833353,8.015107,8.34688,8.680465,9.012237,7.6198816,6.2275267,4.835171,3.442816,2.0504606,2.8898623,3.729264,4.5704784,5.40988,6.249282,5.038223,3.825351,2.612479,1.3996071,0.18673515,0.17223145,0.15772775,0.14322405,0.12690738,0.11240368,1.5101979,2.907992,4.305786,5.7017674,7.0995617,5.9700856,4.84061,3.7093215,2.5798457,1.4503701,1.4902552,1.5301404,1.5700256,1.6099107,1.649796,2.0649643,2.4801328,2.8953013,3.3104696,3.7256382,6.2547207,8.785617,11.314699,13.845595,16.374678,13.127662,9.880646,6.6318173,3.3848011,0.13778515,0.12328146,0.10696479,0.092461094,0.07795739,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.21030366,0.42060733,0.630911,0.83940166,1.0497054,1.2944553,1.5392052,1.7857682,2.030518,2.275268,2.034144,1.794833,1.5555218,1.3143979,1.0750868,1.1276628,1.1802386,1.2328146,1.2853905,1.3379664,1.6226015,1.9072367,2.1918716,2.47832,2.762955,3.2107568,3.6567454,4.1045475,4.552349,5.0001507,4.7173285,4.4345064,4.1516843,3.870675,3.587853,3.3775494,3.1672456,2.956942,2.7466383,2.5381477,2.6723068,2.808279,2.9424384,3.0784104,3.2125697,2.5997884,1.987007,1.3742256,0.76325727,0.15047589,0.6744221,1.2001812,1.7241274,2.2498865,2.7756457,4.102734,5.429823,6.7569118,8.0858135,9.412902,10.520622,11.628342,12.734249,13.8419695,14.94969,13.992445,13.035201,12.077957,11.120712,10.161655,9.046683,7.931711,6.816739,5.7017674,4.5867953,4.0102735,3.4319382,2.855416,2.277081,1.7005589,1.5247015,1.3506571,1.1747998,1.0007553,0.824898,0.6653573,0.5058166,0.3444629,0.18492219,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.1794833,0.36077955,0.5402629,0.7197462,0.89922947,0.9246109,0.9499924,0.97537386,1.0007553,1.0243238,0.88291276,0.73968875,0.5982776,0.4550536,0.31182957,0.25018883,0.18673515,0.12509441,0.06164073,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.26831847,0.43511102,0.60190356,0.7705091,0.93730164,0.7850128,0.6327239,0.48043507,0.32814622,0.17585737,0.18492219,0.19579996,0.20486477,0.21574254,0.22480737,0.1794833,0.13415924,0.09064813,0.045324065,0.0,0.027194439,0.054388877,0.08339628,0.11059072,0.13778515,0.13959812,0.14322405,0.14503701,0.14684997,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.09064813,0.06707962,0.045324065,0.02175555,0.0,0.08339628,0.16497959,0.24837588,0.32995918,0.41335547,0.32995918,0.24837588,0.16497959,0.08339628,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.1794833,0.17223145,0.16497959,0.15772775,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.0,0.0,0.0,0.0,0.0,0.018129626,0.034446288,0.052575916,0.07070554,0.0870222,2.907992,5.727149,8.548119,11.367275,14.188245,13.54283,12.897416,12.252001,11.606586,10.962985,12.242936,13.522888,14.802839,16.08279,17.362743,18.305483,19.248224,20.189152,21.131891,22.074633,19.766731,17.460642,15.152741,12.84484,10.536939,9.840761,9.142771,8.444779,7.746789,7.0506115,5.9465175,4.844236,3.7419548,2.6396735,1.5373923,1.5373923,1.5373923,1.5373923,1.5373923,1.5373923,1.4394923,1.3434052,1.2455053,1.1476053,1.0497054,1.0478923,1.0442665,1.0424535,1.0406405,1.0370146,1.017072,0.99712944,0.97718686,0.9572442,0.93730164,0.90829426,0.8774739,0.8466535,0.81764615,0.7868258,0.7179332,0.64722764,0.57833505,0.5076295,0.43692398,0.34990177,0.26287958,0.17585737,0.0870222,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14503701,0.29007402,0.43511102,0.58014804,0.72518504,1.647983,2.570781,3.491766,4.4145637,5.337362,6.2746634,7.211965,8.149267,9.086569,10.025683,10.085511,10.145339,10.205167,10.264994,10.324821,10.701918,11.080828,11.457924,11.83502,12.212116,11.615651,11.017374,10.419096,9.822631,9.224354,11.7969475,14.369541,16.942135,19.514729,22.087322,20.660522,19.231907,17.805105,16.378304,14.94969,14.715817,14.480132,14.244447,14.010575,13.77489,13.637105,13.499319,13.363347,13.225562,13.087777,12.164979,11.242181,10.319383,9.398398,8.4756,9.195346,9.915092,10.634838,11.354585,12.07433,10.779876,9.48542,8.189152,6.8946967,5.600241,5.4026284,5.2050157,5.0074024,4.8097897,4.612177,5.8323007,7.0524244,8.272549,9.492672,10.712796,10.145339,9.577881,9.010424,8.442966,7.8755093,8.39039,8.9052725,9.420154,9.935035,10.449916,12.400664,12.387974,12.375282,12.362592,12.349901,12.337211,10.903157,9.467291,8.033237,6.5973706,5.163317,6.096993,7.0324817,7.9679704,8.901647,9.837135,11.135216,12.433297,13.729566,15.027647,16.325727,15.326786,14.329657,13.332527,12.335398,11.338268,10.689227,10.042,9.394773,8.747544,8.100317,8.161958,8.225411,8.287052,8.350506,8.412147,6.9200783,5.42801,3.9341288,2.4420607,0.9499924,0.91735905,0.88472575,0.8520924,0.8194591,0.7868258,1.114972,1.4431182,1.7694515,2.0975976,2.4257438,3.5479677,4.670192,5.7924156,6.9146395,8.036863,7.1267557,6.2166486,5.3083544,4.3982472,3.48814,2.810092,2.132044,1.455809,0.7777609,0.099712946,0.45324063,0.80495536,1.1566701,1.5101979,1.8619126,2.2426348,2.6233568,3.002266,3.3829882,3.7618973,3.1708715,2.5780327,1.9851941,1.3923552,0.7995165,1.1657349,1.5301404,1.8945459,2.2607644,2.6251698,2.5599031,2.4946365,2.42937,2.3641033,2.3006494,2.327844,2.3550384,2.382233,2.4094272,2.4366217,2.0178273,1.5972201,1.1766127,0.75781834,0.33721104,0.27013144,0.2030518,0.13415924,0.06707962,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.13053331,0.2229944,0.3154555,0.40791658,0.50037766,0.69255173,0.88472575,1.0768998,1.2708868,1.4630609,1.8002719,2.137483,2.474694,2.811905,3.149116,3.7655232,4.3801174,4.994712,5.6093063,6.2257137,7.4675927,8.709473,9.953164,11.195044,12.436923,11.089892,9.742861,8.39583,7.0469856,5.6999545,7.059676,8.419398,9.780933,11.1406555,12.500377,11.035503,9.570629,8.105756,6.640882,5.1741953,4.6375585,4.099108,3.5624714,3.0258346,2.4873846,5.6800117,8.872639,12.065266,15.257894,18.45052,16.38193,14.315152,12.246562,10.179785,8.113008,8.334189,8.557183,8.780178,9.003172,9.224354,7.7848616,6.345369,4.9040637,3.4645715,2.0250793,3.2832751,4.539658,5.7978544,7.0542374,8.312433,6.70071,5.087173,3.4754493,1.8619126,0.25018883,0.23024625,0.21030366,0.19036107,0.17041849,0.15047589,1.7676386,3.3848011,5.0019636,6.6209393,8.238102,6.8602505,5.482399,4.1045475,2.7266958,1.3506571,1.5192627,1.6896812,1.8600996,2.030518,2.1991236,2.1447346,2.0903459,2.034144,1.9797552,1.9253663,5.5531044,9.179029,12.806767,16.434505,20.062244,16.08279,12.103338,8.122072,4.1426196,0.16316663,0.14322405,0.12328146,0.10333887,0.08339628,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.13053331,0.25925365,0.38978696,0.52032024,0.6508536,0.9481794,1.2455053,1.5428312,1.840157,2.137483,1.8546607,1.5718386,1.2908293,1.0080072,0.72518504,0.75781834,0.7904517,0.823085,0.8557183,0.8883517,1.3669738,1.8474089,2.327844,2.808279,3.2869012,3.9558845,4.6230545,5.290225,5.957395,6.624565,6.189454,5.754343,5.319232,4.8841214,4.4508233,4.157123,3.8652363,3.5733492,3.2796493,2.9877625,2.7303216,2.472881,2.2154403,1.9579996,1.7005589,1.3742256,1.0497054,0.72518504,0.40066472,0.07433146,0.7995165,1.5247015,2.2498865,2.9750717,3.7002566,5.3446136,6.9907837,8.63514,10.279498,11.925668,13.209246,14.494636,15.780026,17.065416,18.350807,16.503399,14.654177,12.806767,10.959359,9.11195,8.01692,6.921891,5.826862,4.7318325,3.636803,3.0802233,2.521831,1.9652514,1.4068589,0.85027945,0.76325727,0.6744221,0.5873999,0.50037766,0.41335547,0.33177215,0.2520018,0.17223145,0.092461094,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.09064813,0.1794833,0.27013144,0.36077955,0.44961473,0.4749962,0.50037766,0.52575916,0.5493277,0.5747091,0.53482395,0.4949388,0.4550536,0.41516843,0.37528324,0.2991388,0.22480737,0.15047589,0.07433146,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.29007402,0.5293851,0.7705091,1.0098201,1.2491312,1.017072,0.7850128,0.5529536,0.3208944,0.0870222,0.13053331,0.17223145,0.21574254,0.2574407,0.2991388,0.23931105,0.1794833,0.11965553,0.059827764,0.0,0.032633327,0.065266654,0.09789998,0.13053331,0.16316663,0.14503701,0.12690738,0.11059072,0.092461094,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.11059072,0.21936847,0.32995918,0.4405499,0.5493277,0.4405499,0.32995918,0.21936847,0.11059072,0.0,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,0.23931105,0.23024625,0.21936847,0.21030366,0.19942589,0.15954071,0.11965553,0.07977036,0.03988518,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,3.7600844,7.4440246,11.129777,14.81553,18.49947,17.553104,16.604925,15.656745,14.710379,13.762199,15.45188,17.143373,18.833055,20.522736,22.212418,22.440851,22.66747,22.895905,23.122524,23.349146,21.340382,19.329807,17.319231,15.310469,13.299893,12.52032,11.740746,10.959359,10.179785,9.400211,7.9298983,6.4595857,4.989273,3.5207734,2.0504606,2.0504606,2.0504606,2.0504606,2.0504606,2.0504606,1.9199274,1.789394,1.6606737,1.5301404,1.3996071,1.3923552,1.3851035,1.3778516,1.3705997,1.3633479,1.2654479,1.167548,1.0696479,0.97174793,0.87566096,0.88472575,0.89560354,0.90466833,0.9155461,0.9246109,0.8520924,0.7795739,0.7070554,0.6345369,0.5620184,0.44961473,0.33721104,0.22480737,0.11240368,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.072518505,0.14503701,0.21755551,0.29007402,0.36259252,1.3180238,2.2716422,3.2270734,4.1825047,5.137936,5.612932,6.0879283,6.5629244,7.037921,7.512917,7.7794223,8.047741,8.314246,8.582565,8.8508835,9.708415,10.564133,11.421664,12.279196,13.136727,12.757817,12.377095,11.998186,11.617464,11.236742,12.717933,14.19731,15.676687,17.157877,18.637255,16.954826,15.272397,13.589968,11.907538,10.225109,10.620335,11.015561,11.410787,11.804199,12.199425,12.375282,12.549327,12.725184,12.899229,13.075087,12.206677,11.340081,10.471672,9.605076,8.736667,9.873394,11.008308,12.143224,13.278138,14.413053,12.877473,11.341894,9.808127,8.272549,6.736969,5.9827766,5.2267714,4.4725785,3.7183862,2.962381,3.8978696,4.8333583,5.767034,6.7025228,7.6380115,7.6216946,7.607191,7.592687,7.5781837,7.5618668,8.582565,9.603263,10.622148,11.642846,12.661731,10.625773,10.536939,10.449916,10.362894,10.275872,10.1870365,8.325124,6.4632115,4.599486,2.7375734,0.87566096,2.1882458,3.5008307,4.8134155,6.1241875,7.4367723,9.324066,11.213174,13.100468,14.9877615,16.875055,15.863422,14.849977,13.838344,12.824898,11.813264,11.088079,10.362894,9.637709,8.912524,8.187339,8.299743,8.412147,8.52455,8.636953,8.749357,7.224656,5.6999545,4.175253,2.6505513,1.1258497,0.9499924,0.774135,0.6000906,0.42423326,0.25018883,0.7995165,1.3506571,1.8999848,2.4493124,3.000453,4.2368937,5.475147,6.7134004,7.949841,9.188094,8.125698,7.063302,5.999093,4.936697,3.874301,3.1255474,2.374981,1.6244144,0.87566096,0.12509441,0.48768693,0.85027945,1.2128719,1.5754645,1.938057,2.2245052,2.5127661,2.7992141,3.0874753,3.3757362,2.7992141,2.2245052,1.649796,1.0750868,0.50037766,0.9119202,1.3252757,1.7368182,2.1501737,2.561716,2.5000753,2.4366217,2.374981,2.3133402,2.2498865,2.2879589,2.324218,2.3622901,2.4003625,2.4366217,2.0250793,1.6117238,1.2001812,0.7868258,0.37528324,0.2991388,0.22480737,0.15047589,0.07433146,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.12509441,0.25018883,0.37528324,0.50037766,0.62547207,0.7868258,0.9499924,1.1131591,1.2745126,1.4376793,1.7495089,2.0631514,2.374981,2.6868105,3.000453,3.1618068,3.3249733,3.48814,3.6494937,3.8126602,5.4008155,6.987158,8.575313,10.161655,11.74981,10.51337,9.275117,8.036863,6.8004227,5.562169,7.462154,9.362139,11.262123,13.162108,15.062093,13.162108,11.262123,9.362139,7.462154,5.562169,4.5632267,3.5624714,2.561716,1.5627737,0.5620184,4.9131284,9.262425,13.613536,17.962833,22.31213,19.62532,16.936697,14.249886,11.563075,8.874452,8.9868555,9.099259,9.211663,9.325879,9.438283,7.949841,6.4632115,4.974769,3.48814,1.9996977,3.6748753,5.3500524,7.02523,8.700407,10.375585,8.363196,6.350808,4.3366065,2.324218,0.31182957,0.28826106,0.26287958,0.2374981,0.21211663,0.18673515,2.0250793,3.8616104,5.6999545,7.5382986,9.374829,7.750415,6.1241875,4.499773,2.8753586,1.2491312,1.550083,1.8492218,2.1501737,2.4493124,2.7502642,2.2245052,1.7005589,1.1747998,0.6508536,0.12509441,4.8496747,9.574255,14.300649,19.025229,23.74981,19.03792,14.326031,9.612328,4.900438,0.18673515,0.16316663,0.13778515,0.11240368,0.0870222,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,0.6000906,0.9499924,1.2998942,1.649796,1.9996977,1.6751775,1.3506571,1.0243238,0.69980353,0.37528324,0.387974,0.40066472,0.41335547,0.42423326,0.43692398,1.1131591,1.7875811,2.4620032,3.1382382,3.8126602,4.699199,5.5875506,6.4759026,7.362441,8.2507925,7.663393,7.07418,6.48678,5.89938,5.3119802,4.936697,4.5632267,4.1879435,3.8126602,3.437377,2.7883365,2.137483,1.4866294,0.8375887,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.9246109,1.8492218,2.7756457,3.7002566,4.6248674,6.588306,8.549932,10.51337,12.474996,14.436621,15.899682,17.362743,18.825804,20.287052,21.750113,19.012539,16.274965,13.537392,10.799818,8.062244,6.987158,5.9120708,4.836984,3.7618973,2.6868105,2.1501737,1.6117238,1.0750868,0.53663695,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.18673515,0.25018883,0.31182957,0.37528324,0.43692398,0.34990177,0.26287958,0.17585737,0.0870222,0.0,0.0,0.0,0.0,0.0,0.0,0.31182957,0.62547207,0.93730164,1.2491312,1.5627737,1.2491312,0.93730164,0.62547207,0.31182957,0.0,0.07433146,0.15047589,0.22480737,0.2991388,0.37528324,0.2991388,0.22480737,0.15047589,0.07433146,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.13778515,0.2755703,0.41335547,0.5493277,0.6871128,0.5493277,0.41335547,0.2755703,0.13778515,0.0,0.06164073,0.12509441,0.18673515,0.25018883,0.31182957,0.2991388,0.28826106,0.2755703,0.26287958,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,4.612177,9.162713,13.713249,18.261972,22.812508,21.561563,20.312433,19.063301,17.812357,16.563227,18.662638,20.762047,22.863272,24.962683,27.062092,26.574406,26.08672,25.600845,25.113157,24.625471,22.912222,21.200785,19.487535,17.774284,16.062849,15.199879,14.336908,13.475751,12.612781,11.74981,9.91328,8.074935,6.2365913,4.40006,2.561716,2.561716,2.561716,2.561716,2.561716,2.561716,2.4003625,2.2371957,2.0758421,1.9126755,1.7495089,1.7368182,1.7241274,1.7132497,1.7005589,1.6878681,1.5120108,1.3379664,1.162109,0.9880646,0.8122072,0.8629702,0.9119202,0.96268314,1.0116332,1.062396,0.9880646,0.9119202,0.8375887,0.76325727,0.6871128,0.5493277,0.41335547,0.2755703,0.13778515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.9880646,1.9743162,2.962381,3.9504454,4.936697,4.949388,4.9620786,4.974769,4.98746,5.0001507,5.475147,5.9501433,6.4251394,6.9001355,7.3751316,8.713099,10.049252,11.3872175,12.725184,14.06315,13.899984,13.736817,13.575464,13.412297,13.24913,13.637105,14.025079,14.413053,14.799213,15.187187,13.24913,11.312886,9.374829,7.4367723,5.5005283,6.5248523,7.550989,8.575313,9.599637,10.625773,11.111648,11.599335,12.087022,12.574709,13.062395,12.250188,11.437981,10.625773,9.811753,8.999546,10.549629,12.099712,13.649796,15.199879,16.749962,14.975071,13.200181,11.42529,9.6504,7.8755093,6.5629244,5.2503395,3.9377546,2.6251698,1.3125849,1.9634385,2.612479,3.2633326,3.9123733,4.5632267,5.0998635,5.638314,6.1749506,6.7115874,7.250037,8.774739,10.29944,11.8241415,13.3506565,14.875358,10.049252,10.074633,10.100015,10.125396,10.150778,10.174346,8.375887,6.5756154,4.7753434,2.9750717,1.1747998,2.231757,3.290527,4.347484,5.4044414,6.4632115,8.033237,9.603263,11.173288,12.743314,14.313339,13.682428,13.05333,12.42242,11.793322,11.162411,10.326634,9.492672,8.656897,7.8229337,6.987158,7.12313,7.2572894,7.3932614,7.5274205,7.66158,6.48678,5.3119802,4.137181,2.962381,1.7875811,1.4703126,1.1530442,0.83577573,0.5166943,0.19942589,0.69073874,1.1802386,1.6697385,2.1592383,2.6505513,3.8471067,5.045475,6.24203,7.440398,8.636953,7.9081426,7.177519,6.446895,5.718084,4.98746,4.1897564,3.392053,2.5943494,1.7966459,1.0007553,1.209246,1.4195497,1.6298534,1.840157,2.0504606,2.2516994,2.4547513,2.657803,2.8608549,3.0620937,2.6795588,2.2970235,1.9144884,1.5319533,1.1494182,1.4648738,1.7803292,2.0957847,2.4094272,2.7248828,2.6016014,2.4801328,2.3568513,2.2353828,2.1121013,2.1519866,2.1918716,2.231757,2.2716422,2.3133402,1.9308052,1.54827,1.1657349,0.78319985,0.40066472,0.3208944,0.23931105,0.15954071,0.07977036,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.099712946,0.19942589,0.2991388,0.40066472,0.50037766,0.67986095,0.85934424,1.0406405,1.2201238,1.3996071,1.6896812,1.9797552,2.269829,2.5599031,2.8499773,3.2016919,3.5552197,3.9069343,4.2604623,4.612177,5.906632,7.2029004,8.497355,9.791811,11.088079,10.060129,9.03218,8.00423,6.978093,5.9501433,7.8102427,9.670342,11.530442,13.390542,15.250641,13.377851,11.50506,9.63227,7.75948,5.8866897,5.0799212,4.273153,3.4645715,2.657803,1.8492218,5.18326,8.515485,11.847711,15.179935,18.512161,16.893185,15.272397,13.651608,12.032633,10.411844,9.864329,9.316814,8.7693,8.221786,7.6742706,6.7532854,5.8304877,4.9076896,3.9848917,3.0620937,4.274966,5.487838,6.70071,7.911769,9.12464,7.3497505,5.57486,3.7999697,2.0250793,0.25018883,0.26287958,0.2755703,0.28826106,0.2991388,0.31182957,2.3641033,4.41819,6.4704633,8.5227375,10.57501,8.714911,6.8548117,4.994712,3.1346123,1.2745126,1.6896812,2.1048496,2.520018,2.9351864,3.350355,2.8282216,2.3042755,1.7821422,1.260009,0.73787576,4.7118897,8.6877165,12.661731,16.637558,20.611572,16.699198,12.786825,8.874452,4.9620786,1.0497054,1.4775645,1.9054236,2.333283,2.759329,3.1871881,2.5798457,1.9725033,1.3651608,0.75781834,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.058014803,0.11421664,0.17223145,0.23024625,0.28826106,0.5982776,0.90829426,1.2183108,1.5283275,1.8383441,1.789394,1.742257,1.69512,1.647983,1.6008459,1.6171626,1.6352923,1.6534219,1.6697385,1.6878681,2.268016,2.8481643,3.4283123,4.006647,4.5867953,5.199577,5.812358,6.4251394,7.037921,7.650702,7.130382,6.6100616,6.089741,5.569421,5.049101,4.7554007,4.459888,4.164375,3.870675,3.5751622,3.4301252,3.2850883,3.1400511,2.9950142,2.8499773,3.247016,3.6458678,4.0429068,4.439945,4.836984,5.772473,6.7079616,7.6434503,8.577126,9.512614,10.781689,12.052575,13.3234625,14.592536,15.863422,16.21695,16.57229,16.927631,17.282972,17.6365,15.399304,13.162108,10.924912,8.6877165,6.450521,5.5893636,4.7300196,3.870675,3.009518,2.1501737,1.7549478,1.3597219,0.9644961,0.56927025,0.17585737,0.13959812,0.10515183,0.07070554,0.034446288,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.15047589,0.19942589,0.25018883,0.2991388,0.34990177,0.35171473,0.35534066,0.35715362,0.36077955,0.36259252,0.29007402,0.21755551,0.14503701,0.072518505,0.0,0.25018883,0.50037766,0.7505665,1.0007553,1.2491312,1.0025684,0.7541924,0.5076295,0.25925365,0.012690738,0.0870222,0.16316663,0.2374981,0.31182957,0.387974,0.3100166,0.23205921,0.15410182,0.07795739,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07977036,0.15954071,0.23931105,0.3208944,0.40066472,0.42060733,0.4405499,0.4604925,0.48043507,0.50037766,0.42423326,0.34990177,0.2755703,0.19942589,0.12509441,0.21936847,0.3154555,0.40972954,0.5058166,0.6000906,0.48587397,0.36984438,0.25562772,0.13959812,0.025381476,0.07795739,0.13053331,0.18310922,0.23568514,0.28826106,0.27013144,0.2520018,0.23568514,0.21755551,0.19942589,0.43329805,0.6653573,0.8974165,1.1294757,1.3633479,1.0895905,0.81764615,0.54570174,0.27194437,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,3.9395678,7.7304726,11.519565,15.310469,19.099562,18.011784,16.92582,15.838041,14.750263,13.662486,15.417434,17.172382,18.92733,20.682278,22.437225,21.967669,21.49811,21.02674,20.557182,20.087626,19.097748,18.10787,17.117992,16.128115,15.138238,14.730321,14.322405,13.914488,13.508384,13.100468,11.624716,10.150778,8.675026,7.1992745,5.7253356,5.5367875,5.3500524,5.163317,4.974769,4.788034,4.421816,4.0574102,3.6930048,3.3267863,2.962381,2.9424384,2.9224956,2.902553,2.8826106,2.8626678,2.6233568,2.382233,2.1429217,1.9017978,1.6624867,1.5591478,1.4576219,1.3542831,1.2527572,1.1494182,1.0424535,0.9354887,0.82671094,0.7197462,0.61278135,0.51306844,0.41335547,0.31182957,0.21211663,0.11240368,0.09064813,0.06707962,0.045324065,0.02175555,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.032633327,0.027194439,0.02175555,0.018129626,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.7904517,1.5790904,2.3695421,3.159994,3.9504454,3.9867048,4.024777,4.062849,4.099108,4.137181,4.5251546,4.9131284,5.2992897,5.6872635,6.0752378,7.124943,8.174648,9.224354,10.274059,11.325577,11.334642,11.34552,11.354585,11.365462,11.374527,11.969179,12.565643,13.1602955,13.754947,14.349599,12.76507,11.18054,9.594198,8.009668,6.4251394,6.929143,7.4349594,7.9407763,8.444779,8.950596,9.407463,9.864329,10.323009,10.779876,11.236742,10.529687,9.822631,9.115576,8.406708,7.699652,8.917963,10.13446,11.352772,12.569269,13.7875805,12.712494,11.637406,10.56232,9.487233,8.412147,7.132195,5.8522434,4.572292,3.29234,2.0123885,2.5127661,3.0131438,3.5117085,4.0120864,4.512464,4.9620786,5.411693,5.863121,6.3127356,6.7623506,8.013294,9.262425,10.51337,11.762501,13.011633,9.474543,9.612328,9.750113,9.8878975,10.025683,10.161655,8.424837,6.688019,4.949388,3.2125697,1.4757515,2.277081,3.0802233,3.8833659,4.6846952,5.487838,6.740595,7.993352,9.244296,10.497053,11.74981,11.503247,11.254871,11.008308,10.7599325,10.51337,9.567003,8.62245,7.6778965,6.733343,5.7869763,5.9447045,6.1024323,6.26016,6.4178877,6.5756154,5.750717,4.9258194,4.099108,3.2742105,2.4493124,1.9906329,1.5301404,1.0696479,0.6091554,0.15047589,0.58014804,1.0098201,1.4394923,1.8691645,2.3006494,3.4573197,4.615803,5.772473,6.929143,8.087626,7.690587,7.2917356,6.8946967,6.497658,6.1006193,5.2557783,4.410938,3.5642843,2.7194438,1.8746033,1.9326181,1.9906329,2.0468347,2.1048496,2.1628644,2.280707,2.3967366,2.514579,2.6324217,2.7502642,2.5599031,2.3695421,2.179181,1.9906329,1.8002719,2.0178273,2.2353828,2.4529383,2.6704938,2.8880494,2.70494,2.521831,2.3405347,2.1574254,1.9743162,2.0178273,2.0595255,2.1030366,2.1447346,2.1882458,1.8347181,1.4830034,1.1294757,0.7777609,0.42423326,0.34083697,0.25562772,0.17041849,0.08520924,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07433146,0.15047589,0.22480737,0.2991388,0.37528324,0.5728962,0.7705091,0.968122,1.1657349,1.3633479,1.6298534,1.8981718,2.1646774,2.4329958,2.6995013,3.24339,3.785466,4.327542,4.8696175,5.411693,6.414262,7.41683,8.419398,9.421967,10.424535,9.606889,8.789243,7.9715962,7.155763,6.338117,8.158332,9.976733,11.7969475,13.617162,15.437376,13.591781,11.747997,9.902402,8.056806,6.2130227,5.5966153,4.9820213,4.367427,3.7528327,3.1382382,5.4515786,7.7667317,10.081885,12.397038,14.712192,14.159238,13.608097,13.055143,12.50219,11.949236,10.741803,9.53437,8.326937,7.119504,5.9120708,5.5549173,5.197764,4.84061,4.4816437,4.12449,4.8750563,5.6256227,6.3743763,7.124943,7.8755093,6.338117,4.800725,3.2633326,1.7241274,0.18673515,0.2374981,0.28826106,0.33721104,0.387974,0.43692398,2.70494,4.972956,7.2409725,9.507175,11.775192,9.679407,7.5854354,5.4896507,3.395679,1.2998942,1.8292793,2.3604772,2.8898623,3.4192474,3.9504454,3.4301252,2.909805,2.3894846,1.8691645,1.3506571,4.574105,7.799365,11.024626,14.249886,17.475147,14.362289,11.249433,8.136576,5.0255322,1.9126755,2.7919624,3.673062,4.552349,5.431636,6.3127356,5.1107416,3.9069343,2.70494,1.502946,0.2991388,0.23931105,0.1794833,0.11965553,0.059827764,0.0,0.065266654,0.13053331,0.19579996,0.25925365,0.3245203,0.5946517,0.86478317,1.1349145,1.405046,1.6751775,1.9054236,2.13567,2.3659163,2.5943494,2.8245957,2.8481643,2.8699198,2.8916752,2.9152439,2.9369993,3.4228733,3.9069343,4.3928084,4.876869,5.3627434,5.6999545,6.037165,6.3743763,6.7134004,7.0506115,6.5973706,6.14413,5.6927023,5.239462,4.788034,4.572292,4.358362,4.1426196,3.926877,3.7129474,4.071914,4.4326935,4.7916603,5.1524396,5.5132194,6.345369,7.177519,8.009668,8.841819,9.675781,10.620335,11.564888,12.509441,13.455809,14.400362,14.976884,15.555219,16.13174,16.710075,17.288412,16.534218,15.781839,15.02946,14.277081,13.524701,11.787883,10.049252,8.312433,6.5756154,4.836984,4.1915693,3.5479677,2.902553,2.2571385,1.6117238,1.3597219,1.1077201,0.8557183,0.60190356,0.34990177,0.27919623,0.21030366,0.13959812,0.07070554,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.11240368,0.15047589,0.18673515,0.22480737,0.26287958,0.35534066,0.44780177,0.5402629,0.6327239,0.72518504,0.58014804,0.43511102,0.29007402,0.14503701,0.0,0.18673515,0.37528324,0.5620184,0.7505665,0.93730164,0.7541924,0.5728962,0.38978696,0.20667773,0.025381476,0.099712946,0.17585737,0.25018883,0.3245203,0.40066472,0.3208944,0.23931105,0.15954071,0.07977036,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.09064813,0.06707962,0.045324065,0.02175555,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.15954071,0.3208944,0.48043507,0.6399758,0.7995165,0.8031424,0.80495536,0.80676836,0.8103943,0.8122072,0.69980353,0.5873999,0.4749962,0.36259252,0.25018883,0.30276474,0.35534066,0.40791658,0.4604925,0.51306844,0.42060733,0.32814622,0.23568514,0.14322405,0.05076295,0.092461094,0.13415924,0.17767033,0.21936847,0.26287958,0.23931105,0.21755551,0.19579996,0.17223145,0.15047589,0.6653573,1.1802386,1.69512,2.2100015,2.7248828,2.179181,1.6352923,1.0895905,0.54570174,0.0,0.047137026,0.09427405,0.14322405,0.19036107,0.2374981,3.2669585,6.298232,9.327692,12.357153,15.386614,14.462003,13.537392,12.612781,11.6881695,10.761745,12.172231,13.582716,14.9932,16.401873,17.812357,17.359118,16.907688,16.454449,16.003021,15.54978,15.283275,15.014956,14.746637,14.480132,14.211814,14.260764,14.3079,14.355038,14.402175,14.449312,13.337966,12.224807,11.111648,10.000301,8.887142,8.511859,8.138389,7.763106,7.3878226,7.0125394,6.445082,5.8776245,5.3101673,4.74271,4.175253,4.1480584,4.120864,4.0918565,4.064662,4.0374675,3.73289,3.4283123,3.1219215,2.817344,2.5127661,2.2571385,2.0033236,1.7476959,1.4920682,1.2382535,1.0968424,0.9572442,0.81764615,0.678048,0.53663695,0.4749962,0.41335547,0.34990177,0.28826106,0.22480737,0.1794833,0.13415924,0.09064813,0.045324065,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.065266654,0.054388877,0.045324065,0.034446288,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.59283876,1.1856775,1.7767034,2.3695421,2.962381,3.0258346,3.0874753,3.149116,3.2125697,3.2742105,3.5751622,3.874301,4.175253,4.4743915,4.7753434,5.5367875,6.300045,7.063302,7.8247466,8.588004,8.7693,8.952409,9.135518,9.316814,9.499924,10.303066,11.104396,11.907538,12.710681,13.512011,12.279196,11.048194,9.815379,8.582565,7.3497505,7.3352466,7.320743,7.304426,7.2899227,7.2754188,7.703278,8.129324,8.557183,8.985043,9.412902,8.809185,8.207282,7.605378,7.0016613,6.399758,7.2844834,8.1692095,9.055748,9.940474,10.825199,10.449916,10.074633,9.699349,9.325879,8.950596,7.703278,6.454147,5.2068286,3.9595103,2.712192,3.0620937,3.4119956,3.7618973,4.1117992,4.461701,4.8242936,5.186886,5.5494785,5.9120708,6.2746634,7.250037,8.225411,9.200785,10.174346,11.14972,8.899834,9.1500225,9.400211,9.6504,9.900589,10.150778,8.4756,6.8004227,5.125245,3.4500678,1.7748904,2.322405,2.8699198,3.4174345,3.9649491,4.512464,5.4479527,6.3816285,7.317117,8.252605,9.188094,9.322253,9.458226,9.592385,9.728357,9.862516,8.807372,7.752228,6.697084,5.6419396,4.5867953,4.7680917,4.947575,5.127058,5.3083544,5.487838,5.0128417,4.537845,4.062849,3.587853,3.1128569,2.5091403,1.9072367,1.305333,0.7016165,0.099712946,0.46955732,0.83940166,1.209246,1.5809034,1.9507477,3.0675328,4.1843176,5.3029156,6.4197006,7.5382986,7.473032,7.407765,7.3424983,7.2772317,7.211965,6.319988,5.42801,4.5342193,3.6422417,2.7502642,2.6541772,2.5599031,2.465629,2.3695421,2.275268,2.3079014,2.3405347,2.373168,2.4058013,2.4366217,2.4402475,2.4420607,2.4456866,2.4474995,2.4493124,2.570781,2.6904364,2.810092,2.9297476,3.049403,2.808279,2.565342,2.322405,2.079468,1.8383441,1.8818551,1.9271792,1.9725033,2.0178273,2.0631514,1.7404441,1.4177368,1.0950294,0.77232206,0.44961473,0.36077955,0.27013144,0.1794833,0.09064813,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,0.46411842,0.67986095,0.89560354,1.1095331,1.3252757,1.5700256,1.8147756,2.0595255,2.3042755,2.5508385,3.2832751,4.0157123,4.748149,5.480586,6.2130227,6.921891,7.6325727,8.343254,9.052122,9.762803,9.155461,8.548119,7.9407763,7.3316207,6.7242785,8.504607,10.284937,12.065266,13.845595,15.624111,13.807523,11.990934,10.172533,8.354132,6.5375433,6.115123,5.6927023,5.2702823,4.847862,4.4254417,5.7217097,7.019791,8.317872,9.6141405,10.912222,11.427103,11.941984,12.456866,12.971747,13.486629,11.619277,9.751925,7.8845744,6.017223,4.1498713,4.358362,4.5650396,4.7717175,4.9802084,5.186886,5.475147,5.7615952,6.049856,6.338117,6.624565,5.3246713,4.024777,2.7248828,1.4249886,0.12509441,0.21211663,0.2991388,0.387974,0.4749962,0.5620184,3.045777,5.527723,8.009668,10.493427,12.975373,10.645717,8.314246,5.9845896,3.6549325,1.3252757,1.9706904,2.6142921,3.2597067,3.9051213,4.550536,4.0320287,3.5153344,2.9968271,2.4801328,1.9616255,4.4381323,6.9128265,9.38752,11.862214,14.336908,12.025381,9.712041,7.400513,5.087173,2.7756457,4.1081734,5.4407005,6.773228,8.105756,9.438283,7.6398244,5.8431783,4.0447197,2.2480736,0.44961473,0.36077955,0.27013144,0.1794833,0.09064813,0.0,0.072518505,0.14503701,0.21755551,0.29007402,0.36259252,0.59283876,0.823085,1.0533313,1.2817645,1.5120108,2.0196402,2.5272698,3.0348995,3.5425289,4.0501585,4.077353,4.1045475,4.1317415,4.160749,4.1879435,4.5777307,4.9675174,5.3573046,5.7470913,6.1368785,6.200332,6.261973,6.3254266,6.3870673,6.450521,6.0643597,5.6800117,5.295664,4.9095025,4.5251546,4.3891826,4.255023,4.120864,3.9848917,3.8507326,4.7155156,5.580299,6.445082,7.309865,8.174648,9.441909,10.70917,11.978244,13.245504,14.512766,15.468197,16.421816,17.377247,18.332678,19.288109,19.17208,19.057863,18.941833,18.827616,18.711586,16.8533,14.9932,13.1331005,11.273002,9.412902,8.174648,6.9382076,5.6999545,4.461701,3.2252605,2.7955883,2.3659163,1.9344311,1.504759,1.0750868,0.9644961,0.8557183,0.7451276,0.6345369,0.52575916,0.42060733,0.3154555,0.21030366,0.10515183,0.0,0.0,0.0,0.0,0.0,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.09064813,0.06707962,0.045324065,0.02175555,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.07433146,0.099712946,0.12509441,0.15047589,0.17585737,0.35715362,0.5402629,0.72337204,0.90466833,1.0877775,0.87022203,0.6526665,0.43511102,0.21755551,0.0,0.12509441,0.25018883,0.37528324,0.50037766,0.62547207,0.5076295,0.38978696,0.27194437,0.15410182,0.038072214,0.11240368,0.18673515,0.26287958,0.33721104,0.41335547,0.32995918,0.24837588,0.16497959,0.08339628,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.23931105,0.48043507,0.7197462,0.96087015,1.2001812,1.1856775,1.1693609,1.1548572,1.1403534,1.1258497,0.97537386,0.824898,0.6744221,0.52575916,0.37528324,0.38434806,0.39522585,0.40429065,0.41516843,0.42423326,0.35534066,0.28463513,0.21574254,0.14503701,0.07433146,0.10696479,0.13959812,0.17223145,0.20486477,0.2374981,0.21030366,0.18310922,0.15410182,0.12690738,0.099712946,0.8974165,1.69512,2.4928236,3.290527,4.0882306,3.2705846,2.4529383,1.6352923,0.81764615,0.0,0.065266654,0.13053331,0.19579996,0.25925365,0.3245203,2.5943494,4.8641787,7.135821,9.40565,11.675479,10.912222,10.150778,9.38752,8.624263,7.8628187,8.927028,9.99305,11.057259,12.123281,13.1874895,12.752378,12.317267,11.882156,11.447045,11.011934,11.466989,11.922042,12.377095,12.8321495,13.287203,13.789393,14.291584,14.795588,15.297778,15.799969,15.049402,14.300649,13.550082,12.799516,12.050762,11.486931,10.924912,10.362894,9.800876,9.237044,8.466536,7.6978393,6.92733,6.156821,5.388125,5.351866,5.317419,5.282973,5.2467136,5.2122674,4.842423,4.4725785,4.102734,3.73289,3.3630457,2.955129,2.5472124,2.1392958,1.7331922,1.3252757,1.1530442,0.9808127,0.80676836,0.6345369,0.46230546,0.43692398,0.41335547,0.387974,0.36259252,0.33721104,0.27013144,0.2030518,0.13415924,0.06707962,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.09789998,0.08339628,0.06707962,0.052575916,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.39522585,0.7904517,1.1856775,1.5790904,1.9743162,2.0631514,2.1501737,2.2371957,2.324218,2.4130533,2.6251698,2.8372865,3.049403,3.2633326,3.4754493,3.9504454,4.4254417,4.900438,5.375434,5.8504305,6.205771,6.5592985,6.9146395,7.26998,7.6253204,8.63514,9.644961,10.654781,11.664601,12.674421,11.795135,10.914035,10.034748,9.155461,8.274362,7.7395372,7.2047133,6.6698895,6.1350656,5.600241,5.99728,6.394319,6.793171,7.1902094,7.5872483,7.0904965,6.591932,6.09518,5.5984282,5.0998635,5.6528172,6.205771,6.7569118,7.309865,7.8628187,8.187339,8.511859,8.838193,9.162713,9.487233,8.272549,7.057863,5.8431783,4.6266804,3.4119956,3.6132345,3.8126602,4.0120864,4.213325,4.4127507,4.688321,4.9620786,5.237649,5.5132194,5.7869763,6.48678,7.1883965,7.8882003,8.588004,9.287807,8.325124,8.6877165,9.050309,9.412902,9.775495,10.138086,8.52455,6.9128265,5.2992897,3.6875658,2.0758421,2.3677292,2.659616,2.953316,3.245203,3.53709,4.15531,4.7717175,5.389938,6.008158,6.624565,7.1430726,7.6597667,8.178274,8.694968,9.211663,8.047741,6.882006,5.718084,4.552349,3.386614,3.589666,3.7927177,3.9957695,4.1970086,4.40006,4.274966,4.1498713,4.024777,3.8996825,3.774588,3.0294604,2.2843328,1.5392052,0.79589057,0.05076295,0.36077955,0.67079616,0.9808127,1.2908293,1.6008459,2.6777458,3.7546456,4.8333583,5.910258,6.987158,7.2554765,7.5219817,7.7903004,8.056806,8.325124,7.3841968,6.445082,5.504154,4.5650396,3.6241121,3.3775494,3.1291735,2.8826106,2.6342347,2.3876717,2.335096,2.2825198,2.229944,2.1773682,2.124792,2.3205922,2.514579,2.7103791,2.904366,3.100166,3.1219215,3.1454902,3.1672456,3.1908143,3.2125697,2.909805,2.6070402,2.3042755,2.0033236,1.7005589,1.7476959,1.794833,1.84197,1.889107,1.938057,1.6443571,1.35247,1.0605831,0.7668832,0.4749962,0.38072214,0.28463513,0.19036107,0.09427405,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.35715362,0.58921283,0.823085,1.0551442,1.2872034,1.5101979,1.7331922,1.9543737,2.1773682,2.4003625,3.3231604,4.2441454,5.1669436,6.089741,7.0125394,7.4295206,7.8483152,8.265296,8.682278,9.099259,8.70222,8.3051815,7.9081426,7.509291,7.112252,8.852696,10.593141,12.331772,14.072216,15.812659,14.023266,12.232059,10.442664,8.653271,6.8620634,6.6318173,6.4033837,6.1731377,5.942891,5.712645,5.9918413,6.2728505,6.552047,6.833056,7.112252,8.694968,10.277685,11.860401,13.443117,15.025834,12.496751,9.969481,7.4422116,4.914942,2.3876717,3.159994,3.9323158,4.704638,5.47696,6.249282,6.0752378,5.89938,5.7253356,5.5494785,5.375434,4.313038,3.2506418,2.1882458,1.1258497,0.06164073,0.18673515,0.31182957,0.43692398,0.5620184,0.6871128,3.3848011,6.0824895,8.780178,11.477866,14.175554,11.610212,9.04487,6.4795284,3.9141862,1.3506571,2.1102884,2.8699198,3.6295512,4.3891826,5.1506267,4.6357455,4.120864,3.6041696,3.0892882,2.5744069,4.3003473,6.0244746,7.750415,9.474543,11.200482,9.686659,8.174648,6.6626377,5.1506267,3.636803,5.422571,7.208339,8.992294,10.778063,12.562017,10.17072,7.7776093,5.384499,2.9932013,0.6000906,0.48043507,0.36077955,0.23931105,0.11965553,0.0,0.07977036,0.15954071,0.23931105,0.3208944,0.40066472,0.58921283,0.7795739,0.969935,1.1602961,1.3506571,2.13567,2.9206827,3.7056956,4.4907084,5.275721,5.3083544,5.3391747,5.371808,5.4044414,5.4370747,5.732588,6.0281005,6.3218007,6.6173134,6.9128265,6.70071,6.48678,6.2746634,6.0625467,5.8504305,5.5331616,5.2158933,4.896812,4.5795436,4.262275,4.207886,4.1516843,4.0972953,4.0429068,3.9867048,5.3573046,6.7279043,8.096691,9.467291,10.837891,12.540262,14.242634,15.945006,17.647377,19.34975,20.314245,21.280556,22.24505,23.209547,24.175856,23.367275,22.560507,21.751925,20.945156,20.138388,17.170568,14.202749,11.234929,8.267109,5.2992897,4.5632267,3.825351,3.0874753,2.3495996,1.6117238,1.3977941,1.1820517,0.968122,0.7523795,0.53663695,0.56927025,0.60190356,0.6345369,0.6671702,0.69980353,0.56020546,0.42060733,0.27919623,0.13959812,0.0,0.0,0.0,0.0,0.0,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.038072214,0.05076295,0.06164073,0.07433146,0.0870222,0.36077955,0.6327239,0.90466833,1.1766127,1.4503701,1.1602961,0.87022203,0.58014804,0.29007402,0.0,0.06164073,0.12509441,0.18673515,0.25018883,0.31182957,0.25925365,0.20667773,0.15410182,0.10333887,0.05076295,0.12509441,0.19942589,0.2755703,0.34990177,0.42423326,0.34083697,0.25562772,0.17041849,0.08520924,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.3208944,0.6399758,0.96087015,1.2799516,1.6008459,1.5682126,1.5355793,1.502946,1.4703126,1.4376793,1.2491312,1.062396,0.87566096,0.6871128,0.50037766,0.46774435,0.43511102,0.40247768,0.36984438,0.33721104,0.29007402,0.24293698,0.19579996,0.14684997,0.099712946,0.12328146,0.14503701,0.16679256,0.19036107,0.21211663,0.1794833,0.14684997,0.11421664,0.08339628,0.05076295,1.1294757,2.2100015,3.290527,4.36924,5.4497657,4.360175,3.2705846,2.179181,1.0895905,0.0,0.08339628,0.16497959,0.24837588,0.32995918,0.41335547,1.9217403,3.4319382,4.942136,6.452334,7.9625316,7.362441,6.7623506,6.16226,5.562169,4.9620786,5.6818247,6.401571,7.12313,7.842876,8.562622,8.145641,7.7268467,7.309865,6.892884,6.474089,7.652515,8.829127,10.007553,11.184166,12.362592,13.319836,14.277081,15.234324,16.193382,17.150625,16.762651,16.374678,15.986704,15.600543,15.212569,14.462003,13.713249,12.962683,12.212116,11.463363,10.489801,9.518054,8.544493,7.572745,6.599184,6.5574856,6.5157876,6.472276,6.430578,6.3870673,5.9519563,5.516845,5.081734,4.646623,4.213325,3.6531196,3.092914,2.5327086,1.9725033,1.4122978,1.2074331,1.0025684,0.79770356,0.59283876,0.387974,0.40066472,0.41335547,0.42423326,0.43692398,0.44961473,0.36077955,0.27013144,0.1794833,0.09064813,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.13053331,0.11059072,0.09064813,0.07070554,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.19761293,0.39522585,0.59283876,0.7904517,0.9880646,1.1004683,1.2128719,1.3252757,1.4376793,1.550083,1.6751775,1.8002719,1.9253663,2.0504606,2.175555,2.3622901,2.5508385,2.7375734,2.9243085,3.1128569,3.6404288,4.168001,4.695573,5.223145,5.750717,6.967215,8.185526,9.402024,10.620335,11.836833,11.30926,10.781689,10.254116,9.728357,9.200785,8.145641,7.0904965,6.035352,4.9802084,3.925064,4.2930956,4.6593137,5.027345,5.3953767,5.7615952,5.369995,4.976582,4.5849824,4.1933823,3.7999697,4.019338,4.2405195,4.459888,4.6792564,4.900438,5.924762,6.9508986,7.9752226,8.999546,10.025683,8.841819,7.6597667,6.4777155,5.295664,4.1117992,4.162562,4.213325,4.262275,4.313038,4.361988,4.550536,4.7372713,4.9258194,5.1125546,5.2992897,5.7253356,6.149569,6.5756154,6.9998484,7.424082,7.750415,8.225411,8.700407,9.175404,9.6504,10.125396,8.575313,7.02523,5.475147,3.925064,2.374981,2.4130533,2.4493124,2.4873846,2.525457,2.561716,2.8626678,3.1618068,3.4627585,3.7618973,4.062849,4.9620786,5.863121,6.7623506,7.663393,8.562622,7.28811,6.011784,4.7372713,3.4627585,2.1882458,2.4130533,2.6378605,2.8626678,3.0874753,3.3122826,3.53709,3.7618973,3.9867048,4.213325,4.4381323,3.5497808,2.663242,1.7748904,0.8883517,0.0,0.25018883,0.50037766,0.7505665,1.0007553,1.2491312,2.2879589,3.3249733,4.361988,5.4008155,6.43783,7.037921,7.6380115,8.238102,8.838193,9.438283,8.450218,7.462154,6.474089,5.487838,4.499773,4.099108,3.7002566,3.299592,2.9007401,2.5000753,2.3622901,2.2245052,2.08672,1.9507477,1.8129625,2.1991236,2.5870976,2.9750717,3.3630457,3.7492065,3.6748753,3.6005437,3.5243993,3.4500678,3.3757362,3.0131438,2.6505513,2.2879589,1.9253663,1.5627737,1.6117238,1.6624867,1.7132497,1.7621996,1.8129625,1.550083,1.2872034,1.0243238,0.76325727,0.50037766,0.40066472,0.2991388,0.19942589,0.099712946,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.25018883,0.50037766,0.7505665,1.0007553,1.2491312,1.4503701,1.649796,1.8492218,2.0504606,2.2498865,3.3630457,4.4743915,5.5875506,6.70071,7.8120556,7.93715,8.062244,8.187339,8.312433,8.437528,8.2507925,8.062244,7.8755093,7.686961,7.500226,9.200785,10.899531,12.60009,14.300649,15.999394,14.237195,12.474996,10.712796,8.950596,7.1883965,7.1503243,7.112252,7.07418,7.037921,6.9998484,6.261973,5.52591,4.788034,4.0501585,3.3122826,5.962834,8.611572,11.262123,13.912675,16.563227,13.374225,10.1870365,6.9998484,3.8126602,0.62547207,1.9616255,3.299592,4.6375585,5.975525,7.311678,6.6753283,6.037165,5.4008155,4.762653,4.12449,3.299592,2.474694,1.649796,0.824898,0.0,0.16316663,0.3245203,0.48768693,0.6508536,0.8122072,3.7256382,6.637256,9.550687,12.462305,15.375735,12.574709,9.775495,6.9744673,4.175253,1.3742256,2.2498865,3.1255474,3.9993954,4.8750563,5.750717,5.237649,4.7245803,4.213325,3.7002566,3.1871881,4.162562,5.137936,6.11331,7.0868707,8.062244,7.3497505,6.637256,5.924762,5.2122674,4.499773,6.736969,8.974165,11.213174,13.45037,15.687565,12.699803,9.712041,6.7242785,3.738329,0.7505665,0.6000906,0.44961473,0.2991388,0.15047589,0.0,0.0870222,0.17585737,0.26287958,0.34990177,0.43692398,0.5873999,0.73787576,0.8883517,1.0370146,1.1874905,2.2498865,3.3122826,4.3746786,5.4370747,6.4994707,6.5375433,6.5756154,6.6118746,6.6499467,6.688019,6.887445,7.0868707,7.28811,7.4875355,7.686961,7.1992745,6.7134004,6.2257137,5.7380266,5.2503395,5.0001507,4.749962,4.499773,4.249584,3.9993954,4.024777,4.0501585,4.07554,4.099108,4.12449,5.999093,7.8755093,9.750113,11.624716,13.499319,15.636803,17.774284,19.911768,22.049252,24.186733,25.162107,26.137482,27.112856,28.08823,29.06179,27.56247,26.06315,24.562017,23.062696,21.563377,17.487837,13.412297,9.336758,5.2630305,1.1874905,0.9499924,0.7124943,0.4749962,0.2374981,0.0,0.0,0.0,0.0,0.0,0.0,0.17585737,0.34990177,0.52575916,0.69980353,0.87566096,0.69980353,0.52575916,0.34990177,0.17585737,0.0,0.0,0.0,0.0,0.0,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.36259252,0.72518504,1.0877775,1.4503701,1.8129625,1.4503701,1.0877775,0.72518504,0.36259252,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.13778515,0.21211663,0.28826106,0.36259252,0.43692398,0.34990177,0.26287958,0.17585737,0.0870222,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.40066472,0.7995165,1.2001812,1.6008459,1.9996977,1.9507477,1.8999848,1.8492218,1.8002719,1.7495089,1.5247015,1.2998942,1.0750868,0.85027945,0.62547207,0.5493277,0.4749962,0.40066472,0.3245203,0.25018883,0.22480737,0.19942589,0.17585737,0.15047589,0.12509441,0.13778515,0.15047589,0.16316663,0.17585737,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,1.3633479,2.7248828,4.0882306,5.4497657,6.813113,5.4497657,4.0882306,2.7248828,1.3633479,0.0,0.099712946,0.19942589,0.2991388,0.40066472,0.50037766,1.2509441,1.9996977,2.7502642,3.5008307,4.249584,3.8126602,3.3757362,2.9369993,2.5000753,2.0631514,2.4366217,2.811905,3.1871881,3.5624714,3.9377546,3.53709,3.1382382,2.7375734,2.3369088,1.938057,3.8380418,5.7380266,7.6380115,9.537996,11.437981,12.850279,14.262577,15.674874,17.087172,18.49947,18.475903,18.45052,18.425138,18.399757,18.374376,17.437075,16.499773,15.56247,14.625169,13.687867,12.513068,11.338268,10.161655,8.9868555,7.8120556,7.763106,7.7123427,7.663393,7.61263,7.5618668,7.063302,6.5629244,6.0625467,5.562169,5.0617914,4.349297,3.636803,2.9243085,2.2118144,1.49932,1.261822,1.0243238,0.7868258,0.5493277,0.31182957,0.36259252,0.41335547,0.46230546,0.51306844,0.5620184,0.44961473,0.33721104,0.22480737,0.11240368,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.16316663,0.13778515,0.11240368,0.0870222,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13778515,0.2755703,0.41335547,0.5493277,0.6871128,0.72518504,0.76325727,0.7995165,0.8375887,0.87566096,0.774135,0.6744221,0.5747091,0.4749962,0.37528324,1.0750868,1.7748904,2.474694,3.1744974,3.874301,5.2992897,6.7242785,8.149267,9.574255,10.999244,10.825199,10.649343,10.475298,10.29944,10.125396,8.549932,6.9744673,5.4008155,3.825351,2.2498865,2.5870976,2.9243085,3.2633326,3.6005437,3.9377546,3.6494937,3.3630457,3.0747845,2.7883365,2.5000753,2.3876717,2.275268,2.1628644,2.0504606,1.938057,3.6621845,5.388125,7.112252,8.838193,10.56232,9.412902,8.26167,7.112252,5.962834,4.8116026,4.7118897,4.612177,4.512464,4.4127507,4.313038,4.4127507,4.512464,4.612177,4.7118897,4.8116026,4.9620786,5.1125546,5.2630305,5.411693,5.562169,7.9244595,8.207282,8.490104,8.772926,9.055748,9.336758,8.067683,6.796797,5.527723,4.256836,2.9877625,3.3666716,3.7473936,4.1281157,4.507025,4.8877473,5.132497,5.377247,5.621997,5.866747,6.11331,6.985345,7.85738,8.729415,9.603263,10.475298,9.284182,8.094878,6.9055743,5.714458,4.5251546,4.4925213,4.459888,4.4272547,4.3946214,4.361988,4.465327,4.5668526,4.670192,4.7717175,4.8750563,4.064662,3.254268,2.4456866,1.6352923,0.824898,0.85934424,0.89560354,0.9300498,0.9644961,1.0007553,1.9507477,2.9007401,3.8507326,4.800725,5.750717,6.352621,6.9545245,7.558241,8.160145,8.762048,7.902704,7.0433598,6.1822023,5.3228583,4.461701,4.1299286,3.7981565,3.4645715,3.1327994,2.7992141,2.6233568,2.4456866,2.268016,2.0903459,1.9126755,2.2154403,2.518205,2.819157,3.1219215,3.4246864,3.3666716,3.3104696,3.2524548,3.1944401,3.1382382,2.817344,2.4982624,2.1773682,1.8582866,1.5373923,1.5718386,1.6080978,1.6425442,1.6769904,1.7132497,1.5192627,1.3270886,1.1349145,0.94274056,0.7505665,0.6073425,0.46411842,0.32270733,0.1794833,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.26287958,0.52575916,0.7868258,1.0497054,1.3125849,1.4431182,1.5718386,1.7023718,1.8329052,1.9616255,2.902553,3.8416677,4.782595,5.7217097,6.6626377,7.0143523,7.36788,7.7195945,8.073122,8.424837,8.096691,7.7703576,7.4422116,7.115878,6.787732,8.285239,9.782746,11.280253,12.7777605,14.275268,12.754191,11.234929,9.715667,8.194591,6.6753283,6.740595,6.8058615,6.869315,6.9345818,6.9998484,6.167699,5.335549,4.501586,3.6694362,2.8372865,5.047288,7.2572894,9.467291,11.677292,13.887294,11.445232,9.003172,6.5592985,4.117238,1.6751775,2.6704938,3.6658103,4.6593137,5.65463,6.6499467,5.9918413,5.335549,4.6774435,4.019338,3.3630457,2.8826106,2.4021754,1.9217403,1.4431182,0.96268314,1.3307146,1.696933,2.0649643,2.4329958,2.7992141,4.699199,6.599184,8.499168,10.399154,12.299138,10.31757,8.334189,6.352621,4.36924,2.3876717,2.8300345,3.2723975,3.7147603,4.157123,4.599486,4.255023,3.9105604,3.5642843,3.2198215,2.8753586,3.6458678,4.4145637,5.185073,5.955582,6.7242785,6.987158,7.250037,7.512917,7.7757964,8.036863,10.3502035,12.661731,14.975071,17.288412,19.59994,17.176008,14.750263,12.32452,9.900589,7.474845,6.7859187,6.09518,5.4044414,4.7155156,4.024777,4.0555973,4.0846047,4.115425,4.1444325,4.175253,4.160749,4.1444325,4.1299286,4.115425,4.100921,4.934884,5.77066,6.604623,7.440398,8.274362,8.0858135,7.895452,7.705091,7.51473,7.324369,7.5346723,7.744976,7.95528,8.165584,8.375887,7.850128,7.324369,6.8004227,6.2746634,5.750717,5.582112,5.4153194,5.2467136,5.0799212,4.9131284,5.315606,5.718084,6.1205616,6.5230393,6.925517,8.285239,9.644961,11.004683,12.364405,13.724127,15.179935,16.635744,18.08974,19.54555,20.999546,21.481794,21.96404,22.448103,22.930351,23.4126,22.179785,20.94697,19.714155,18.483154,17.25034,13.990632,10.730926,7.4694057,4.209699,0.9499924,0.75963134,0.56927025,0.38072214,0.19036107,0.0,0.0,0.0,0.0,0.0,0.0,0.13959812,0.27919623,0.42060733,0.56020546,0.69980353,0.56020546,0.42060733,0.27919623,0.13959812,0.0,0.0,0.0,0.0,0.0,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.29007402,0.58014804,0.87022203,1.1602961,1.4503701,1.162109,0.87566096,0.5873999,0.2991388,0.012690738,0.047137026,0.08339628,0.11784257,0.15228885,0.18673515,0.16497959,0.14322405,0.11965553,0.09789998,0.07433146,0.3154555,0.55476654,0.79589057,1.0352017,1.2745126,1.0478923,0.8194591,0.59283876,0.36440548,0.13778515,0.11059072,0.08339628,0.054388877,0.027194439,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.48587397,0.969935,1.455809,1.93987,2.4257438,2.2607644,2.0957847,1.9308052,1.7658255,1.6008459,1.455809,1.310772,1.1657349,1.020698,0.87566096,0.75963134,0.64541465,0.5293851,0.41516843,0.2991388,0.26469254,0.23024625,0.19579996,0.15954071,0.12509441,0.13234627,0.13959812,0.14684997,0.15410182,0.16316663,0.19761293,0.23205921,0.26831847,0.30276474,0.33721104,1.5319533,2.7266958,3.923251,5.1179934,6.3127356,5.069043,3.827164,2.5852847,1.3415923,0.099712946,0.35534066,0.6091554,0.86478317,1.1204109,1.3742256,1.8981718,2.420305,2.9424384,3.4645715,3.9867048,3.5497808,3.1128569,2.6741197,2.2371957,1.8002719,2.0704033,2.3405347,2.610666,2.8807976,3.149116,2.8318477,2.514579,2.1973107,1.8800422,1.5627737,3.245203,4.9276323,6.6100616,8.292491,9.97492,11.050007,12.125093,13.200181,14.275268,15.350354,15.257894,15.165432,15.072971,14.98051,14.888049,14.231756,13.577277,12.922797,12.268318,11.612025,10.754494,9.896963,9.039432,8.1819,7.324369,7.3570023,7.3896356,7.422269,7.454902,7.4875355,7.0071006,6.526665,6.0480433,5.567608,5.087173,4.5269675,3.966762,3.4083695,2.8481643,2.2879589,1.9851941,1.6824293,1.3796645,1.0768998,0.774135,0.7541924,0.73424983,0.71430725,0.69436467,0.6744221,0.5475147,0.42060733,0.291887,0.16497959,0.038072214,0.059827764,0.08339628,0.10515183,0.12690738,0.15047589,0.13053331,0.11059072,0.09064813,0.07070554,0.05076295,0.054388877,0.059827764,0.065266654,0.07070554,0.07433146,0.092461094,0.11059072,0.12690738,0.14503701,0.16316663,0.13053331,0.09789998,0.065266654,0.032633327,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.12328146,0.23205921,0.34264994,0.45324063,0.5620184,0.61459434,0.6671702,0.7197462,0.77232206,0.824898,0.7469406,0.67079616,0.59283876,0.5148814,0.43692398,1.0025684,1.5682126,2.132044,2.6976883,3.2633326,4.505212,5.7470913,6.9907837,8.232663,9.474543,9.27693,9.079316,8.881703,8.684091,8.488291,7.2373466,5.9882154,4.7372713,3.48814,2.2371957,2.4620032,2.6868105,2.911618,3.1382382,3.3630457,3.1708715,2.9768846,2.7847104,2.5925364,2.4003625,2.333283,2.2643902,2.1973107,2.1302311,2.0631514,3.529838,4.9983377,6.4650245,7.931711,9.400211,8.415772,7.4295206,6.445082,5.4606433,4.4743915,4.4127507,4.349297,4.2876563,4.2242026,4.162562,4.195195,4.227829,4.2604623,4.2930956,4.325729,4.3982472,4.4707656,4.5432844,4.615803,4.688321,8.100317,8.189152,8.2798,8.370448,8.459284,8.549932,7.560054,6.5701766,5.580299,4.590421,3.6005437,4.322103,5.045475,5.767034,6.490406,7.211965,7.402326,7.592687,7.783048,7.9734097,8.161958,9.006798,9.851639,10.698292,11.543133,12.387974,11.282066,10.177972,9.072064,7.9679704,6.8620634,6.5719895,6.281915,5.9918413,5.7017674,5.411693,5.391751,5.371808,5.351866,5.331923,5.3119802,4.5795436,3.8471067,3.1146698,2.382233,1.649796,1.4703126,1.2908293,1.1095331,0.9300498,0.7505665,1.6117238,2.474694,3.3376641,4.2006345,5.0617914,5.667321,6.2728505,6.87838,7.4820967,8.087626,7.3551893,6.622752,5.8903155,5.1578784,4.4254417,4.160749,3.8942437,3.6295512,3.3648586,3.100166,2.8826106,2.665055,2.4474995,2.229944,2.0123885,2.229944,2.4474995,2.665055,2.8826106,3.100166,3.0602808,3.0203958,2.9805105,2.9406252,2.9007401,2.6233568,2.3441606,2.0667772,1.789394,1.5120108,1.5319533,1.551896,1.5718386,1.5917811,1.6117238,1.4902552,1.3669738,1.2455053,1.1222239,1.0007553,0.81583315,0.630911,0.44417584,0.25925365,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.2755703,0.5493277,0.824898,1.1004683,1.3742256,1.4358664,1.4956942,1.5555218,1.6153497,1.6751775,2.4420607,3.2107568,3.97764,4.744523,5.5132194,6.093367,6.6717024,7.25185,7.8319983,8.412147,7.944402,7.476658,7.0107265,6.542982,6.0752378,7.369693,8.664148,9.960417,11.254871,12.549327,11.273002,9.994863,8.716724,7.440398,6.16226,6.3308654,6.497658,6.6644506,6.833056,6.9998484,6.071612,5.145188,4.216951,3.290527,2.3622901,4.1317415,5.903006,7.6724577,9.441909,11.213174,9.514427,7.817495,6.1205616,4.421816,2.7248828,3.3775494,4.0302157,4.6828823,5.335549,5.9882154,5.3101673,4.632119,3.9540713,3.2778363,2.5997884,2.465629,2.3296568,2.1954978,2.0595255,1.9253663,2.4982624,3.0693457,3.6422417,4.215138,4.788034,5.674573,6.5629244,7.4494634,8.337815,9.224354,8.0604315,6.8946967,5.730775,4.5650396,3.3993049,3.4101827,3.4192474,3.4301252,3.43919,3.4500678,3.2723975,3.094727,2.9170568,2.7393866,2.561716,3.1273603,3.6930048,4.256836,4.8224807,5.388125,6.624565,7.8628187,9.099259,10.337513,11.575767,13.961625,16.349297,18.736969,21.12464,23.512312,21.650398,19.788486,17.92476,16.062849,14.200936,12.969934,11.740746,10.509744,9.280556,8.049554,8.02236,7.995165,7.9679704,7.9407763,7.911769,7.7322855,7.552802,7.3733187,7.192023,7.0125394,7.6198816,8.227224,8.834567,9.441909,10.049252,9.63227,9.215289,8.798307,8.379513,7.9625316,8.1819,8.403082,8.62245,8.841819,9.063,8.499168,7.93715,7.3751316,6.813113,6.249282,6.165886,6.0806766,5.995467,5.910258,5.825049,6.604623,7.3841968,8.165584,8.945157,9.724731,10.5695715,11.4144125,12.259253,13.1059065,13.9507475,14.723069,15.495391,16.267714,17.040035,17.812357,17.803293,17.792416,17.78335,17.772472,17.761595,16.797098,15.8326025,14.868106,13.901797,12.937301,10.491614,8.047741,5.6020546,3.1581807,0.7124943,0.56927025,0.42785916,0.28463513,0.14322405,0.0,0.0,0.0,0.0,0.0,0.0,0.10515183,0.21030366,0.3154555,0.42060733,0.52575916,0.42060733,0.3154555,0.21030366,0.10515183,0.0,0.0,0.0,0.0,0.0,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.09064813,0.06707962,0.045324065,0.02175555,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.21755551,0.43511102,0.6526665,0.87022203,1.0877775,0.87566096,0.66173136,0.44961473,0.2374981,0.025381476,0.09427405,0.16497959,0.23568514,0.3045777,0.37528324,0.31726846,0.25925365,0.2030518,0.14503701,0.0870222,0.49312583,0.8974165,1.3017071,1.7078108,2.1121013,1.745883,1.3778516,1.0098201,0.6417888,0.2755703,0.21936847,0.16497959,0.11059072,0.054388877,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.56927025,1.1403534,1.7096237,2.280707,2.8499773,2.570781,2.2897718,2.0105755,1.7295663,1.4503701,1.3851035,1.3198367,1.2545701,1.1893034,1.1258497,0.969935,0.81583315,0.65991837,0.5058166,0.34990177,0.3045777,0.25925365,0.21574254,0.17041849,0.12509441,0.12690738,0.13053331,0.13234627,0.13415924,0.13778515,0.24474995,0.35171473,0.4604925,0.56745726,0.6744221,1.7023718,2.7303216,3.7582715,4.784408,5.812358,4.690134,3.5679104,2.4456866,1.3216497,0.19942589,0.6091554,1.020698,1.4304274,1.840157,2.2498865,2.5453994,2.8390994,3.1346123,3.4301252,3.7256382,3.2869012,2.8499773,2.4130533,1.9743162,1.5373923,1.7023718,1.8673514,2.032331,2.1973107,2.3622901,2.126605,1.892733,1.6570477,1.4231756,1.1874905,2.6523643,4.117238,5.582112,7.0469856,8.511859,9.249735,9.987611,10.725487,11.463363,12.199425,12.039885,11.880343,11.720803,11.559449,11.399909,11.028252,10.654781,10.283124,9.909654,9.537996,8.997733,8.457471,7.9172077,7.3769445,6.836682,6.9527116,7.066928,7.1829576,7.2971745,7.413204,6.9527116,6.492219,6.0317264,5.573047,5.1125546,4.704638,4.2967215,3.8906176,3.482701,3.0747845,2.7067533,2.3405347,1.9725033,1.6044719,1.2382535,1.1476053,1.0569572,0.968122,0.8774739,0.7868258,0.64541465,0.50219065,0.36077955,0.21755551,0.07433146,0.08339628,0.09064813,0.09789998,0.10515183,0.11240368,0.09789998,0.08339628,0.06707962,0.052575916,0.038072214,0.059827764,0.08339628,0.10515183,0.12690738,0.15047589,0.18492219,0.21936847,0.25562772,0.29007402,0.3245203,0.25925365,0.19579996,0.13053331,0.065266654,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.10696479,0.19036107,0.27194437,0.35534066,0.43692398,0.5058166,0.5728962,0.6399758,0.7070554,0.774135,0.7197462,0.6653573,0.6091554,0.55476654,0.50037766,0.9300498,1.3597219,1.789394,2.2190661,2.6505513,3.7093215,4.7699046,5.8304877,6.889258,7.949841,7.7304726,7.509291,7.2899227,7.0705543,6.849373,5.924762,5.0001507,4.07554,3.150929,2.2245052,2.3369088,2.4493124,2.561716,2.6741197,2.7883365,2.6904364,2.5925364,2.4946365,2.3967366,2.3006494,2.277081,2.2553256,2.231757,2.2100015,2.1882458,3.397492,4.608551,5.8177967,7.027043,8.238102,7.41683,6.5973706,5.7779117,4.9584527,4.137181,4.1117992,4.0882306,4.062849,4.0374675,4.0120864,3.97764,3.9431937,3.9069343,3.872488,3.8380418,3.832603,3.827164,3.8217251,3.8180993,3.8126602,8.274362,8.172835,8.069496,7.9679704,7.8646317,7.763106,7.0524244,6.341743,5.632875,4.9221935,4.213325,5.277534,6.341743,7.407765,8.471974,9.537996,9.672155,9.808127,9.9422865,10.078259,10.212419,11.030065,11.847711,12.665357,13.483003,14.300649,13.279951,12.259253,11.240368,10.21967,9.200785,8.653271,8.105756,7.558241,7.0107265,6.4632115,6.319988,6.1767635,6.035352,5.8921285,5.750717,5.0944247,4.439945,3.785466,3.1291735,2.474694,2.079468,1.6842422,1.2908293,0.89560354,0.50037766,1.2745126,2.0504606,2.8245957,3.6005437,4.3746786,4.9820213,5.5893636,6.1967063,6.8058615,7.413204,6.8076744,6.202145,5.5966153,4.992899,4.3873696,4.1897564,3.9921436,3.7945306,3.5969179,3.3993049,3.141864,2.8844235,2.6269827,2.3695421,2.1121013,2.2444477,2.3767939,2.5091403,2.6432993,2.7756457,2.752077,2.7303216,2.7067533,2.6849976,2.663242,2.427557,2.1918716,1.9579996,1.7223145,1.4866294,1.4920682,1.4975071,1.502946,1.5083848,1.5120108,1.4594349,1.4068589,1.3542831,1.3017071,1.2491312,1.0225109,0.79589057,0.56745726,0.34083697,0.11240368,0.09064813,0.06707962,0.045324065,0.02175555,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.28826106,0.5747091,0.8629702,1.1494182,1.4376793,1.4268016,1.4177368,1.4068589,1.3977941,1.3869164,1.983381,2.5780327,3.1726844,3.7673361,4.361988,5.1705694,5.977338,6.7859187,7.592687,8.399456,7.7921133,7.1847706,6.5774283,5.9700856,5.3627434,6.454147,7.5473633,8.640579,9.731983,10.825199,9.789998,8.754796,7.7195945,6.684393,5.6491914,5.919323,6.189454,6.4595857,6.7297173,6.9998484,5.977338,4.954827,3.9323158,2.909805,1.887294,3.2180085,4.5469103,5.8776245,7.208339,8.537241,7.5854354,6.6318173,5.6800117,4.7282066,3.774588,4.0846047,4.3946214,4.704638,5.0146546,5.3246713,4.6266804,3.930503,3.2325122,2.5345216,1.8383441,2.0468347,2.2571385,2.467442,2.6777458,2.8880494,3.6658103,4.441758,5.219519,5.99728,6.775041,6.6499467,6.5248523,6.399758,6.2746634,6.149569,5.803293,5.4552045,5.1071157,4.76084,4.4127507,3.9903307,3.5679104,3.1454902,2.72307,2.3006494,2.2897718,2.280707,2.269829,2.2607644,2.2498865,2.610666,2.9696326,3.3304121,3.6893787,4.0501585,6.261973,8.4756,10.687414,12.899229,15.112856,17.57486,20.036863,22.500679,24.962683,27.424685,26.12479,24.824896,23.525002,22.22511,20.925215,19.155762,17.384499,15.6150465,13.845595,12.07433,11.989121,11.9057255,11.820516,11.735307,11.650098,11.3056345,10.959359,10.614896,10.270433,9.924157,10.304879,10.685601,11.06451,11.445232,11.8241415,11.18054,10.535126,9.88971,9.244296,8.600695,8.829127,9.059374,9.28962,9.519867,9.750113,9.1500225,8.549932,7.949841,7.3497505,6.7496595,6.7478466,6.7442207,6.742408,6.740595,6.736969,7.895452,9.052122,10.210606,11.367275,12.525759,12.855718,13.185677,13.515636,13.845595,14.175554,14.26439,14.355038,14.445685,14.534521,14.625169,14.122978,13.620788,13.116784,12.6145935,12.112403,11.4144125,10.718235,10.020245,9.322253,8.624263,6.9944096,5.3645563,3.7347028,2.1048496,0.4749962,0.38072214,0.28463513,0.19036107,0.09427405,0.0,0.0,0.0,0.0,0.0,0.0,0.07070554,0.13959812,0.21030366,0.27919623,0.34990177,0.27919623,0.21030366,0.13959812,0.07070554,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.14503701,0.29007402,0.43511102,0.58014804,0.72518504,0.5873999,0.44961473,0.31182957,0.17585737,0.038072214,0.14322405,0.24837588,0.35171473,0.45686656,0.5620184,0.46955732,0.3770962,0.28463513,0.19217403,0.099712946,0.67079616,1.2400664,1.8093367,2.38042,2.94969,2.4420607,1.9344311,1.4268016,0.91917205,0.41335547,0.32995918,0.24837588,0.16497959,0.08339628,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.6544795,1.310772,1.9652514,2.619731,3.2742105,2.8807976,2.4855716,2.0903459,1.69512,1.2998942,1.3143979,1.3307146,1.3452182,1.3597219,1.3742256,1.1802386,0.98443866,0.7904517,0.5946517,0.40066472,0.3444629,0.29007402,0.23568514,0.1794833,0.12509441,0.12328146,0.11965553,0.11784257,0.11421664,0.11240368,0.291887,0.47318324,0.6526665,0.8321498,1.0116332,1.8727903,2.7321346,3.5932918,4.4526362,5.3119802,4.309412,3.3068438,2.3042755,1.3017071,0.2991388,0.86478317,1.4304274,1.9942589,2.5599031,3.1255474,3.1926272,3.2597067,3.3267863,3.395679,3.4627585,3.0258346,2.5870976,2.1501737,1.7132497,1.2745126,1.3343405,1.3941683,1.455809,1.5156367,1.5754645,1.4231756,1.2708868,1.1167849,0.9644961,0.8122072,2.0595255,3.3068438,4.554162,5.803293,7.0506115,7.4494634,7.850128,8.2507925,8.649645,9.050309,8.821876,8.595256,8.366822,8.140202,7.911769,7.8229337,7.7322855,7.6416373,7.552802,7.462154,7.2391596,7.017978,6.794984,6.5719895,6.350808,6.548421,6.7442207,6.9418335,7.1394467,7.3370595,6.8983226,6.4577727,6.017223,5.576673,5.137936,4.882308,4.6266804,4.3728657,4.117238,3.8616104,3.4301252,2.9968271,2.565342,2.132044,1.7005589,1.5392052,1.3796645,1.2201238,1.0605831,0.89922947,0.7433147,0.5855869,0.42785916,0.27013144,0.11240368,0.10515183,0.09789998,0.09064813,0.08339628,0.07433146,0.065266654,0.054388877,0.045324065,0.034446288,0.025381476,0.065266654,0.10515183,0.14503701,0.18492219,0.22480737,0.27738327,0.32995918,0.3825351,0.43511102,0.48768693,0.38978696,0.291887,0.19579996,0.09789998,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.092461094,0.14684997,0.2030518,0.2574407,0.31182957,0.39522585,0.47680917,0.56020546,0.6417888,0.72518504,0.69255173,0.65991837,0.62728506,0.5946517,0.5620184,0.8575313,1.1530442,1.4467441,1.742257,2.03777,2.9152439,3.7927177,4.670192,5.5476656,6.4251394,6.1822023,5.9392653,5.6981416,5.4552045,5.2122674,4.612177,4.0120864,3.4119956,2.811905,2.2118144,2.2118144,2.2118144,2.2118144,2.2118144,2.2118144,2.2100015,2.2081885,2.2045624,2.2027495,2.1991236,2.222692,2.2444477,2.268016,2.2897718,2.3133402,3.2651455,4.216951,5.1705694,6.1223745,7.07418,6.4197006,5.765221,5.1107416,4.454449,3.7999697,3.8126602,3.825351,3.8380418,3.8507326,3.8616104,3.7600844,3.6567454,3.5552197,3.4518807,3.350355,3.2669585,3.1853752,3.101979,3.0203958,2.9369993,8.450218,8.154706,7.859193,7.5654926,7.26998,6.9744673,6.544795,6.115123,5.6854506,5.2557783,4.8242936,6.2329655,7.6398244,9.046683,10.455356,11.862214,11.941984,12.021755,12.103338,12.183108,12.262879,13.05333,13.8419695,14.632421,15.422873,16.213324,15.277836,14.342347,13.406858,12.473183,11.537694,10.7327385,9.927783,9.122828,8.317872,7.512917,7.2482243,6.981719,6.717026,6.452334,6.187641,5.6093063,5.032784,4.454449,3.877927,3.299592,2.6904364,2.079468,1.4703126,0.85934424,0.25018883,0.93730164,1.6244144,2.3133402,3.000453,3.6875658,4.2967215,4.9076896,5.516845,6.1278133,6.736969,6.26016,5.7833505,5.3047285,4.8279195,4.349297,4.220577,4.0900435,3.9595103,3.83079,3.7002566,3.4029307,3.105605,2.808279,2.5091403,2.2118144,2.2607644,2.3079014,2.3550384,2.4021754,2.4493124,2.4456866,2.4402475,2.4348087,2.42937,2.4257438,2.231757,2.039583,1.8474089,1.6552348,1.4630609,1.452183,1.4431182,1.4322405,1.4231756,1.4122978,1.4304274,1.4467441,1.4648738,1.4830034,1.49932,1.2291887,0.96087015,0.69073874,0.42060733,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.2991388,0.6000906,0.89922947,1.2001812,1.49932,1.4195497,1.3397794,1.260009,1.1802386,1.1004683,1.5228885,1.9453088,2.3677292,2.7901495,3.2125697,4.2477713,5.282973,6.3181744,7.3533764,8.386765,7.6398244,6.892884,6.14413,5.3971896,4.650249,5.540414,6.430578,7.320743,8.209095,9.099259,8.306994,7.51473,6.722465,5.9302006,5.137936,5.5095935,5.883064,6.2547207,6.628191,6.9998484,5.883064,4.764466,3.6476808,2.5290828,1.4122978,2.3024626,3.1926272,4.082792,4.972956,5.863121,5.65463,5.4479527,5.239462,5.032784,4.8242936,4.7916603,4.76084,4.7282066,4.695573,4.6629395,3.9450066,3.2270734,2.5091403,1.79302,1.0750868,1.6298534,2.18462,2.7393866,3.294153,3.8507326,4.8333583,5.814171,6.796797,7.7794223,8.762048,7.6253204,6.48678,5.3500524,4.213325,3.0747845,3.5443418,4.0157123,4.4852695,4.954827,5.424384,4.5704784,3.7147603,2.8608549,2.0051367,1.1494182,1.3071461,1.4648738,1.6226015,1.7803292,1.938057,2.0921588,2.2480736,2.4021754,2.5580902,2.712192,5.89938,9.086569,12.27557,15.462758,18.649946,21.188093,23.724428,26.262575,28.800724,31.337059,30.599182,29.86312,29.125244,28.387367,27.649492,25.339779,23.030064,20.72035,18.410635,16.100922,15.957697,15.814472,15.673061,15.529838,15.388427,14.877171,14.367728,13.858286,13.347031,12.837588,12.989877,13.142166,13.294455,13.446743,13.600845,12.726997,11.854962,10.982927,10.110892,9.237044,9.4781685,9.71748,9.956791,10.197914,10.437225,9.800876,9.162713,8.52455,7.8882003,7.250037,7.3298078,7.409578,7.4893484,7.569119,7.650702,9.184468,10.720048,12.255627,13.789393,15.324973,15.140051,14.955129,14.770206,14.585284,14.400362,13.807523,13.2146845,12.621845,12.03082,11.437981,10.442664,9.447348,8.452031,7.456715,6.4632115,6.0317264,5.6020546,5.1723824,4.74271,4.313038,3.4972048,2.6831846,1.8673514,1.0533313,0.2374981,0.19036107,0.14322405,0.09427405,0.047137026,0.0,0.0,0.0,0.0,0.0,0.0,0.034446288,0.07070554,0.10515183,0.13959812,0.17585737,0.13959812,0.10515183,0.07070554,0.034446288,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.072518505,0.14503701,0.21755551,0.29007402,0.36259252,0.2991388,0.2374981,0.17585737,0.11240368,0.05076295,0.19036107,0.32995918,0.46955732,0.6091554,0.7505665,0.62184614,0.4949388,0.3680314,0.23931105,0.11240368,0.8466535,1.5827163,2.3169663,3.053029,3.787279,3.1400511,2.4928236,1.845596,1.1983683,0.5493277,0.4405499,0.32995918,0.21936847,0.11059072,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.73968875,1.4793775,2.220879,2.960568,3.7002566,3.1908143,2.6795588,2.1701162,1.6606737,1.1494182,1.2455053,1.3397794,1.4358664,1.5301404,1.6244144,1.3905423,1.1548572,0.91917205,0.6852999,0.44961473,0.38434806,0.3208944,0.25562772,0.19036107,0.12509441,0.11784257,0.11059072,0.10333887,0.09427405,0.0870222,0.34083697,0.59283876,0.8448406,1.0968424,1.3506571,2.0432088,2.7357605,3.4283123,4.120864,4.8116026,3.930503,3.04759,2.1646774,1.2817645,0.40066472,1.1204109,1.840157,2.5599031,3.2796493,3.9993954,3.8398547,3.680314,3.5207734,3.3594196,3.199879,2.762955,2.324218,1.887294,1.4503701,1.0116332,0.968122,0.922798,0.8774739,0.8321498,0.7868258,0.7179332,0.64722764,0.57833505,0.5076295,0.43692398,1.4666867,2.4982624,3.5280252,4.557788,5.5875506,5.6491914,5.712645,5.774286,5.8377395,5.89938,5.6056805,5.3101673,5.0146546,4.7191415,4.4254417,4.6176157,4.8097897,5.0019636,5.1941376,5.388125,5.482399,5.576673,5.67276,5.767034,5.863121,6.1423173,6.4233265,6.7025228,6.981719,7.262728,6.8421206,6.4233265,6.002719,5.582112,5.163317,5.0599785,4.95664,4.855114,4.751775,4.650249,4.1516843,3.6549325,3.1581807,2.659616,2.1628644,1.9326181,1.7023718,1.4721256,1.2418793,1.0116332,0.83940166,0.6671702,0.4949388,0.32270733,0.15047589,0.12690738,0.10515183,0.08339628,0.059827764,0.038072214,0.032633327,0.027194439,0.02175555,0.018129626,0.012690738,0.07070554,0.12690738,0.18492219,0.24293698,0.2991388,0.36984438,0.4405499,0.5094425,0.58014804,0.6508536,0.52032024,0.38978696,0.25925365,0.13053331,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.07795739,0.10515183,0.13234627,0.15954071,0.18673515,0.28463513,0.3825351,0.48043507,0.57833505,0.6744221,0.6653573,0.6544795,0.64541465,0.6345369,0.62547207,0.7850128,0.9445535,1.1040943,1.2654479,1.4249886,2.1193533,2.8155308,3.5098956,4.2042603,4.900438,4.6357455,4.36924,4.1045475,3.8398547,3.5751622,3.299592,3.0258346,2.7502642,2.474694,2.1991236,2.08672,1.9743162,1.8619126,1.7495089,1.6371052,1.7295663,1.8220274,1.9144884,2.0069497,2.0994108,2.1683033,2.2353828,2.3024626,2.3695421,2.4366217,3.1327994,3.827164,4.5233417,5.217706,5.9120708,5.422571,4.933071,4.441758,3.9522583,3.4627585,3.5117085,3.5624714,3.6132345,3.6621845,3.7129474,3.5425289,3.3721104,3.2016919,3.0330863,2.8626678,2.7031271,2.5417736,2.382233,2.222692,2.0631514,8.624263,8.138389,7.650702,7.1630154,6.6753283,6.187641,6.037165,5.8866897,5.7380266,5.5875506,5.4370747,7.1865835,8.937905,10.687414,12.436923,14.188245,14.211814,14.237195,14.262577,14.287958,14.313339,15.074784,15.838041,16.599485,17.362743,18.124187,17.27572,16.425442,15.575162,14.724882,13.874602,12.812206,11.74981,10.687414,9.625018,8.562622,8.174648,7.7866745,7.400513,7.0125394,6.624565,6.1241875,5.6256227,5.125245,4.6248674,4.12449,3.299592,2.474694,1.649796,0.824898,0.0,0.6000906,1.2001812,1.8002719,2.4003625,3.000453,3.6132345,4.2242026,4.836984,5.4497657,6.0625467,5.712645,5.3627434,5.0128417,4.6629395,4.313038,4.249584,4.1879435,4.12449,4.062849,3.9993954,3.6621845,3.3249733,2.9877625,2.6505513,2.3133402,2.275268,2.2371957,2.1991236,2.1628644,2.124792,2.137483,2.1501737,2.1628644,2.175555,2.1882458,2.03777,1.887294,1.7368182,1.5881553,1.4376793,1.4122978,1.3869164,1.3633479,1.3379664,1.3125849,1.3996071,1.4866294,1.5754645,1.6624867,1.7495089,1.4376793,1.1258497,0.8122072,0.50037766,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.31182957,0.62547207,0.93730164,1.2491312,1.5627737,1.4122978,1.261822,1.1131591,0.96268314,0.8122072,1.062396,1.3125849,1.5627737,1.8129625,2.0631514,3.3249733,4.5867953,5.8504305,7.112252,8.375887,7.4875355,6.599184,5.712645,4.8242936,3.9377546,4.6248674,5.3119802,6.000906,6.688019,7.3751316,6.825804,6.2746634,5.7253356,5.1741953,4.6248674,5.0998635,5.57486,6.049856,6.5248523,6.9998484,5.7869763,4.5759177,3.3630457,2.1501737,0.93730164,1.3869164,1.8383441,2.2879589,2.7375734,3.1871881,3.7256382,4.262275,4.800725,5.337362,5.8758116,5.5005283,5.125245,4.749962,4.3746786,3.9993954,3.2633326,2.525457,1.7875811,1.0497054,0.31182957,1.2128719,2.1121013,3.0131438,3.9123733,4.8116026,5.999093,7.1865835,8.375887,9.563377,10.750868,8.600695,6.450521,4.3003473,2.1501737,0.0,1.2872034,2.5744069,3.8634233,5.1506267,6.43783,5.1506267,3.8634233,2.5744069,1.2872034,0.0,0.3245203,0.6508536,0.97537386,1.2998942,1.6244144,1.5754645,1.5247015,1.4757515,1.4249886,1.3742256,5.5367875,9.699349,13.861912,18.024473,22.187037,24.799515,27.411995,30.024473,32.63695,35.24943,35.075386,34.89953,34.725487,34.54963,34.375584,31.525606,28.675629,25.825651,22.975676,20.125698,19.92446,19.725033,19.525606,19.324368,19.124943,18.45052,17.774284,17.099863,16.425442,15.749206,15.674874,15.600543,15.524399,15.4500675,15.375735,14.275268,13.174799,12.07433,10.975676,9.875207,10.125396,10.375585,10.625773,10.874149,11.124338,10.449916,9.775495,9.099259,8.424837,7.750415,7.911769,8.074935,8.238102,8.399456,8.562622,10.475298,12.387974,14.300649,16.213324,18.124187,17.424383,16.72458,16.024776,15.324973,14.625169,13.3506565,12.07433,10.799818,9.525306,8.2507925,6.7623506,5.275721,3.787279,2.3006494,0.8122072,0.6508536,0.48768693,0.3245203,0.16316663,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.2374981,0.41335547,0.5873999,0.76325727,0.93730164,0.774135,0.61278135,0.44961473,0.28826106,0.12509441,1.0243238,1.9253663,2.8245957,3.7256382,4.6248674,3.8380418,3.049403,2.2625773,1.4757515,0.6871128,0.5493277,0.41335547,0.2755703,0.13778515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.824898,1.649796,2.474694,3.299592,4.12449,3.5008307,2.8753586,2.2498865,1.6244144,1.0007553,1.1747998,1.3506571,1.5247015,1.7005589,1.8746033,1.6008459,1.3252757,1.0497054,0.774135,0.50037766,0.42423326,0.34990177,0.2755703,0.19942589,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.387974,0.7124943,1.0370146,1.3633479,1.6878681,2.2118144,2.7375734,3.2633326,3.787279,4.313038,3.5497808,2.7883365,2.0250793,1.261822,0.50037766,1.3742256,2.2498865,3.1255474,3.9993954,4.8750563,4.4870825,4.099108,3.7129474,3.3249733,2.9369993,2.5000753,2.0631514,1.6244144,1.1874905,0.7505665,0.6000906,0.44961473,0.2991388,0.15047589,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.87566096,1.6878681,2.5000753,3.3122826,4.12449,3.8507326,3.5751622,3.299592,3.0258346,2.7502642,2.3876717,2.0250793,1.6624867,1.2998942,0.93730164,1.4122978,1.887294,2.3622901,2.8372865,3.3122826,3.7256382,4.137181,4.550536,4.9620786,5.375434,5.7380266,6.1006193,6.4632115,6.825804,7.1883965,6.787732,6.3870673,5.9882154,5.5875506,5.186886,5.237649,5.2865987,5.337362,5.388125,5.4370747,4.8750563,4.313038,3.7492065,3.1871881,2.6251698,2.324218,2.0250793,1.7241274,1.4249886,1.1258497,0.93730164,0.7505665,0.5620184,0.37528324,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.0,0.0,0.0,0.0,0.0,0.07433146,0.15047589,0.22480737,0.2991388,0.37528324,0.46230546,0.5493277,0.63816285,0.72518504,0.8122072,0.6508536,0.48768693,0.3245203,0.16316663,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.17585737,0.28826106,0.40066472,0.51306844,0.62547207,0.63816285,0.6508536,0.66173136,0.6744221,0.6871128,0.7124943,0.73787576,0.76325727,0.7868258,0.8122072,1.3252757,1.8383441,2.3495996,2.8626678,3.3757362,3.0874753,2.7992141,2.5127661,2.2245052,1.938057,1.987007,2.03777,2.08672,2.137483,2.1882458,1.9616255,1.7368182,1.5120108,1.2872034,1.062396,1.2491312,1.4376793,1.6244144,1.8129625,1.9996977,2.1121013,2.2245052,2.3369088,2.4493124,2.561716,3.000453,3.437377,3.874301,4.313038,4.749962,4.4254417,4.099108,3.774588,3.4500678,3.1255474,3.2125697,3.299592,3.386614,3.4754493,3.5624714,3.3249733,3.0874753,2.8499773,2.612479,2.374981,2.137483,1.8999848,1.6624867,1.4249886,1.1874905,8.52455,7.9842873,7.4458375,6.9055743,6.3653116,5.825049,5.718084,5.6093063,5.5023413,5.3953767,5.2865987,6.735156,8.1819,9.630457,11.077202,12.525759,12.567456,12.609155,12.652666,12.694364,12.737875,13.68968,14.643299,15.595104,16.54691,17.500528,16.36924,15.239763,14.110288,12.980812,11.849524,11.080828,10.310318,9.539809,8.7693,8.000604,7.574558,7.1503243,6.7242785,6.300045,5.8758116,5.371808,4.8696175,4.367427,3.8652363,3.3630457,2.7176309,2.0722163,1.4268016,0.78319985,0.13778515,0.6200332,1.1022812,1.5845293,2.0667772,2.5508385,3.0983531,3.6458678,4.1933823,4.740897,5.2865987,5.1107416,4.933071,4.7554007,4.5777307,4.40006,4.441758,4.4852695,4.5269675,4.5704784,4.612177,4.1480584,3.682127,3.2180085,2.752077,2.2879589,2.18462,2.0830941,1.9797552,1.8782293,1.7748904,1.8147756,1.8546607,1.8945459,1.9344311,1.9743162,1.8655385,1.7549478,1.6443571,1.5355793,1.4249886,1.4177368,1.4104849,1.403233,1.3941683,1.3869164,1.4141108,1.4431182,1.4703126,1.4975071,1.5247015,1.2491312,0.97537386,0.69980353,0.42423326,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.027194439,0.054388877,0.08339628,0.11059072,0.13778515,0.43692398,0.73787576,1.0370146,1.3379664,1.6371052,1.5228885,1.4068589,1.2926424,1.1766127,1.062396,1.2527572,1.4431182,1.6316663,1.8220274,2.0123885,3.2016919,4.3928084,5.582112,6.773228,7.9625316,6.9998484,6.037165,5.0744824,4.1117992,3.149116,3.7002566,4.249584,4.800725,5.3500524,5.89938,5.565795,5.230397,4.894999,4.559601,4.2242026,4.550536,4.8750563,5.199577,5.524097,5.8504305,4.98746,4.12449,3.2633326,2.4003625,1.5373923,2.039583,2.5417736,3.045777,3.5479677,4.0501585,4.273153,4.494334,4.7173285,4.940323,5.163317,5.6981416,6.2329655,6.7677894,7.3026133,7.837437,6.735156,5.632875,4.5305934,3.4283123,2.324218,2.8445382,3.3648586,3.8851788,4.405499,4.9258194,5.814171,6.7043357,7.5945,8.484665,9.374829,7.590874,5.805106,4.019338,2.2353828,0.44961473,1.4630609,2.474694,3.48814,4.499773,5.5132194,4.41819,3.3231604,2.228131,1.1331016,0.038072214,0.29732585,0.55839247,0.81764615,1.0768998,1.3379664,1.2908293,1.2418793,1.1947423,1.1476053,1.1004683,4.9294453,8.760235,12.589212,16.420002,20.250792,22.069193,23.889408,25.709621,27.529837,29.350052,29.712645,30.075235,30.437828,30.80042,31.163013,28.202446,25.241879,22.283123,19.322556,16.361988,16.757214,17.15244,17.547665,17.94289,18.338116,17.513218,16.68832,15.861609,15.036712,14.211814,14.064963,13.918114,13.769451,13.622601,13.475751,12.516694,11.559449,10.602205,9.644961,8.6877165,8.749357,8.812811,8.874452,8.937905,8.999546,8.479226,7.9607186,7.440398,6.9200783,6.399758,6.5701766,6.740595,6.9092,7.079619,7.250037,8.832754,10.41547,11.998186,13.57909,15.161806,14.554463,13.947122,13.339779,12.732436,12.125093,11.019187,9.915092,8.809185,7.705091,6.599184,5.40988,4.220577,3.0294604,1.840157,0.6508536,0.533011,0.41516843,0.29732585,0.1794833,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.047137026,0.09427405,0.14322405,0.19036107,0.2374981,0.21030366,0.18310922,0.15410182,0.12690738,0.099712946,0.10333887,0.10515183,0.10696479,0.11059072,0.11240368,0.17585737,0.2374981,0.2991388,0.36259252,0.42423326,0.34990177,0.2755703,0.19942589,0.12509441,0.05076295,0.19036107,0.32995918,0.46955732,0.6091554,0.7505665,1.6697385,2.5907235,3.5098956,4.4308805,5.3500524,5.040036,4.7300196,4.420003,4.1099863,3.7999697,3.1817493,2.565342,1.9471219,1.3307146,0.7124943,0.6200332,0.5275721,0.43511102,0.34264994,0.25018883,0.2955129,0.34083697,0.38434806,0.42967212,0.4749962,0.38072214,0.28463513,0.19036107,0.09427405,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.11784257,0.23568514,0.35171473,0.46955732,0.5873999,1.2056202,1.8220274,2.4402475,3.056655,3.6748753,3.2869012,2.9007401,2.5127661,2.124792,1.7368182,1.7096237,1.6824293,1.6552348,1.6280404,1.6008459,1.3597219,1.1204109,0.8792868,0.6399758,0.40066472,0.34264994,0.28463513,0.22662032,0.17041849,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.05076295,0.31182957,0.5747091,0.8375887,1.1004683,1.3633479,1.938057,2.5127661,3.0874753,3.6621845,4.2368937,4.0356545,3.832603,3.6295512,3.4283123,3.2252605,4.1281157,5.029158,5.9320135,6.834869,7.7377243,7.0868707,6.43783,5.7869763,5.137936,4.4870825,4.0320287,3.576975,3.1219215,2.666868,2.2118144,1.8691645,1.5283275,1.1856775,0.8430276,0.50037766,0.48768693,0.4749962,0.46230546,0.44961473,0.43692398,1.0732739,1.7078108,2.3423476,2.9768846,3.6132345,3.3304121,3.04759,2.764768,2.4819458,2.1991236,1.9108626,1.6207886,1.3307146,1.0406405,0.7505665,1.1294757,1.5101979,1.889107,2.269829,2.6505513,2.9805105,3.3104696,3.6404288,3.9703882,4.3003473,4.590421,4.880495,5.1705694,5.4606433,5.750717,5.429823,5.1107416,4.7898474,4.4707656,4.1498713,4.1897564,4.229642,4.269527,4.309412,4.349297,4.022964,3.6948178,3.3666716,3.0403383,2.712192,2.7466383,2.7828975,2.817344,2.8517902,2.8880494,2.6251698,2.3622901,2.0994108,1.8383441,1.5754645,1.3851035,1.1947423,1.0043813,0.81583315,0.62547207,0.50219065,0.38072214,0.2574407,0.13415924,0.012690738,0.24837588,0.48224804,0.7179332,0.95180535,1.1874905,1.3307146,1.4721256,1.6153497,1.7567607,1.8999848,1.5954071,1.2908293,0.98443866,0.67986095,0.37528324,0.2991388,0.22480737,0.15047589,0.07433146,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.072518505,0.07070554,0.06707962,0.065266654,0.06164073,0.15047589,0.2374981,0.3245203,0.41335547,0.50037766,0.5094425,0.52032024,0.5293851,0.5402629,0.5493277,0.56927025,0.58921283,0.6091554,0.629098,0.6508536,1.2545701,1.8600996,2.465629,3.0693457,3.6748753,3.2597067,2.8445382,2.42937,2.0142014,1.6008459,1.7078108,1.8147756,1.9217403,2.030518,2.137483,1.987007,1.8383441,1.6878681,1.5373923,1.3869164,1.4358664,1.4830034,1.5301404,1.5772774,1.6244144,1.8474089,2.0704033,2.2933977,2.514579,2.7375734,3.0892882,3.442816,3.7945306,4.1480584,4.499773,4.2894692,4.079166,3.870675,3.6603715,3.4500678,3.5570326,3.6658103,3.7727752,3.87974,3.9867048,3.720199,3.4518807,3.1853752,2.9170568,2.6505513,2.6849976,2.7194438,2.7557032,2.7901495,2.8245957,8.424837,7.8319983,7.2391596,6.6481338,6.055295,5.462456,5.3971896,5.331923,5.2666564,5.2032027,5.137936,6.281915,7.4277077,8.571687,9.71748,10.863272,10.9230995,10.982927,11.042755,11.102583,11.162411,12.304577,13.446743,14.590723,15.732889,16.875055,15.464571,14.055899,12.645414,11.234929,9.824444,9.347635,8.870826,8.392203,7.915395,7.4367723,6.9744673,6.5121617,6.049856,5.5875506,5.125245,4.6194286,4.115425,3.6096084,3.105605,2.5997884,2.13567,1.6697385,1.2056202,0.73968875,0.2755703,0.6399758,1.0043813,1.3705997,1.7350051,2.0994108,2.5816586,3.0657198,3.5479677,4.0302157,4.512464,4.507025,4.503399,4.49796,4.4925213,4.4870825,4.6357455,4.782595,4.9294453,5.0781083,5.224958,4.632119,4.0392804,3.4482548,2.855416,2.2625773,2.0957847,1.9271792,1.7603867,1.5917811,1.4249886,1.4920682,1.5591478,1.6280404,1.69512,1.7621996,1.693307,1.6226015,1.551896,1.4830034,1.4122978,1.4231756,1.4322405,1.4431182,1.452183,1.4630609,1.4304274,1.3977941,1.3651608,1.3325275,1.2998942,1.062396,0.824898,0.5873999,0.34990177,0.11240368,0.09064813,0.06707962,0.045324065,0.02175555,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.054388877,0.11059072,0.16497959,0.21936847,0.2755703,0.5620184,0.85027945,1.1367276,1.4249886,1.7132497,1.6316663,1.551896,1.4721256,1.3923552,1.3125849,1.4431182,1.5718386,1.7023718,1.8329052,1.9616255,3.0802233,4.1970086,5.315606,6.432391,7.549176,6.5121617,5.475147,4.4381323,3.3993049,2.3622901,2.7756457,3.1871881,3.6005437,4.0120864,4.4254417,4.305786,4.1843176,4.064662,3.9450066,3.825351,3.9993954,4.175253,4.349297,4.5251546,4.699199,4.1879435,3.6748753,3.1618068,2.6505513,2.137483,2.6922495,3.247016,3.8017826,4.358362,4.9131284,4.8206677,4.7282066,4.6357455,4.5432844,4.4508233,5.8957543,7.3406854,8.785617,10.230548,11.675479,10.20698,8.740293,7.271793,5.805106,4.3384194,4.478018,4.6176157,4.7572136,4.896812,5.038223,5.6292486,6.2220874,6.814926,7.407765,8.000604,6.5792413,5.1596913,3.7401419,2.3205922,0.89922947,1.6371052,2.374981,3.1128569,3.8507326,4.5867953,3.6857529,2.7828975,1.8800422,0.97718686,0.07433146,0.27013144,0.46411842,0.65991837,0.8557183,1.0497054,1.0043813,0.96087015,0.9155461,0.87022203,0.824898,4.322103,7.819308,11.318325,14.81553,18.312735,19.340685,20.366821,21.394772,22.422722,23.45067,24.349901,25.24913,26.150173,27.049402,27.950443,24.879286,21.80994,18.740595,15.6694355,12.60009,13.589968,14.579845,15.569723,16.5596,17.549479,16.574104,15.600543,14.625169,13.649796,12.674421,12.455053,12.235684,12.0145035,11.795135,11.575767,10.7599325,9.945912,9.130079,8.314246,7.500226,7.3751316,7.250037,7.124943,6.9998484,6.874754,6.510349,6.14413,5.7797246,5.4153194,5.049101,5.2267714,5.4044414,5.582112,5.7597823,5.9374523,7.1902094,8.442966,9.695724,10.946668,12.199425,11.684544,11.169662,10.654781,10.139899,9.625018,8.689529,7.755854,6.8203654,5.8848767,4.949388,4.0574102,3.1654327,2.2716422,1.3796645,0.48768693,0.41516843,0.34264994,0.27013144,0.19761293,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.09427405,0.19036107,0.28463513,0.38072214,0.4749962,0.39522585,0.3154555,0.23568514,0.15410182,0.07433146,0.10515183,0.13415924,0.16497959,0.19579996,0.22480737,0.34990177,0.4749962,0.6000906,0.72518504,0.85027945,0.6871128,0.52575916,0.36259252,0.19942589,0.038072214,0.14322405,0.24837588,0.35171473,0.45686656,0.5620184,2.565342,4.5668526,6.5701766,8.571687,10.57501,9.055748,7.5346723,6.01541,4.494334,2.9750717,2.5272698,2.079468,1.6316663,1.1856775,0.73787576,0.69073874,0.6417888,0.5946517,0.5475147,0.50037766,0.58921283,0.67986095,0.7705091,0.85934424,0.9499924,0.75963134,0.56927025,0.38072214,0.19036107,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.23568514,0.46955732,0.70524246,0.93911463,1.1747998,1.5845293,1.9942589,2.4058013,2.8155308,3.2252605,3.0747845,2.9243085,2.7756457,2.6251698,2.474694,2.2444477,2.0142014,1.7857682,1.5555218,1.3252757,1.1204109,0.9155461,0.7106813,0.5058166,0.2991388,0.25925365,0.21936847,0.1794833,0.13959812,0.099712946,0.0870222,0.07433146,0.06164073,0.05076295,0.038072214,0.2374981,0.43692398,0.63816285,0.8375887,1.0370146,1.6624867,2.2879589,2.911618,3.53709,4.162562,4.519716,4.876869,5.235836,5.5929894,5.9501433,6.880193,7.8102427,8.740293,9.670342,10.600392,9.686659,8.774739,7.8628187,6.9508986,6.037165,5.565795,5.092612,4.6194286,4.1480584,3.6748753,3.1400511,2.6052272,2.0704033,1.5355793,1.0007553,0.96268314,0.9246109,0.8883517,0.85027945,0.8122072,1.2708868,1.7277533,2.18462,2.6432993,3.100166,2.810092,2.520018,2.229944,1.93987,1.649796,1.4322405,1.214685,0.99712944,0.7795739,0.5620184,0.8466535,1.1331016,1.4177368,1.7023718,1.987007,2.2353828,2.4819458,2.7303216,2.9768846,3.2252605,3.442816,3.6603715,3.877927,4.0954823,4.313038,4.071914,3.832603,3.5932918,3.3521678,3.1128569,3.141864,3.1726844,3.2016919,3.2325122,3.2633326,3.1708715,3.0765975,2.9841363,2.8916752,2.7992141,3.1708715,3.540716,3.9105604,4.2804046,4.650249,4.313038,3.975827,3.636803,3.299592,2.962381,2.619731,2.277081,1.9344311,1.5917811,1.2491312,1.0043813,0.75963134,0.5148814,0.27013144,0.025381476,0.42060733,0.81583315,1.209246,1.6044719,1.9996977,2.1973107,2.3949237,2.5925364,2.7901495,2.9877625,2.5399606,2.0921588,1.6443571,1.1983683,0.7505665,0.6000906,0.44961473,0.2991388,0.15047589,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.018129626,0.034446288,0.052575916,0.07070554,0.0870222,0.08339628,0.07795739,0.072518505,0.06707962,0.06164073,0.12509441,0.18673515,0.25018883,0.31182957,0.37528324,0.3825351,0.38978696,0.39703882,0.40429065,0.41335547,0.42785916,0.44236287,0.45686656,0.47318324,0.48768693,1.1856775,1.8818551,2.5798457,3.2778363,3.975827,3.4319382,2.8898623,2.3477864,1.8057107,1.261822,1.4268016,1.5917811,1.7567607,1.9217403,2.08672,2.0123885,1.938057,1.8619126,1.7875811,1.7132497,1.6207886,1.5283275,1.4358664,1.3434052,1.2491312,1.5827163,1.9144884,2.2480736,2.5798457,2.911618,3.1799364,3.4482548,3.7147603,3.9830787,4.249584,4.15531,4.059223,3.9649491,3.870675,3.774588,3.9033084,4.0302157,4.157123,4.2858434,4.4127507,4.115425,3.8180993,3.5207734,3.2216346,2.9243085,3.2325122,3.540716,3.8471067,4.15531,4.461701,8.325124,7.6797094,7.0342946,6.390693,5.7452784,5.0998635,5.0781083,5.0545397,5.032784,5.009216,4.98746,5.8304877,6.6717024,7.51473,8.357758,9.200785,9.27693,9.354887,9.432844,9.510801,9.5869465,10.919474,12.252001,13.584529,14.917056,16.249584,14.559902,12.870221,11.18054,9.490859,7.799365,7.614443,7.4295206,7.2445984,7.059676,6.874754,6.3743763,5.8758116,5.375434,4.8750563,4.3746786,3.8670492,3.3594196,2.8517902,2.3441606,1.8383441,1.551896,1.2672608,0.9826257,0.6979906,0.41335547,0.65991837,0.90829426,1.1548572,1.403233,1.649796,2.0667772,2.4855716,2.902553,3.3195345,3.738329,3.9051213,4.071914,4.2405195,4.407312,4.574105,4.8279195,5.0799212,5.331923,5.5857377,5.8377395,5.1179934,4.3982472,3.6766882,2.956942,2.2371957,2.0051367,1.7730774,1.5392052,1.3071461,1.0750868,1.1693609,1.2654479,1.3597219,1.455809,1.550083,1.5192627,1.4902552,1.4594349,1.4304274,1.3996071,1.4268016,1.455809,1.4830034,1.5101979,1.5373923,1.4449311,1.35247,1.260009,1.167548,1.0750868,0.87566096,0.6744221,0.4749962,0.2755703,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08339628,0.16497959,0.24837588,0.32995918,0.41335547,0.6871128,0.96268314,1.2382535,1.5120108,1.7875811,1.742257,1.696933,1.651609,1.6080978,1.5627737,1.6316663,1.7023718,1.7730774,1.84197,1.9126755,2.956942,4.0030212,5.047288,6.093367,7.137634,6.0244746,4.9131284,3.7999697,2.6868105,1.5754645,1.8492218,2.124792,2.4003625,2.6741197,2.94969,3.045777,3.1400511,3.2343252,3.3304121,3.4246864,3.4500678,3.4754493,3.5008307,3.5243993,3.5497808,3.386614,3.2252605,3.0620937,2.9007401,2.7375734,3.3449159,3.9522583,4.559601,5.1669436,5.774286,5.368182,4.9602656,4.552349,4.1444325,3.738329,6.093367,8.446592,10.803444,13.15667,15.511708,13.680615,11.847711,10.014805,8.1819,6.350808,6.109684,5.870373,5.6292486,5.389938,5.1506267,5.4443264,5.7398396,6.035352,6.3308654,6.624565,5.569421,4.514277,3.4591327,2.4058013,1.3506571,1.8129625,2.275268,2.7375734,3.199879,3.6621845,2.953316,2.2426348,1.5319533,0.823085,0.11240368,0.24293698,0.37165734,0.50219065,0.6327239,0.76325727,0.7197462,0.678048,0.6345369,0.59283876,0.5493277,3.7147603,6.880193,10.045626,13.209246,16.374678,16.610363,16.844234,17.07992,17.315605,17.549479,18.987158,20.424837,21.862516,23.300196,24.737875,21.557938,18.378002,15.198066,12.018129,8.838193,10.422722,12.007251,13.591781,15.1781225,16.762651,15.636803,14.512766,13.386916,12.262879,11.137029,10.845142,10.553255,10.259555,9.967669,9.675781,9.003172,8.330563,7.6579537,6.985345,6.3127356,6.000906,5.6872635,5.375434,5.0617914,4.749962,4.539658,4.329355,4.120864,3.9105604,3.7002566,3.8851788,4.070101,4.255023,4.439945,4.6248674,5.5476656,6.4704633,7.3932614,8.314246,9.237044,8.814624,8.392203,7.9697833,7.5473633,7.124943,6.359873,5.5948024,4.8297324,4.064662,3.299592,2.70494,2.1102884,1.5156367,0.91917205,0.3245203,0.29732585,0.27013144,0.24293698,0.21574254,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14322405,0.28463513,0.42785916,0.56927025,0.7124943,0.58014804,0.44780177,0.3154555,0.18310922,0.05076295,0.10696479,0.16497959,0.2229944,0.27919623,0.33721104,0.52575916,0.7124943,0.89922947,1.0877775,1.2745126,1.0243238,0.774135,0.52575916,0.2755703,0.025381476,0.09427405,0.16497959,0.23568514,0.3045777,0.37528324,3.4609456,6.544795,9.630457,12.714307,15.799969,13.069647,10.339326,7.609004,4.880495,2.1501737,1.8727903,1.5954071,1.3180238,1.0406405,0.76325727,0.75963134,0.75781834,0.7541924,0.7523795,0.7505665,0.88472575,1.020698,1.1548572,1.2908293,1.4249886,1.1403534,0.8557183,0.56927025,0.28463513,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.35171473,0.70524246,1.0569572,1.4104849,1.7621996,1.9652514,2.1683033,2.3695421,2.572594,2.7756457,2.8626678,2.94969,3.0367124,3.1255474,3.2125697,2.7792716,2.3477864,1.9144884,1.4830034,1.0497054,0.8792868,0.7106813,0.5402629,0.36984438,0.19942589,0.17767033,0.15410182,0.13234627,0.11059072,0.0870222,0.07433146,0.06164073,0.05076295,0.038072214,0.025381476,0.16316663,0.2991388,0.43692398,0.5747091,0.7124943,1.3869164,2.0631514,2.7375734,3.4119956,4.0882306,5.0055895,5.922949,6.8403077,7.757667,8.675026,9.63227,10.589515,11.546759,12.5058155,13.46306,12.28826,11.111648,9.936848,8.762048,7.5872483,7.0977483,6.6082487,6.1169357,5.6274357,5.137936,4.409125,3.682127,2.955129,2.228131,1.49932,1.4376793,1.3742256,1.3125849,1.2491312,1.1874905,1.4666867,1.7476959,2.0268922,2.3079014,2.5870976,2.2897718,1.9924458,1.69512,1.3977941,1.1004683,0.9554313,0.8103943,0.6653573,0.52032024,0.37528324,0.5656443,0.7541924,0.9445535,1.1349145,1.3252757,1.4902552,1.6552348,1.8202144,1.9851941,2.1501737,2.2952106,2.4402475,2.5852847,2.7303216,2.8753586,2.715818,2.5544643,2.3949237,2.2353828,2.0758421,2.0957847,2.1157274,2.13567,2.1556125,2.175555,2.3169663,2.4601903,2.6016014,2.7448254,2.8880494,3.5932918,4.2967215,5.0019636,5.7072062,6.412449,5.999093,5.5875506,5.1741953,4.762653,4.349297,3.8543584,3.3594196,2.864481,2.3695421,1.8746033,1.5065719,1.1403534,0.77232206,0.40429065,0.038072214,0.59283876,1.1476053,1.7023718,2.2571385,2.811905,3.0657198,3.3177216,3.5697234,3.8217251,4.07554,3.484514,2.8953013,2.3042755,1.7150626,1.1258497,0.89922947,0.6744221,0.44961473,0.22480737,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.092461094,0.08520924,0.07795739,0.07070554,0.06164073,0.099712946,0.13778515,0.17585737,0.21211663,0.25018883,0.25562772,0.25925365,0.26469254,0.27013144,0.2755703,0.28463513,0.2955129,0.3045777,0.3154555,0.3245203,1.114972,1.9054236,2.6958754,3.484514,4.274966,3.6041696,2.9351864,2.2643902,1.5954071,0.9246109,1.1476053,1.3705997,1.5917811,1.8147756,2.03777,2.03777,2.03777,2.03777,2.03777,2.03777,1.8057107,1.5718386,1.3397794,1.1077201,0.87566096,1.3180238,1.7603867,2.2027495,2.6451125,3.0874753,3.2705846,3.4518807,3.63499,3.8180993,3.9993954,4.019338,4.0392804,4.059223,4.079166,4.099108,4.2477713,4.3946214,4.5432844,4.690134,4.836984,4.510651,4.1825047,3.8543584,3.5280252,3.199879,3.780027,4.360175,4.940323,5.520471,6.1006193,8.225411,7.5274205,6.82943,6.1332526,5.4352617,4.7372713,4.7572136,4.7771564,4.797099,4.8170414,4.836984,5.377247,5.91751,6.4577727,6.9980354,7.5382986,7.6325727,7.7268467,7.8229337,7.9172077,8.013294,9.53437,11.057259,12.580148,14.103036,15.624111,13.655234,11.684544,9.715667,7.744976,5.774286,5.883064,5.9900284,6.096993,6.205771,6.3127356,5.774286,5.237649,4.699199,4.162562,3.6241121,3.1146698,2.6052272,2.0957847,1.5845293,1.0750868,0.969935,0.86478317,0.75963134,0.6544795,0.5493277,0.67986095,0.8103943,0.93911463,1.0696479,1.2001812,1.551896,1.9054236,2.2571385,2.610666,2.962381,3.303218,3.6422417,3.9830787,4.322103,4.6629395,5.0200934,5.377247,5.7344007,6.093367,6.450521,5.6020546,4.7554007,3.9069343,3.0602808,2.2118144,1.9144884,1.6171626,1.3198367,1.0225109,0.72518504,0.8466535,0.969935,1.0932164,1.214685,1.3379664,1.3470312,1.357909,1.3669738,1.3778516,1.3869164,1.4322405,1.4775645,1.5228885,1.5682126,1.6117238,1.4594349,1.3071461,1.1548572,1.0025684,0.85027945,0.6871128,0.52575916,0.36259252,0.19942589,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.11059072,0.21936847,0.32995918,0.4405499,0.5493277,0.8122072,1.0750868,1.3379664,1.6008459,1.8619126,1.8528478,1.84197,1.8329052,1.8220274,1.8129625,1.8220274,1.8329052,1.84197,1.8528478,1.8619126,2.8354735,3.8072214,4.780782,5.75253,6.7242785,5.5367875,4.349297,3.1618068,1.9743162,0.7868258,0.9246109,1.062396,1.2001812,1.3379664,1.4757515,1.7857682,2.0957847,2.4058013,2.715818,3.0258346,2.9007401,2.7756457,2.6505513,2.525457,2.4003625,2.5870976,2.7756457,2.962381,3.149116,3.3376641,3.9975824,4.6575007,5.317419,5.977338,6.637256,5.915697,5.1923246,4.4707656,3.7473936,3.0258346,6.2891674,9.554313,12.819458,16.084604,19.34975,17.15244,14.955129,12.757817,10.560507,8.363196,7.743163,7.12313,6.5030966,5.883064,5.2630305,5.2594047,5.2575917,5.2557783,5.2521524,5.2503395,4.559601,3.870675,3.1799364,2.4891977,1.8002719,1.987007,2.175555,2.3622901,2.5508385,2.7375734,2.220879,1.7023718,1.1856775,0.6671702,0.15047589,0.21574254,0.27919623,0.3444629,0.40972954,0.4749962,0.43511102,0.39522585,0.35534066,0.3154555,0.2755703,3.1074178,5.9392653,8.772926,11.6047735,14.436621,13.880041,13.321649,12.76507,12.206677,11.650098,13.6244135,15.600543,17.57486,19.549175,21.525305,18.234777,14.94425,11.655537,8.365009,5.0744824,7.2554765,9.434657,11.615651,13.794832,15.975826,14.699501,13.424988,12.1504755,10.874149,9.599637,9.235231,8.870826,8.504607,8.140202,7.7757964,7.2445984,6.7152133,6.185828,5.65463,5.125245,4.6248674,4.12449,3.6241121,3.1255474,2.6251698,2.570781,2.514579,2.4601903,2.4058013,2.3495996,2.5417736,2.7357605,2.9279346,3.1201086,3.3122826,3.9051213,4.49796,5.090799,5.6818247,6.2746634,5.9447045,5.614745,5.2847857,4.954827,4.6248674,4.0302157,3.435564,2.8390994,2.2444477,1.649796,1.35247,1.0551442,0.75781834,0.4604925,0.16316663,0.1794833,0.19761293,0.21574254,0.23205921,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.19036107,0.38072214,0.56927025,0.75963134,0.9499924,0.7650702,0.58014804,0.39522585,0.21030366,0.025381476,0.11059072,0.19579996,0.27919623,0.36440548,0.44961473,0.69980353,0.9499924,1.2001812,1.4503701,1.7005589,1.3633479,1.0243238,0.6871128,0.34990177,0.012690738,0.047137026,0.08339628,0.11784257,0.15228885,0.18673515,4.3547363,8.5227375,12.690738,16.856926,21.024927,17.08536,13.145792,9.2044115,5.2648435,1.3252757,1.2183108,1.1095331,1.0025684,0.89560354,0.7868258,0.83033687,0.872035,0.9155461,0.9572442,1.0007553,1.1802386,1.3597219,1.5392052,1.7205015,1.8999848,1.5192627,1.1403534,0.75963134,0.38072214,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.46955732,0.93911463,1.4104849,1.8800422,2.3495996,2.3441606,2.3405347,2.335096,2.3296568,2.324218,2.6505513,2.9750717,3.299592,3.6241121,3.9504454,3.3140955,2.6795588,2.0450218,1.4104849,0.774135,0.6399758,0.5058166,0.36984438,0.23568514,0.099712946,0.09427405,0.09064813,0.08520924,0.07977036,0.07433146,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0870222,0.16316663,0.2374981,0.31182957,0.387974,1.1131591,1.8383441,2.561716,3.2869012,4.0120864,5.4896507,6.967215,8.444779,9.922344,11.399909,12.384347,13.370599,14.355038,15.339477,16.325727,14.888049,13.45037,12.012691,10.57501,9.137331,8.629702,8.122072,7.614443,7.1068134,6.599184,5.6800117,4.76084,3.8398547,2.9206827,1.9996977,1.9126755,1.8256533,1.7368182,1.649796,1.5627737,1.6642996,1.7676386,1.8691645,1.9725033,2.0758421,1.7694515,1.4648738,1.1602961,0.8557183,0.5493277,0.47680917,0.40429065,0.33177215,0.25925365,0.18673515,0.28282216,0.3770962,0.47318324,0.56745726,0.66173136,0.7451276,0.82671094,0.9101072,0.9916905,1.0750868,1.1476053,1.2201238,1.2926424,1.3651608,1.4376793,1.357909,1.2781386,1.1983683,1.1167849,1.0370146,1.0478923,1.0569572,1.067835,1.0768998,1.0877775,1.4648738,1.84197,2.220879,2.5979755,2.9750717,4.0157123,5.0545397,6.09518,7.135821,8.174648,7.686961,7.1992745,6.7134004,6.2257137,5.7380266,5.090799,4.441758,3.7945306,3.147303,2.5000753,2.0105755,1.5192627,1.0297627,0.5402629,0.05076295,0.7650702,1.4793775,2.1954978,2.909805,3.6241121,3.9323158,4.2405195,4.5469103,4.855114,5.163317,4.4290676,3.6966307,2.9641938,2.231757,1.49932,1.2001812,0.89922947,0.6000906,0.2991388,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.10333887,0.092461094,0.08339628,0.072518505,0.06164073,0.07433146,0.0870222,0.099712946,0.11240368,0.12509441,0.12690738,0.13053331,0.13234627,0.13415924,0.13778515,0.14322405,0.14684997,0.15228885,0.15772775,0.16316663,1.0442665,1.9271792,2.810092,3.6930048,4.574105,3.778214,2.9805105,2.182807,1.3851035,0.5873999,0.8684091,1.1476053,1.4268016,1.7078108,1.987007,2.0631514,2.137483,2.2118144,2.2879589,2.3622901,1.9906329,1.6171626,1.2455053,0.872035,0.50037766,1.0533313,1.6044719,2.1574254,2.7103791,3.2633326,3.3594196,3.4573197,3.5552197,3.6531196,3.7492065,3.8851788,4.019338,4.15531,4.2894692,4.4254417,4.592234,4.76084,4.9276323,5.0944247,5.2630305,4.9058766,4.5469103,4.1897564,3.832603,3.4754493,4.327542,5.179634,6.0317264,6.885632,7.7377243,8.125698,7.3751316,6.624565,5.8758116,5.125245,4.3746786,4.4381323,4.499773,4.5632267,4.6248674,4.688321,4.9258194,5.163317,5.4008155,5.638314,5.8758116,5.9882154,6.1006193,6.2130227,6.3254266,6.43783,8.149267,9.862516,11.575767,13.287203,15.000452,12.750566,10.500679,8.2507925,5.999093,3.7492065,4.1498713,4.550536,4.949388,5.3500524,5.750717,5.1741953,4.599486,4.024777,3.4500678,2.8753586,2.3622901,1.8492218,1.3379664,0.824898,0.31182957,0.387974,0.46230546,0.53663695,0.61278135,0.6871128,0.69980353,0.7124943,0.72518504,0.73787576,0.7505665,1.0370146,1.3252757,1.6117238,1.8999848,2.1882458,2.6995013,3.2125697,3.7256382,4.2368937,4.749962,5.2122674,5.674573,6.1368785,6.599184,7.063302,6.0879283,5.1125546,4.137181,3.1618068,2.1882458,1.8256533,1.4630609,1.1004683,0.73787576,0.37528324,0.52575916,0.6744221,0.824898,0.97537386,1.1258497,1.1747998,1.2255627,1.2745126,1.3252757,1.3742256,1.4376793,1.49932,1.5627737,1.6244144,1.6878681,1.4757515,1.261822,1.0497054,0.8375887,0.62547207,0.50037766,0.37528324,0.25018883,0.12509441,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13778515,0.2755703,0.41335547,0.5493277,0.6871128,0.93730164,1.1874905,1.4376793,1.6878681,1.938057,1.9616255,1.987007,2.0123885,2.03777,2.0631514,2.0123885,1.9616255,1.9126755,1.8619126,1.8129625,2.712192,3.6132345,4.512464,5.411693,6.3127356,5.050914,3.787279,2.525457,1.261822,0.0,0.0,0.0,0.0,0.0,0.0,0.52575916,1.0497054,1.5754645,2.0994108,2.6251698,2.3495996,2.0758421,1.8002719,1.5247015,1.2491312,1.7875811,2.324218,2.8626678,3.3993049,3.9377546,4.650249,5.3627434,6.0752378,6.787732,7.500226,6.4632115,5.424384,4.3873696,3.350355,2.3133402,6.48678,10.662033,14.837286,19.012539,23.187792,20.624262,18.062546,15.499017,12.937301,10.375585,9.374829,8.375887,7.3751316,6.3743763,5.375434,5.0744824,4.7753434,4.4743915,4.175253,3.874301,3.5497808,3.2252605,2.9007401,2.5744069,2.2498865,2.1628644,2.0758421,1.987007,1.8999848,1.8129625,1.4866294,1.162109,0.8375887,0.51306844,0.18673515,0.18673515,0.18673515,0.18673515,0.18673515,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,2.5000753,5.0001507,7.500226,10.000301,12.500377,11.14972,9.800876,8.450218,7.0995617,5.750717,8.26167,10.774437,13.287203,15.799969,18.312735,14.91343,11.512312,8.113008,4.7118897,1.3125849,4.0882306,6.8620634,9.637709,12.413355,15.187187,13.762199,12.337211,10.912222,9.487233,8.062244,7.6253204,7.1883965,6.7496595,6.3127356,5.8758116,5.487838,5.0998635,4.7118897,4.325729,3.9377546,3.2506418,2.561716,1.8746033,1.1874905,0.50037766,0.6000906,0.69980353,0.7995165,0.89922947,1.0007553,1.2001812,1.3996071,1.6008459,1.8002719,1.9996977,2.2625773,2.525457,2.7883365,3.049403,3.3122826,3.0747845,2.8372865,2.5997884,2.3622901,2.124792,1.7005589,1.2745126,0.85027945,0.42423326,0.0,0.0,0.0,0.0,0.0,0.0,0.06164073,0.12509441,0.18673515,0.25018883,0.31182957,0.25018883,0.18673515,0.12509441,0.06164073,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.2374981,0.4749962,0.7124943,0.9499924,1.1874905,0.9499924,0.7124943,0.4749962,0.2374981,0.0,0.11240368,0.22480737,0.33721104,0.44961473,0.5620184,0.87566096,1.1874905,1.49932,1.8129625,2.124792,1.7005589,1.2745126,0.85027945,0.42423326,0.0,0.0,0.0,0.0,0.0,0.0,5.2503395,10.500679,15.751019,20.999546,26.249886,21.099258,15.950445,10.799818,5.6491914,0.50037766,0.5620184,0.62547207,0.6871128,0.7505665,0.8122072,0.89922947,0.9880646,1.0750868,1.162109,1.2491312,1.4757515,1.7005589,1.9253663,2.1501737,2.374981,1.8999848,1.4249886,0.9499924,0.4749962,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.5873999,1.1747998,1.7621996,2.3495996,2.9369993,2.7248828,2.5127661,2.3006494,2.08672,1.8746033,2.4384346,3.000453,3.5624714,4.12449,4.688321,3.8507326,3.0131438,2.175555,1.3379664,0.50037766,0.40066472,0.2991388,0.19942589,0.099712946,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.8375887,1.6117238,2.3876717,3.1618068,3.9377546,5.975525,8.013294,10.049252,12.087022,14.124791,15.138238,16.14987,17.163317,18.17495,19.188396,17.487837,15.787278,14.0867195,12.387974,10.687414,10.161655,9.637709,9.11195,8.588004,8.062244,6.9490857,5.8377395,4.7245803,3.6132345,2.5000753,2.3876717,2.275268,2.1628644,2.0504606,1.938057,1.8619126,1.7875811,1.7132497,1.6371052,1.5627737,1.2491312,0.93730164,0.62547207,0.31182957,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.61278135,1.2255627,1.8383441,2.4493124,3.0620937,4.4381323,5.812358,7.1883965,8.562622,9.936848,9.374829,8.812811,8.2507925,7.686961,7.124943,6.3254266,5.52591,4.7245803,3.925064,3.1255474,2.5127661,1.8999848,1.2872034,0.6744221,0.06164073,0.93730164,1.8129625,2.6868105,3.5624714,4.4381323,4.800725,5.163317,5.52591,5.8866897,6.249282,5.375434,4.499773,3.6241121,2.7502642,1.8746033,1.49932,1.1258497,0.7505665,0.37528324,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.97537386,1.9507477,2.9243085,3.8996825,4.8750563,3.9504454,3.0240216,2.0994108,1.1747998,0.25018883,0.5873999,0.9246109,1.261822,1.6008459,1.938057,2.08672,2.2371957,2.3876717,2.5381477,2.6868105,2.175555,1.6624867,1.1494182,0.63816285,0.12509441,0.7868258,1.4503701,2.1121013,2.7756457,3.437377,3.4500678,3.4627585,3.4754493,3.48814,3.5008307,3.7492065,3.9993954,4.249584,4.499773,4.749962,4.936697,5.125245,5.3119802,5.5005283,5.6872635,5.2992897,4.9131284,4.5251546,4.137181,3.7492065,4.8750563,6.000906,7.124943,8.2507925,9.374829,7.462154,6.784106,6.107871,5.429823,4.751775,4.07554,4.137181,4.2006345,4.262275,4.325729,4.3873696,4.6792564,4.972956,5.2648435,5.5567303,5.8504305,5.9519563,6.055295,6.156821,6.26016,6.3616858,7.690587,9.017676,10.344765,11.671853,13.000754,11.530442,10.060129,8.589817,7.119504,5.6510043,5.6927023,5.7344007,5.7779117,5.81961,5.863121,5.2702823,4.6774435,4.0846047,3.491766,2.9007401,2.5816586,2.2643902,1.9471219,1.6298534,1.3125849,1.4177368,1.5228885,1.6280404,1.7331922,1.8383441,1.7150626,1.5917811,1.4703126,1.3470312,1.2255627,1.3542831,1.4848163,1.6153497,1.745883,1.8746033,2.5345216,3.1944401,3.8543584,4.514277,5.1741953,5.669134,6.165886,6.6608243,7.155763,7.650702,6.816739,5.9845896,5.1524396,4.3202896,3.48814,3.1817493,2.8771715,2.572594,2.268016,1.9634385,2.030518,2.0975976,2.1646774,2.231757,2.3006494,2.2607644,2.220879,2.179181,2.1392958,2.0994108,2.0994108,2.0994108,2.0994108,2.0994108,2.0994108,1.7966459,1.4956942,1.1929294,0.8901646,0.5873999,0.46955732,0.35171473,0.23568514,0.11784257,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.2374981,0.41335547,0.5873999,0.76325727,0.93730164,1.79302,2.6469254,3.5026438,4.358362,5.2122674,4.9783955,4.74271,4.507025,4.273153,4.0374675,3.874301,3.7129474,3.5497808,3.388427,3.2252605,3.8108473,4.3946214,4.9802084,5.565795,6.149569,4.942136,3.7347028,2.5272698,1.3198367,0.11240368,0.21211663,0.31182957,0.41335547,0.51306844,0.61278135,1.0569572,1.502946,1.9471219,2.3931105,2.8372865,2.520018,2.2027495,1.8854811,1.5682126,1.2491312,1.6552348,2.0595255,2.465629,2.8699198,3.2742105,3.8199122,4.365614,4.9095025,5.4552045,5.999093,5.864934,5.730775,5.5948024,5.4606433,5.3246713,8.158332,10.990179,13.822026,16.655687,19.487535,17.322857,15.15818,12.99169,10.827013,8.662335,7.8483152,7.0324817,6.2166486,5.4026284,4.5867953,4.3003473,4.0120864,3.7256382,3.437377,3.149116,3.0367124,2.9243085,2.811905,2.6995013,2.5870976,2.4801328,2.373168,2.2643902,2.1574254,2.0504606,1.693307,1.3343405,0.97718686,0.6200332,0.26287958,0.2755703,0.28826106,0.2991388,0.31182957,0.3245203,0.4550536,0.5855869,0.71430725,0.8448406,0.97537386,3.4119956,5.8504305,8.287052,10.725487,13.162108,12.717933,12.271944,11.827768,11.383592,10.937603,13.211059,15.4827,17.756155,20.027798,22.29944,19.5945,16.889559,14.184619,11.479679,8.774739,10.466233,12.155914,13.845595,15.535276,17.224958,15.218008,13.209246,11.202296,9.195346,7.1865835,6.816739,6.446895,6.0770507,5.7072062,5.337362,4.9983377,4.6575007,4.3166637,3.97764,3.636803,2.9932013,2.3477864,1.7023718,1.0569572,0.41335547,0.62184614,0.8321498,1.0424535,1.2527572,1.4630609,1.5917811,1.7223145,1.8528478,1.983381,2.1121013,2.220879,2.327844,2.4348087,2.5417736,2.6505513,2.4601903,2.269829,2.079468,1.889107,1.7005589,1.3597219,1.020698,0.67986095,0.34083697,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.059827764,0.10696479,0.15410182,0.2030518,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.065266654,0.13053331,0.19579996,0.25925365,0.3245203,0.27919623,0.23568514,0.19036107,0.14503701,0.099712946,0.27013144,0.4405499,0.6091554,0.7795739,0.9499924,0.75963134,0.56927025,0.38072214,0.19036107,0.0,0.09064813,0.1794833,0.27013144,0.36077955,0.44961473,0.69980353,0.9499924,1.2001812,1.4503701,1.7005589,1.3597219,1.020698,0.67986095,0.34083697,0.0,0.06164073,0.12509441,0.18673515,0.25018883,0.31182957,4.4526362,8.59163,12.732436,16.87143,21.012236,17.346426,13.682428,10.016619,6.352621,2.6868105,2.5127661,2.3369088,2.1628644,1.987007,1.8129625,1.6570477,1.502946,1.3470312,1.1929294,1.0370146,1.2291887,1.4231756,1.6153497,1.8075237,1.9996977,1.6008459,1.2001812,0.7995165,0.40066472,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.10515183,0.08520924,0.065266654,0.045324065,0.025381476,0.03988518,0.054388877,0.07070554,0.08520924,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0870222,0.17585737,0.26287958,0.34990177,0.43692398,0.41516843,0.3934129,0.36984438,0.3480888,0.3245203,1.0098201,1.69512,2.38042,3.0657198,3.7492065,3.5171473,3.2850883,3.053029,2.819157,2.5870976,2.8245957,3.0620937,3.299592,3.53709,3.774588,3.100166,2.4257438,1.7495089,1.0750868,0.40066472,0.3208944,0.23931105,0.15954071,0.07977036,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.13053331,0.13415924,0.13959812,0.14503701,0.15047589,0.20486477,0.25925365,0.3154555,0.36984438,0.42423326,1.5083848,2.5907235,3.673062,4.7554007,5.8377395,7.0342946,8.232663,9.429218,10.627586,11.8241415,12.750566,13.675177,14.599788,15.524399,16.449009,15.20713,13.965251,12.721559,11.479679,10.2378,9.976733,9.71748,9.458226,9.197159,8.937905,8.113008,7.28811,6.4632115,5.638314,4.8134155,4.461701,4.1117992,3.7618973,3.4119956,3.0620937,2.8681068,2.6723068,2.47832,2.2825198,2.08672,1.7767034,1.4666867,1.1566701,0.8466535,0.53663695,0.47318324,0.40791658,0.34264994,0.27738327,0.21211663,0.2755703,0.33721104,0.40066472,0.46230546,0.52575916,0.7505665,0.97537386,1.2001812,1.4249886,1.649796,1.8347181,2.0196402,2.2045624,2.3894846,2.5744069,2.1102884,1.6443571,1.1802386,0.71430725,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.4894999,0.9808127,1.4703126,1.9598125,2.4493124,3.5932918,4.7354584,5.8776245,7.019791,8.161958,7.9226465,7.6833353,7.4422116,7.2029004,6.9617763,6.24203,5.522284,4.802538,4.082792,3.3630457,2.7031271,2.0432088,1.3832904,0.72337204,0.06164073,0.7795739,1.4975071,2.2154403,2.9315605,3.6494937,3.9703882,4.2894692,4.610364,4.9294453,5.2503395,4.5632267,3.874301,3.1871881,2.5000753,1.8129625,1.452183,1.0932164,0.7324369,0.37165734,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.072518505,0.13234627,0.19217403,0.2520018,0.31182957,0.27194437,0.23205921,0.19217403,0.15228885,0.11240368,0.17223145,0.23205921,0.291887,0.35171473,0.41335547,0.33721104,0.26287958,0.18673515,0.11240368,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.81764615,1.6226015,2.427557,3.2325122,4.0374675,3.3721104,2.7067533,2.0432088,1.3778516,0.7124943,0.91735905,1.1222239,1.3270886,1.5319533,1.7368182,1.9144884,2.0921588,2.269829,2.4474995,2.6251698,2.1628644,1.7005589,1.2382535,0.774135,0.31182957,0.83033687,1.3470312,1.8655385,2.382233,2.9007401,2.9351864,2.9696326,3.004079,3.0403383,3.0747845,3.3829882,3.6893787,3.9975824,4.305786,4.612177,4.7554007,4.896812,5.040036,5.18326,5.3246713,4.9294453,4.5342193,4.1408067,3.7455807,3.350355,4.2767787,5.2050157,6.1332526,7.059676,7.987913,6.8004227,6.1948934,5.5893636,4.985647,4.3801174,3.774588,3.8380418,3.8996825,3.9631362,4.024777,4.0882306,4.4345064,4.782595,5.130684,5.47696,5.825049,5.91751,6.009971,6.1024323,6.1948934,6.2873545,7.230095,8.172835,9.115576,10.058316,10.999244,10.310318,9.619579,8.930654,8.239915,7.549176,7.2355337,6.9200783,6.604623,6.2891674,5.975525,5.3645563,4.7554007,4.1444325,3.5352771,2.9243085,2.8028402,2.6795588,2.5580902,2.4348087,2.3133402,2.4474995,2.5816586,2.7176309,2.8517902,2.9877625,2.7303216,2.472881,2.2154403,1.9579996,1.7005589,1.6733645,1.6443571,1.6171626,1.5899682,1.5627737,2.3695421,3.1781235,3.9848917,4.7916603,5.600241,6.1278133,6.6553855,7.1829576,7.71053,8.238102,7.5473633,6.8566246,6.167699,5.47696,4.788034,4.539658,4.2930956,4.0447197,3.7981565,3.5497808,3.5352771,3.5207734,3.5044568,3.489953,3.4754493,3.3449159,3.2143826,3.0856624,2.955129,2.8245957,2.762955,2.6995013,2.6378605,2.5744069,2.5127661,2.1193533,1.7277533,1.3343405,0.94274056,0.5493277,0.4405499,0.32995918,0.21936847,0.11059072,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.33721104,0.5493277,0.76325727,0.97537386,1.1874905,2.6469254,4.1081734,5.567608,7.027043,8.488291,7.991539,7.4966,7.0016613,6.506723,6.011784,5.7380266,5.462456,5.186886,4.9131284,4.6375585,4.9076896,5.177821,5.4479527,5.718084,5.9882154,4.835171,3.682127,2.5290828,1.3778516,0.22480737,0.42423326,0.62547207,0.824898,1.0243238,1.2255627,1.5899682,1.9543737,2.3205922,2.6849976,3.049403,2.6904364,2.3296568,1.9706904,1.6099107,1.2491312,1.5228885,1.794833,2.0667772,2.3405347,2.612479,2.9895754,3.3666716,3.7455807,4.122677,4.499773,5.2666564,6.035352,6.8022356,7.569119,8.337815,9.82807,11.318325,12.806767,14.297023,15.787278,14.01964,12.252001,10.484363,8.716724,6.9508986,6.319988,5.6908894,5.0599785,4.4308805,3.7999697,3.5243993,3.2506418,2.9750717,2.6995013,2.4257438,2.525457,2.6251698,2.7248828,2.8245957,2.9243085,2.7974012,2.6704938,2.5417736,2.4148662,2.2879589,1.8981718,1.5083848,1.1167849,0.726998,0.33721104,0.36259252,0.387974,0.41335547,0.43692398,0.46230546,0.75963134,1.0569572,1.3542831,1.651609,1.9507477,4.325729,6.70071,9.07569,11.450671,13.825653,14.284332,14.744824,15.2053175,15.663997,16.124489,18.15682,20.189152,22.223295,24.255627,26.287958,24.277382,22.266806,20.258043,18.247469,16.236893,16.842422,17.447952,18.051668,18.657198,19.262728,16.672005,14.083094,11.49237,8.901647,6.3127356,6.009971,5.7072062,5.4044414,5.101677,4.800725,4.507025,4.215138,3.923251,3.6295512,3.3376641,2.7357605,2.132044,1.5301404,0.92823684,0.3245203,0.64541465,0.9644961,1.2853905,1.6044719,1.9253663,1.9851941,2.0450218,2.1048496,2.1646774,2.2245052,2.1773682,2.1302311,2.0830941,2.034144,1.987007,1.845596,1.7023718,1.5591478,1.4177368,1.2745126,1.020698,0.7650702,0.5094425,0.25562772,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.058014803,0.09064813,0.12328146,0.15410182,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13053331,0.25925365,0.38978696,0.52032024,0.6508536,0.56020546,0.46955732,0.38072214,0.29007402,0.19942589,0.30276474,0.40429065,0.5076295,0.6091554,0.7124943,0.56927025,0.42785916,0.28463513,0.14322405,0.0,0.06707962,0.13415924,0.2030518,0.27013144,0.33721104,0.52575916,0.7124943,0.89922947,1.0877775,1.2745126,1.020698,0.7650702,0.5094425,0.25562772,0.0,0.12509441,0.25018883,0.37528324,0.50037766,0.62547207,3.6549325,6.684393,9.715667,12.745127,15.774588,13.595407,11.4144125,9.235231,7.0542374,4.8750563,4.461701,4.0501585,3.636803,3.2252605,2.811905,2.4148662,2.0178273,1.6207886,1.2219368,0.824898,0.98443866,1.1457924,1.305333,1.4648738,1.6244144,1.2998942,0.97537386,0.6508536,0.3245203,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,0.21030366,0.17041849,0.13053331,0.09064813,0.05076295,0.054388877,0.059827764,0.065266654,0.07070554,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.17585737,0.34990177,0.52575916,0.69980353,0.87566096,0.83033687,0.7850128,0.73968875,0.69436467,0.6508536,1.4322405,2.2154403,2.9968271,3.780027,4.5632267,4.309412,4.0574102,3.8054085,3.5515938,3.299592,3.2125697,3.1255474,3.0367124,2.94969,2.8626678,2.3495996,1.8383441,1.3252757,0.8122072,0.2991388,0.23931105,0.1794833,0.11965553,0.059827764,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.21030366,0.23205921,0.25562772,0.27738327,0.2991388,0.39703882,0.4949388,0.59283876,0.69073874,0.7868258,2.1773682,3.5679104,4.95664,6.347182,7.7377243,8.094878,8.452031,8.809185,9.168152,9.525306,10.362894,11.200482,12.038072,12.87566,13.713249,12.928236,12.143224,11.358211,10.573197,9.788185,9.791811,9.79725,9.802689,9.808127,9.811753,9.275117,8.736667,8.200029,7.66158,7.124943,6.5375433,5.9501433,5.3627434,4.7753434,4.1879435,3.872488,3.5570326,3.2415771,2.9279346,2.612479,2.3042755,1.9978848,1.6896812,1.3832904,1.0750868,0.9445535,0.81583315,0.6852999,0.55476654,0.42423326,0.5493277,0.6744221,0.7995165,0.9246109,1.0497054,1.49932,1.9507477,2.4003625,2.8499773,3.299592,3.6694362,4.0392804,4.409125,4.780782,5.1506267,4.220577,3.290527,2.3604772,1.4304274,0.50037766,0.40066472,0.2991388,0.19942589,0.099712946,0.0,0.3680314,0.73424983,1.1022812,1.4703126,1.8383441,2.7484512,3.6567454,4.5668526,5.47696,6.3870673,6.4704633,6.552047,6.635443,6.717026,6.8004227,6.1604466,5.520471,4.880495,4.2405195,3.6005437,2.8916752,2.18462,1.4775645,0.7705091,0.06164073,0.62184614,1.1820517,1.742257,2.3024626,2.8626678,3.1400511,3.4174345,3.6948178,3.972201,4.249584,3.7492065,3.2506418,2.7502642,2.2498865,1.7495089,1.405046,1.0605831,0.71430725,0.36984438,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.14503701,0.26469254,0.38434806,0.5058166,0.62547207,0.52032024,0.41516843,0.3100166,0.20486477,0.099712946,0.23205921,0.36440548,0.49675176,0.629098,0.76325727,0.62547207,0.48768693,0.34990177,0.21211663,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.65991837,1.2944553,1.9308052,2.565342,3.199879,2.7955883,2.3894846,1.9851941,1.5809034,1.1747998,1.2473183,1.3198367,1.3923552,1.4648738,1.5373923,1.742257,1.9471219,2.1519866,2.3568513,2.561716,2.1501737,1.7368182,1.3252757,0.9119202,0.50037766,0.872035,1.2455053,1.6171626,1.9906329,2.3622901,2.420305,2.47832,2.5345216,2.5925364,2.6505513,3.0149567,3.3793623,3.7455807,4.1099863,4.4743915,4.572292,4.670192,4.7680917,4.8641787,4.9620786,4.559601,4.157123,3.7546456,3.3521678,2.94969,3.680314,4.410938,5.139749,5.870373,6.599184,6.1368785,5.6056805,5.0726695,4.539658,4.006647,3.4754493,3.53709,3.6005437,3.6621845,3.7256382,3.787279,4.1897564,4.592234,4.994712,5.3971896,5.7996674,5.883064,5.964647,6.0480433,6.1296263,6.2130227,6.7696023,7.327995,7.8845744,8.442966,8.999546,9.090195,9.180842,9.269678,9.360326,9.449161,8.778365,8.105756,7.4331465,6.7605376,6.0879283,5.4606433,4.8333583,4.2042603,3.576975,2.94969,3.0222087,3.094727,3.1672456,3.2397642,3.3122826,3.4772623,3.6422417,3.8072214,3.972201,4.137181,3.7455807,3.3521678,2.960568,2.5671551,2.175555,1.9906329,1.8057107,1.6207886,1.4358664,1.2491312,2.2045624,3.159994,4.115425,5.0708566,6.0244746,6.58468,7.1448855,7.705091,8.265296,8.825501,8.2779875,7.7304726,7.1829576,6.635443,6.0879283,5.8975673,5.7072062,5.516845,5.328297,5.137936,5.040036,4.942136,4.844236,4.748149,4.650249,4.4308805,4.209699,3.9903307,3.7691493,3.5497808,3.4246864,3.299592,3.1744974,3.049403,2.9243085,2.4420607,1.9598125,1.4775645,0.99531645,0.51306844,0.40972954,0.30820364,0.20486477,0.10333887,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.43692398,0.6871128,0.93730164,1.1874905,1.4376793,3.5026438,5.567608,7.6325727,9.697536,11.762501,11.008308,10.252303,9.498111,8.7421055,7.987913,7.5999393,7.211965,6.825804,6.43783,6.049856,6.004532,5.959208,5.915697,5.870373,5.825049,4.7282066,3.6295512,2.5327086,1.4358664,0.33721104,0.63816285,0.93730164,1.2382535,1.5373923,1.8383441,2.1229792,2.4076142,2.6922495,2.9768846,3.2633326,2.8608549,2.4583774,2.0540867,1.651609,1.2491312,1.3905423,1.5301404,1.6697385,1.8093367,1.9507477,2.1592383,2.3695421,2.5798457,2.7901495,3.000453,4.670192,6.33993,8.009668,9.679407,11.350959,11.497808,11.644659,11.793322,11.940171,12.087022,10.718235,9.347635,7.9770355,6.6082487,5.237649,4.7916603,4.347484,3.9033084,3.4573197,3.0131438,2.7502642,2.4873846,2.2245052,1.9616255,1.7005589,2.0123885,2.324218,2.6378605,2.94969,3.2633326,3.1146698,2.9678197,2.819157,2.6723068,2.525457,2.1030366,1.6806163,1.258196,0.83577573,0.41335547,0.44961473,0.48768693,0.52575916,0.5620184,0.6000906,1.064209,1.5301404,1.9942589,2.4601903,2.9243085,5.237649,7.549176,9.862516,12.175857,14.487384,15.852545,17.217705,18.582867,19.948027,21.313189,23.104395,24.897415,26.690435,28.483456,30.274662,28.960264,27.645866,26.329655,25.015257,23.70086,23.220425,22.73999,22.259554,21.780933,21.300497,18.127813,14.955129,11.782444,8.609759,5.4370747,5.2032027,4.9675174,4.7318325,4.49796,4.262275,4.017525,3.7727752,3.5280252,3.2832751,3.0367124,2.47832,1.9181144,1.357909,0.79770356,0.2374981,0.6671702,1.0968424,1.5283275,1.9579996,2.3876717,2.3767939,2.3677292,2.3568513,2.3477864,2.3369088,2.13567,1.9326181,1.7295663,1.5283275,1.3252757,1.2291887,1.1349145,1.0406405,0.9445535,0.85027945,0.67986095,0.5094425,0.34083697,0.17041849,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.054388877,0.072518505,0.09064813,0.10696479,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.19579996,0.38978696,0.5855869,0.7795739,0.97537386,0.83940166,0.70524246,0.56927025,0.43511102,0.2991388,0.33539808,0.36984438,0.40429065,0.4405499,0.4749962,0.38072214,0.28463513,0.19036107,0.09427405,0.0,0.045324065,0.09064813,0.13415924,0.1794833,0.22480737,0.34990177,0.4749962,0.6000906,0.72518504,0.85027945,0.67986095,0.5094425,0.34083697,0.17041849,0.0,0.18673515,0.37528324,0.5620184,0.7505665,0.93730164,2.857229,4.7771564,6.697084,8.617011,10.536939,9.842574,9.14821,8.452031,7.757667,7.063302,6.412449,5.763408,5.1125546,4.461701,3.8126602,3.1726844,2.5327086,1.892733,1.2527572,0.61278135,0.73968875,0.8665961,0.99531645,1.1222239,1.2491312,1.0007553,0.7505665,0.50037766,0.25018883,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.07433146,0.15047589,0.22480737,0.2991388,0.37528324,0.3154555,0.25562772,0.19579996,0.13415924,0.07433146,0.07070554,0.065266654,0.059827764,0.054388877,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.26287958,0.52575916,0.7868258,1.0497054,1.3125849,1.2455053,1.1766127,1.1095331,1.0424535,0.97537386,1.8546607,2.7357605,3.6150475,4.494334,5.375434,5.101677,4.8297324,4.557788,4.2858434,4.0120864,3.6005437,3.1871881,2.7756457,2.3622901,1.9507477,1.6008459,1.2491312,0.89922947,0.5493277,0.19942589,0.15954071,0.11965553,0.07977036,0.03988518,0.0,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,0.29007402,0.32995918,0.36984438,0.40972954,0.44961473,0.58921283,0.7306239,0.87022203,1.0098201,1.1494182,2.8481643,4.5450974,6.24203,7.9407763,9.637709,9.155461,8.673213,8.189152,7.706904,7.224656,7.9752226,8.725789,9.474543,10.225109,10.975676,10.64753,10.319383,9.99305,9.664904,9.336758,9.606889,9.87702,10.147152,10.417283,10.687414,10.437225,10.1870365,9.936848,9.686659,9.438283,8.613385,7.7884874,6.9617763,6.1368785,5.3119802,4.876869,4.441758,4.006647,3.5733492,3.1382382,2.8318477,2.5272698,2.222692,1.9181144,1.6117238,1.4177368,1.2219368,1.0279498,0.8321498,0.63816285,0.824898,1.0116332,1.2001812,1.3869164,1.5754645,2.2498865,2.9243085,3.6005437,4.274966,4.949388,5.505967,6.060734,6.6155005,7.170267,7.7250338,6.3308654,4.934884,3.540716,2.1447346,0.7505665,0.6000906,0.44961473,0.2991388,0.15047589,0.0,0.24474995,0.4894999,0.73424983,0.9808127,1.2255627,1.9017978,2.5798457,3.2578938,3.9341288,4.612177,5.0182805,5.422571,5.826862,6.2329655,6.637256,6.0770507,5.516845,4.95664,4.3982472,3.8380418,3.0820365,2.327844,1.5718386,0.81764615,0.06164073,0.46411842,0.8665961,1.2708868,1.6715515,2.0758421,2.3097143,2.5453994,2.7792716,3.0149567,3.2506418,2.9369993,2.6251698,2.3133402,1.9996977,1.6878681,1.357909,1.0279498,0.6979906,0.3680314,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.21755551,0.39703882,0.57833505,0.75781834,0.93730164,0.7668832,0.5982776,0.42785916,0.2574407,0.0870222,0.291887,0.49675176,0.7016165,0.90829426,1.1131591,0.9119202,0.7124943,0.51306844,0.31182957,0.11240368,0.09064813,0.06707962,0.045324065,0.02175555,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.50219065,0.968122,1.4322405,1.8981718,2.3622901,2.2172532,2.0722163,1.9271792,1.7821422,1.6371052,1.5772774,1.5174497,1.4576219,1.3977941,1.3379664,1.5700256,1.8020848,2.034144,2.268016,2.5000753,2.137483,1.7748904,1.4122978,1.0497054,0.6871128,0.9155461,1.1421664,1.3705997,1.5972201,1.8256533,1.9054236,1.9851941,2.0649643,2.1447346,2.2245052,2.6469254,3.0693457,3.491766,3.9141862,4.3366065,4.3891826,4.441758,4.494334,4.5469103,4.599486,4.1897564,3.780027,3.3702974,2.960568,2.5508385,3.0820365,3.6150475,4.1480584,4.6792564,5.2122674,5.475147,5.0146546,4.554162,4.0954823,3.63499,3.1744974,3.2379513,3.299592,3.3630457,3.4246864,3.48814,3.9450066,4.401873,4.860553,5.317419,5.774286,5.846804,5.919323,5.9918413,6.0643597,6.1368785,6.3091097,6.4831543,6.6553855,6.827617,6.9998484,7.8700705,8.740293,9.610515,10.480737,11.349146,10.319383,9.28962,8.259857,7.230095,6.200332,5.5549173,4.9095025,4.264088,3.6204863,2.9750717,3.24339,3.5098956,3.778214,4.0447197,4.313038,4.507025,4.702825,4.896812,5.092612,5.2884116,4.76084,4.233268,3.7056956,3.1781235,2.6505513,2.3079014,1.9652514,1.6226015,1.2799516,0.93730164,2.039583,3.141864,4.2441454,5.3482394,6.450521,7.0433598,7.6343856,8.227224,8.820063,9.412902,9.006798,8.602508,8.198216,7.7921133,7.3878226,7.2554765,7.12313,6.9907837,6.8566246,6.7242785,6.544795,6.3653116,6.185828,6.004532,5.825049,5.5150323,5.2050157,4.894999,4.5849824,4.274966,4.0882306,3.8996825,3.7129474,3.5243993,3.3376641,2.764768,2.1918716,1.6207886,1.0478923,0.4749962,0.38072214,0.28463513,0.19036107,0.09427405,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,0.53663695,0.824898,1.1131591,1.3996071,1.6878681,4.358362,7.027043,9.697536,12.368031,15.036712,14.023266,13.008006,11.992747,10.9774885,9.96223,9.461852,8.963287,8.46291,7.9625316,7.462154,7.1031876,6.742408,6.3816285,6.0226617,5.661882,4.6194286,3.576975,2.5345216,1.4920682,0.44961473,0.85027945,1.2491312,1.649796,2.0504606,2.4493124,2.6541772,2.8608549,3.0657198,3.2705846,3.4754493,3.0294604,2.5852847,2.1392958,1.69512,1.2491312,1.258196,1.2654479,1.2726997,1.2799516,1.2872034,1.3307146,1.3724127,1.4141108,1.4576219,1.49932,4.071914,6.644508,9.217102,11.789696,14.362289,13.167547,11.972805,10.778063,9.583321,8.386765,7.415017,6.4432693,5.469708,4.49796,3.5243993,3.2651455,3.005892,2.7448254,2.4855716,2.2245052,1.9743162,1.7241274,1.4757515,1.2255627,0.97537386,1.49932,2.0250793,2.5508385,3.0747845,3.6005437,3.4319382,3.2651455,3.0983531,2.9297476,2.762955,2.3079014,1.8528478,1.3977941,0.94274056,0.48768693,0.53663695,0.5873999,0.63816285,0.6871128,0.73787576,1.3705997,2.0033236,2.6342347,3.2669585,3.8996825,6.149569,8.399456,10.649343,12.899229,15.149116,17.420757,19.690586,21.960415,24.230246,26.500074,28.05197,29.605679,31.157576,32.709473,34.26318,33.643147,33.023113,32.40308,31.783047,31.163013,29.598427,28.032028,26.467442,24.902855,23.338266,19.581808,15.827164,12.072517,8.317872,4.5632267,4.3946214,4.227829,4.059223,3.8924308,3.7256382,3.5280252,3.3304121,3.1327994,2.9351864,2.7375734,2.220879,1.7023718,1.1856775,0.6671702,0.15047589,0.69073874,1.2291887,1.7694515,2.3097143,2.8499773,2.770207,2.6904364,2.610666,2.5308957,2.4493124,2.0921588,1.7350051,1.3778516,1.020698,0.66173136,0.61459434,0.56745726,0.52032024,0.47318324,0.42423326,0.34083697,0.25562772,0.17041849,0.08520924,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.052575916,0.054388877,0.058014803,0.059827764,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.25925365,0.52032024,0.7795739,1.0406405,1.2998942,1.1204109,0.93911463,0.75963134,0.58014804,0.40066472,0.3680314,0.33539808,0.30276474,0.27013144,0.2374981,0.19036107,0.14322405,0.09427405,0.047137026,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.17585737,0.2374981,0.2991388,0.36259252,0.42423326,0.34083697,0.25562772,0.17041849,0.08520924,0.0,0.25018883,0.50037766,0.7505665,1.0007553,1.2491312,2.0595255,2.8699198,3.680314,4.4907084,5.2992897,6.089741,6.880193,7.6706448,8.459284,9.249735,8.363196,7.474845,6.588306,5.6999545,4.8134155,3.930503,3.04759,2.1646774,1.2817645,0.40066472,0.4949388,0.58921283,0.6852999,0.7795739,0.87566096,0.69980353,0.52575916,0.34990177,0.17585737,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.099712946,0.19942589,0.2991388,0.40066472,0.50037766,0.42060733,0.34083697,0.25925365,0.1794833,0.099712946,0.08520924,0.07070554,0.054388877,0.03988518,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.34990177,0.69980353,1.0497054,1.3996071,1.7495089,1.6606737,1.5700256,1.4793775,1.3905423,1.2998942,2.277081,3.254268,4.233268,5.2104545,6.187641,5.8957543,5.6020546,5.3101673,5.0182805,4.7245803,3.9867048,3.2506418,2.5127661,1.7748904,1.0370146,0.85027945,0.66173136,0.4749962,0.28826106,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.06164073,0.12509441,0.18673515,0.25018883,0.31182957,0.36984438,0.42785916,0.48587397,0.5420758,0.6000906,0.78319985,0.9644961,1.1476053,1.3307146,1.5120108,3.5171473,5.522284,7.5274205,9.5325575,11.537694,10.2142315,8.892582,7.569119,6.247469,4.9258194,5.5875506,6.249282,6.9128265,7.574558,8.238102,8.366822,8.497355,8.627889,8.756609,8.887142,9.421967,9.956791,10.493427,11.028252,11.563075,11.599335,11.637406,11.675479,11.711739,11.74981,10.687414,9.625018,8.562622,7.500226,6.43783,5.883064,5.328297,4.7717175,4.216951,3.6621845,3.3594196,3.056655,2.7557032,2.4529383,2.1501737,1.889107,1.6298534,1.3705997,1.1095331,0.85027945,1.1004683,1.3506571,1.6008459,1.8492218,2.0994108,3.000453,3.8996825,4.800725,5.6999545,6.599184,7.3406854,8.080374,8.820063,9.5597515,10.29944,8.439341,6.5792413,4.7191415,2.8608549,1.0007553,0.7995165,0.6000906,0.40066472,0.19942589,0.0,0.12328146,0.24474995,0.3680314,0.4894999,0.61278135,1.0569572,1.502946,1.9471219,2.3931105,2.8372865,3.5642843,4.2930956,5.0200934,5.7470913,6.4759026,5.995467,5.5150323,5.034597,4.554162,4.07554,3.2723975,2.469255,1.6679256,0.86478317,0.06164073,0.30820364,0.5529536,0.79770356,1.0424535,1.2872034,1.4793775,1.6733645,1.8655385,2.0577126,2.2498865,2.124792,1.9996977,1.8746033,1.7495089,1.6244144,1.310772,0.99531645,0.67986095,0.36440548,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.29007402,0.5293851,0.7705091,1.0098201,1.2491312,1.015259,0.7795739,0.54570174,0.3100166,0.07433146,0.35171473,0.629098,0.90829426,1.1856775,1.4630609,1.2001812,0.93730164,0.6744221,0.41335547,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.3444629,0.6399758,0.9354887,1.2291887,1.5247015,1.6407311,1.7549478,1.8691645,1.9851941,2.0994108,1.9072367,1.7150626,1.5228885,1.3307146,1.1367276,1.3977941,1.6570477,1.9181144,2.1773682,2.4366217,2.124792,1.8129625,1.49932,1.1874905,0.87566096,0.9572442,1.0406405,1.1222239,1.2056202,1.2872034,1.3905423,1.4920682,1.5954071,1.696933,1.8002719,2.280707,2.759329,3.2397642,3.720199,4.2006345,4.207886,4.215138,4.2223897,4.229642,4.2368937,3.8199122,3.4029307,2.9841363,2.5671551,2.1501737,2.4855716,2.819157,3.1545548,3.489953,3.825351,4.8116026,4.4254417,4.0374675,3.6494937,3.2633326,2.8753586,2.9369993,3.000453,3.0620937,3.1255474,3.1871881,3.7002566,4.213325,4.7245803,5.237649,5.750717,5.812358,5.8758116,5.9374523,6.000906,6.0625467,5.8504305,5.638314,5.424384,5.2122674,5.0001507,6.6499467,8.299743,9.949538,11.599335,13.24913,11.862214,10.475298,9.086569,7.699652,6.3127356,5.6491914,4.98746,4.325729,3.6621845,3.000453,3.4627585,3.925064,4.3873696,4.8496747,5.3119802,5.5367875,5.7615952,5.9882154,6.2130227,6.43783,5.774286,5.1125546,4.4508233,3.787279,3.1255474,2.6251698,2.124792,1.6244144,1.1258497,0.62547207,1.8746033,3.1255474,4.3746786,5.6256227,6.874754,7.500226,8.125698,8.749357,9.374829,10.000301,9.737422,9.474543,9.211663,8.950596,8.6877165,8.613385,8.537241,8.46291,8.386765,8.312433,8.049554,7.7866745,7.5256076,7.262728,6.9998484,6.599184,6.200332,5.7996674,5.4008155,5.0001507,4.749962,4.499773,4.249584,3.9993954,3.7492065,3.0874753,2.4257438,1.7621996,1.1004683,0.43692398,0.34990177,0.26287958,0.17585737,0.0870222,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06164073,0.12509441,0.18673515,0.25018883,0.31182957,0.63816285,0.96268314,1.2872034,1.6117238,1.938057,5.2122674,8.488291,11.762501,15.036712,18.312735,17.038223,15.761897,14.487384,13.212872,11.938358,11.325577,10.712796,10.100015,9.487233,8.874452,8.200029,7.5256076,6.849373,6.1749506,5.5005283,4.512464,3.5243993,2.5381477,1.550083,0.5620184,1.062396,1.5627737,2.0631514,2.561716,3.0620937,3.1871881,3.3122826,3.437377,3.5624714,3.6875658,3.199879,2.712192,2.2245052,1.7368182,1.2491312,1.1258497,1.0007553,0.87566096,0.7505665,0.62547207,0.50037766,0.37528324,0.25018883,0.12509441,0.0,3.4754493,6.9490857,10.424535,13.899984,17.375433,14.837286,12.300951,9.762803,7.224656,4.688321,4.1117992,3.53709,2.962381,2.3876717,1.8129625,1.7368182,1.6624867,1.5881553,1.5120108,1.4376793,1.2001812,0.96268314,0.72518504,0.48768693,0.25018883,0.9880646,1.7241274,2.4620032,3.199879,3.9377546,3.7492065,3.5624714,3.3757362,3.1871881,3.000453,2.5127661,2.0250793,1.5373923,1.0497054,0.5620184,0.62547207,0.6871128,0.7505665,0.8122072,0.87566096,1.6751775,2.474694,3.2742105,4.07554,4.8750563,7.063302,9.249735,11.437981,13.6244135,15.812659,18.987158,22.161655,25.337965,28.512463,31.68696,32.999546,34.31213,35.624714,36.937298,38.249886,38.324215,38.40036,38.474693,38.550835,38.625168,35.974617,33.32588,30.675327,28.024776,25.374224,21.037619,16.701012,12.362592,8.024173,3.6875658,3.587853,3.48814,3.386614,3.2869012,3.1871881,3.0367124,2.8880494,2.7375734,2.5870976,2.4366217,1.9616255,1.4866294,1.0116332,0.53663695,0.06164073,0.7124943,1.3633479,2.0123885,2.663242,3.3122826,3.1618068,3.0131438,2.8626678,2.712192,2.561716,2.0504606,1.5373923,1.0243238,0.51306844,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.3245203,0.6508536,0.97537386,1.2998942,1.6244144,1.3996071,1.1747998,0.9499924,0.72518504,0.50037766,0.40066472,0.2991388,0.19942589,0.099712946,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.31182957,0.62547207,0.93730164,1.2491312,1.5627737,1.261822,0.96268314,0.66173136,0.36259252,0.06164073,2.3369088,4.612177,6.887445,9.162713,11.437981,10.312131,9.188094,8.062244,6.9382076,5.812358,4.688321,3.5624714,2.4366217,1.3125849,0.18673515,0.25018883,0.31182957,0.37528324,0.43692398,0.50037766,0.40066472,0.2991388,0.19942589,0.099712946,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.12509441,0.25018883,0.37528324,0.50037766,0.62547207,0.52575916,0.42423326,0.3245203,0.22480737,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.43692398,0.87566096,1.3125849,1.7495089,2.1882458,2.0758421,1.9616255,1.8492218,1.7368182,1.6244144,2.6995013,3.774588,4.8496747,5.924762,6.9998484,6.688019,6.3743763,6.0625467,5.750717,5.4370747,4.3746786,3.3122826,2.2498865,1.1874905,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.07433146,0.15047589,0.22480737,0.2991388,0.37528324,0.44961473,0.52575916,0.6000906,0.6744221,0.7505665,0.97537386,1.2001812,1.4249886,1.649796,1.8746033,4.1879435,6.4994707,8.812811,11.124338,13.437678,11.274815,9.11195,6.9490857,4.788034,2.6251698,3.199879,3.774588,4.349297,4.9258194,5.5005283,6.0879283,6.6753283,7.262728,7.850128,8.437528,9.237044,10.038374,10.837891,11.637406,12.436923,12.763257,13.087777,13.412297,13.736817,14.06315,12.763257,11.463363,10.161655,8.861761,7.5618668,6.887445,6.2130227,5.5367875,4.8623657,4.1879435,3.8869917,3.587853,3.2869012,2.9877625,2.6868105,2.3622901,2.03777,1.7132497,1.3869164,1.062396,1.3742256,1.6878681,1.9996977,2.3133402,2.6251698,3.7492065,4.8750563,6.000906,7.124943,8.2507925,9.175404,10.100015,11.024626,11.949236,12.87566,10.549629,8.225411,5.89938,3.5751622,1.2491312,1.0007553,0.7505665,0.50037766,0.25018883,0.0,0.0,0.0,0.0,0.0,0.0,0.21211663,0.42423326,0.63816285,0.85027945,1.062396,2.1121013,3.1618068,4.213325,5.2630305,6.3127356,5.9120708,5.5132194,5.1125546,4.7118897,4.313038,3.4627585,2.612479,1.7621996,0.9119202,0.06164073,0.15047589,0.2374981,0.3245203,0.41335547,0.50037766,0.6508536,0.7995165,0.9499924,1.1004683,1.2491312,1.3125849,1.3742256,1.4376793,1.49932,1.5627737,1.261822,0.96268314,0.66173136,0.36259252,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.36259252,0.66173136,0.96268314,1.261822,1.5627737,1.261822,0.96268314,0.66173136,0.36259252,0.06164073,0.41335547,0.76325727,1.1131591,1.4630609,1.8129625,1.4866294,1.162109,0.8375887,0.51306844,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.18673515,0.31182957,0.43692398,0.5620184,0.6871128,1.062396,1.4376793,1.8129625,2.1882458,2.561716,2.2371957,1.9126755,1.5881553,1.261822,0.93730164,1.2255627,1.5120108,1.8002719,2.08672,2.374981,2.1121013,1.8492218,1.5881553,1.3252757,1.062396,1.0007553,0.93730164,0.87566096,0.8122072,0.7505665,0.87566096,1.0007553,1.1258497,1.2491312,1.3742256,1.9126755,2.4493124,2.9877625,3.5243993,4.062849,4.024777,3.9867048,3.9504454,3.9123733,3.874301,3.4500678,3.0258346,2.5997884,2.175555,1.7495089,1.887294,2.0250793,2.1628644,2.3006494,2.4366217,4.4508233,4.157123,3.8652363,3.5733492,3.2796493,2.9877625,3.009518,3.0330863,3.054842,3.0765975,3.100166,3.5806012,4.059223,4.539658,5.0200934,5.5005283,5.667321,5.8341136,6.002719,6.169512,6.338117,6.3254266,6.3127356,6.300045,6.2873545,6.2746634,7.6398244,9.004985,10.370146,11.735307,13.100468,11.952863,10.805257,9.657652,8.510046,7.362441,6.9055743,6.446895,5.9900284,5.5331616,5.0744824,5.3083544,5.540414,5.772473,6.004532,6.2384043,6.3743763,6.5121617,6.6499467,6.787732,6.925517,6.4051967,5.8848767,5.3645563,4.844236,4.325729,3.9830787,3.6404288,3.2977788,2.955129,2.612479,3.4228733,4.233268,5.041849,5.8522434,6.6626377,7.135821,7.607191,8.080374,8.551744,9.024928,9.11195,9.200785,9.287807,9.374829,9.461852,9.262425,9.063,8.861761,8.662335,8.46291,8.212721,7.9625316,7.7123427,7.462154,7.211965,6.9128265,6.6118746,6.3127356,6.011784,5.712645,5.3119802,4.9131284,4.512464,4.1117992,3.7129474,3.1908143,2.666868,2.1447346,1.6226015,1.1004683,0.9445535,0.7904517,0.6345369,0.48043507,0.3245203,0.28282216,0.23931105,0.19761293,0.15591478,0.11240368,0.11059072,0.10696479,0.10515183,0.10333887,0.099712946,0.11965553,0.13959812,0.15954071,0.1794833,0.19942589,0.23568514,0.27013144,0.3045777,0.34083697,0.37528324,0.61278135,0.85027945,1.0877775,1.3252757,1.5627737,4.4526362,7.3424983,10.232361,13.122223,16.012085,14.951503,13.892733,12.8321495,11.771566,10.712796,10.419096,10.127209,9.835322,9.541622,9.249735,8.404895,7.560054,6.7152133,5.870373,5.0255322,4.2767787,3.529838,2.7828975,2.034144,1.2872034,1.8020848,2.3169663,2.8318477,3.346729,3.8634233,3.8978696,3.9323158,3.966762,4.0030212,4.0374675,3.6041696,3.1726844,2.7393866,2.3079014,1.8746033,1.6008459,1.3252757,1.0497054,0.774135,0.50037766,0.8448406,1.1893034,1.5355793,1.8800422,2.2245052,4.7898474,7.3551893,9.920531,12.48406,15.049402,12.908294,10.765372,8.62245,6.4795284,4.3366065,3.7890918,3.24339,2.6940625,2.1483607,1.6008459,1.9308052,2.2607644,2.5907235,2.9206827,3.2506418,2.6396735,2.030518,1.4195497,0.8103943,0.19942589,0.7904517,1.3796645,1.9706904,2.5599031,3.149116,3.0675328,2.9841363,2.902553,2.819157,2.7375734,2.3967366,2.0577126,1.7168756,1.3778516,1.0370146,1.5228885,2.0069497,2.4928236,2.9768846,3.4627585,3.8996825,4.3384194,4.7753434,5.2122674,5.6491914,7.0524244,8.455658,9.857078,11.26031,12.661731,15.199879,17.738026,20.27436,22.812508,25.348843,26.452936,27.555218,28.6575,29.75978,30.862062,30.901947,30.941832,30.981718,31.021603,31.061487,29.065416,27.067532,25.069647,23.071762,21.073877,17.487837,13.899984,10.312131,6.7242785,3.1382382,3.0330863,2.9279346,2.8227828,2.7176309,2.612479,2.4819458,2.3532255,2.222692,2.0921588,1.9616255,1.5790904,1.1983683,0.81583315,0.43329805,0.05076295,0.56927025,1.0895905,1.6099107,2.1302311,2.6505513,2.5290828,2.4094272,2.2897718,2.1701162,2.0504606,1.6407311,1.2291887,0.8194591,0.40972954,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.047137026,0.07070554,0.092461094,0.11421664,0.13778515,0.19942589,0.26287958,0.3245203,0.387974,0.44961473,0.3825351,0.3154555,0.24837588,0.1794833,0.11240368,0.37528324,0.63816285,0.89922947,1.162109,1.4249886,1.2201238,1.015259,0.8103943,0.6055295,0.40066472,0.3208944,0.23931105,0.15954071,0.07977036,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.33177215,0.61459434,0.8974165,1.1802386,1.4630609,1.1929294,0.922798,0.6526665,0.3825351,0.11240368,1.9344311,3.7582715,5.580299,7.402326,9.224354,8.486478,7.750415,7.0125394,6.2746634,5.5367875,4.459888,3.3829882,2.3042755,1.2273756,0.15047589,0.19942589,0.25018883,0.2991388,0.34990177,0.40066472,0.33721104,0.2755703,0.21211663,0.15047589,0.0870222,0.07070554,0.052575916,0.034446288,0.018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.19579996,0.38978696,0.5855869,0.7795739,0.97537386,0.8792868,0.7850128,0.69073874,0.5946517,0.50037766,0.42060733,0.34083697,0.25925365,0.1794833,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.07795739,0.15410182,0.23205921,0.3100166,0.387974,0.70342946,1.017072,1.3325275,1.647983,1.9616255,1.8292793,1.696933,1.5645868,1.4322405,1.2998942,2.1646774,3.0294604,3.8942437,4.76084,5.6256227,5.369995,5.1143675,4.860553,4.604925,4.349297,3.4990177,2.6505513,1.8002719,0.9499924,0.099712946,0.08339628,0.065266654,0.047137026,0.030820364,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.13053331,0.24837588,0.36440548,0.48224804,0.6000906,0.9644961,1.3307146,1.69512,2.0595255,2.4257438,2.6795588,2.9351864,3.1908143,3.444629,3.7002566,5.230397,6.7605376,8.290678,9.820818,11.349146,9.867955,8.384952,6.9019485,5.4207582,3.9377546,4.40006,4.8623657,5.3246713,5.7869763,6.249282,6.4269524,6.604623,6.782293,6.9599633,7.137634,7.9770355,8.81825,9.657652,10.497053,11.338268,11.512312,11.6881695,11.862214,12.038072,12.212116,10.991992,9.771869,8.551744,7.3316207,6.11331,5.562169,5.0128417,4.461701,3.9123733,3.3630457,3.247016,3.1327994,3.0167696,2.902553,2.7883365,2.4003625,2.0123885,1.6244144,1.2382535,0.85027945,1.1004683,1.3506571,1.6008459,1.8492218,2.0994108,3.000453,3.8996825,4.800725,5.6999545,6.599184,7.3406854,8.080374,8.820063,9.5597515,10.29944,8.539054,6.78048,5.0200934,3.2597067,1.49932,1.2799516,1.0605831,0.83940166,0.6200332,0.40066472,0.3208944,0.23931105,0.15954071,0.07977036,0.0,0.17585737,0.34990177,0.52575916,0.69980353,0.87566096,1.7621996,2.6505513,3.53709,4.4254417,5.3119802,5.045475,4.7771564,4.510651,4.2423325,3.975827,3.245203,2.514579,1.7857682,1.0551442,0.3245203,0.3444629,0.36440548,0.38434806,0.40429065,0.42423326,0.69436467,0.9644961,1.2346275,1.504759,1.7748904,1.7368182,1.7005589,1.6624867,1.6244144,1.5881553,1.5247015,1.4630609,1.3996071,1.3379664,1.2745126,1.3143979,1.3542831,1.3959812,1.4358664,1.4757515,1.7132497,1.9507477,2.1882458,2.4257438,2.663242,2.1701162,1.6769904,1.1856775,0.69255173,0.19942589,0.44961473,0.69980353,0.9499924,1.2001812,1.4503701,1.1893034,0.9300498,0.67079616,0.40972954,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.032633327,0.065266654,0.09789998,0.13053331,0.16316663,0.3045777,0.44780177,0.58921283,0.7324369,0.87566096,1.1222239,1.3705997,1.6171626,1.8655385,2.1121013,1.8945459,1.6769904,1.4594349,1.2418793,1.0243238,1.258196,1.4902552,1.7223145,1.9543737,2.1882458,1.9507477,1.7132497,1.4757515,1.2382535,1.0007553,1.0116332,1.0243238,1.0370146,1.0497054,1.062396,1.1457924,1.2273756,1.310772,1.3923552,1.4757515,1.8673514,2.2607644,2.6523643,3.045777,3.437377,3.4482548,3.4573197,3.4681973,3.4772623,3.48814,3.1744974,2.8626678,2.5508385,2.2371957,1.9253663,2.0432088,2.1592383,2.277081,2.3949237,2.5127661,4.0882306,3.8906176,3.6930048,3.4953918,3.2977788,3.100166,3.0820365,3.0657198,3.04759,3.0294604,3.0131438,3.4591327,3.9069343,4.3547363,4.802538,5.2503395,5.522284,5.7942286,6.0679855,6.33993,6.6118746,6.8004227,6.987158,7.175706,7.362441,7.549176,8.629702,9.710228,10.790753,11.869466,12.949992,12.0416975,11.135216,10.226922,9.32044,8.412147,8.160145,7.9081426,7.654328,7.402326,7.1503243,7.1521373,7.155763,7.157576,7.159389,7.1630154,7.211965,7.262728,7.311678,7.362441,7.413204,7.0342946,6.6571984,6.2801023,5.903006,5.524097,5.3391747,5.1542525,4.9693303,4.784408,4.599486,4.9693303,5.3391747,5.710832,6.0806766,6.450521,6.7696023,7.0904965,7.409578,7.7304726,8.049554,8.488291,8.925215,9.362139,9.800876,10.2378,9.91328,9.5869465,9.262425,8.937905,8.613385,8.375887,8.138389,7.900891,7.663393,7.4258947,7.224656,7.02523,6.825804,6.624565,6.4251394,5.8758116,5.3246713,4.7753434,4.2242026,3.6748753,3.29234,2.909805,2.5272698,2.1447346,1.7621996,1.5392052,1.3180238,1.0950294,0.872035,0.6508536,0.5656443,0.48043507,0.39522585,0.3100166,0.22480737,0.21936847,0.21574254,0.21030366,0.20486477,0.19942589,0.23931105,0.27919623,0.3208944,0.36077955,0.40066472,0.40791658,0.41516843,0.4224203,0.42967212,0.43692398,0.5873999,0.73787576,0.8883517,1.0370146,1.1874905,3.6930048,6.1967063,8.70222,11.207735,13.713249,12.868408,12.021755,11.176914,10.332074,9.487233,9.514427,9.541622,9.570629,9.597824,9.625018,8.609759,7.5945,6.5792413,5.565795,4.550536,4.0429068,3.5352771,3.0276475,2.520018,2.0123885,2.5417736,3.0729716,3.6023567,4.1317415,4.6629395,4.606738,4.552349,4.49796,4.441758,4.3873696,4.0102735,3.633177,3.254268,2.8771715,2.5000753,2.0758421,1.649796,1.2255627,0.7995165,0.37528324,1.1893034,2.0051367,2.819157,3.63499,4.4508233,6.104245,7.75948,9.414715,11.069949,12.725184,10.9774885,9.229793,7.4820967,5.7344007,3.9867048,3.4681973,2.9478772,2.427557,1.9072367,1.3869164,2.1229792,2.857229,3.5932918,4.327542,5.0617914,4.079166,3.0983531,2.1157274,1.1331016,0.15047589,0.59283876,1.0352017,1.4775645,1.9199274,2.3622901,2.3858588,2.4076142,2.42937,2.4529383,2.474694,2.2825198,2.0903459,1.8981718,1.7041848,1.5120108,2.420305,3.3267863,4.2350807,5.141562,6.049856,6.1241875,6.200332,6.2746634,6.350808,6.4251394,7.0433598,7.6597667,8.2779875,8.894395,9.512614,11.4126,13.312584,15.212569,17.112555,19.012539,19.904516,20.798307,21.690285,22.582262,23.476053,23.47968,23.485117,23.490557,23.495995,23.49962,22.154404,20.810997,19.465778,18.120562,16.775343,13.938056,11.10077,8.26167,5.424384,2.5870976,2.47832,2.3677292,2.2571385,2.1483607,2.03777,1.9271792,1.8184015,1.7078108,1.5972201,1.4866294,1.1983683,0.90829426,0.61822027,0.32814622,0.038072214,0.42785916,0.81764615,1.2074331,1.5972201,1.987007,1.8981718,1.8075237,1.7168756,1.6280404,1.5373923,1.2291887,0.922798,0.61459434,0.30820364,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.09427405,0.13959812,0.18492219,0.23024625,0.2755703,0.40066472,0.52575916,0.6508536,0.774135,0.89922947,0.7650702,0.629098,0.4949388,0.36077955,0.22480737,0.42423326,0.62547207,0.824898,1.0243238,1.2255627,1.0406405,0.8557183,0.67079616,0.48587397,0.2991388,0.23931105,0.1794833,0.11965553,0.059827764,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.35171473,0.6055295,0.8575313,1.1095331,1.3633479,1.1222239,0.88291276,0.6417888,0.40247768,0.16316663,1.5319533,2.902553,4.273153,5.6419396,7.0125394,6.6626377,6.3127356,5.962834,5.612932,5.2630305,4.233268,3.2016919,2.1719291,1.1421664,0.11240368,0.15047589,0.18673515,0.22480737,0.26287958,0.2991388,0.2755703,0.25018883,0.22480737,0.19942589,0.17585737,0.13959812,0.10515183,0.07070554,0.034446288,0.0,0.0,0.0,0.0,0.0,0.0,0.38978696,0.7795739,1.1693609,1.5591478,1.9507477,1.6352923,1.3198367,1.0043813,0.69073874,0.37528324,0.3154555,0.25562772,0.19579996,0.13415924,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.15410182,0.3100166,0.46411842,0.6200332,0.774135,0.968122,1.1602961,1.35247,1.5446441,1.7368182,1.5845293,1.4322405,1.2799516,1.1276628,0.97537386,1.6298534,2.2843328,2.9406252,3.5951047,4.249584,4.0519714,3.8543584,3.6567454,3.4591327,3.2633326,2.6251698,1.987007,1.3506571,0.7124943,0.07433146,0.065266654,0.054388877,0.045324065,0.034446288,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.18492219,0.3444629,0.5058166,0.6653573,0.824898,1.4793775,2.13567,2.7901495,3.444629,4.099108,4.3855567,4.670192,4.954827,5.239462,5.524097,6.2728505,7.019791,7.7667317,8.515485,9.262425,8.459284,7.6579537,6.8548117,6.051669,5.2503395,5.600241,5.9501433,6.300045,6.6499467,6.9998484,6.7677894,6.53573,6.301858,6.069799,5.8377395,6.717026,7.5981264,8.477413,9.3567,10.2378,10.263181,10.28675,10.312131,10.337513,10.362894,9.222541,8.082188,6.9418335,5.803293,4.6629395,4.2368937,3.8126602,3.386614,2.962381,2.5381477,2.6070402,2.6777458,2.7466383,2.817344,2.8880494,2.4366217,1.987007,1.5373923,1.0877775,0.63816285,0.824898,1.0116332,1.2001812,1.3869164,1.5754645,2.2498865,2.9243085,3.6005437,4.274966,4.949388,5.505967,6.060734,6.6155005,7.170267,7.7250338,6.530291,5.335549,4.1408067,2.9442513,1.7495089,1.5591478,1.3705997,1.1802386,0.9898776,0.7995165,0.6399758,0.48043507,0.3208944,0.15954071,0.0,0.13778515,0.2755703,0.41335547,0.5493277,0.6871128,1.4122978,2.137483,2.8626678,3.587853,4.313038,4.177066,4.0429068,3.9069343,3.7727752,3.636803,3.0276475,2.4166791,1.8075237,1.1983683,0.5873999,0.5402629,0.49312583,0.44417584,0.39703882,0.34990177,0.73968875,1.1294757,1.5192627,1.9108626,2.3006494,2.1628644,2.0250793,1.887294,1.7495089,1.6117238,1.7875811,1.9616255,2.137483,2.3133402,2.4873846,2.5671551,2.6469254,2.7266958,2.808279,2.8880494,3.0620937,3.2379513,3.4119956,3.587853,3.7618973,3.0765975,2.3931105,1.7078108,1.0225109,0.33721104,0.48768693,0.63816285,0.7868258,0.93730164,1.0877775,0.8919776,0.6979906,0.50219065,0.30820364,0.11240368,0.09064813,0.06707962,0.045324065,0.02175555,0.0,0.052575916,0.10515183,0.15772775,0.21030366,0.26287958,0.4224203,0.581961,0.7433147,0.90285534,1.062396,1.1820517,1.3017071,1.4231756,1.5428312,1.6624867,1.551896,1.4431182,1.3325275,1.2219368,1.1131591,1.2908293,1.4666867,1.6443571,1.8220274,1.9996977,1.7875811,1.5754645,1.3633479,1.1494182,0.93730164,1.0243238,1.1131591,1.2001812,1.2872034,1.3742256,1.4141108,1.455809,1.4956942,1.5355793,1.5754645,1.8220274,2.0704033,2.3169663,2.565342,2.811905,2.8699198,2.9279346,2.9841363,3.0421512,3.100166,2.9007401,2.6995013,2.5000753,2.3006494,2.0994108,2.1973107,2.2952106,2.3931105,2.4891977,2.5870976,3.7256382,3.6222992,3.5207734,3.4174345,3.3140955,3.2125697,3.1545548,3.0983531,3.0403383,2.9823234,2.9243085,3.339477,3.7546456,4.169814,4.5849824,5.0001507,5.377247,5.754343,6.1332526,6.510349,6.887445,7.2754188,7.663393,8.049554,8.437528,8.825501,9.619579,10.41547,11.209548,12.005438,12.799516,12.132345,11.465176,10.798005,10.130835,9.461852,9.414715,9.367578,9.32044,9.273304,9.224354,8.997733,8.7693,8.54268,8.314246,8.087626,8.049554,8.013294,7.9752226,7.93715,7.900891,7.665206,7.4295206,7.1956487,6.9599633,6.7242785,6.697084,6.6698895,6.642695,6.6155005,6.588306,6.5176005,6.446895,6.378002,6.3072968,6.2365913,6.4051967,6.5719895,6.740595,6.9073873,7.07418,7.8628187,8.649645,9.438283,10.225109,11.011934,10.56232,10.112705,9.663091,9.211663,8.762048,8.537241,8.312433,8.087626,7.8628187,7.6380115,7.5382986,7.4367723,7.3370595,7.2373466,7.137634,6.43783,5.7380266,5.038223,4.3366065,3.636803,3.395679,3.152742,2.909805,2.666868,2.4257438,2.13567,1.845596,1.5555218,1.2654479,0.97537386,0.8466535,0.7197462,0.59283876,0.46411842,0.33721104,0.32995918,0.32270733,0.3154555,0.30820364,0.2991388,0.36077955,0.42060733,0.48043507,0.5402629,0.6000906,0.58014804,0.56020546,0.5402629,0.52032024,0.50037766,0.5620184,0.62547207,0.6871128,0.7505665,0.8122072,2.9315605,5.0527267,7.17208,9.293246,11.4126,10.781689,10.152591,9.52168,8.892582,8.26167,8.609759,8.957849,9.304124,9.652213,10.000301,8.814624,7.6307597,6.445082,5.2594047,4.07554,3.8072214,3.540716,3.2723975,3.005892,2.7375734,3.2832751,3.827164,4.3728657,4.9167547,5.462456,5.317419,5.1723824,5.027345,4.882308,4.7372713,4.4145637,4.0918565,3.7691493,3.4482548,3.1255474,2.5508385,1.9743162,1.3996071,0.824898,0.25018883,1.5355793,2.819157,4.1045475,5.389938,6.6753283,7.420456,8.165584,8.910711,9.655839,10.399154,9.046683,7.6942134,6.341743,4.989273,3.636803,3.1454902,2.6523643,2.1592383,1.6679256,1.1747998,2.3151531,3.4555066,4.59586,5.7344007,6.874754,5.520471,4.164375,2.810092,1.455809,0.099712946,0.39522585,0.69073874,0.98443866,1.2799516,1.5754645,1.7023718,1.8292793,1.9579996,2.084907,2.2118144,2.1683033,2.1229792,2.077655,2.032331,1.987007,3.3177216,4.646623,5.977338,7.308052,8.636953,8.350506,8.062244,7.7757964,7.4875355,7.1992745,7.0324817,6.8656893,6.697084,6.530291,6.3616858,7.6253204,8.887142,10.150778,11.4126,12.674421,13.357908,14.039582,14.723069,15.404743,16.086416,16.05741,16.026588,15.9975815,15.966762,15.937754,15.245202,14.55265,13.860099,13.167547,12.474996,10.388275,8.299743,6.2130227,4.12449,2.03777,1.9217403,1.8075237,1.693307,1.5772774,1.4630609,1.3724127,1.2817645,1.1929294,1.1022812,1.0116332,0.81583315,0.61822027,0.42060733,0.2229944,0.025381476,0.28463513,0.54570174,0.80495536,1.064209,1.3252757,1.2654479,1.2056202,1.1457924,1.0841516,1.0243238,0.8194591,0.61459434,0.40972954,0.20486477,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.14322405,0.21030366,0.27738327,0.3444629,0.41335547,0.6000906,0.7868258,0.97537386,1.162109,1.3506571,1.1476053,0.9445535,0.7433147,0.5402629,0.33721104,0.4749962,0.61278135,0.7505665,0.8883517,1.0243238,0.85934424,0.69436467,0.5293851,0.36440548,0.19942589,0.15954071,0.11965553,0.07977036,0.03988518,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.37165734,0.5946517,0.81764615,1.0406405,1.261822,1.0533313,0.8430276,0.6327239,0.4224203,0.21211663,1.1294757,2.0468347,2.9641938,3.8833659,4.800725,4.836984,4.8750563,4.9131284,4.949388,4.98746,4.004834,3.0222087,2.039583,1.0569572,0.07433146,0.099712946,0.12509441,0.15047589,0.17585737,0.19942589,0.21211663,0.22480737,0.2374981,0.25018883,0.26287958,0.21030366,0.15772775,0.10515183,0.052575916,0.0,0.0,0.0,0.0,0.0,0.0,0.5855869,1.1693609,1.7549478,2.3405347,2.9243085,2.3894846,1.8546607,1.3198367,0.7850128,0.25018883,0.21030366,0.17041849,0.13053331,0.09064813,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.23205921,0.46411842,0.6979906,0.9300498,1.162109,1.2328146,1.3017071,1.3724127,1.4431182,1.5120108,1.3397794,1.167548,0.99531645,0.823085,0.6508536,1.0950294,1.5392052,1.9851941,2.42937,2.8753586,2.7357605,2.5943494,2.4547513,2.3151531,2.175555,1.7495089,1.3252757,0.89922947,0.4749962,0.05076295,0.047137026,0.045324065,0.04169814,0.03988518,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.23931105,0.44236287,0.64541465,0.8466535,1.0497054,1.9942589,2.9406252,3.8851788,4.8297324,5.774286,6.089741,6.4051967,6.720652,7.0342946,7.3497505,7.315304,7.2808576,7.2445984,7.210152,7.175706,7.0524244,6.929143,6.8076744,6.684393,6.5629244,6.8004227,7.037921,7.2754188,7.512917,7.750415,7.1068134,6.4650245,5.823236,5.179634,4.537845,5.4570174,6.378002,7.2971745,8.21816,9.137331,9.012237,8.887142,8.762048,8.636953,8.511859,7.453089,6.392506,5.331923,4.273153,3.2125697,2.911618,2.612479,2.3133402,2.0123885,1.7132497,1.9670644,2.222692,2.47832,2.7321346,2.9877625,2.474694,1.9616255,1.4503701,0.93730164,0.42423326,0.5493277,0.6744221,0.7995165,0.9246109,1.0497054,1.49932,1.9507477,2.4003625,2.8499773,3.299592,3.6694362,4.0392804,4.409125,4.780782,5.1506267,4.519716,3.8906176,3.2597067,2.6306088,1.9996977,1.840157,1.6806163,1.5192627,1.3597219,1.2001812,0.96087015,0.7197462,0.48043507,0.23931105,0.0,0.099712946,0.19942589,0.2991388,0.40066472,0.50037766,1.062396,1.6244144,2.1882458,2.7502642,3.3122826,3.3104696,3.3068438,3.3050308,3.303218,3.299592,2.810092,2.3205922,1.8292793,1.3397794,0.85027945,0.73424983,0.6200332,0.5058166,0.38978696,0.2755703,0.7850128,1.2944553,1.8057107,2.3151531,2.8245957,2.5870976,2.3495996,2.1121013,1.8746033,1.6371052,2.0504606,2.4620032,2.8753586,3.2869012,3.7002566,3.8199122,3.9395678,4.059223,4.1806917,4.3003473,4.4127507,4.5251546,4.6375585,4.749962,4.8623657,3.9848917,3.1074178,2.229944,1.35247,0.4749962,0.52575916,0.5747091,0.62547207,0.6744221,0.72518504,0.5946517,0.46411842,0.33539808,0.20486477,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.072518505,0.14503701,0.21755551,0.29007402,0.36259252,0.5402629,0.7179332,0.89560354,1.0732739,1.2491312,1.2418793,1.2346275,1.2273756,1.2201238,1.2128719,1.209246,1.2074331,1.2056202,1.2019942,1.2001812,1.3216497,1.4449311,1.5682126,1.6896812,1.8129625,1.6244144,1.4376793,1.2491312,1.062396,0.87566096,1.0370146,1.2001812,1.3633479,1.5247015,1.6878681,1.6842422,1.6824293,1.6806163,1.6769904,1.6751775,1.7767034,1.8800422,1.983381,2.084907,2.1882458,2.2915847,2.3967366,2.5018883,2.6070402,2.712192,2.6251698,2.5381477,2.4493124,2.3622901,2.275268,2.3532255,2.42937,2.5073273,2.5852847,2.663242,3.3630457,3.3557937,3.346729,3.339477,3.3322253,3.3249733,3.2270734,3.1291735,3.0330863,2.9351864,2.8372865,3.2198215,3.6023567,3.9848917,4.367427,4.749962,5.23221,5.714458,6.1967063,6.680767,7.1630154,7.750415,8.337815,8.925215,9.512614,10.100015,10.609457,11.120712,11.630155,12.139598,12.650853,12.222994,11.795135,11.367275,10.939416,10.51337,10.669285,10.827013,10.98474,11.142468,11.300196,10.843329,10.384649,9.927783,9.470917,9.012237,8.887142,8.762048,8.636953,8.511859,8.386765,8.294304,8.201842,8.109382,8.01692,7.9244595,8.054993,8.185526,8.314246,8.444779,8.575313,8.06587,7.554615,7.0451727,6.53573,6.0244746,6.0407915,6.055295,6.069799,6.0843024,6.1006193,7.2373466,8.374074,9.512614,10.649343,11.787883,11.213174,10.636651,10.061942,9.487233,8.912524,8.700407,8.488291,8.274362,8.062244,7.850128,7.850128,7.850128,7.850128,7.850128,7.850128,6.9998484,6.149569,5.2992897,4.4508233,3.6005437,3.4972048,3.395679,3.29234,3.1908143,3.0874753,2.7303216,2.373168,2.0142014,1.6570477,1.2998942,1.1294757,0.96087015,0.7904517,0.6200332,0.44961473,0.4405499,0.42967212,0.42060733,0.40972954,0.40066472,0.48043507,0.56020546,0.6399758,0.7197462,0.7995165,0.7523795,0.70524246,0.65810543,0.6091554,0.5620184,0.53663695,0.51306844,0.48768693,0.46230546,0.43692398,2.1719291,3.9069343,5.6419396,7.3769445,9.11195,8.696781,8.281613,7.8682575,7.453089,7.037921,7.705091,8.372261,9.039432,9.708415,10.375585,9.019489,7.665206,6.3091097,4.954827,3.6005437,3.5733492,3.5443418,3.5171473,3.489953,3.4627585,4.022964,4.5831695,5.143375,5.7017674,6.261973,6.0281005,5.7924156,5.5567303,5.3228583,5.087173,4.8206677,4.552349,4.2858434,4.017525,3.7492065,3.0258346,2.3006494,1.5754645,0.85027945,0.12509441,1.8800422,3.63499,5.389938,7.1448855,8.899834,8.734854,8.569874,8.404895,8.239915,8.074935,7.117691,6.1604466,5.2032027,4.2441454,3.2869012,2.8227828,2.3568513,1.892733,1.4268016,0.96268314,2.5073273,4.0519714,5.5984282,7.1430726,8.6877165,6.9599633,5.23221,3.5044568,1.7767034,0.05076295,0.19761293,0.3444629,0.49312583,0.6399758,0.7868258,1.020698,1.2527572,1.4848163,1.7168756,1.9507477,2.0522738,2.1556125,2.2571385,2.3604772,2.4620032,4.215138,5.9682727,7.7195945,9.47273,11.225864,10.57501,9.924157,9.275117,8.624263,7.9752226,7.023417,6.069799,5.1179934,4.164375,3.2125697,3.8380418,4.461701,5.087173,5.712645,6.338117,6.8094873,7.2826705,7.754041,8.227224,8.700407,8.63514,8.569874,8.504607,8.439341,8.374074,8.334189,8.294304,8.254418,8.214534,8.174648,6.836682,5.5005283,4.162562,2.8245957,1.4866294,1.3669738,1.2473183,1.1276628,1.0080072,0.8883517,0.81764615,0.7469406,0.678048,0.6073425,0.53663695,0.43329805,0.32814622,0.2229944,0.11784257,0.012690738,0.14322405,0.27194437,0.40247768,0.533011,0.66173136,0.6327239,0.60190356,0.5728962,0.5420758,0.51306844,0.40972954,0.30820364,0.20486477,0.10333887,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.19036107,0.27919623,0.36984438,0.4604925,0.5493277,0.7995165,1.0497054,1.2998942,1.550083,1.8002719,1.5301404,1.260009,0.9898776,0.7197462,0.44961473,0.52575916,0.6000906,0.6744221,0.7505665,0.824898,0.67986095,0.53482395,0.38978696,0.24474995,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03988518,0.07977036,0.11965553,0.15954071,0.19942589,0.3934129,0.5855869,0.7777609,0.969935,1.162109,0.9826257,0.8031424,0.62184614,0.44236287,0.26287958,0.726998,1.1929294,1.6570477,2.1229792,2.5870976,3.0131438,3.437377,3.8616104,4.2876563,4.7118897,3.778214,2.8427253,1.9072367,0.97174793,0.038072214,0.05076295,0.06164073,0.07433146,0.0870222,0.099712946,0.15047589,0.19942589,0.25018883,0.2991388,0.34990177,0.27919623,0.21030366,0.13959812,0.07070554,0.0,0.0,0.0,0.0,0.0,0.0,0.7795739,1.5591478,2.3405347,3.1201086,3.8996825,3.1454902,2.3894846,1.6352923,0.8792868,0.12509441,0.10515183,0.08520924,0.065266654,0.045324065,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.3100166,0.6200332,0.9300498,1.2400664,1.550083,1.4975071,1.4449311,1.3923552,1.3397794,1.2872034,1.0950294,0.90285534,0.7106813,0.5166943,0.3245203,0.56020546,0.79407763,1.0297627,1.2654479,1.49932,1.4177368,1.3343405,1.2527572,1.1693609,1.0877775,0.87566096,0.66173136,0.44961473,0.2374981,0.025381476,0.030820364,0.034446288,0.03988518,0.045324065,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.2955129,0.5402629,0.7850128,1.0297627,1.2745126,2.5109532,3.7455807,4.9802084,6.2148356,7.4494634,7.795739,8.140202,8.484665,8.829127,9.175404,8.357758,7.5401115,6.722465,5.904819,5.087173,5.6455655,6.202145,6.7605376,7.317117,7.8755093,8.000604,8.125698,8.2507925,8.375887,8.499168,7.4476504,6.394319,5.3428006,4.2894692,3.2379513,4.1970086,5.1578784,6.1169357,7.077806,8.036863,7.763106,7.4875355,7.211965,6.9382076,6.6626377,5.6818247,4.702825,3.7220123,2.7430124,1.7621996,1.5881553,1.4122978,1.2382535,1.062396,0.8883517,1.3270886,1.7676386,2.2081885,2.6469254,3.0874753,2.5127661,1.938057,1.3633479,0.7868258,0.21211663,0.2755703,0.33721104,0.40066472,0.46230546,0.52575916,0.7505665,0.97537386,1.2001812,1.4249886,1.649796,1.8347181,2.0196402,2.2045624,2.3894846,2.5744069,2.5091403,2.4456866,2.38042,2.3151531,2.2498865,2.1193533,1.9906329,1.8600996,1.7295663,1.6008459,1.2799516,0.96087015,0.6399758,0.3208944,0.0,0.06164073,0.12509441,0.18673515,0.25018883,0.31182957,0.7124943,1.1131591,1.5120108,1.9126755,2.3133402,2.4420607,2.572594,2.7031271,2.8318477,2.962381,2.5925364,2.222692,1.8528478,1.4830034,1.1131591,0.9300498,0.7469406,0.5656443,0.3825351,0.19942589,0.83033687,1.4594349,2.0903459,2.7194438,3.350355,3.0131438,2.6741197,2.3369088,1.9996977,1.6624867,2.3133402,2.962381,3.6132345,4.262275,4.9131284,5.0726695,5.23221,5.391751,5.5531044,5.712645,5.763408,5.812358,5.863121,5.9120708,5.962834,4.893186,3.8217251,2.752077,1.6824293,0.61278135,0.5620184,0.51306844,0.46230546,0.41335547,0.36259252,0.29732585,0.23205921,0.16679256,0.10333887,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.092461094,0.18492219,0.27738327,0.36984438,0.46230546,0.65810543,0.8520924,1.0478923,1.2418793,1.4376793,1.3017071,1.167548,1.0333886,0.8974165,0.76325727,0.8665961,0.97174793,1.0768998,1.1820517,1.2872034,1.3542831,1.4231756,1.4902552,1.5573349,1.6244144,1.4630609,1.2998942,1.1367276,0.97537386,0.8122072,1.0497054,1.2872034,1.5247015,1.7621996,1.9996977,1.9543737,1.9108626,1.8655385,1.8202144,1.7748904,1.7331922,1.6896812,1.647983,1.6044719,1.5627737,1.7150626,1.8673514,2.0196402,2.1719291,2.324218,2.3495996,2.374981,2.4003625,2.4257438,2.4493124,2.5073273,2.565342,2.6233568,2.6795588,2.7375734,3.000453,3.0874753,3.1744974,3.2633326,3.350355,3.437377,3.299592,3.1618068,3.0258346,2.8880494,2.7502642,3.100166,3.4500678,3.7999697,4.1498713,4.499773,5.087173,5.674573,6.261973,6.849373,7.4367723,8.225411,9.012237,9.800876,10.587702,11.374527,11.599335,11.8241415,12.050762,12.27557,12.500377,12.311829,12.125093,11.938358,11.74981,11.563075,11.925668,12.28826,12.650853,13.011633,13.374225,12.687112,11.999999,11.312886,10.625773,9.936848,9.724731,9.512614,9.300498,9.088382,8.874452,8.925215,8.974165,9.024928,9.07569,9.12464,9.412902,9.699349,9.987611,10.275872,10.56232,9.612328,8.662335,7.7123427,6.7623506,5.812358,5.674573,5.5367875,5.4008155,5.2630305,5.125245,6.6118746,8.100317,9.5869465,11.075388,12.562017,11.862214,11.162411,10.462607,9.762803,9.063,8.861761,8.662335,8.46291,8.26167,8.062244,8.161958,8.26167,8.363196,8.46291,8.562622,7.5618668,6.5629244,5.562169,4.5632267,3.5624714,3.6005437,3.636803,3.6748753,3.7129474,3.7492065,3.3249733,2.9007401,2.474694,2.0504606,1.6244144,1.4122978,1.2001812,0.9880646,0.774135,0.5620184,0.5493277,0.53663695,0.52575916,0.51306844,0.50037766,0.6000906,0.69980353,0.7995165,0.89922947,1.0007553,0.9246109,0.85027945,0.774135,0.69980353,0.62547207,0.51306844,0.40066472,0.28826106,0.17585737,0.06164073,1.4122978,2.762955,4.1117992,5.462456,6.813113,6.6118746,6.412449,6.2130227,6.011784,5.812358,6.8004227,7.7866745,8.774739,9.762803,10.750868,9.224354,7.699652,6.1749506,4.650249,3.1255474,3.3376641,3.5497808,3.7618973,3.975827,4.1879435,4.762653,5.337362,5.9120708,6.48678,7.063302,6.736969,6.412449,6.0879283,5.7615952,5.4370747,5.224958,5.0128417,4.800725,4.5867953,4.3746786,3.5008307,2.6251698,1.7495089,0.87566096,0.0,2.2245052,4.4508233,6.6753283,8.899834,11.124338,10.049252,8.974165,7.899078,6.825804,5.750717,5.186886,4.6248674,4.062849,3.5008307,2.9369993,2.5000753,2.0631514,1.6244144,1.1874905,0.7505665,2.6995013,4.650249,6.599184,8.549932,10.500679,8.399456,6.300045,4.2006345,2.0994108,0.0,0.0,0.0,0.0,0.0,0.0,0.33721104,0.6744221,1.0116332,1.3506571,1.6878681,1.938057,2.1882458,2.4366217,2.6868105,2.9369993,5.1125546,7.28811,9.461852,11.637406,13.812962,12.799516,11.787883,10.774437,9.762803,8.749357,7.0125394,5.275721,3.53709,1.8002719,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.26287958,0.52575916,0.7868258,1.0497054,1.3125849,1.2128719,1.1131591,1.0116332,0.9119202,0.8122072,1.4249886,2.03777,2.6505513,3.2633326,3.874301,3.2869012,2.6995013,2.1121013,1.5247015,0.93730164,0.8122072,0.6871128,0.5620184,0.43692398,0.31182957,0.26287958,0.21211663,0.16316663,0.11240368,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.2374981,0.34990177,0.46230546,0.5747091,0.6871128,1.0007553,1.3125849,1.6244144,1.938057,2.2498865,1.9126755,1.5754645,1.2382535,0.89922947,0.5620184,0.5747091,0.5873999,0.6000906,0.61278135,0.62547207,0.50037766,0.37528324,0.25018883,0.12509441,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,0.41335547,0.5747091,0.73787576,0.89922947,1.062396,0.9119202,0.76325727,0.61278135,0.46230546,0.31182957,0.3245203,0.33721104,0.34990177,0.36259252,0.37528324,1.1874905,1.9996977,2.811905,3.6241121,4.4381323,3.5497808,2.663242,1.7748904,0.8883517,0.0,0.0,0.0,0.0,0.0,0.0,0.0870222,0.17585737,0.26287958,0.34990177,0.43692398,0.34990177,0.26287958,0.17585737,0.0870222,0.0,0.0,0.0,0.0,0.0,0.0,0.97537386,1.9507477,2.9243085,3.8996825,4.8750563,3.8996825,2.9243085,1.9507477,0.97537386,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.387974,0.774135,1.162109,1.550083,1.938057,1.7621996,1.5881553,1.4122978,1.2382535,1.062396,0.85027945,0.63816285,0.42423326,0.21211663,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.34990177,0.63816285,0.9246109,1.2128719,1.49932,3.0258346,4.550536,6.0752378,7.5999393,9.12464,9.499924,9.875207,10.25049,10.625773,10.999244,9.400211,7.799365,6.200332,4.599486,3.000453,4.2368937,5.475147,6.7134004,7.949841,9.188094,9.200785,9.211663,9.224354,9.237044,9.249735,7.7866745,6.3254266,4.8623657,3.3993049,1.938057,2.9369993,3.9377546,4.936697,5.9374523,6.9382076,6.5121617,6.0879283,5.661882,5.237649,4.8116026,3.9123733,3.0131438,2.1121013,1.2128719,0.31182957,0.26287958,0.21211663,0.16316663,0.11240368,0.06164073,0.6871128,1.3125849,1.938057,2.561716,3.1871881,2.5508385,1.9126755,1.2745126,0.63816285,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.50037766,1.0007553,1.49932,1.9996977,2.5000753,2.4003625,2.3006494,2.1991236,2.0994108,1.9996977,1.6008459,1.2001812,0.7995165,0.40066472,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.36259252,0.6000906,0.8375887,1.0750868,1.3125849,1.5754645,1.8383441,2.0994108,2.3622901,2.6251698,2.374981,2.124792,1.8746033,1.6244144,1.3742256,1.1258497,0.87566096,0.62547207,0.37528324,0.12509441,0.87566096,1.6244144,2.374981,3.1255474,3.874301,3.437377,3.000453,2.561716,2.124792,1.6878681,2.5744069,3.4627585,4.349297,5.237649,6.1241875,6.3254266,6.5248523,6.7242785,6.925517,7.124943,7.112252,7.0995617,7.0868707,7.07418,7.063302,5.7996674,4.537845,3.2742105,2.0123885,0.7505665,0.6000906,0.44961473,0.2991388,0.15047589,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.11240368,0.22480737,0.33721104,0.44961473,0.5620184,0.774135,0.9880646,1.2001812,1.4122978,1.6244144,1.3633479,1.1004683,0.8375887,0.5747091,0.31182957,0.52575916,0.73787576,0.9499924,1.162109,1.3742256,1.3869164,1.3996071,1.4122978,1.4249886,1.4376793,1.2998942,1.162109,1.0243238,0.8883517,0.7505665,1.062396,1.3742256,1.6878681,1.9996977,2.3133402,2.2245052,2.137483,2.0504606,1.9616255,1.8746033,1.6878681,1.49932,1.3125849,1.1258497,0.93730164,1.1367276,1.3379664,1.5373923,1.7368182,1.938057,2.0758421,2.2118144,2.3495996,2.4873846,2.6251698,2.663242,2.6995013,2.7375734,2.7756457,2.811905,2.6378605,2.9007401,3.1618068,3.4246864,3.6875658,3.9504454,3.7075086,3.4645715,3.2216346,2.9805105,2.7375734,3.000453,3.2633326,3.5243993,3.787279,4.0501585,4.6303062,5.2104545,5.7906027,6.3707504,6.9490857,7.6180687,8.285239,8.952409,9.619579,10.28675,10.475298,10.662033,10.850581,11.037316,11.224051,11.111648,10.999244,10.88684,10.774437,10.662033,10.937603,11.213174,11.486931,11.762501,12.038072,11.514126,10.991992,10.469859,9.947725,9.425592,9.425592,9.425592,9.425592,9.425592,9.425592,9.3150015,9.2044115,9.0956335,8.985043,8.874452,9.177217,9.479981,9.782746,10.085511,10.388275,9.567003,8.747544,7.9280853,7.1068134,6.2873545,6.189454,6.093367,5.995467,5.8975673,5.7996674,7.166641,8.535428,9.902402,11.269376,12.638163,11.854962,11.071762,10.290376,9.507175,8.725789,8.529989,8.334189,8.140202,7.944402,7.750415,7.757667,7.764919,7.7721705,7.7794223,7.7866745,7.0542374,6.3218007,5.5893636,4.856927,4.12449,3.9903307,3.8543584,3.720199,3.584227,3.4500678,3.198066,2.9442513,2.6922495,2.4402475,2.1882458,1.9453088,1.7023718,1.4594349,1.2183108,0.97537386,0.94274056,0.9101072,0.8774739,0.8448406,0.8122072,0.96268314,1.1131591,1.261822,1.4122978,1.5627737,1.3796645,1.1983683,1.015259,0.8321498,0.6508536,0.6417888,0.6345369,0.62728506,0.6200332,0.61278135,1.7857682,2.956942,4.1299286,5.3029156,6.474089,6.450521,6.4251394,6.399758,6.3743763,6.350808,7.17208,7.995165,8.81825,9.639522,10.462607,9.373016,8.283426,7.192023,6.1024323,5.0128417,5.038223,5.0617914,5.087173,5.1125546,5.137936,5.4171324,5.6981416,5.977338,6.258347,6.5375433,6.1749506,5.812358,5.4497657,5.087173,4.7245803,4.690134,4.655688,4.6194286,4.5849824,4.550536,3.9051213,3.2597067,2.6142921,1.9706904,1.3252757,2.8826106,4.439945,5.99728,7.554615,9.11195,8.477413,7.842876,7.208339,6.5719895,5.9374523,5.235836,4.5324063,3.83079,3.1273603,2.4257438,2.1429217,1.8600996,1.5772774,1.2944553,1.0116332,2.6777458,4.3420453,6.008158,7.6724577,9.336758,7.4694057,5.6020546,3.7347028,1.8673514,0.0,0.06707962,0.13415924,0.2030518,0.27013144,0.33721104,0.5402629,0.7433147,0.9445535,1.1476053,1.3506571,1.550083,1.7495089,1.9507477,2.1501737,2.3495996,4.1045475,5.859495,7.614443,9.3693905,11.124338,10.489801,9.855265,9.220728,8.584378,7.949841,6.604623,5.2594047,3.9141862,2.570781,1.2255627,1.1403534,1.0551442,0.969935,0.88472575,0.7995165,0.9808127,1.1602961,1.3397794,1.5192627,1.7005589,1.6769904,1.6552348,1.6316663,1.6099107,1.5881553,2.0957847,2.6034143,3.1092308,3.6168604,4.12449,3.4700103,2.8155308,2.1592383,1.504759,0.85027945,0.7324369,0.61459434,0.49675176,0.38072214,0.26287958,0.21936847,0.17767033,0.13415924,0.092461094,0.05076295,0.054388877,0.059827764,0.065266654,0.07070554,0.07433146,0.065266654,0.054388877,0.045324065,0.034446288,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.17223145,0.15772775,0.14322405,0.12690738,0.11240368,0.25562772,0.39703882,0.5402629,0.68167394,0.824898,1.167548,1.5101979,1.8528478,2.1954978,2.5381477,2.220879,1.9017978,1.5845293,1.2672608,0.9499924,0.8883517,0.824898,0.76325727,0.69980353,0.63816285,0.5094425,0.3825351,0.25562772,0.12690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.06707962,0.11059072,0.15228885,0.19579996,0.2374981,0.36259252,0.48768693,0.61278135,0.73787576,0.8629702,0.7433147,0.62184614,0.50219065,0.3825351,0.26287958,0.27738327,0.291887,0.30820364,0.32270733,0.33721104,0.9808127,1.6226015,2.2643902,2.907992,3.5497808,2.8390994,2.1302311,1.4195497,0.7106813,0.0,0.0,0.0,0.0,0.0,0.0,0.38978696,0.7795739,1.1693609,1.5609608,1.9507477,1.7078108,1.4648738,1.2219368,0.9808127,0.73787576,0.59283876,0.44780177,0.30276474,0.15772775,0.012690738,0.7904517,1.5682126,2.3441606,3.1219215,3.8996825,3.1201086,2.3405347,1.5591478,0.7795739,0.0,0.20486477,0.40972954,0.61459434,0.8194591,1.0243238,0.8448406,0.6653573,0.48587397,0.3045777,0.12509441,0.40972954,0.69436467,0.9808127,1.2654479,1.550083,1.4122978,1.2745126,1.1367276,1.0007553,0.8629702,1.1820517,1.502946,1.8220274,2.1429217,2.4620032,1.9996977,1.5373923,1.0750868,0.61278135,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.054388877,0.08520924,0.11421664,0.14503701,0.17585737,0.46230546,0.7505665,1.0370146,1.3252757,1.6117238,1.6153497,1.6171626,1.6207886,1.6226015,1.6244144,2.8717327,4.119051,5.368182,6.6155005,7.8628187,8.363196,8.861761,9.362139,9.862516,10.362894,9.046683,7.7322855,6.4178877,5.101677,3.787279,4.64481,5.5023413,6.359873,7.217404,8.074935,7.9679704,7.859193,7.752228,7.645263,7.5382986,6.3616858,5.186886,4.0120864,2.8372865,1.6624867,2.4402475,3.2180085,3.9957695,4.7717175,5.5494785,5.2104545,4.8696175,4.5305934,4.1897564,3.8507326,3.1291735,2.4094272,1.6896812,0.969935,0.25018883,0.21030366,0.17041849,0.13053331,0.09064813,0.05076295,0.5493277,1.0497054,1.550083,2.0504606,2.5508385,2.039583,1.5301404,1.020698,0.5094425,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.41516843,0.83033687,1.2455053,1.6606737,2.0758421,2.0722163,2.0704033,2.0667772,2.0649643,2.0631514,1.7621996,1.4630609,1.162109,0.8629702,0.5620184,0.8774739,1.1929294,1.5083848,1.8220274,2.137483,2.1628644,2.1882458,2.2118144,2.2371957,2.2625773,2.5417736,2.8227828,3.101979,3.3829882,3.6621845,3.442816,3.2234476,3.002266,2.7828975,2.561716,2.1628644,1.7621996,1.3633479,0.96268314,0.5620184,1.2654479,1.9670644,2.6704938,3.3721104,4.07554,3.5479677,3.0203958,2.4928236,1.9652514,1.4376793,2.4384346,3.437377,4.4381323,5.4370747,6.43783,6.6553855,6.872941,7.0904965,7.308052,7.5256076,7.3424983,7.159389,6.978093,6.794984,6.6118746,5.4606433,4.307599,3.1545548,2.0033236,0.85027945,0.75963134,0.67079616,0.58014804,0.4894999,0.40066472,0.3245203,0.25018883,0.17585737,0.099712946,0.025381476,0.054388877,0.08520924,0.11421664,0.14503701,0.17585737,0.26469254,0.35534066,0.44417584,0.53482395,0.62547207,0.79226464,0.96087015,1.1276628,1.2944553,1.4630609,1.2382535,1.0116332,0.7868258,0.5620184,0.33721104,0.61459434,0.8919776,1.1693609,1.4467441,1.7241274,1.6280404,1.5301404,1.4322405,1.3343405,1.2382535,1.1947423,1.1530442,1.1095331,1.067835,1.0243238,1.310772,1.5954071,1.8800422,2.1646774,2.4493124,2.374981,2.3006494,2.2245052,2.1501737,2.0758421,1.8746033,1.6751775,1.4757515,1.2745126,1.0750868,1.2473183,1.4195497,1.5917811,1.7658255,1.938057,2.084907,2.231757,2.38042,2.5272698,2.6741197,2.7502642,2.8245957,2.9007401,2.9750717,3.049403,2.275268,2.712192,3.149116,3.587853,4.024777,4.461701,4.115425,3.7673361,3.4192474,3.0729716,2.7248828,2.9007401,3.0747845,3.2506418,3.4246864,3.6005437,4.171627,4.744523,5.317419,5.8903155,6.4632115,7.0107265,7.558241,8.105756,8.653271,9.200785,9.349448,9.499924,9.6504,9.800876,9.949538,9.91328,9.875207,9.837135,9.800876,9.762803,9.949538,10.138086,10.324821,10.51337,10.700105,10.342952,9.985798,9.626831,9.269678,8.912524,9.12464,9.336758,9.550687,9.762803,9.97492,9.704789,9.434657,9.164526,8.894395,8.624263,8.943344,9.2606125,9.577881,9.89515,10.212419,9.52168,8.832754,8.1420145,7.453089,6.7623506,6.7043357,6.6481338,6.590119,6.532104,6.474089,7.723221,8.970539,10.217857,11.465176,12.712494,11.847711,10.982927,10.118144,9.253361,8.386765,8.198216,8.007855,7.817495,7.6271334,7.4367723,7.3533764,7.268167,7.1829576,7.0977483,7.0125394,6.548421,6.0824895,5.618371,5.1524396,4.688321,4.3801174,4.071914,3.7655232,3.4573197,3.149116,3.0693457,2.9895754,2.909805,2.8300345,2.7502642,2.47832,2.2045624,1.9326181,1.6606737,1.3869164,1.3343405,1.2817645,1.2291887,1.1766127,1.1258497,1.3252757,1.5247015,1.7241274,1.9253663,2.124792,1.8347181,1.5446441,1.2545701,0.9644961,0.6744221,0.77232206,0.87022203,0.968122,1.064209,1.162109,2.1574254,3.152742,4.1480584,5.143375,6.1368785,6.2873545,6.43783,6.588306,6.736969,6.887445,7.5455503,8.201842,8.859948,9.518054,10.174346,9.519867,8.865387,8.209095,7.554615,6.9001355,6.736969,6.5756154,6.412449,6.249282,6.0879283,6.071612,6.057108,6.0426044,6.0281005,6.011784,5.612932,5.2122674,4.8116026,4.4127507,4.0120864,4.15531,4.2967215,4.439945,4.5831695,4.7245803,4.309412,3.8942437,3.4790752,3.0657198,2.6505513,3.540716,4.4290676,5.319232,6.209397,7.0995617,6.9055743,6.7097745,6.5157876,6.319988,6.1241875,5.282973,4.439945,3.5969179,2.7557032,1.9126755,1.7857682,1.6570477,1.5301404,1.403233,1.2745126,2.6541772,4.0356545,5.4153194,6.794984,8.174648,6.539356,4.9058766,3.2705846,1.6352923,0.0,0.13415924,0.27013144,0.40429065,0.5402629,0.6744221,0.7433147,0.8103943,0.8774739,0.9445535,1.0116332,1.162109,1.3125849,1.4630609,1.6117238,1.7621996,3.0983531,4.4326935,5.767034,7.1031876,8.437528,8.180087,7.9226465,7.665206,7.407765,7.1503243,6.1967063,5.2449007,4.2930956,3.339477,2.3876717,2.229944,2.0722163,1.9144884,1.7567607,1.6008459,1.696933,1.794833,1.892733,1.9906329,2.08672,2.1429217,2.1973107,2.2516994,2.3079014,2.3622901,2.764768,3.1672456,3.5697234,3.972201,4.3746786,3.6531196,2.9297476,2.2081885,1.4848163,0.76325727,0.6526665,0.5420758,0.43329805,0.32270733,0.21211663,0.17767033,0.14322405,0.10696479,0.072518505,0.038072214,0.059827764,0.08339628,0.10515183,0.12690738,0.15047589,0.13053331,0.11059072,0.09064813,0.07070554,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.07433146,0.15047589,0.22480737,0.2991388,0.37528324,0.3208944,0.26469254,0.21030366,0.15410182,0.099712946,0.27194437,0.44417584,0.61822027,0.7904517,0.96268314,1.3343405,1.7078108,2.079468,2.4529383,2.8245957,2.5272698,2.229944,1.9326181,1.6352923,1.3379664,1.2001812,1.062396,0.9246109,0.7868258,0.6508536,0.52032024,0.38978696,0.25925365,0.13053331,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.08520924,0.11965553,0.15410182,0.19036107,0.22480737,0.31182957,0.40066472,0.48768693,0.5747091,0.66173136,0.5728962,0.48224804,0.39159992,0.30276474,0.21211663,0.23024625,0.24837588,0.26469254,0.28282216,0.2991388,0.77232206,1.2455053,1.7168756,2.1900587,2.663242,2.1302311,1.5972201,1.064209,0.533011,0.0,0.0,0.0,0.0,0.0,0.0,0.69255173,1.3851035,2.077655,2.770207,3.4627585,3.0657198,2.666868,2.269829,1.8727903,1.4757515,1.1856775,0.89560354,0.6055295,0.3154555,0.025381476,0.6055295,1.1856775,1.7658255,2.3441606,2.9243085,2.3405347,1.7549478,1.1693609,0.5855869,0.0,0.40972954,0.8194591,1.2291887,1.6407311,2.0504606,1.6896812,1.3307146,0.969935,0.6091554,0.25018883,0.43329805,0.61459434,0.79770356,0.9808127,1.162109,1.062396,0.96268314,0.8629702,0.76325727,0.66173136,1.5156367,2.3677292,3.2198215,4.071914,4.9258194,3.974014,3.0258346,2.0758421,1.1258497,0.17585737,0.13959812,0.10515183,0.07070554,0.034446288,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.09789998,0.14503701,0.19217403,0.23931105,0.28826106,0.8629702,1.4376793,2.0123885,2.5870976,3.1618068,2.8807976,2.5979755,2.3151531,2.032331,1.7495089,2.7194438,3.6893787,4.6593137,5.6292486,6.599184,7.224656,7.850128,8.4756,9.099259,9.724731,8.694968,7.665206,6.635443,5.6056805,4.574105,5.0527267,5.529536,6.008158,6.484967,6.9617763,6.735156,6.506723,6.2801023,6.051669,5.825049,4.936697,4.0501585,3.1618068,2.275268,1.3869164,1.9416829,2.4982624,3.053029,3.6077955,4.162562,3.9069343,3.6531196,3.397492,3.141864,2.8880494,2.3477864,1.8075237,1.2672608,0.726998,0.18673515,0.15772775,0.12690738,0.09789998,0.06707962,0.038072214,0.41335547,0.7868258,1.162109,1.5373923,1.9126755,1.5301404,1.1476053,0.7650702,0.3825351,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.32995918,0.65991837,0.9898776,1.3198367,1.649796,1.745883,1.840157,1.9344311,2.030518,2.124792,1.9253663,1.7241274,1.5247015,1.3252757,1.1258497,1.7295663,2.335096,2.9406252,3.5443418,4.1498713,3.9631362,3.774588,3.587853,3.3993049,3.2125697,3.5098956,3.8072214,4.1045475,4.401873,4.699199,4.510651,4.3202896,4.1299286,3.9395678,3.7492065,3.199879,2.6505513,2.0994108,1.550083,1.0007553,1.6552348,2.3097143,2.9641938,3.6204863,4.274966,3.6567454,3.0403383,2.422118,1.8057107,1.1874905,2.3006494,3.4119956,4.5251546,5.638314,6.7496595,6.985345,7.219217,7.454902,7.690587,7.9244595,7.572745,7.219217,6.867502,6.5157876,6.16226,5.1198063,4.077353,3.0348995,1.9924458,0.9499924,0.91917205,0.8901646,0.85934424,0.83033687,0.7995165,0.6508536,0.50037766,0.34990177,0.19942589,0.05076295,0.11059072,0.17041849,0.23024625,0.29007402,0.34990177,0.4169814,0.48587397,0.5529536,0.6200332,0.6871128,0.8103943,0.9318628,1.0551442,1.1766127,1.2998942,1.1131591,0.9246109,0.73787576,0.5493277,0.36259252,0.70524246,1.0478923,1.3905423,1.7331922,2.0758421,1.8673514,1.6606737,1.452183,1.2455053,1.0370146,1.0895905,1.1421664,1.1947423,1.2473183,1.2998942,1.5573349,1.8147756,2.0722163,2.3296568,2.5870976,2.525457,2.4620032,2.4003625,2.3369088,2.275268,2.0631514,1.8492218,1.6371052,1.4249886,1.2128719,1.357909,1.502946,1.647983,1.79302,1.938057,2.0957847,2.2516994,2.4094272,2.5671551,2.7248828,2.8372865,2.94969,3.0620937,3.1744974,3.2869012,1.9126755,2.525457,3.1382382,3.7492065,4.361988,4.974769,4.5233417,4.070101,3.6168604,3.1654327,2.712192,2.7992141,2.8880494,2.9750717,3.0620937,3.149116,3.7147603,4.2804046,4.844236,5.40988,5.975525,6.401571,6.82943,7.2572894,7.6851482,8.113008,8.225411,8.337815,8.450218,8.562622,8.675026,8.713099,8.749357,8.78743,8.825501,8.861761,8.963287,9.063,9.162713,9.262425,9.362139,9.169965,8.977791,8.785617,8.59163,8.399456,8.825501,9.249735,9.675781,10.100015,10.524248,10.094576,9.664904,9.235231,8.805559,8.375887,8.70766,9.039432,9.373016,9.704789,10.038374,9.4781685,8.917963,8.357758,7.797552,7.2373466,7.219217,7.2029004,7.1847706,7.166641,7.1503243,8.2779875,9.40565,10.533313,11.6591625,12.786825,11.840459,10.89228,9.944099,8.997733,8.049554,7.8646317,7.6797094,7.494787,7.309865,7.124943,6.947273,6.7696023,6.591932,6.414262,6.2365913,6.0407915,5.8431783,5.6455655,5.4479527,5.2503395,4.7699046,4.2894692,3.8108473,3.3304121,2.8499773,2.9424384,3.0348995,3.1273603,3.2198215,3.3122826,3.009518,2.7067533,2.4058013,2.1030366,1.8002719,1.7277533,1.6552348,1.5827163,1.5101979,1.4376793,1.6878681,1.938057,2.1882458,2.4366217,2.6868105,2.2897718,1.892733,1.4956942,1.0968424,0.69980353,0.90285534,1.1059072,1.3071461,1.5101979,1.7132497,2.5308957,3.346729,4.164375,4.9820213,5.7996674,6.1241875,6.450521,6.775041,7.0995617,7.4258947,7.9172077,8.410334,8.901647,9.394773,9.8878975,9.666717,9.447348,9.22798,9.006798,8.78743,8.437528,8.087626,7.7377243,7.3878226,7.037921,6.7279043,6.4178877,6.107871,5.7978544,5.487838,5.049101,4.612177,4.175253,3.738329,3.299592,3.6204863,3.9395678,4.2604623,4.5795436,4.900438,4.7155156,4.5305934,4.345671,4.160749,3.975827,4.1970086,4.420003,4.6429973,4.8641787,5.087173,5.331923,5.576673,5.823236,6.0679855,6.3127356,5.33011,4.347484,3.3648586,2.382233,1.3996071,1.4268016,1.455809,1.4830034,1.5101979,1.5373923,2.6324217,3.727451,4.8224807,5.91751,7.0125394,5.6093063,4.207886,2.8046532,1.403233,0.0,0.2030518,0.40429065,0.6073425,0.8103943,1.0116332,0.9445535,0.8774739,0.8103943,0.7433147,0.6744221,0.774135,0.87566096,0.97537386,1.0750868,1.1747998,2.0903459,3.004079,3.919625,4.835171,5.750717,5.870373,5.9900284,6.109684,6.2293396,6.350808,5.7906027,5.230397,4.670192,4.1099863,3.5497808,3.3195345,3.0892882,2.8608549,2.6306088,2.4003625,2.4148662,2.42937,2.4456866,2.4601903,2.474694,2.6070402,2.7393866,2.8717327,3.005892,3.1382382,3.435564,3.73289,4.0302157,4.327542,4.6248674,3.834416,3.045777,2.2553256,1.4648738,0.6744221,0.5728962,0.46955732,0.3680314,0.26469254,0.16316663,0.13415924,0.10696479,0.07977036,0.052575916,0.025381476,0.065266654,0.10515183,0.14503701,0.18492219,0.22480737,0.19579996,0.16497959,0.13415924,0.10515183,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.11240368,0.22480737,0.33721104,0.44961473,0.5620184,0.46774435,0.37165734,0.27738327,0.18310922,0.0870222,0.29007402,0.49312583,0.69436467,0.8974165,1.1004683,1.502946,1.9054236,2.3079014,2.7103791,3.1128569,2.8354735,2.5580902,2.280707,2.0033236,1.7241274,1.5120108,1.2998942,1.0877775,0.87566096,0.66173136,0.5293851,0.39703882,0.26469254,0.13234627,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.07433146,0.07433146,0.07433146,0.07433146,0.07433146,0.10333887,0.13053331,0.15772775,0.18492219,0.21211663,0.26287958,0.31182957,0.36259252,0.41335547,0.46230546,0.40247768,0.34264994,0.28282216,0.2229944,0.16316663,0.18310922,0.2030518,0.2229944,0.24293698,0.26287958,0.5656443,0.8665961,1.1693609,1.4721256,1.7748904,1.4195497,1.064209,0.7106813,0.35534066,0.0,0.0,0.0,0.0,0.0,0.0,0.99531645,1.9906329,2.9859493,3.9794528,4.974769,4.421816,3.870675,3.3177216,2.764768,2.2118144,1.7767034,1.3434052,0.90829426,0.47318324,0.038072214,0.42060733,0.8031424,1.1856775,1.5682126,1.9507477,1.5591478,1.1693609,0.7795739,0.38978696,0.0,0.61459434,1.2291887,1.845596,2.4601903,3.0747845,2.5345216,1.9942589,1.455809,0.9155461,0.37528324,0.4550536,0.53482395,0.61459434,0.69436467,0.774135,0.7124943,0.6508536,0.5873999,0.52575916,0.46230546,1.8474089,3.2325122,4.6176157,6.002719,7.3878226,5.9501433,4.512464,3.0747845,1.6371052,0.19942589,0.15954071,0.11965553,0.07977036,0.03988518,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.13959812,0.20486477,0.27013144,0.33539808,0.40066472,1.261822,2.124792,2.9877625,3.8507326,4.7118897,4.1444325,3.576975,3.009518,2.4420607,1.8746033,2.5671551,3.2597067,3.9522583,4.64481,5.337362,6.0879283,6.836682,7.5872483,8.337815,9.088382,8.343254,7.5981264,6.8529987,6.107871,5.3627434,5.4606433,5.5567303,5.65463,5.75253,5.8504305,5.5023413,5.1542525,4.8079767,4.459888,4.1117992,3.5117085,2.911618,2.3133402,1.7132497,1.1131591,1.4449311,1.7767034,2.1102884,2.4420607,2.7756457,2.6052272,2.4348087,2.2643902,2.0957847,1.9253663,1.5645868,1.2056202,0.8448406,0.48587397,0.12509441,0.10515183,0.08520924,0.065266654,0.045324065,0.025381476,0.2755703,0.52575916,0.774135,1.0243238,1.2745126,1.020698,0.7650702,0.5094425,0.25562772,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.24474995,0.4894999,0.73424983,0.9808127,1.2255627,1.4177368,1.6099107,1.8020848,1.9942589,2.1882458,2.08672,1.987007,1.887294,1.7875811,1.6878681,2.5834718,3.4772623,4.3728657,5.2684693,6.16226,5.763408,5.3627434,4.9620786,4.5632267,4.162562,4.478018,4.7916603,5.1071157,5.422571,5.7380266,5.576673,5.4171324,5.2575917,5.0980506,4.936697,4.2368937,3.53709,2.8372865,2.137483,1.4376793,2.0450218,2.6523643,3.2597067,3.8670492,4.4743915,3.7673361,3.0602808,2.3532255,1.6443571,0.93730164,2.1628644,3.386614,4.612177,5.8377395,7.063302,7.315304,7.567306,7.819308,8.073122,8.325124,7.802991,7.2808576,6.7569118,6.2347784,5.712645,4.780782,3.8471067,2.9152439,1.983381,1.0497054,1.0805258,1.1095331,1.1403534,1.1693609,1.2001812,0.97537386,0.7505665,0.52575916,0.2991388,0.07433146,0.16497959,0.25562772,0.3444629,0.43511102,0.52575916,0.56927025,0.61459434,0.65991837,0.70524246,0.7505665,0.82671094,0.90466833,0.9826257,1.0605831,1.1367276,0.9880646,0.8375887,0.6871128,0.53663695,0.387974,0.79589057,1.2019942,1.6099107,2.0178273,2.4257438,2.1066625,1.789394,1.4721256,1.1548572,0.8375887,0.98443866,1.1331016,1.2799516,1.4268016,1.5754645,1.8057107,2.034144,2.2643902,2.4946365,2.7248828,2.6741197,2.6251698,2.5744069,2.525457,2.474694,2.2498865,2.0250793,1.8002719,1.5754645,1.3506571,1.4666867,1.5845293,1.7023718,1.8202144,1.938057,2.1048496,2.2716422,2.4402475,2.6070402,2.7756457,2.9243085,3.0747845,3.2252605,3.3757362,3.5243993,1.550083,2.3369088,3.1255474,3.9123733,4.699199,5.487838,4.9294453,4.3728657,3.8144734,3.2578938,2.6995013,2.6995013,2.6995013,2.6995013,2.6995013,2.6995013,3.2578938,3.8144734,4.3728657,4.9294453,5.487838,5.7942286,6.1024323,6.4106355,6.717026,7.02523,7.0995617,7.175706,7.250037,7.324369,7.400513,7.512917,7.6253204,7.7377243,7.850128,7.9625316,7.9752226,7.987913,8.000604,8.013294,8.024173,7.996978,7.9697833,7.9425893,7.915395,7.8882003,8.52455,9.162713,9.800876,10.437225,11.075388,10.484363,9.89515,9.304124,8.714911,8.125698,8.471974,8.820063,9.168152,9.514427,9.862516,9.432844,9.003172,8.571687,8.1420145,7.7123427,7.7359114,7.757667,7.7794223,7.802991,7.8247466,8.832754,9.840761,10.846955,11.854962,12.862969,11.833207,10.801631,9.771869,8.7421055,7.7123427,7.5328593,7.3533764,7.17208,6.9925966,6.813113,6.542982,6.2728505,6.002719,5.732588,5.462456,5.5331616,5.6020546,5.67276,5.7416525,5.812358,5.1596913,4.507025,3.8543584,3.2016919,2.5508385,2.8155308,3.0802233,3.3449159,3.6096084,3.874301,3.5425289,3.2107568,2.8771715,2.5453994,2.2118144,2.1193533,2.0268922,1.9344311,1.84197,1.7495089,2.0504606,2.3495996,2.6505513,2.94969,3.2506418,2.7448254,2.2408218,1.7350051,1.2291887,0.72518504,1.0333886,1.3397794,1.647983,1.9543737,2.2625773,2.902553,3.5425289,4.1825047,4.8224807,5.462456,5.962834,6.4632115,6.9617763,7.462154,7.9625316,8.290678,8.617011,8.945157,9.273304,9.599637,9.815379,10.029309,10.245051,10.460794,10.674724,10.138086,9.599637,9.063,8.52455,7.987913,7.382384,6.776854,6.1731377,5.567608,4.9620786,4.4870825,4.0120864,3.53709,3.0620937,2.5870976,3.0856624,3.5824142,4.079166,4.5777307,5.0744824,5.1198063,5.1651306,5.2104545,5.2557783,5.2992897,4.855114,4.409125,3.9649491,3.5207734,3.0747845,3.7600844,4.445384,5.130684,5.814171,6.4994707,5.377247,4.255023,3.1327994,2.0105755,0.8883517,1.0696479,1.2527572,1.4358664,1.6171626,1.8002719,2.610666,3.4192474,4.229642,5.040036,5.8504305,4.6792564,3.5098956,2.3405347,1.1693609,0.0,0.27013144,0.5402629,0.8103943,1.0805258,1.3506571,1.1476053,0.9445535,0.7433147,0.5402629,0.33721104,0.387974,0.43692398,0.48768693,0.53663695,0.5873999,1.0823387,1.5772774,2.0722163,2.5671551,3.0620937,3.5606585,4.0574102,4.554162,5.0527267,5.5494785,5.382686,5.2158933,5.047288,4.880495,4.7118897,4.409125,4.1081734,3.8054085,3.5026438,3.199879,3.1327994,3.0657198,2.9968271,2.9297476,2.8626678,3.0729716,3.2832751,3.491766,3.7020695,3.9123733,4.1045475,4.2967215,4.4907084,4.6828823,4.8750563,4.017525,3.159994,2.3024626,1.4449311,0.5873999,0.49312583,0.39703882,0.30276474,0.20667773,0.11240368,0.092461094,0.072518505,0.052575916,0.032633327,0.012690738,0.07070554,0.12690738,0.18492219,0.24293698,0.2991388,0.25925365,0.21936847,0.1794833,0.13959812,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.15047589,0.2991388,0.44961473,0.6000906,0.7505665,0.61459434,0.48043507,0.3444629,0.21030366,0.07433146,0.30820364,0.5402629,0.77232206,1.0043813,1.2382535,1.6697385,2.1030366,2.5345216,2.9678197,3.3993049,3.141864,2.8844235,2.6269827,2.3695421,2.1121013,1.8256533,1.5373923,1.2491312,0.96268314,0.6744221,0.5402629,0.40429065,0.27013144,0.13415924,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.099712946,0.099712946,0.099712946,0.099712946,0.099712946,0.11965553,0.13959812,0.15954071,0.1794833,0.19942589,0.21211663,0.22480737,0.2374981,0.25018883,0.26287958,0.23205921,0.2030518,0.17223145,0.14322405,0.11240368,0.13415924,0.15772775,0.1794833,0.2030518,0.22480737,0.35715362,0.4894999,0.62184614,0.7541924,0.8883517,0.7106813,0.533011,0.35534066,0.17767033,0.0,0.0,0.0,0.0,0.0,0.0,1.2980812,2.5943494,3.8924308,5.1905117,6.48678,5.7797246,5.0726695,4.365614,3.6567454,2.94969,2.3695421,1.789394,1.209246,0.629098,0.05076295,0.23568514,0.42060733,0.6055295,0.7904517,0.97537386,0.7795739,0.5855869,0.38978696,0.19579996,0.0,0.8194591,1.6407311,2.4601903,3.2796493,4.100921,3.3793623,2.659616,1.93987,1.2201238,0.50037766,0.47680917,0.4550536,0.43329805,0.40972954,0.387974,0.36259252,0.33721104,0.31182957,0.28826106,0.26287958,2.180994,4.0972953,6.01541,7.931711,9.849826,7.9244595,6.000906,4.07554,2.1501737,0.22480737,0.1794833,0.13415924,0.09064813,0.045324065,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.18310922,0.26469254,0.3480888,0.42967212,0.51306844,1.6624867,2.811905,3.9631362,5.1125546,6.261973,5.40988,4.557788,3.7056956,2.8517902,1.9996977,2.4148662,2.8300345,3.245203,3.6603715,4.07554,4.949388,5.825049,6.70071,7.574558,8.450218,7.989726,7.5292335,7.0705543,6.6100616,6.149569,5.866747,5.5857377,5.3029156,5.0200934,4.7372713,4.269527,3.8017826,3.3358512,2.8681068,2.4003625,2.08672,1.7748904,1.4630609,1.1494182,0.8375887,0.9481794,1.0569572,1.167548,1.2781386,1.3869164,1.3017071,1.2183108,1.1331016,1.0478923,0.96268314,0.78319985,0.60190356,0.4224203,0.24293698,0.06164073,0.052575916,0.04169814,0.032633327,0.02175555,0.012690738,0.13778515,0.26287958,0.387974,0.51306844,0.63816285,0.5094425,0.3825351,0.25562772,0.12690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.15954071,0.3208944,0.48043507,0.6399758,0.7995165,1.0895905,1.3796645,1.6697385,1.9598125,2.2498865,2.2498865,2.2498865,2.2498865,2.2498865,2.2498865,3.435564,4.6194286,5.805106,6.9907837,8.174648,7.5618668,6.9508986,6.338117,5.7253356,5.1125546,5.4443264,5.7779117,6.109684,6.4432693,6.775041,6.644508,6.5157876,6.3852544,6.2547207,6.1241875,5.275721,4.4254417,3.5751622,2.7248828,1.8746033,2.4348087,2.9950142,3.5552197,4.115425,4.6756306,3.877927,3.0802233,2.2825198,1.4848163,0.6871128,2.0250793,3.3630457,4.699199,6.037165,7.3751316,7.645263,7.915395,8.185526,8.455658,8.725789,8.033237,7.3406854,6.6481338,5.955582,5.2630305,4.439945,3.6168604,2.7955883,1.9725033,1.1494182,1.2400664,1.3307146,1.4195497,1.5101979,1.6008459,1.2998942,1.0007553,0.69980353,0.40066472,0.099712946,0.21936847,0.34083697,0.4604925,0.58014804,0.69980353,0.72337204,0.7451276,0.7668832,0.7904517,0.8122072,0.8448406,0.8774739,0.9101072,0.94274056,0.97537386,0.8629702,0.7505665,0.63816285,0.52575916,0.41335547,0.88472575,1.357909,1.8292793,2.3024626,2.7756457,2.3477864,1.9199274,1.4920682,1.064209,0.63816285,0.8792868,1.1222239,1.3651608,1.6080978,1.8492218,2.0522738,2.2553256,2.4583774,2.659616,2.8626678,2.8245957,2.7883365,2.7502642,2.712192,2.6741197,2.4366217,2.1991236,1.9616255,1.7241274,1.4866294,1.5772774,1.6679256,1.7567607,1.8474089,1.938057,2.1157274,2.2933977,2.469255,2.6469254,2.8245957,3.0131438,3.199879,3.386614,3.5751622,3.7618973,1.1874905,2.1501737,3.1128569,4.07554,5.038223,6.000906,5.337362,4.6756306,4.0120864,3.350355,2.6868105,2.5997884,2.5127661,2.4257438,2.3369088,2.2498865,2.7992141,3.350355,3.8996825,4.4508233,5.0001507,5.186886,5.375434,5.562169,5.750717,5.9374523,5.975525,6.011784,6.049856,6.0879283,6.1241875,6.3127356,6.4994707,6.688019,6.874754,7.063302,6.987158,6.9128265,6.836682,6.7623506,6.688019,6.825804,6.9617763,7.0995617,7.2373466,7.3751316,8.225411,9.07569,9.924157,10.774437,11.624716,10.874149,10.125396,9.374829,8.624263,7.8755093,8.238102,8.600695,8.963287,9.325879,9.686659,9.38752,9.088382,8.78743,8.488291,8.187339,8.2507925,8.312433,8.375887,8.437528,8.499168,9.38752,10.275872,11.162411,12.050762,12.937301,11.8241415,10.712796,9.599637,8.488291,7.3751316,7.1992745,7.02523,6.849373,6.6753283,6.4994707,6.1368785,5.774286,5.411693,5.049101,4.688321,5.0255322,5.3627434,5.6999545,6.037165,6.3743763,5.5494785,4.7245803,3.8996825,3.0747845,2.2498865,2.6868105,3.1255474,3.5624714,3.9993954,4.4381323,4.07554,3.7129474,3.350355,2.9877625,2.6251698,2.5127661,2.4003625,2.2879589,2.175555,2.0631514,2.4130533,2.762955,3.1128569,3.4627585,3.8126602,3.199879,2.5870976,1.9743162,1.3633479,0.7505665,1.162109,1.5754645,1.987007,2.4003625,2.811905,3.2742105,3.738329,4.2006345,4.6629395,5.125245,5.7996674,6.474089,7.1503243,7.8247466,8.499168,8.662335,8.825501,8.9868555,9.1500225,9.313189,9.96223,10.613083,11.262123,11.912977,12.562017,11.836833,11.111648,10.388275,9.663091,8.937905,8.036863,7.137634,6.2365913,5.337362,4.4381323,3.925064,3.4119956,2.9007401,2.3876717,1.8746033,2.5508385,3.2252605,3.8996825,4.574105,5.2503395,5.524097,5.7996674,6.0752378,6.350808,6.624565,5.5132194,4.40006,3.2869012,2.175555,1.062396,2.1882458,3.3122826,4.4381323,5.562169,6.688019,5.424384,4.162562,2.9007401,1.6371052,0.37528324,0.7124943,1.0497054,1.3869164,1.7241274,2.0631514,2.5870976,3.1128569,3.636803,4.162562,4.688321,3.7492065,2.811905,1.8746033,0.93730164,0.0,0.33721104,0.6744221,1.0116332,1.3506571,1.6878681,1.3506571,1.0116332,0.6744221,0.33721104,0.0,0.0,0.0,0.0,0.0,0.0,0.07433146,0.15047589,0.22480737,0.2991388,0.37528324,1.2491312,2.124792,3.000453,3.874301,4.749962,4.974769,5.199577,5.424384,5.6491914,5.8758116,5.5005283,5.125245,4.749962,4.3746786,3.9993954,3.8507326,3.7002566,3.5497808,3.3993049,3.2506418,3.53709,3.825351,4.1117992,4.40006,4.688321,4.7753434,4.8623657,4.949388,5.038223,5.125245,4.2006345,3.2742105,2.3495996,1.4249886,0.50037766,0.41335547,0.3245203,0.2374981,0.15047589,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.07433146,0.15047589,0.22480737,0.2991388,0.37528324,0.3245203,0.2755703,0.22480737,0.17585737,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.18673515,0.37528324,0.5620184,0.7505665,0.93730164,0.76325727,0.5873999,0.41335547,0.2374981,0.06164073,0.3245203,0.5873999,0.85027945,1.1131591,1.3742256,1.8383441,2.3006494,2.762955,3.2252605,3.6875658,3.4500678,3.2125697,2.9750717,2.7375734,2.5000753,2.137483,1.7748904,1.4122978,1.0497054,0.6871128,0.5493277,0.41335547,0.2755703,0.13778515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.13778515,0.15047589,0.16316663,0.17585737,0.18673515,0.16316663,0.13778515,0.11240368,0.0870222,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.0870222,0.11240368,0.13778515,0.16316663,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.6008459,3.199879,4.800725,6.399758,8.000604,7.137634,6.2746634,5.411693,4.550536,3.6875658,2.962381,2.2371957,1.5120108,0.7868258,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,1.0243238,2.0504606,3.0747845,4.100921,5.125245,4.2242026,3.3249733,2.4257438,1.5247015,0.62547207,0.50037766,0.37528324,0.25018883,0.12509441,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,2.5127661,4.9620786,7.413204,9.862516,12.311829,9.900589,7.4875355,5.0744824,2.663242,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.22480737,0.3245203,0.42423326,0.52575916,0.62547207,2.0631514,3.5008307,4.936697,6.3743763,7.8120556,6.6753283,5.5367875,4.40006,3.2633326,2.124792,2.2625773,2.4003625,2.5381477,2.6741197,2.811905,3.8126602,4.8116026,5.812358,6.813113,7.8120556,7.6380115,7.462154,7.28811,7.112252,6.9382076,6.2746634,5.612932,4.949388,4.2876563,3.6241121,3.0367124,2.4493124,1.8619126,1.2745126,0.6871128,0.66173136,0.63816285,0.61278135,0.5873999,0.5620184,0.44961473,0.33721104,0.22480737,0.11240368,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07433146,0.15047589,0.22480737,0.2991388,0.37528324,0.76325727,1.1494182,1.5373923,1.9253663,2.3133402,2.4130533,2.5127661,2.612479,2.712192,2.811905,4.2876563,5.7615952,7.2373466,8.713099,10.1870365,9.362139,8.537241,7.7123427,6.887445,6.0625467,6.412449,6.7623506,7.112252,7.462154,7.8120556,7.7123427,7.61263,7.512917,7.413204,7.311678,6.3127356,5.3119802,4.313038,3.3122826,2.3133402,2.8245957,3.3376641,3.8507326,4.361988,4.8750563,3.9867048,3.100166,2.2118144,1.3252757,0.43692398,1.887294,3.3376641,4.788034,6.2365913,7.686961,7.9752226,8.26167,8.549932,8.838193,9.12464,8.26167,7.400513,6.5375433,5.674573,4.8116026,4.099108,3.388427,2.6741197,1.9634385,1.2491312,1.3996071,1.550083,1.7005589,1.8492218,1.9996977,1.6244144,1.2491312,0.87566096,0.50037766,0.12509441,0.2755703,0.42423326,0.5747091,0.72518504,0.87566096,0.87566096,0.87566096,0.87566096,0.87566096,0.87566096,0.8629702,0.85027945,0.8375887,0.824898,0.8122072,0.73787576,0.66173136,0.5873999,0.51306844,0.43692398,0.97537386,1.5120108,2.0504606,2.5870976,3.1255474,2.5870976,2.0504606,1.5120108,0.97537386,0.43692398,0.774135,1.1131591,1.4503701,1.7875811,2.124792,2.3006494,2.474694,2.6505513,2.8245957,3.000453,2.9750717,2.94969,2.9243085,2.9007401,2.8753586,2.6251698,2.374981,2.124792,1.8746033,1.6244144,1.6878681,1.7495089,1.8129625,1.8746033,1.938057,2.124792,2.3133402,2.5000753,2.6868105,2.8753586,3.100166,3.3249733,3.5497808,3.774588,3.9993954,2.374981,3.0784104,3.780027,4.4816437,5.185073,5.8866897,5.3047285,4.7227674,4.1408067,3.5570326,2.9750717,2.8844235,2.7955883,2.70494,2.6142921,2.525457,2.9406252,3.3557937,3.7691493,4.1843176,4.599486,4.7898474,4.9802084,5.1705694,5.3591175,5.5494785,5.667321,5.7851634,5.903006,6.0208488,6.1368785,6.3725634,6.6082487,6.8421206,7.077806,7.311678,7.2772317,7.2427855,7.208339,7.17208,7.137634,7.0850577,7.0324817,6.979906,6.92733,6.874754,7.817495,8.760235,9.702975,10.645717,11.586644,10.926725,10.266808,9.606889,8.94697,8.287052,8.629702,8.972352,9.3150015,9.657652,10.000301,9.768243,9.53437,9.302311,9.070251,8.838193,8.747544,8.656897,8.568061,8.477413,8.386765,9.030367,9.672155,10.315757,10.957546,11.599335,10.749055,9.900589,9.050309,8.200029,7.3497505,7.228282,7.1050005,6.981719,6.8602505,6.736969,6.3653116,5.9918413,5.620184,5.2467136,4.8750563,5.0998635,5.3246713,5.5494785,5.774286,5.999093,5.2648435,4.5305934,3.7945306,3.0602808,2.324218,2.6904364,3.054842,3.4192474,3.785466,4.1498713,3.7981565,3.444629,3.092914,2.7393866,2.3876717,2.2716422,2.1574254,2.0432088,1.9271792,1.8129625,2.0649643,2.3169663,2.570781,2.8227828,3.0747845,2.5798457,2.084907,1.5899682,1.0950294,0.6000906,0.99531645,1.3905423,1.7857682,2.179181,2.5744069,3.1726844,3.7691493,4.367427,4.9657044,5.562169,5.8522434,6.1423173,6.432391,6.722465,7.0125394,7.4966,7.9824743,8.4683485,8.952409,9.438283,9.880646,10.323009,10.765372,11.207735,11.650098,11.253058,10.854207,10.457169,10.060129,9.663091,8.569874,7.476658,6.3852544,5.292038,4.2006345,3.6930048,3.1853752,2.6777458,2.1701162,1.6624867,2.2371957,2.811905,3.386614,3.9631362,4.537845,4.7717175,5.0074024,5.243088,5.47696,5.712645,4.860553,4.006647,3.1545548,2.3024626,1.4503701,2.759329,4.070101,5.3808727,6.6898317,8.000604,6.542982,5.08536,3.6277382,2.1701162,0.7124943,0.9119202,1.1131591,1.3125849,1.5120108,1.7132497,2.1193533,2.5272698,2.9351864,3.343103,3.7492065,3.000453,2.2498865,1.49932,0.7505665,0.0,0.27013144,0.5402629,0.8103943,1.0805258,1.3506571,1.0805258,0.8103943,0.5402629,0.27013144,0.0,0.0,0.0,0.0,0.0,0.0,0.059827764,0.11965553,0.1794833,0.23931105,0.2991388,1.0007553,1.7005589,2.4003625,3.100166,3.7999697,3.9794528,4.160749,4.3402324,4.519716,4.699199,4.401873,4.1045475,3.8072214,3.5098956,3.2125697,3.2343252,3.2578938,3.2796493,3.303218,3.3249733,3.531651,3.7401419,3.9468195,4.15531,4.361988,4.3347936,4.307599,4.2804046,4.25321,4.2242026,3.5153344,2.8046532,2.0957847,1.3851035,0.6744221,0.6073425,0.5402629,0.47318324,0.40429065,0.33721104,0.34990177,0.36259252,0.37528324,0.387974,0.40066472,0.40972954,0.42060733,0.42967212,0.4405499,0.44961473,0.40791658,0.36440548,0.32270733,0.27919623,0.2374981,0.2030518,0.16679256,0.13234627,0.09789998,0.06164073,0.10696479,0.15228885,0.19761293,0.24293698,0.28826106,0.24293698,0.19761293,0.15228885,0.10696479,0.06164073,0.052575916,0.04169814,0.032633327,0.02175555,0.012690738,0.01994259,0.027194439,0.034446288,0.04169814,0.05076295,0.04169814,0.034446288,0.027194439,0.01994259,0.012690738,0.25925365,0.5076295,0.7541924,1.0025684,1.2491312,1.0352017,0.8194591,0.6055295,0.38978696,0.17585737,0.36077955,0.54570174,0.7306239,0.9155461,1.1004683,1.4703126,1.840157,2.2100015,2.5798457,2.94969,2.759329,2.570781,2.38042,2.1900587,1.9996977,1.7096237,1.4195497,1.1294757,0.83940166,0.5493277,0.44236287,0.33539808,0.22662032,0.11965553,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.099712946,0.099712946,0.099712946,0.099712946,0.099712946,0.11059072,0.11965553,0.13053331,0.13959812,0.15047589,0.13053331,0.11059072,0.09064813,0.07070554,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.07070554,0.09064813,0.11059072,0.13053331,0.15047589,0.20667773,0.26469254,0.32270733,0.38072214,0.43692398,0.44236287,0.44780177,0.45324063,0.45686656,0.46230546,0.37165734,0.28282216,0.19217403,0.10333887,0.012690738,1.2908293,2.5671551,3.8452935,5.121619,6.399758,5.709019,5.0200934,4.329355,3.6404288,2.94969,2.3695421,1.789394,1.209246,0.629098,0.05076295,0.0870222,0.12509441,0.16316663,0.19942589,0.2374981,0.5402629,0.8430276,1.1457924,1.4467441,1.7495089,2.570781,3.39024,4.209699,5.030971,5.8504305,4.802538,3.7546456,2.7067533,1.6606737,0.61278135,0.49312583,0.37165734,0.2520018,0.13234627,0.012690738,0.2755703,0.53663695,0.7995165,1.062396,1.3252757,3.141864,4.9602656,6.776854,8.595256,10.411844,8.437528,6.4632115,4.4870825,2.5127661,0.53663695,0.52032024,0.50219065,0.48587397,0.46774435,0.44961473,0.40066472,0.34990177,0.2991388,0.25018883,0.19942589,0.5148814,0.83033687,1.1457924,1.4594349,1.7748904,2.6904364,3.6041696,4.519716,5.4352617,6.350808,5.422571,4.494334,3.5679104,2.6396735,1.7132497,1.93987,2.1683033,2.3949237,2.6233568,2.8499773,3.7220123,4.59586,5.467895,6.33993,7.211965,6.9001355,6.588306,6.2746634,5.962834,5.6491914,5.0998635,4.550536,3.9993954,3.4500678,2.9007401,2.47832,2.0540867,1.6316663,1.209246,0.7868258,0.87022203,0.95180535,1.0352017,1.1167849,1.2001812,0.96087015,0.7197462,0.48043507,0.23931105,0.0,0.092461094,0.18492219,0.27738327,0.36984438,0.46230546,0.36984438,0.27738327,0.18492219,0.092461094,0.0,0.16679256,0.33539808,0.50219065,0.67079616,0.8375887,0.7668832,0.6979906,0.62728506,0.55839247,0.48768693,0.43329805,0.3770962,0.32270733,0.26831847,0.21211663,0.33539808,0.45686656,0.58014804,0.70342946,0.824898,0.6653573,0.5058166,0.3444629,0.18492219,0.025381476,0.038072214,0.05076295,0.06164073,0.07433146,0.0870222,0.15954071,0.23205921,0.3045777,0.3770962,0.44961473,0.9318628,1.4141108,1.8981718,2.38042,2.8626678,2.9841363,3.1074178,3.2306993,3.3521678,3.4754493,4.6846952,5.8957543,7.1050005,8.314246,9.525306,8.94697,8.370448,7.7921133,7.215591,6.637256,6.8403077,7.0433598,7.2445984,7.4476504,7.650702,7.560054,7.4694057,7.380571,7.2899227,7.1992745,6.454147,5.710832,4.9657044,4.220577,3.4754493,3.7401419,4.004834,4.269527,4.5342193,4.800725,4.4381323,4.07554,3.7129474,3.350355,2.9877625,3.7056956,4.421816,5.139749,5.857682,6.5756154,6.73153,6.889258,7.0469856,7.2047133,7.362441,6.94546,6.526665,6.109684,5.6927023,5.275721,4.514277,3.7546456,2.9950142,2.2353828,1.4757515,1.5228885,1.5700256,1.6171626,1.6642996,1.7132497,1.3923552,1.0732739,0.7523795,0.43329805,0.11240368,0.2374981,0.36259252,0.48768693,0.61278135,0.73787576,0.78319985,0.82671094,0.872035,0.91735905,0.96268314,0.90829426,0.8520924,0.79770356,0.7433147,0.6871128,0.6327239,0.57833505,0.52213323,0.46774435,0.41335547,0.88472575,1.357909,1.8292793,2.3024626,2.7756457,2.3641033,1.9543737,1.5446441,1.1349145,0.72518504,0.97537386,1.2255627,1.4757515,1.7241274,1.9743162,2.1175404,2.2607644,2.4021754,2.5453994,2.6868105,2.7919624,2.8971143,3.002266,3.1074178,3.2125697,2.9895754,2.7683938,2.5453994,2.322405,2.0994108,2.1973107,2.2952106,2.3931105,2.4891977,2.5870976,2.8354735,3.0820365,3.3304121,3.576975,3.825351,4.1045475,4.3855567,4.664753,4.945762,5.224958,3.5624714,4.004834,4.4471974,4.88956,5.331923,5.774286,5.272095,4.7699046,4.267714,3.7655232,3.2633326,3.1708715,3.0765975,2.9841363,2.8916752,2.7992141,3.0802233,3.3594196,3.6404288,3.919625,4.2006345,4.3928084,4.5849824,4.7771564,4.9693303,5.163317,5.3591175,5.5567303,5.754343,5.9519563,6.149569,6.432391,6.7152133,6.9980354,7.2808576,7.5618668,7.567306,7.572745,7.5781837,7.5818095,7.5872483,7.344311,7.1031876,6.8602505,6.6173134,6.3743763,7.409578,8.444779,9.479981,10.515183,11.5503845,10.979301,10.410031,9.840761,9.269678,8.700407,9.023115,9.345822,9.666717,9.989424,10.312131,10.147152,9.982172,9.817192,9.652213,9.487233,9.244296,9.003172,8.760235,8.517298,8.274362,8.673213,9.070251,9.467291,9.864329,10.263181,9.675781,9.088382,8.499168,7.911769,7.324369,7.2554765,7.1847706,7.115878,7.0451727,6.9744673,6.591932,6.209397,5.826862,5.4443264,5.0617914,5.1741953,5.2865987,5.4008155,5.5132194,5.6256227,4.9802084,4.3347936,3.6893787,3.045777,2.4003625,2.6922495,2.9841363,3.2778363,3.5697234,3.8616104,3.5207734,3.1781235,2.8354735,2.4928236,2.1501737,2.032331,1.9144884,1.7966459,1.6806163,1.5627737,1.7168756,1.8727903,2.0268922,2.182807,2.3369088,1.9598125,1.5827163,1.2056202,0.82671094,0.44961473,0.82671094,1.2056202,1.5827163,1.9598125,2.3369088,3.0693457,3.8017826,4.5342193,5.2666564,5.999093,5.904819,5.810545,5.714458,5.620184,5.52591,6.3326783,7.1394467,7.948028,8.754796,9.563377,9.79725,10.032935,10.266808,10.502492,10.738177,10.667472,10.596766,10.527874,10.457169,10.388275,9.102885,7.817495,6.532104,5.2467136,3.9631362,3.4591327,2.956942,2.4547513,1.9525607,1.4503701,1.9253663,2.4003625,2.8753586,3.350355,3.825351,4.019338,4.215138,4.410938,4.604925,4.800725,4.207886,3.6150475,3.0222087,2.42937,1.8383441,3.3322253,4.8279195,6.3218007,7.817495,9.313189,7.6597667,6.008158,4.3547363,2.7031271,1.0497054,1.1131591,1.1747998,1.2382535,1.2998942,1.3633479,1.651609,1.9416829,2.231757,2.521831,2.811905,2.2498865,1.6878681,1.1258497,0.5620184,0.0,0.2030518,0.40429065,0.6073425,0.8103943,1.0116332,0.8103943,0.6073425,0.40429065,0.2030518,0.0,0.0,0.0,0.0,0.0,0.0,0.045324065,0.09064813,0.13415924,0.1794833,0.22480737,0.7505665,1.2745126,1.8002719,2.324218,2.8499773,2.9841363,3.1201086,3.254268,3.39024,3.5243993,3.3050308,3.0856624,2.864481,2.6451125,2.4257438,2.619731,2.8155308,3.009518,3.2053177,3.3993049,3.5280252,3.6549325,3.7818398,3.9105604,4.0374675,3.8942437,3.7528327,3.6096084,3.4681973,3.3249733,2.8300345,2.335096,1.840157,1.3452182,0.85027945,0.8031424,0.7541924,0.7070554,0.65991837,0.61278135,0.6508536,0.6871128,0.72518504,0.76325727,0.7995165,0.7451276,0.69073874,0.6345369,0.58014804,0.52575916,0.4894999,0.4550536,0.42060733,0.38434806,0.34990177,0.3045777,0.25925365,0.21574254,0.17041849,0.12509441,0.21574254,0.3045777,0.39522585,0.48587397,0.5747091,0.47318324,0.36984438,0.26831847,0.16497959,0.06164073,0.054388877,0.047137026,0.03988518,0.032633327,0.025381476,0.027194439,0.030820364,0.032633327,0.034446288,0.038072214,0.034446288,0.032633327,0.030820364,0.027194439,0.025381476,0.33177215,0.6399758,0.9481794,1.2545701,1.5627737,1.3071461,1.0533313,0.79770356,0.5420758,0.28826106,0.39522585,0.50219065,0.6091554,0.7179332,0.824898,1.1022812,1.3796645,1.6570477,1.9344311,2.2118144,2.0704033,1.9271792,1.7857682,1.6425442,1.49932,1.2817645,1.064209,0.8466535,0.629098,0.41335547,0.33539808,0.2574407,0.1794833,0.10333887,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.07433146,0.07433146,0.07433146,0.07433146,0.07433146,0.08339628,0.09064813,0.09789998,0.10515183,0.11240368,0.09789998,0.08339628,0.06707962,0.052575916,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.052575916,0.06707962,0.08339628,0.09789998,0.11240368,0.26469254,0.4169814,0.56927025,0.72337204,0.87566096,0.88472575,0.89560354,0.90466833,0.9155461,0.9246109,0.7451276,0.5656443,0.38434806,0.20486477,0.025381476,0.9808127,1.9344311,2.8898623,3.8452935,4.800725,4.2822175,3.7655232,3.247016,2.7303216,2.2118144,1.7767034,1.3434052,0.90829426,0.47318324,0.038072214,0.12509441,0.21211663,0.2991388,0.387974,0.4749962,1.0805258,1.6842422,2.2897718,2.8953013,3.5008307,4.115425,4.7300196,5.3446136,5.959208,6.5756154,5.37906,4.1843176,2.9895754,1.794833,0.6000906,0.48587397,0.36984438,0.25562772,0.13959812,0.025381476,0.53663695,1.0497054,1.5627737,2.0758421,2.5870976,3.7727752,4.95664,6.1423173,7.327995,8.511859,6.9744673,5.4370747,3.8996825,2.3622901,0.824898,0.83940166,0.8557183,0.87022203,0.88472575,0.89922947,0.774135,0.6508536,0.52575916,0.40066472,0.2755703,0.80495536,1.3343405,1.8655385,2.3949237,2.9243085,3.3177216,3.7093215,4.102734,4.494334,4.8877473,4.169814,3.4518807,2.7357605,2.0178273,1.2998942,1.6171626,1.9344311,2.2516994,2.570781,2.8880494,3.633177,4.3783045,5.123432,5.866747,6.6118746,6.16226,5.712645,5.2630305,4.8134155,4.361988,3.925064,3.48814,3.049403,2.612479,2.175555,1.9181144,1.6606737,1.403233,1.1457924,0.8883517,1.0768998,1.2672608,1.4576219,1.647983,1.8383441,1.4703126,1.1022812,0.73424983,0.3680314,0.0,0.18492219,0.36984438,0.55476654,0.73968875,0.9246109,0.73968875,0.55476654,0.36984438,0.18492219,0.0,0.33539808,0.67079616,1.0043813,1.3397794,1.6751775,1.5355793,1.3941683,1.2545701,1.114972,0.97537386,0.86478317,0.7541924,0.64541465,0.53482395,0.42423326,0.67079616,0.9155461,1.1602961,1.405046,1.649796,1.3307146,1.0098201,0.69073874,0.36984438,0.05076295,0.07433146,0.099712946,0.12509441,0.15047589,0.17585737,0.24474995,0.3154555,0.38434806,0.4550536,0.52575916,1.1022812,1.6806163,2.2571385,2.8354735,3.4119956,3.5570326,3.7020695,3.8471067,3.9921436,4.137181,5.081734,6.0281005,6.972654,7.9172077,8.861761,8.531802,8.201842,7.8718834,7.5419245,7.211965,7.268167,7.322556,7.3769445,7.4331465,7.4875355,7.407765,7.327995,7.2482243,7.166641,7.0868707,6.5973706,6.107871,5.618371,5.127058,4.6375585,4.655688,4.6720047,4.690134,4.708264,4.7245803,4.8877473,5.049101,5.2122674,5.375434,5.5367875,5.522284,5.5077806,5.4932766,5.47696,5.462456,5.4896507,5.516845,5.5458527,5.573047,5.600241,5.6274357,5.65463,5.6818247,5.710832,5.7380266,4.9294453,4.122677,3.3140955,2.5073273,1.7005589,1.6443571,1.5899682,1.5355793,1.4793775,1.4249886,1.1602961,0.89560354,0.629098,0.36440548,0.099712946,0.19942589,0.2991388,0.40066472,0.50037766,0.6000906,0.69073874,0.7795739,0.87022203,0.96087015,1.0497054,0.95180535,0.8557183,0.75781834,0.65991837,0.5620184,0.5275721,0.49312583,0.45686656,0.4224203,0.387974,0.79589057,1.2019942,1.6099107,2.0178273,2.4257438,2.1429217,1.8600996,1.5772774,1.2944553,1.0116332,1.1747998,1.3379664,1.49932,1.6624867,1.8256533,1.9344311,2.0450218,2.1556125,2.2643902,2.374981,2.610666,2.8445382,3.0802233,3.3140955,3.5497808,3.3557937,3.159994,2.9641938,2.770207,2.5744069,2.7067533,2.8390994,2.9732587,3.105605,3.2379513,3.5443418,3.8525455,4.160749,4.4671397,4.7753434,5.1107416,5.4443264,5.7797246,6.115123,6.450521,4.749962,4.933071,5.1143675,5.297477,5.480586,5.661882,5.239462,4.8170414,4.3946214,3.972201,3.5497808,3.4555066,3.3594196,3.2651455,3.1708715,3.0747845,3.2198215,3.3648586,3.5098956,3.6549325,3.7999697,3.9957695,4.1897564,4.3855567,4.5795436,4.7753434,5.0527267,5.33011,5.6074934,5.8848767,6.16226,6.492219,6.8221784,7.1521373,7.4820967,7.8120556,7.85738,7.902704,7.948028,7.993352,8.036863,7.605378,7.17208,6.740595,6.3072968,5.8758116,7.0016613,8.129324,9.256987,10.384649,11.512312,11.0318775,10.553255,10.07282,9.592385,9.11195,9.414715,9.71748,10.020245,10.323009,10.625773,10.527874,10.429974,10.332074,10.234174,10.138086,9.742861,9.347635,8.952409,8.557183,8.161958,8.314246,8.4683485,8.620637,8.772926,8.925215,8.600695,8.274362,7.949841,7.6253204,7.3008003,7.2826705,7.264541,7.2482243,7.230095,7.211965,6.8203654,6.4269524,6.035352,5.6419396,5.2503395,5.2503395,5.2503395,5.2503395,5.2503395,5.2503395,4.695573,4.1408067,3.584227,3.0294604,2.474694,2.6958754,2.9152439,3.1346123,3.3557937,3.5751622,3.24339,2.909805,2.5780327,2.2444477,1.9126755,1.79302,1.6733645,1.551896,1.4322405,1.3125849,1.3705997,1.4268016,1.4848163,1.5428312,1.6008459,1.3397794,1.0805258,0.8194591,0.56020546,0.2991388,0.65991837,1.020698,1.3796645,1.7404441,2.0994108,2.9678197,3.834416,4.702825,5.569421,6.43783,5.957395,5.47696,4.9983377,4.517903,4.0374675,5.1669436,6.298232,7.4277077,8.557183,9.686659,9.715667,9.742861,9.770056,9.79725,9.824444,10.081885,10.339326,10.596766,10.854207,11.111648,9.635896,8.158332,6.680767,5.2032027,3.7256382,3.2270734,2.7303216,2.231757,1.7350051,1.2382535,1.6117238,1.987007,2.3622901,2.7375734,3.1128569,3.2669585,3.4228733,3.576975,3.73289,3.8869917,3.5552197,3.2216346,2.8898623,2.5580902,2.2245052,3.9051213,5.5857377,7.264541,8.945157,10.625773,8.778365,6.930956,5.081734,3.2343252,1.3869164,1.3125849,1.2382535,1.162109,1.0877775,1.0116332,1.1856775,1.357909,1.5301404,1.7023718,1.8746033,1.49932,1.1258497,0.7505665,0.37528324,0.0,0.13415924,0.27013144,0.40429065,0.5402629,0.6744221,0.5402629,0.40429065,0.27013144,0.13415924,0.0,0.0,0.0,0.0,0.0,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.50037766,0.85027945,1.2001812,1.550083,1.8999848,1.9906329,2.079468,2.1701162,2.2607644,2.3495996,2.2081885,2.0649643,1.9217403,1.7803292,1.6371052,2.0051367,2.373168,2.7393866,3.1074178,3.4754493,3.5225863,3.5697234,3.6168604,3.6658103,3.7129474,3.4555066,3.198066,2.9406252,2.6831846,2.4257438,2.1447346,1.8655385,1.5845293,1.305333,1.0243238,0.99712944,0.969935,0.94274056,0.9155461,0.8883517,0.9499924,1.0116332,1.0750868,1.1367276,1.2001812,1.0805258,0.96087015,0.83940166,0.7197462,0.6000906,0.5728962,0.54570174,0.5166943,0.4894999,0.46230546,0.40791658,0.35171473,0.29732585,0.24293698,0.18673515,0.32270733,0.45686656,0.59283876,0.726998,0.8629702,0.7016165,0.5420758,0.3825351,0.2229944,0.06164073,0.058014803,0.052575916,0.047137026,0.04169814,0.038072214,0.034446288,0.032633327,0.030820364,0.027194439,0.025381476,0.027194439,0.030820364,0.032633327,0.034446288,0.038072214,0.40429065,0.77232206,1.1403534,1.5083848,1.8746033,1.5809034,1.2853905,0.9898776,0.69436467,0.40066472,0.42967212,0.4604925,0.4894999,0.52032024,0.5493277,0.73424983,0.91917205,1.1040943,1.2908293,1.4757515,1.3796645,1.2853905,1.1893034,1.0950294,1.0007553,0.8557183,0.7106813,0.5656443,0.42060733,0.2755703,0.22662032,0.1794833,0.13234627,0.08520924,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.054388877,0.059827764,0.065266654,0.07070554,0.07433146,0.065266654,0.054388877,0.045324065,0.034446288,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.034446288,0.045324065,0.054388877,0.065266654,0.07433146,0.32270733,0.56927025,0.81764615,1.064209,1.3125849,1.3270886,1.3434052,1.357909,1.3724127,1.3869164,1.1167849,0.8466535,0.57833505,0.30820364,0.038072214,0.67079616,1.3017071,1.9344311,2.5671551,3.199879,2.855416,2.5091403,2.1646774,1.8202144,1.4757515,1.1856775,0.89560354,0.6055295,0.3154555,0.025381476,0.16316663,0.2991388,0.43692398,0.5747091,0.7124943,1.6207886,2.5272698,3.435564,4.3420453,5.2503395,5.660069,6.069799,6.4795284,6.889258,7.3008003,5.957395,4.615803,3.2723975,1.9308052,0.5873999,0.47680917,0.3680314,0.2574407,0.14684997,0.038072214,0.7995165,1.5627737,2.324218,3.0874753,3.8507326,4.401873,4.954827,5.5077806,6.060734,6.6118746,5.5132194,4.4127507,3.3122826,2.2118144,1.1131591,1.1602961,1.2074331,1.2545701,1.3017071,1.3506571,1.1494182,0.9499924,0.7505665,0.5493277,0.34990177,1.0950294,1.840157,2.5852847,3.3304121,4.07554,3.9450066,3.8144734,3.6857529,3.5552197,3.4246864,2.9170568,2.4094272,1.9017978,1.3941683,0.8883517,1.2944553,1.7023718,2.1102884,2.518205,2.9243085,3.5425289,4.160749,4.7771564,5.3953767,6.011784,5.424384,4.836984,4.249584,3.6621845,3.0747845,2.7502642,2.4257438,2.0994108,1.7748904,1.4503701,1.357909,1.2654479,1.1729867,1.0805258,0.9880646,1.2853905,1.5827163,1.8800422,2.1773682,2.474694,1.9797552,1.4848163,0.9898776,0.4949388,0.0,0.27738327,0.55476654,0.8321498,1.1095331,1.3869164,1.1095331,0.8321498,0.55476654,0.27738327,0.0,0.50219065,1.0043813,1.5083848,2.0105755,2.5127661,2.3024626,2.0921588,1.8818551,1.6733645,1.4630609,1.2980812,1.1331016,0.968122,0.8031424,0.63816285,1.0043813,1.3724127,1.7404441,2.1066625,2.474694,1.9942589,1.5156367,1.0352017,0.55476654,0.07433146,0.11240368,0.15047589,0.18673515,0.22480737,0.26287958,0.32995918,0.39703882,0.46411842,0.533011,0.6000906,1.2726997,1.9453088,2.617918,3.290527,3.9631362,4.1299286,4.2967215,4.465327,4.632119,4.800725,5.480586,6.1604466,6.8403077,7.520169,8.200029,8.116633,8.03505,7.951654,7.8700705,7.7866745,7.6942134,7.6017523,7.509291,7.41683,7.324369,7.2554765,7.1847706,7.115878,7.0451727,6.9744673,6.740595,6.5049095,6.2692246,6.035352,5.7996674,5.569421,5.3391747,5.1107416,4.880495,4.650249,5.337362,6.0244746,6.7134004,7.400513,8.087626,7.3406854,6.591932,5.844991,5.0980506,4.349297,4.2477713,4.1444325,4.0429068,3.9395678,3.8380418,4.309412,4.782595,5.2557783,5.727149,6.200332,5.3446136,4.4907084,3.63499,2.7792716,1.9253663,1.7676386,1.6099107,1.452183,1.2944553,1.1367276,0.92823684,0.7179332,0.5076295,0.29732585,0.0870222,0.16316663,0.2374981,0.31182957,0.387974,0.46230546,0.5982776,0.7324369,0.8684091,1.0025684,1.1367276,0.99712944,0.8575313,0.7179332,0.57833505,0.43692398,0.4224203,0.40791658,0.39159992,0.3770962,0.36259252,0.70524246,1.0478923,1.3905423,1.7331922,2.0758421,1.9199274,1.7658255,1.6099107,1.455809,1.2998942,1.3742256,1.4503701,1.5247015,1.6008459,1.6751775,1.7531348,1.8292793,1.9072367,1.9851941,2.0631514,2.427557,2.7919624,3.1581807,3.5225863,3.8869917,3.720199,3.5515938,3.3848011,3.2180085,3.049403,3.2180085,3.3848011,3.5534067,3.720199,3.8869917,4.255023,4.6230545,4.989273,5.3573046,5.7253356,6.115123,6.5049095,6.8946967,7.2844834,7.6742706,5.9374523,5.859495,5.7833505,5.7053933,5.6274357,5.5494785,5.2068286,4.8641787,4.5233417,4.1806917,3.8380418,3.7401419,3.6422417,3.5443418,3.4482548,3.350355,3.3594196,3.3702974,3.3793623,3.39024,3.3993049,3.5969179,3.7945306,3.9921436,4.1897564,4.3873696,4.744523,5.101677,5.4606433,5.8177967,6.1749506,6.552047,6.929143,7.308052,7.6851482,8.062244,8.147454,8.232663,8.317872,8.403082,8.488291,7.8646317,7.2427855,6.6191263,5.99728,5.375434,6.5955577,7.8156815,9.035806,10.254116,11.47424,11.084454,10.694666,10.304879,9.915092,9.525306,9.808127,10.089137,10.371959,10.654781,10.937603,10.906783,10.877775,10.846955,10.817947,10.7871275,10.239613,9.692098,9.144584,8.597069,8.049554,7.957093,7.8646317,7.7721705,7.6797094,7.5872483,7.5256076,7.462154,7.400513,7.3370595,7.2754188,7.309865,7.344311,7.380571,7.415017,7.4494634,7.0469856,6.644508,6.24203,5.8395524,5.4370747,5.3246713,5.2122674,5.0998635,4.98746,4.8750563,4.409125,3.9450066,3.4808881,3.0149567,2.5508385,2.6976883,2.8445382,2.9932013,3.1400511,3.2869012,2.9641938,2.6432993,2.3205922,1.9978848,1.6751775,1.551896,1.4304274,1.3071461,1.1856775,1.062396,1.0225109,0.9826257,0.94274056,0.90285534,0.8629702,0.7197462,0.57833505,0.43511102,0.291887,0.15047589,0.49312583,0.83577573,1.1766127,1.5192627,1.8619126,2.864481,3.8670492,4.8696175,5.8721857,6.874754,6.009971,5.145188,4.2804046,3.4156215,2.5508385,4.0030212,5.4552045,6.9073873,8.3595705,9.811753,9.63227,9.452786,9.273304,9.092008,8.912524,9.498111,10.081885,10.667472,11.253058,11.836833,10.167094,8.497355,6.827617,5.1578784,3.48814,2.9950142,2.5018883,2.0105755,1.5174497,1.0243238,1.2998942,1.5754645,1.8492218,2.124792,2.4003625,2.514579,2.6306088,2.7448254,2.8608549,2.9750717,2.902553,2.8300345,2.7575161,2.6849976,2.612479,4.478018,6.341743,8.207282,10.07282,11.938358,9.89515,7.851941,5.810545,3.7673361,1.7241274,1.5120108,1.2998942,1.0877775,0.87566096,0.66173136,0.7179332,0.77232206,0.82671094,0.88291276,0.93730164,0.7505665,0.5620184,0.37528324,0.18673515,0.0,0.06707962,0.13415924,0.2030518,0.27013144,0.33721104,0.27013144,0.2030518,0.13415924,0.06707962,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.25018883,0.42423326,0.6000906,0.774135,0.9499924,0.99531645,1.0406405,1.0841516,1.1294757,1.1747998,1.1095331,1.0442665,0.9808127,0.9155461,0.85027945,1.3905423,1.9308052,2.469255,3.009518,3.5497808,3.5171473,3.484514,3.4518807,3.4192474,3.386614,3.0149567,2.6432993,2.269829,1.8981718,1.5247015,1.4594349,1.3941683,1.3307146,1.2654479,1.2001812,1.1929294,1.1856775,1.1766127,1.1693609,1.162109,1.2491312,1.3379664,1.4249886,1.5120108,1.6008459,1.4141108,1.2291887,1.0442665,0.85934424,0.6744221,0.6544795,0.6345369,0.61459434,0.5946517,0.5747091,0.5094425,0.44417584,0.38072214,0.3154555,0.25018883,0.42967212,0.6091554,0.7904517,0.969935,1.1494182,0.9318628,0.71430725,0.49675176,0.27919623,0.06164073,0.059827764,0.058014803,0.054388877,0.052575916,0.05076295,0.04169814,0.034446288,0.027194439,0.01994259,0.012690738,0.01994259,0.027194439,0.034446288,0.04169814,0.05076295,0.47680917,0.90466833,1.3325275,1.7603867,2.1882458,1.8528478,1.5174497,1.1820517,0.8466535,0.51306844,0.46411842,0.4169814,0.36984438,0.32270733,0.2755703,0.3680314,0.4604925,0.5529536,0.64541465,0.73787576,0.69073874,0.6417888,0.5946517,0.5475147,0.50037766,0.42785916,0.35534066,0.28282216,0.21030366,0.13778515,0.11965553,0.10333887,0.08520924,0.06707962,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.027194439,0.030820364,0.032633327,0.034446288,0.038072214,0.032633327,0.027194439,0.02175555,0.018129626,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.018129626,0.02175555,0.027194439,0.032633327,0.038072214,0.38072214,0.72337204,1.064209,1.4068589,1.7495089,1.7694515,1.789394,1.8093367,1.8292793,1.8492218,1.4902552,1.1294757,0.7705091,0.40972954,0.05076295,0.36077955,0.67079616,0.9808127,1.2908293,1.6008459,1.4268016,1.2545701,1.0823387,0.9101072,0.73787576,0.59283876,0.44780177,0.30276474,0.15772775,0.012690738,0.19942589,0.387974,0.5747091,0.76325727,0.9499924,2.1592383,3.3702974,4.5795436,5.7906027,6.9998484,7.2047133,7.409578,7.614443,7.819308,8.024173,6.53573,5.045475,3.5552197,2.0649643,0.5747091,0.46955732,0.36440548,0.25925365,0.15410182,0.05076295,1.062396,2.0758421,3.0874753,4.100921,5.1125546,5.032784,4.953014,4.8732433,4.7916603,4.7118897,4.0501585,3.386614,2.7248828,2.0631514,1.3996071,1.4793775,1.5591478,1.6407311,1.7205015,1.8002719,1.5247015,1.2491312,0.97537386,0.69980353,0.42423326,1.3851035,2.3441606,3.3050308,4.265901,5.224958,4.572292,3.919625,3.2669585,2.6142921,1.9616255,1.6642996,1.3669738,1.0696479,0.77232206,0.4749962,0.97174793,1.4703126,1.9670644,2.465629,2.962381,3.4518807,3.9431937,4.4326935,4.9221935,5.411693,4.688321,3.9631362,3.2379513,2.5127661,1.7875811,1.5754645,1.3633479,1.1494182,0.93730164,0.72518504,0.79770356,0.87022203,0.94274056,1.015259,1.0877775,1.4920682,1.8981718,2.3024626,2.7067533,3.1128569,2.4891977,1.8673514,1.2455053,0.62184614,0.0,0.36984438,0.73968875,1.1095331,1.4793775,1.8492218,1.4793775,1.1095331,0.73968875,0.36984438,0.0,0.67079616,1.3397794,2.0105755,2.6795588,3.350355,3.0693457,2.7901495,2.5091403,2.229944,1.9507477,1.7295663,1.5101979,1.2908293,1.0696479,0.85027945,1.3397794,1.8292793,2.3205922,2.810092,3.299592,2.659616,2.0196402,1.3796645,0.73968875,0.099712946,0.15047589,0.19942589,0.25018883,0.2991388,0.34990177,0.41516843,0.48043507,0.54570174,0.6091554,0.6744221,1.4431182,2.2100015,2.9768846,3.7455807,4.512464,4.702825,4.893186,5.081734,5.272095,5.462456,5.8776245,6.2927933,6.7079616,7.12313,7.5382986,7.703278,7.8682575,8.033237,8.198216,8.363196,8.122072,7.8827615,7.6416373,7.402326,7.1630154,7.1031876,7.0433598,6.981719,6.921891,6.8620634,6.882006,6.9019485,6.921891,6.9418335,6.9617763,6.484967,6.008158,5.529536,5.0527267,4.574105,5.7869763,6.9998484,8.212721,9.425592,10.636651,9.157274,7.6778965,6.1967063,4.7173285,3.2379513,3.004079,2.7720199,2.5399606,2.3079014,2.0758421,2.9932013,3.9105604,4.8279195,5.7452784,6.6626377,5.7597823,4.856927,3.9540713,3.053029,2.1501737,1.889107,1.6298534,1.3705997,1.1095331,0.85027945,0.69436467,0.5402629,0.38434806,0.23024625,0.07433146,0.12509441,0.17585737,0.22480737,0.2755703,0.3245203,0.5058166,0.6852999,0.86478317,1.0442665,1.2255627,1.0424535,0.85934424,0.678048,0.4949388,0.31182957,0.31726846,0.32270733,0.32814622,0.33177215,0.33721104,0.61459434,0.8919776,1.1693609,1.4467441,1.7241274,1.696933,1.6697385,1.6425442,1.6153497,1.5881553,1.5754645,1.5627737,1.550083,1.5373923,1.5247015,1.5700256,1.6153497,1.6606737,1.7041848,1.7495089,2.2444477,2.7393866,3.2343252,3.729264,4.2242026,4.0846047,3.9450066,3.8054085,3.6658103,3.5243993,3.727451,3.930503,4.1317415,4.3347936,4.537845,4.9657044,5.391751,5.81961,6.247469,6.6753283,7.119504,7.5654926,8.009668,8.455658,8.899834,7.124943,6.787732,6.450521,6.11331,5.774286,5.4370747,5.1741953,4.9131284,4.650249,4.3873696,4.12449,4.024777,3.925064,3.825351,3.7256382,3.6241121,3.5008307,3.3757362,3.2506418,3.1255474,3.000453,3.199879,3.3993049,3.6005437,3.7999697,3.9993954,4.4381323,4.8750563,5.3119802,5.750717,6.187641,6.6118746,7.037921,7.462154,7.8882003,8.312433,8.437528,8.562622,8.6877165,8.812811,8.937905,8.125698,7.311678,6.4994707,5.6872635,4.8750563,6.187641,7.500226,8.812811,10.125396,11.437981,11.137029,10.837891,10.536939,10.2378,9.936848,10.199727,10.462607,10.725487,10.988366,11.249433,11.287505,11.325577,11.361836,11.399909,11.437981,10.738177,10.038374,9.336758,8.636953,7.93715,7.5999393,7.262728,6.925517,6.588306,6.249282,6.450521,6.6499467,6.849373,7.0506115,7.250037,7.3370595,7.4258947,7.512917,7.5999393,7.686961,7.2754188,6.8620634,6.450521,6.037165,5.6256227,5.4008155,5.1741953,4.949388,4.7245803,4.499773,4.12449,3.7492065,3.3757362,3.000453,2.6251698,2.6995013,2.7756457,2.8499773,2.9243085,3.000453,2.6868105,2.374981,2.0631514,1.7495089,1.4376793,1.3125849,1.1874905,1.062396,0.93730164,0.8122072,0.6744221,0.53663695,0.40066472,0.26287958,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.3245203,0.6508536,0.97537386,1.2998942,1.6244144,2.762955,3.8996825,5.038223,6.1749506,7.311678,6.0625467,4.8134155,3.5624714,2.3133402,1.062396,2.8372865,4.612177,6.3870673,8.161958,9.936848,9.550687,9.162713,8.774739,8.386765,8.000604,8.912524,9.824444,10.738177,11.650098,12.562017,10.700105,8.838193,6.9744673,5.1125546,3.2506418,2.762955,2.275268,1.7875811,1.2998942,0.8122072,0.9880646,1.162109,1.3379664,1.5120108,1.6878681,1.7621996,1.8383441,1.9126755,1.987007,2.0631514,2.2498865,2.4366217,2.6251698,2.811905,3.000453,5.049101,7.0995617,9.1500225,11.200482,13.24913,11.011934,8.774739,6.5375433,4.3003473,2.0631514,1.7132497,1.3633479,1.0116332,0.66173136,0.31182957,0.25018883,0.18673515,0.12509441,0.06164073,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.774135,1.4866294,2.1991236,2.911618,3.6241121,3.5117085,3.3993049,3.2869012,3.1744974,3.0620937,2.5744069,2.08672,1.6008459,1.1131591,0.62547207,0.774135,0.9246109,1.0750868,1.2255627,1.3742256,1.3869164,1.3996071,1.4122978,1.4249886,1.4376793,1.550083,1.6624867,1.7748904,1.887294,1.9996977,1.7495089,1.49932,1.2491312,1.0007553,0.7505665,0.73787576,0.72518504,0.7124943,0.69980353,0.6871128,0.61278135,0.53663695,0.46230546,0.387974,0.31182957,0.53663695,0.76325727,0.9880646,1.2128719,1.4376793,1.162109,0.8883517,0.61278135,0.33721104,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.5493277,1.0370146,1.5247015,2.0123885,2.5000753,2.124792,1.7495089,1.3742256,1.0007553,0.62547207,0.50037766,0.37528324,0.25018883,0.12509441,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.43692398,0.87566096,1.3125849,1.7495089,2.1882458,2.2118144,2.2371957,2.2625773,2.2879589,2.3133402,1.8619126,1.4122978,0.96268314,0.51306844,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.2374981,0.4749962,0.7124943,0.9499924,1.1874905,2.6995013,4.213325,5.7253356,7.2373466,8.749357,8.749357,8.749357,8.749357,8.749357,8.749357,7.112252,5.475147,3.8380418,2.1991236,0.5620184,0.46230546,0.36259252,0.26287958,0.16316663,0.06164073,1.3252757,2.5870976,3.8507326,5.1125546,6.3743763,5.661882,4.949388,4.2368937,3.5243993,2.811905,2.5870976,2.3622901,2.137483,1.9126755,1.6878681,1.8002719,1.9126755,2.0250793,2.137483,2.2498865,1.8999848,1.550083,1.2001812,0.85027945,0.50037766,1.6751775,2.8499773,4.024777,5.199577,6.3743763,5.199577,4.024777,2.8499773,1.6751775,0.50037766,0.41335547,0.3245203,0.2374981,0.15047589,0.06164073,0.6508536,1.2382535,1.8256533,2.4130533,3.000453,3.3630457,3.7256382,4.0882306,4.4508233,4.8116026,3.9504454,3.0874753,2.2245052,1.3633479,0.50037766,0.40066472,0.2991388,0.19942589,0.099712946,0.0,0.2374981,0.4749962,0.7124943,0.9499924,1.1874905,1.7005589,2.2118144,2.7248828,3.2379513,3.7492065,3.000453,2.2498865,1.49932,0.7505665,0.0,0.46230546,0.9246109,1.3869164,1.8492218,2.3133402,1.8492218,1.3869164,0.9246109,0.46230546,0.0,0.8375887,1.6751775,2.5127661,3.350355,4.1879435,3.8380418,3.48814,3.1382382,2.7883365,2.4366217,2.1628644,1.887294,1.6117238,1.3379664,1.062396,1.6751775,2.2879589,2.9007401,3.5117085,4.12449,3.3249733,2.525457,1.7241274,0.9246109,0.12509441,0.18673515,0.25018883,0.31182957,0.37528324,0.43692398,0.50037766,0.5620184,0.62547207,0.6871128,0.7505665,1.6117238,2.474694,3.3376641,4.2006345,5.0617914,5.275721,5.487838,5.6999545,5.9120708,6.1241875,6.2746634,6.4251394,6.5756154,6.7242785,6.874754,7.28811,7.699652,8.113008,8.52455,8.937905,8.549932,8.161958,7.7757964,7.3878226,6.9998484,6.9508986,6.9001355,6.849373,6.8004227,6.7496595,7.02523,7.3008003,7.574558,7.850128,8.125698,7.400513,6.6753283,5.9501433,5.224958,4.499773,6.2384043,7.9752226,9.712041,11.450671,13.1874895,10.975676,8.762048,6.550234,4.3384194,2.124792,1.7621996,1.3996071,1.0370146,0.6744221,0.31182957,1.6751775,3.0367124,4.40006,5.7615952,7.124943,6.1749506,5.224958,4.274966,3.3249733,2.374981,2.0123885,1.649796,1.2872034,0.9246109,0.5620184,0.46230546,0.36259252,0.26287958,0.16316663,0.06164073,0.0870222,0.11240368,0.13778515,0.16316663,0.18673515,0.41335547,0.63816285,0.8629702,1.0877775,1.3125849,1.0877775,0.8629702,0.63816285,0.41335547,0.18673515,0.21211663,0.2374981,0.26287958,0.28826106,0.31182957,0.52575916,0.73787576,0.9499924,1.162109,1.3742256,1.4757515,1.5754645,1.6751775,1.7748904,1.8746033,1.7748904,1.6751775,1.5754645,1.4757515,1.3742256,1.3869164,1.3996071,1.4122978,1.4249886,1.4376793,2.0631514,2.6868105,3.3122826,3.9377546,4.5632267,4.4508233,4.3366065,4.2242026,4.1117992,3.9993954,4.2368937,4.4743915,4.7118897,4.949388,5.186886,5.674573,6.16226,6.6499467,7.137634,7.6253204,8.125698,8.624263,9.12464,9.625018,10.125396,8.450218,8.05318,7.654328,7.2572894,6.8602505,6.4632115,6.115123,5.767034,5.4207582,5.0726695,4.7245803,4.5777307,4.4308805,4.2822175,4.135368,3.9867048,3.8126602,3.636803,3.4627585,3.2869012,3.1128569,3.3159087,3.5171473,3.720199,3.923251,4.12449,4.507025,4.88956,5.272095,5.65463,6.037165,6.247469,6.4577727,6.6680765,6.876567,7.0868707,7.3298078,7.572745,7.8156815,8.056806,8.299743,7.705091,7.1104393,6.5157876,5.919323,5.3246713,6.3653116,7.404139,8.444779,9.48542,10.524248,10.274059,10.025683,9.775495,9.525306,9.275117,9.510801,9.744674,9.980359,10.2142315,10.449916,10.468046,10.484363,10.502492,10.520622,10.536939,9.967669,9.396585,8.827314,8.258044,7.686961,7.3769445,7.066928,6.7569118,6.446895,6.1368785,6.3344913,6.532104,6.7297173,6.92733,7.124943,7.170267,7.215591,7.2591023,7.304426,7.3497505,7.0071006,6.6644506,6.3218007,5.979151,5.638314,5.2630305,4.8877473,4.512464,4.137181,3.7618973,3.435564,3.1074178,2.7792716,2.4529383,2.124792,2.1900587,2.2553256,2.3205922,2.3858588,2.4493124,2.1918716,1.9344311,1.6769904,1.4195497,1.162109,1.062396,0.96268314,0.8629702,0.76325727,0.66173136,0.5493277,0.43692398,0.3245203,0.21211663,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.25925365,0.52032024,0.7795739,1.0406405,1.2998942,2.2245052,3.149116,4.07554,5.0001507,5.924762,4.985647,4.0447197,3.105605,2.1646774,1.2255627,2.9152439,4.604925,6.294606,7.9842873,9.675781,9.119202,8.564435,8.009668,7.454902,6.9001355,7.6325727,8.365009,9.097446,9.829884,10.56232,8.970539,7.3769445,5.7851634,4.1915693,2.5997884,2.2118144,1.8256533,1.4376793,1.0497054,0.66173136,1.0098201,1.357909,1.7041848,2.0522738,2.4003625,2.3604772,2.3205922,2.280707,2.2408218,2.1991236,2.427557,2.6541772,2.8826106,3.1092308,3.3376641,4.992899,6.6481338,8.303369,9.956791,11.612025,9.755551,7.897265,6.0407915,4.1825047,2.324218,1.9996977,1.6751775,1.3506571,1.0243238,0.69980353,0.56020546,0.42060733,0.27919623,0.13959812,0.0,0.058014803,0.11421664,0.17223145,0.23024625,0.28826106,0.31726846,0.3480888,0.3770962,0.40791658,0.43692398,0.36077955,0.28282216,0.20486477,0.12690738,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.045324065,0.09064813,0.13415924,0.1794833,0.22480737,0.43692398,0.6508536,0.8629702,1.0750868,1.2872034,1.1856775,1.0823387,0.9808127,0.8774739,0.775948,1.4159238,2.0558996,2.6958754,3.3358512,3.975827,3.8597972,3.7455807,3.6295512,3.5153344,3.3993049,2.8771715,2.3550384,1.8329052,1.310772,0.7868258,0.86478317,0.94274056,1.020698,1.0968424,1.1747998,1.1693609,1.1657349,1.1602961,1.1548572,1.1494182,1.2491312,1.3506571,1.4503701,1.550083,1.649796,1.452183,1.2545701,1.0569572,0.85934424,0.66173136,0.6417888,0.62184614,0.60190356,0.581961,0.5620184,0.50037766,0.43692398,0.37528324,0.31182957,0.25018883,0.42967212,0.6091554,0.7904517,0.969935,1.1494182,0.9554313,0.75963134,0.5656443,0.36984438,0.17585737,0.36440548,0.55476654,0.7451276,0.9354887,1.1258497,0.96268314,0.7995165,0.63816285,0.4749962,0.31182957,0.34990177,0.387974,0.42423326,0.46230546,0.50037766,0.80495536,1.1095331,1.4141108,1.7205015,2.0250793,1.7205015,1.4141108,1.1095331,0.80495536,0.50037766,0.40066472,0.2991388,0.19942589,0.099712946,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.34990177,0.69980353,1.0497054,1.3996071,1.7495089,1.8020848,1.8546607,1.9072367,1.9598125,2.0123885,1.7621996,1.5120108,1.261822,1.0116332,0.76325727,0.67986095,0.5982776,0.5148814,0.43329805,0.34990177,0.30276474,0.25562772,0.20667773,0.15954071,0.11240368,0.40066472,0.6871128,0.97537386,1.261822,1.550083,1.7549478,1.9598125,2.1646774,2.3695421,2.5744069,3.5624714,4.550536,5.5367875,6.5248523,7.512917,7.6724577,7.8319983,7.993352,8.152893,8.312433,6.9073873,5.5023413,4.0972953,2.6922495,1.2872034,1.9652514,2.6432993,3.3195345,3.9975824,4.6756306,4.9584527,5.239462,5.522284,5.805106,6.0879283,5.37906,4.6720047,3.9649491,3.2578938,2.5508385,2.3169663,2.084907,1.8528478,1.6207886,1.3869164,1.5373923,1.6878681,1.8383441,1.987007,2.137483,1.983381,1.8274662,1.6733645,1.5174497,1.3633479,2.2118144,3.0620937,3.9123733,4.762653,5.612932,4.5704784,3.5280252,2.4855716,1.4431182,0.40066472,0.32995918,0.25925365,0.19036107,0.11965553,0.05076295,0.55476654,1.0605831,1.5645868,2.0704033,2.5744069,2.8880494,3.199879,3.5117085,3.825351,4.137181,3.4192474,2.7031271,1.9851941,1.2672608,0.5493277,0.48043507,0.40972954,0.34083697,0.27013144,0.19942589,0.35534066,0.5094425,0.6653573,0.8194591,0.97537386,1.3796645,1.7857682,2.1900587,2.5943494,3.000453,2.4003625,1.8002719,1.2001812,0.6000906,0.0,0.36984438,0.73968875,1.1095331,1.4793775,1.8492218,1.9416829,2.034144,2.128418,2.220879,2.3133402,2.752077,3.1926272,3.633177,4.071914,4.512464,4.2441454,3.97764,3.7093215,3.442816,3.1744974,2.8916752,2.610666,2.327844,2.0450218,1.7621996,2.1900587,2.617918,3.045777,3.4718235,3.8996825,3.159994,2.420305,1.6806163,0.93911463,0.19942589,0.33539808,0.46955732,0.6055295,0.73968875,0.87566096,0.8974165,0.91917205,0.94274056,0.9644961,0.9880646,1.7259403,2.4620032,3.199879,3.9377546,4.6756306,4.8333583,4.989273,5.147001,5.3047285,5.462456,5.612932,5.7615952,5.9120708,6.0625467,6.2130227,6.8094873,7.407765,8.00423,8.602508,9.200785,8.9052725,8.609759,8.314246,8.020547,7.7250338,7.7377243,7.750415,7.763106,7.7757964,7.7866745,8.624263,9.461852,10.29944,11.137029,11.974618,10.370146,8.765674,7.159389,5.5549173,3.9504454,5.2702823,6.590119,7.909956,9.229793,10.549629,8.834567,7.119504,5.4044414,3.6893787,1.9743162,1.9416829,1.9108626,1.8782293,1.845596,1.8129625,2.9732587,4.1317415,5.292038,6.452334,7.61263,6.58468,5.5567303,4.5305934,3.5026438,2.474694,2.077655,1.6806163,1.2817645,0.88472575,0.48768693,0.40066472,0.31182957,0.22480737,0.13778515,0.05076295,0.07070554,0.09064813,0.11059072,0.13053331,0.15047589,0.32995918,0.5094425,0.69073874,0.87022203,1.0497054,0.87022203,0.69073874,0.5094425,0.32995918,0.15047589,0.17041849,0.19036107,0.21030366,0.23024625,0.25018883,0.4405499,0.630911,0.8194591,1.0098201,1.2001812,1.2908293,1.3796645,1.4703126,1.5591478,1.649796,1.6606737,1.6697385,1.6806163,1.6896812,1.7005589,1.69512,1.6896812,1.6842422,1.6806163,1.6751775,2.2371957,2.7992141,3.3630457,3.925064,4.4870825,4.517903,4.5469103,4.5777307,4.606738,4.6375585,4.88956,5.143375,5.3953767,5.6473784,5.89938,6.2801023,6.6608243,7.039734,7.420456,7.799365,8.312433,8.825501,9.336758,9.849826,10.362894,9.775495,9.316814,8.859948,8.403082,7.944402,7.4875355,7.0542374,6.622752,6.189454,5.7579694,5.3246713,5.130684,4.934884,4.7390842,4.5450974,4.349297,4.12449,3.8996825,3.6748753,3.4500678,3.2252605,3.4301252,3.63499,3.8398547,4.0447197,4.249584,4.5777307,4.9058766,5.23221,5.560356,5.8866897,5.883064,5.8776245,5.8721857,5.866747,5.863121,6.2220874,6.582867,6.9418335,7.3026133,7.663393,7.2844834,6.9073873,6.530291,6.153195,5.774286,6.542982,7.309865,8.076748,8.845445,9.612328,9.412902,9.211663,9.012237,8.812811,8.613385,8.820063,9.026741,9.235231,9.441909,9.6504,9.646774,9.644961,9.643148,9.639522,9.637709,9.197159,8.758422,8.317872,7.877322,7.4367723,7.155763,6.872941,6.590119,6.3072968,6.0244746,6.2202744,6.414262,6.6100616,6.8058615,6.9998484,7.0016613,7.0052876,7.0071006,7.0107265,7.0125394,6.740595,6.4668374,6.1948934,5.922949,5.6491914,5.125245,4.599486,4.07554,3.5497808,3.0258346,2.7448254,2.465629,2.18462,1.9054236,1.6244144,1.6806163,1.7350051,1.789394,1.845596,1.8999848,1.696933,1.4956942,1.2926424,1.0895905,0.8883517,0.8122072,0.73787576,0.66173136,0.5873999,0.51306844,0.42423326,0.33721104,0.25018883,0.16316663,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.19579996,0.38978696,0.5855869,0.7795739,0.97537386,1.6878681,2.4003625,3.1128569,3.825351,4.537845,3.9069343,3.2778363,2.6469254,2.0178273,1.3869164,2.9932013,4.597673,6.202145,7.8084297,9.412902,8.689529,7.9679704,7.2445984,6.5230393,5.7996674,6.352621,6.9055743,7.456715,8.009668,8.562622,7.2409725,5.91751,4.59586,3.2723975,1.9507477,1.6624867,1.3742256,1.0877775,0.7995165,0.51306844,1.0333886,1.551896,2.0722163,2.5925364,3.1128569,2.956942,2.8028402,2.6469254,2.4928236,2.3369088,2.6052272,2.8717327,3.1400511,3.4083695,3.6748753,4.934884,6.1948934,7.454902,8.714911,9.97492,8.497355,7.019791,5.542227,4.064662,2.5870976,2.2879589,1.987007,1.6878681,1.3869164,1.0877775,0.87022203,0.6526665,0.43511102,0.21755551,0.0,0.11421664,0.23024625,0.3444629,0.4604925,0.5747091,0.6345369,0.69436467,0.7541924,0.81583315,0.87566096,0.7197462,0.5656443,0.40972954,0.25562772,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0,0.0,0.0,0.0,0.0,0.09064813,0.1794833,0.27013144,0.36077955,0.44961473,0.87566096,1.2998942,1.7241274,2.1501737,2.5744069,2.3568513,2.1392958,1.9217403,1.7041848,1.4866294,2.0540867,2.6233568,3.1908143,3.7582715,4.325729,4.207886,4.0900435,3.972201,3.8543584,3.738329,3.1799364,2.6233568,2.0649643,1.5083848,0.9499924,0.9554313,0.96087015,0.9644961,0.969935,0.97537386,0.95180535,0.9300498,0.90829426,0.88472575,0.8629702,0.9499924,1.0370146,1.1258497,1.2128719,1.2998942,1.1548572,1.0098201,0.86478317,0.7197462,0.5747091,0.5475147,0.52032024,0.49312583,0.46411842,0.43692398,0.387974,0.33721104,0.28826106,0.2374981,0.18673515,0.32270733,0.45686656,0.59283876,0.726998,0.8629702,0.7469406,0.6327239,0.5166943,0.40247768,0.28826106,0.6671702,1.0478923,1.4268016,1.8075237,2.1882458,1.8746033,1.5627737,1.2491312,0.93730164,0.62547207,0.6871128,0.7505665,0.8122072,0.87566096,0.93730164,1.0605831,1.1820517,1.305333,1.4268016,1.550083,1.3143979,1.0805258,0.8448406,0.6091554,0.37528324,0.2991388,0.22480737,0.15047589,0.07433146,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.26287958,0.52575916,0.7868258,1.0497054,1.3125849,1.3923552,1.4721256,1.551896,1.6316663,1.7132497,1.6624867,1.6117238,1.5627737,1.5120108,1.4630609,1.310772,1.1566701,1.0043813,0.8520924,0.69980353,0.6055295,0.5094425,0.41516843,0.3208944,0.22480737,0.7995165,1.3742256,1.9507477,2.525457,3.100166,3.2723975,3.444629,3.6168604,3.7890918,3.9631362,4.4254417,4.8877473,5.3500524,5.812358,6.2746634,6.5955577,6.9146395,7.2355337,7.554615,7.8755093,6.7025228,5.529536,4.358362,3.1853752,2.0123885,3.4681973,4.9221935,6.378002,7.8319983,9.287807,8.589817,7.891826,7.1956487,6.497658,5.7996674,5.0980506,4.3946214,3.6930048,2.9895754,2.2879589,2.0468347,1.8075237,1.5682126,1.3270886,1.0877775,1.2745126,1.4630609,1.649796,1.8383441,2.0250793,2.0649643,2.1048496,2.1447346,2.18462,2.2245052,2.7502642,3.2742105,3.7999697,4.325729,4.8496747,3.9395678,3.0294604,2.1193533,1.209246,0.2991388,0.24837588,0.19579996,0.14322405,0.09064813,0.038072214,0.4604925,0.88291276,1.305333,1.7277533,2.1501737,2.4130533,2.6741197,2.9369993,3.199879,3.4627585,2.8898623,2.3169663,1.745883,1.1729867,0.6000906,0.56020546,0.52032024,0.48043507,0.4405499,0.40066472,0.47318324,0.54570174,0.61822027,0.69073874,0.76325727,1.0605831,1.357909,1.6552348,1.9525607,2.2498865,1.8002719,1.3506571,0.89922947,0.44961473,0.0,0.27738327,0.55476654,0.8321498,1.1095331,1.3869164,2.034144,2.6831846,3.3304121,3.97764,4.6248674,4.666566,4.710077,4.751775,4.795286,4.836984,4.652062,4.4671397,4.2822175,4.0972953,3.9123733,3.6222992,3.3322253,3.0421512,2.752077,2.4620032,2.70494,2.9478772,3.1908143,3.4319382,3.6748753,2.9950142,2.3151531,1.6352923,0.9554313,0.2755703,0.48224804,0.69073874,0.8974165,1.1040943,1.3125849,1.2944553,1.2781386,1.260009,1.2418793,1.2255627,1.8383441,2.4493124,3.0620937,3.6748753,4.2876563,4.3891826,4.4925213,4.59586,4.6973863,4.800725,4.949388,5.0998635,5.2503395,5.4008155,5.5494785,6.3326783,7.115878,7.897265,8.680465,9.461852,9.2606125,9.057561,8.854509,8.653271,8.450218,8.52455,8.600695,8.675026,8.749357,8.825501,10.225109,11.624716,13.024323,14.42393,15.825351,13.339779,10.854207,8.370448,5.8848767,3.3993049,4.3021603,5.2050157,6.107871,7.0107265,7.911769,6.695271,5.47696,4.2604623,3.0421512,1.8256533,2.1229792,2.420305,2.7176309,3.0149567,3.3122826,4.269527,5.2267714,6.185828,7.1430726,8.100317,6.9944096,5.8903155,4.784408,3.680314,2.5744069,2.1429217,1.7096237,1.2781386,0.8448406,0.41335547,0.33721104,0.26287958,0.18673515,0.11240368,0.038072214,0.052575916,0.06707962,0.08339628,0.09789998,0.11240368,0.24837588,0.3825351,0.5166943,0.6526665,0.7868258,0.6526665,0.5166943,0.3825351,0.24837588,0.11240368,0.12690738,0.14322405,0.15772775,0.17223145,0.18673515,0.35534066,0.52213323,0.69073874,0.8575313,1.0243238,1.1059072,1.1856775,1.2654479,1.3452182,1.4249886,1.5446441,1.6642996,1.7857682,1.9054236,2.0250793,2.0033236,1.9797552,1.9579996,1.9344311,1.9126755,2.4130533,2.913431,3.4119956,3.9123733,4.4127507,4.5849824,4.7572136,4.9294453,5.101677,5.275721,5.542227,5.810545,6.0770507,6.345369,6.6118746,6.885632,7.157576,7.4295206,7.703278,7.9752226,8.499168,9.024928,9.550687,10.074633,10.600392,11.10077,10.582263,10.065568,9.547061,9.030367,8.511859,7.995165,7.476658,6.9599633,6.4432693,5.924762,5.6818247,5.4407005,5.197764,4.954827,4.7118897,4.4381323,4.162562,3.8869917,3.6132345,3.3376641,3.5443418,3.7528327,3.9595103,4.168001,4.3746786,4.646623,4.9203806,5.1923246,5.464269,5.7380266,5.516845,5.297477,5.0781083,4.856927,4.6375585,5.1143675,5.5929894,6.069799,6.546608,7.02523,6.8656893,6.7043357,6.544795,6.3852544,6.2257137,6.720652,7.215591,7.71053,8.205468,8.700407,8.549932,8.399456,8.2507925,8.100317,7.949841,8.129324,8.31062,8.490104,8.669587,8.849071,8.827314,8.805559,8.781991,8.760235,8.736667,8.42665,8.116633,7.806617,7.4966,7.1883965,6.932769,6.677141,6.4233265,6.167699,5.9120708,6.104245,6.298232,6.490406,6.68258,6.874754,6.834869,6.794984,6.755099,6.7152133,6.6753283,6.472276,6.2692246,6.0679855,5.864934,5.661882,4.98746,4.313038,3.636803,2.962381,2.2879589,2.0540867,1.8220274,1.5899682,1.357909,1.1258497,1.1693609,1.214685,1.260009,1.305333,1.3506571,1.2019942,1.0551442,0.90829426,0.75963134,0.61278135,0.5620184,0.51306844,0.46230546,0.41335547,0.36259252,0.2991388,0.2374981,0.17585737,0.11240368,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.13053331,0.25925365,0.38978696,0.52032024,0.6508536,1.1494182,1.649796,2.1501737,2.6505513,3.149116,2.8300345,2.5091403,2.1900587,1.8691645,1.550083,3.0693457,4.590421,6.109684,7.6307597,9.1500225,8.259857,7.369693,6.4795284,5.5893636,4.699199,5.0726695,5.4443264,5.8177967,6.189454,6.5629244,5.5095935,4.458075,3.4047437,2.3532255,1.2998942,1.1131591,0.9246109,0.73787576,0.5493277,0.36259252,1.0551442,1.7476959,2.4402475,3.1327994,3.825351,3.5552197,3.2850883,3.0149567,2.7448254,2.474694,2.7828975,3.0892882,3.397492,3.7056956,4.0120864,4.876869,5.7416525,6.6082487,7.473032,8.337815,7.2391596,6.1423173,5.045475,3.9468195,2.8499773,2.5744069,2.3006494,2.0250793,1.7495089,1.4757515,1.1802386,0.88472575,0.58921283,0.2955129,0.0,0.17223145,0.3444629,0.5166943,0.69073874,0.8629702,0.95180535,1.0424535,1.1331016,1.2219368,1.3125849,1.0805258,0.8466535,0.61459434,0.3825351,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.0,0.0,0.0,0.0,0.0,0.13415924,0.27013144,0.40429065,0.5402629,0.6744221,1.3125849,1.9507477,2.5870976,3.2252605,3.8634233,3.529838,3.198066,2.864481,2.5327086,2.1991236,2.6958754,3.1908143,3.6857529,4.1806917,4.6756306,4.554162,4.4345064,4.314851,4.195195,4.07554,3.482701,2.8898623,2.2970235,1.7041848,1.1131591,1.0442665,0.97718686,0.9101072,0.8430276,0.774135,0.73424983,0.69436467,0.6544795,0.61459434,0.5747091,0.6508536,0.72518504,0.7995165,0.87566096,0.9499924,0.8575313,0.7650702,0.6726091,0.58014804,0.48768693,0.45324063,0.4169814,0.3825351,0.3480888,0.31182957,0.2755703,0.2374981,0.19942589,0.16316663,0.12509441,0.21574254,0.3045777,0.39522585,0.48587397,0.5747091,0.5402629,0.5058166,0.46955732,0.43511102,0.40066472,0.969935,1.5392052,2.1102884,2.6795588,3.2506418,2.7883365,2.324218,1.8619126,1.3996071,0.93730164,1.0243238,1.1131591,1.2001812,1.2872034,1.3742256,1.3143979,1.2545701,1.1947423,1.1349145,1.0750868,0.9101072,0.7451276,0.58014804,0.41516843,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.17585737,0.34990177,0.52575916,0.69980353,0.87566096,0.9826257,1.0895905,1.1983683,1.305333,1.4122978,1.5627737,1.7132497,1.8619126,2.0123885,2.1628644,1.93987,1.7168756,1.4956942,1.2726997,1.0497054,0.90829426,0.7650702,0.62184614,0.48043507,0.33721104,1.2001812,2.0631514,2.9243085,3.787279,4.650249,4.7898474,4.9294453,5.0708566,5.2104545,5.3500524,5.2884116,5.224958,5.163317,5.0998635,5.038223,5.516845,5.99728,6.4777155,6.9581504,7.4367723,6.497658,5.5567303,4.6176157,3.6766882,2.7375734,4.9693303,7.2029004,9.434657,11.668227,13.899984,12.222994,10.546003,8.8672,7.1902094,5.5132194,4.8152285,4.117238,3.4192474,2.72307,2.0250793,1.7767034,1.5301404,1.2817645,1.0352017,0.7868258,1.0116332,1.2382535,1.4630609,1.6878681,1.9126755,2.1483607,2.382233,2.617918,2.8517902,3.0874753,3.2869012,3.48814,3.6875658,3.8869917,4.0882306,3.3104696,2.5327086,1.7549478,0.97718686,0.19942589,0.16497959,0.13053331,0.09427405,0.059827764,0.025381476,0.36440548,0.70524246,1.0442665,1.3851035,1.7241274,1.938057,2.1501737,2.3622901,2.5744069,2.7883365,2.3604772,1.9326181,1.504759,1.0768998,0.6508536,0.6399758,0.629098,0.6200332,0.6091554,0.6000906,0.58921283,0.58014804,0.56927025,0.56020546,0.5493277,0.73968875,0.9300498,1.1204109,1.310772,1.49932,1.2001812,0.89922947,0.6000906,0.2991388,0.0,0.18492219,0.36984438,0.55476654,0.73968875,0.9246109,2.128418,3.3304121,4.5324063,5.7344007,6.9382076,6.582867,6.2275267,5.8721857,5.516845,5.163317,5.0599785,4.95664,4.855114,4.751775,4.650249,4.3529234,4.0555973,3.7582715,3.4591327,3.1618068,3.2198215,3.2778363,3.3358512,3.392053,3.4500678,2.8300345,2.2100015,1.5899682,0.969935,0.34990177,0.630911,0.9101072,1.1893034,1.4703126,1.7495089,1.693307,1.6352923,1.5772774,1.5192627,1.4630609,1.9507477,2.4366217,2.9243085,3.4119956,3.8996825,3.9468195,3.9957695,4.0429068,4.0900435,4.137181,4.2876563,4.4381323,4.5867953,4.7372713,4.8877473,5.8558693,6.8221784,7.7903004,8.758422,9.724731,9.6141405,9.5053625,9.394773,9.284182,9.175404,9.313189,9.449161,9.5869465,9.724731,9.862516,11.825955,13.7875805,15.751019,17.712645,19.67427,16.309412,12.944552,9.579695,6.2148356,2.8499773,3.3358512,3.8199122,4.305786,4.7898474,5.275721,4.554162,3.834416,3.1146698,2.3949237,1.6751775,2.3024626,2.9297476,3.5570326,4.1843176,4.8134155,5.567608,6.3218007,7.077806,7.8319983,8.588004,7.404139,6.2220874,5.040036,3.8579843,2.6741197,2.2081885,1.7404441,1.2726997,0.80495536,0.33721104,0.2755703,0.21211663,0.15047589,0.0870222,0.025381476,0.034446288,0.045324065,0.054388877,0.065266654,0.07433146,0.16497959,0.25562772,0.3444629,0.43511102,0.52575916,0.43511102,0.3444629,0.25562772,0.16497959,0.07433146,0.08520924,0.09427405,0.10515183,0.11421664,0.12509441,0.27013144,0.41516843,0.56020546,0.70524246,0.85027945,0.91917205,0.9898776,1.0605831,1.1294757,1.2001812,1.4304274,1.6606737,1.889107,2.1193533,2.3495996,2.3097143,2.269829,2.229944,2.1900587,2.1501737,2.5870976,3.0258346,3.4627585,3.8996825,4.3366065,4.652062,4.9675174,5.282973,5.5966153,5.9120708,6.1948934,6.4777155,6.7605376,7.0433598,7.324369,7.4893484,7.654328,7.819308,7.9842873,8.149267,8.6877165,9.224354,9.762803,10.29944,10.837891,12.4242325,11.847711,11.269376,10.692853,10.114518,9.537996,8.934279,8.3323765,7.7304726,7.1267557,6.5248523,6.2347784,5.9447045,5.65463,5.3645563,5.0744824,4.749962,4.4254417,4.099108,3.774588,3.4500678,3.6603715,3.870675,4.079166,4.2894692,4.499773,4.7173285,4.934884,5.1524396,5.369995,5.5875506,5.1524396,4.7173285,4.2822175,3.8471067,3.4119956,4.006647,4.603112,5.197764,5.7924156,6.3870673,6.445082,6.5030966,6.5592985,6.6173134,6.6753283,6.8983226,7.119504,7.3424983,7.5654926,7.7866745,7.686961,7.5872483,7.4875355,7.3878226,7.28811,7.440398,7.592687,7.744976,7.897265,8.049554,8.007855,7.9643445,7.9226465,7.8791356,7.837437,7.6579537,7.476658,7.2971745,7.117691,6.9382076,6.7097745,6.4831543,6.2547207,6.0281005,5.7996674,5.9900284,6.1803894,6.3707504,6.5592985,6.7496595,6.6680765,6.58468,6.5030966,6.4197006,6.338117,6.205771,6.071612,5.9392653,5.806919,5.674573,4.8496747,4.024777,3.199879,2.374981,1.550083,1.3651608,1.1802386,0.99531645,0.8103943,0.62547207,0.65991837,0.69436467,0.7306239,0.7650702,0.7995165,0.7070554,0.61459434,0.52213323,0.42967212,0.33721104,0.31182957,0.28826106,0.26287958,0.2374981,0.21211663,0.17585737,0.13778515,0.099712946,0.06164073,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.065266654,0.13053331,0.19579996,0.25925365,0.3245203,0.61278135,0.89922947,1.1874905,1.4757515,1.7621996,1.7531348,1.742257,1.7331922,1.7223145,1.7132497,3.147303,4.5831695,6.017223,7.453089,8.887142,7.8301854,6.773228,5.714458,4.6575007,3.6005437,3.7927177,3.9848917,4.177066,4.36924,4.5632267,3.780027,2.9968271,2.2154403,1.4322405,0.6508536,0.5620184,0.4749962,0.387974,0.2991388,0.21211663,1.0768998,1.9416829,2.808279,3.673062,4.537845,4.1516843,3.7673361,3.3829882,2.9968271,2.612479,2.960568,3.3068438,3.6549325,4.0030212,4.349297,4.8206677,5.290225,5.7597823,6.2293396,6.70071,5.9827766,5.2648435,4.5469103,3.83079,3.1128569,2.8626678,2.612479,2.3622901,2.1121013,1.8619126,1.4902552,1.1167849,0.7451276,0.37165734,0.0,0.23024625,0.4604925,0.69073874,0.91917205,1.1494182,1.2708868,1.3905423,1.5101979,1.6298534,1.7495089,1.4394923,1.1294757,0.8194591,0.5094425,0.19942589,0.15954071,0.11965553,0.07977036,0.03988518,0.0,0.0,0.0,0.0,0.0,0.0,0.1794833,0.36077955,0.5402629,0.7197462,0.89922947,1.7495089,2.5997884,3.4500678,4.3003473,5.1506267,4.702825,4.255023,3.8072214,3.3594196,2.911618,3.3358512,3.7582715,4.1806917,4.603112,5.0255322,4.902251,4.780782,4.6575007,4.5342193,4.4127507,3.785466,3.1581807,2.5290828,1.9017978,1.2745126,1.1349145,0.99531645,0.8557183,0.71430725,0.5747091,0.5166943,0.4604925,0.40247768,0.3444629,0.28826106,0.34990177,0.41335547,0.4749962,0.53663695,0.6000906,0.56020546,0.52032024,0.48043507,0.4405499,0.40066472,0.35715362,0.3154555,0.27194437,0.23024625,0.18673515,0.16316663,0.13778515,0.11240368,0.0870222,0.06164073,0.10696479,0.15228885,0.19761293,0.24293698,0.28826106,0.33177215,0.3770962,0.4224203,0.46774435,0.51306844,1.2726997,2.032331,2.7919624,3.5534067,4.313038,3.7002566,3.0874753,2.474694,1.8619126,1.2491312,1.3633479,1.4757515,1.5881553,1.7005589,1.8129625,1.5700256,1.3270886,1.0841516,0.8430276,0.6000906,0.5058166,0.40972954,0.3154555,0.21936847,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0870222,0.17585737,0.26287958,0.34990177,0.43692398,0.5728962,0.7070554,0.8430276,0.97718686,1.1131591,1.4630609,1.8129625,2.1628644,2.5127661,2.8626678,2.570781,2.277081,1.9851941,1.693307,1.3996071,1.209246,1.020698,0.83033687,0.6399758,0.44961473,1.6008459,2.7502642,3.8996825,5.050914,6.200332,6.3072968,6.414262,6.5230393,6.630004,6.736969,6.149569,5.562169,4.974769,4.3873696,3.7999697,4.439945,5.0799212,5.719897,6.359873,6.9998484,6.2927933,5.5857377,4.876869,4.169814,3.4627585,6.472276,9.481794,12.493125,15.502643,18.512161,15.854358,13.198368,10.540565,7.8827615,5.224958,4.5324063,3.8398547,3.147303,2.4547513,1.7621996,1.5083848,1.2527572,0.99712944,0.7433147,0.48768693,0.7505665,1.0116332,1.2745126,1.5373923,1.8002719,2.229944,2.659616,3.0892882,3.5207734,3.9504454,3.825351,3.7002566,3.5751622,3.4500678,3.3249733,2.6795588,2.034144,1.3905423,0.7451276,0.099712946,0.08339628,0.065266654,0.047137026,0.030820364,0.012690738,0.27013144,0.5275721,0.7850128,1.0424535,1.2998942,1.4630609,1.6244144,1.7875811,1.9507477,2.1121013,1.8292793,1.54827,1.2654479,0.9826257,0.69980353,0.7197462,0.73968875,0.75963134,0.7795739,0.7995165,0.7070554,0.61459434,0.52213323,0.42967212,0.33721104,0.42060733,0.50219065,0.5855869,0.6671702,0.7505665,0.6000906,0.44961473,0.2991388,0.15047589,0.0,0.092461094,0.18492219,0.27738327,0.36984438,0.46230546,2.220879,3.97764,5.7344007,7.4929743,9.249735,8.497355,7.744976,6.9925966,6.240217,5.487838,5.467895,5.4479527,5.42801,5.408067,5.388125,5.081734,4.7771564,4.4725785,4.168001,3.8616104,3.7347028,3.6077955,3.4808881,3.3521678,3.2252605,2.665055,2.1048496,1.5446441,0.98443866,0.42423326,0.7777609,1.1294757,1.4830034,1.8347181,2.1882458,2.0903459,1.9924458,1.8945459,1.7966459,1.7005589,2.0631514,2.4257438,2.7883365,3.149116,3.5117085,3.5044568,3.4972048,3.489953,3.482701,3.4754493,3.6241121,3.774588,3.925064,4.07554,4.2242026,5.377247,6.530291,7.6833353,8.834567,9.987611,9.969481,9.953164,9.935035,9.916905,9.900589,10.100015,10.29944,10.500679,10.700105,10.899531,13.424988,15.950445,18.475903,20.999546,23.525002,19.279043,15.034899,10.790753,6.544795,2.3006494,2.3677292,2.4348087,2.5018883,2.570781,2.6378605,2.4148662,2.1918716,1.9706904,1.7476959,1.5247015,2.4819458,3.43919,4.3982472,5.3554916,6.3127356,6.8656893,7.41683,7.9697833,8.5227375,9.07569,7.8156815,6.5556726,5.295664,4.0356545,2.7756457,2.2716422,1.7694515,1.2672608,0.7650702,0.26287958,0.21211663,0.16316663,0.11240368,0.06164073,0.012690738,0.018129626,0.02175555,0.027194439,0.032633327,0.038072214,0.08339628,0.12690738,0.17223145,0.21755551,0.26287958,0.21755551,0.17223145,0.12690738,0.08339628,0.038072214,0.04169814,0.047137026,0.052575916,0.058014803,0.06164073,0.18492219,0.30820364,0.42967212,0.5529536,0.6744221,0.73424983,0.79589057,0.8557183,0.9155461,0.97537386,1.3143979,1.6552348,1.9942589,2.335096,2.6741197,2.617918,2.5599031,2.5018883,2.4456866,2.3876717,2.762955,3.1382382,3.5117085,3.8869917,4.262275,4.7191415,5.177821,5.634688,6.093367,6.550234,6.8475595,7.1448855,7.4422116,7.7395372,8.036863,8.094878,8.152893,8.210908,8.267109,8.325124,8.874452,9.425592,9.97492,10.524248,11.075388,13.749508,13.113158,12.474996,11.836833,11.200482,10.56232,9.875207,9.188094,8.499168,7.8120556,7.124943,6.787732,6.450521,6.11331,5.774286,5.4370747,5.0617914,4.688321,4.313038,3.9377546,3.5624714,3.774588,3.9867048,4.2006345,4.4127507,4.6248674,4.788034,4.949388,5.1125546,5.275721,5.4370747,4.788034,4.137181,3.48814,2.8372865,2.1882458,2.9007401,3.6132345,4.325729,5.038223,5.750717,6.0244746,6.300045,6.5756154,6.849373,7.124943,7.07418,7.02523,6.9744673,6.925517,6.874754,6.825804,6.775041,6.7242785,6.6753283,6.624565,6.7496595,6.874754,6.9998484,7.124943,7.250037,7.1883965,7.124943,7.063302,6.9998484,6.9382076,6.887445,6.836682,6.787732,6.736969,6.688019,6.48678,6.2873545,6.0879283,5.8866897,5.6872635,5.8758116,6.0625467,6.249282,6.43783,6.624565,6.4994707,6.3743763,6.249282,6.1241875,6.000906,5.9374523,5.8758116,5.812358,5.750717,5.6872635,4.7118897,3.738329,2.762955,1.7875811,0.8122072,0.6744221,0.53663695,0.40066472,0.26287958,0.12509441,0.15047589,0.17585737,0.19942589,0.22480737,0.25018883,0.21211663,0.17585737,0.13778515,0.099712946,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07433146,0.15047589,0.22480737,0.2991388,0.37528324,0.6744221,0.97537386,1.2745126,1.5754645,1.8746033,3.2252605,4.574105,5.924762,7.2754188,8.624263,7.400513,6.1749506,4.949388,3.7256382,2.5000753,2.5127661,2.525457,2.5381477,2.5508385,2.561716,2.0504606,1.5373923,1.0243238,0.51306844,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,1.1004683,2.137483,3.1744974,4.213325,5.2503395,4.749962,4.249584,3.7492065,3.2506418,2.7502642,3.1382382,3.5243993,3.9123733,4.3003473,4.688321,4.762653,4.836984,4.9131284,4.98746,5.0617914,4.7245803,4.3873696,4.0501585,3.7129474,3.3757362,3.149116,2.9243085,2.6995013,2.474694,2.2498865,1.8002719,1.3506571,0.89922947,0.44961473,0.0,0.28826106,0.5747091,0.8629702,1.1494182,1.4376793,1.5881553,1.7368182,1.887294,2.03777,2.1882458,1.8002719,1.4122978,1.0243238,0.63816285,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.0,0.0,0.0,0.0,0.0,0.22480737,0.44961473,0.6744221,0.89922947,1.1258497,2.1882458,3.2506418,4.313038,5.375434,6.43783,5.8758116,5.3119802,4.749962,4.1879435,3.6241121,3.975827,4.325729,4.6756306,5.0255322,5.375434,5.2503395,5.125245,5.0001507,4.8750563,4.749962,4.0882306,3.4246864,2.762955,2.0994108,1.4376793,1.2255627,1.0116332,0.7995165,0.5873999,0.37528324,0.2991388,0.22480737,0.15047589,0.07433146,0.0,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,0.26287958,0.2755703,0.28826106,0.2991388,0.31182957,0.26287958,0.21211663,0.16316663,0.11240368,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.12509441,0.25018883,0.37528324,0.50037766,0.62547207,1.5754645,2.525457,3.4754493,4.4254417,5.375434,4.612177,3.8507326,3.0874753,2.324218,1.5627737,1.7005589,1.8383441,1.9743162,2.1121013,2.2498865,1.8256533,1.3996071,0.97537386,0.5493277,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.16316663,0.3245203,0.48768693,0.6508536,0.8122072,1.3633479,1.9126755,2.4620032,3.0131438,3.5624714,3.199879,2.8372865,2.474694,2.1121013,1.7495089,1.5120108,1.2745126,1.0370146,0.7995165,0.5620184,1.9996977,3.437377,4.8750563,6.3127356,7.750415,7.8247466,7.900891,7.9752226,8.049554,8.125698,7.0125394,5.89938,4.788034,3.6748753,2.561716,3.3630457,4.162562,4.9620786,5.763408,6.5629244,6.0879283,5.612932,5.137936,4.6629395,4.1879435,7.9752226,11.762501,15.54978,19.337059,23.124338,19.487535,15.850732,12.212116,8.575313,4.936697,4.249584,3.5624714,2.8753586,2.1882458,1.49932,1.2382535,0.97537386,0.7124943,0.44961473,0.18673515,0.48768693,0.7868258,1.0877775,1.3869164,1.6878681,2.3133402,2.9369993,3.5624714,4.1879435,4.8116026,4.361988,3.9123733,3.4627585,3.0131438,2.561716,2.0504606,1.5373923,1.0243238,0.51306844,0.0,0.0,0.0,0.0,0.0,0.0,0.17585737,0.34990177,0.52575916,0.69980353,0.87566096,0.9880646,1.1004683,1.2128719,1.3252757,1.4376793,1.2998942,1.162109,1.0243238,0.8883517,0.7505665,0.7995165,0.85027945,0.89922947,0.9499924,1.0007553,0.824898,0.6508536,0.4749962,0.2991388,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.3133402,4.6248674,6.9382076,9.249735,11.563075,10.411844,9.262425,8.113008,6.9617763,5.812358,5.8758116,5.9374523,6.000906,6.0625467,6.1241875,5.812358,5.5005283,5.186886,4.8750563,4.5632267,4.249584,3.9377546,3.6241121,3.3122826,3.000453,2.5000753,1.9996977,1.49932,1.0007553,0.50037766,0.9246109,1.3506571,1.7748904,2.1991236,2.6251698,2.4873846,2.3495996,2.2118144,2.0758421,1.938057,2.175555,2.4130533,2.6505513,2.8880494,3.1255474,3.0620937,3.000453,2.9369993,2.8753586,2.811905,2.962381,3.1128569,3.2633326,3.4119956,3.5624714,4.900438,6.2365913,7.574558,8.912524,10.25049,10.324821,10.399154,10.475298,10.549629,10.625773,10.88684,11.14972,11.4126,11.675479,11.938358,15.025834,18.11331,21.200785,24.286448,27.375734,22.25049,17.125244,11.999999,6.874754,1.7495089,1.3996071,1.0497054,0.69980353,0.34990177,0.0,0.2755703,0.5493277,0.824898,1.1004683,1.3742256,2.663242,3.9504454,5.237649,6.5248523,7.8120556,8.161958,8.511859,8.861761,9.211663,9.563377,8.225411,6.887445,5.5494785,4.213325,2.8753586,2.3369088,1.8002719,1.261822,0.72518504,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.099712946,0.19942589,0.2991388,0.40066472,0.50037766,0.5493277,0.6000906,0.6508536,0.69980353,0.7505665,1.2001812,1.649796,2.0994108,2.5508385,3.000453,2.9243085,2.8499773,2.7756457,2.6995013,2.6251698,2.9369993,3.2506418,3.5624714,3.874301,4.1879435,4.788034,5.388125,5.9882154,6.588306,7.1883965,7.500226,7.8120556,8.125698,8.437528,8.749357,8.700407,8.649645,8.600695,8.549932,8.499168,9.063,9.625018,10.1870365,10.750868,11.312886,13.849221,13.044266,12.23931,11.434355,10.629399,9.824444,9.262425,8.700407,8.136576,7.574558,7.0125394,6.9200783,6.827617,6.735156,6.642695,6.550234,6.051669,5.5549173,5.0581656,4.559601,4.062849,4.1480584,4.233268,4.3166637,4.401873,4.4870825,4.6629395,4.836984,5.0128417,5.186886,5.3627434,4.782595,4.2024474,3.6222992,3.0421512,2.4620032,3.0602808,3.6567454,4.255023,4.853301,5.4497657,5.750717,6.049856,6.350808,6.6499467,6.9490857,6.816739,6.684393,6.552047,6.4197006,6.2873545,6.19308,6.096993,6.002719,5.906632,5.812358,5.810545,5.806919,5.805106,5.803293,5.7996674,5.750717,5.6999545,5.6491914,5.600241,5.5494785,5.5567303,5.565795,5.573047,5.580299,5.5875506,5.4044414,5.223145,5.040036,4.856927,4.6756306,4.853301,5.029158,5.2068286,5.384499,5.562169,5.487838,5.411693,5.337362,5.2630305,5.186886,5.1071157,5.027345,4.947575,4.8678045,4.788034,3.9595103,3.1327994,2.3042755,1.4775645,0.6508536,0.5402629,0.42967212,0.3208944,0.21030366,0.099712946,0.11965553,0.13959812,0.15954071,0.1794833,0.19942589,0.17041849,0.13959812,0.11059072,0.07977036,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.18673515,0.37528324,0.5620184,0.7505665,0.93730164,1.1693609,1.403233,1.6352923,1.8673514,2.0994108,3.0602808,4.019338,4.9802084,5.9392653,6.9001355,5.919323,4.940323,3.9595103,2.9805105,1.9996977,2.0105755,2.0196402,2.030518,2.039583,2.0504606,1.6407311,1.2291887,0.8194591,0.40972954,0.0,0.027194439,0.054388877,0.08339628,0.11059072,0.13778515,1.1077201,2.077655,3.04759,4.017525,4.98746,4.554162,4.122677,3.6893787,3.2578938,2.8245957,3.0367124,3.2506418,3.4627585,3.6748753,3.8869917,4.0972953,4.307599,4.517903,4.7282066,4.936697,4.668379,4.3982472,4.1281157,3.8579843,3.587853,3.3376641,3.0874753,2.8372865,2.5870976,2.3369088,1.8782293,1.4177368,0.9572442,0.49675176,0.038072214,0.42967212,0.823085,1.214685,1.6080978,1.9996977,2.2027495,2.4058013,2.6070402,2.810092,3.0131438,2.6723068,2.333283,1.9924458,1.6534219,1.3125849,1.2346275,1.1566701,1.0805258,1.0025684,0.9246109,0.9898776,1.0551442,1.1204109,1.1856775,1.2509441,1.2853905,1.3198367,1.3542831,1.3905423,1.4249886,2.269829,3.1146698,3.9595103,4.804351,5.6491914,5.1578784,4.664753,4.171627,3.680314,3.1871881,3.4101827,3.633177,3.8543584,4.077353,4.3003473,4.2006345,4.099108,3.9993954,3.8996825,3.7999697,3.2705846,2.7393866,2.2100015,1.6806163,1.1494182,0.9808127,0.8103943,0.6399758,0.46955732,0.2991388,0.23931105,0.1794833,0.11965553,0.059827764,0.0,0.03988518,0.07977036,0.11965553,0.15954071,0.19942589,0.21030366,0.21936847,0.23024625,0.23931105,0.25018883,0.21030366,0.17041849,0.13053331,0.09064813,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.10333887,0.20486477,0.30820364,0.40972954,0.51306844,1.2726997,2.032331,2.7919624,3.5515938,4.313038,3.7020695,3.092914,2.4819458,1.8727903,1.261822,1.3705997,1.4775645,1.5845293,1.693307,1.8002719,1.4594349,1.1204109,0.7795739,0.4405499,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.09064813,0.06707962,0.045324065,0.02175555,0.0,0.092461094,0.18492219,0.27738327,0.36984438,0.46230546,0.5420758,0.62184614,0.7016165,0.78319985,0.8629702,1.4467441,2.032331,2.617918,3.2016919,3.787279,3.4681973,3.147303,2.8282216,2.5073273,2.1882458,2.7393866,3.29234,3.8452935,4.3982472,4.949388,5.5984282,6.245656,6.892884,7.5401115,8.187339,7.8682575,7.5473633,7.228282,6.9073873,6.588306,6.3145485,6.0426044,5.77066,5.4969025,5.224958,5.4352617,5.6455655,5.8558693,6.0643597,6.2746634,6.3616858,6.450521,6.5375433,6.624565,6.7134004,9.285995,11.856775,14.429369,17.001963,19.574556,16.570478,13.564586,10.560507,7.554615,4.550536,3.9830787,3.4156215,2.8481643,2.280707,1.7132497,1.6352923,1.5573349,1.4793775,1.403233,1.3252757,1.4648738,1.6044719,1.745883,1.8854811,2.0250793,2.5018883,2.9805105,3.4573197,3.9341288,4.4127507,4.0030212,3.5932918,3.1817493,2.7720199,2.3622901,2.4094272,2.4583774,2.5055144,2.5526514,2.5997884,2.3767939,2.1556125,1.9326181,1.7096237,1.4884423,1.3452182,1.2019942,1.0605831,0.91735905,0.774135,0.85027945,0.9246109,1.0007553,1.0750868,1.1494182,1.0732739,0.99531645,0.91735905,0.83940166,0.76325727,0.7777609,0.79226464,0.80676836,0.823085,0.8375887,0.69073874,0.5420758,0.39522585,0.24837588,0.099712946,0.07977036,0.059827764,0.03988518,0.01994259,0.0,0.32814622,0.6544795,0.9826257,1.310772,1.6371052,1.5156367,1.3923552,1.2708868,1.1476053,1.0243238,2.7792716,4.5342193,6.2891674,8.044115,9.799063,8.887142,7.9752226,7.063302,6.149569,5.237649,5.7470913,6.258347,6.7677894,7.2772317,7.7884874,7.2554765,6.722465,6.189454,5.658256,5.125245,4.8170414,4.510651,4.2024474,3.8942437,3.587853,3.1074178,2.6269827,2.1483607,1.6679256,1.1874905,1.6751775,2.1628644,2.6505513,3.1382382,3.625925,3.392053,3.159994,2.9279346,2.6958754,2.4620032,2.8282216,3.1926272,3.5570326,3.923251,4.2876563,4.314851,4.3420453,4.36924,4.3982472,4.4254417,4.9294453,5.4352617,5.941078,6.445082,6.9508986,8.488291,10.025683,11.563075,13.100468,14.63786,14.418491,14.19731,13.9779415,13.758573,13.537392,13.397794,13.258195,13.116784,12.977186,12.837588,14.995013,17.15244,19.309864,21.46729,23.624716,19.407764,15.190813,10.97205,6.755099,2.5381477,2.0595255,1.5827163,1.1059072,0.62728506,0.15047589,0.43329805,0.71430725,0.99712944,1.2799516,1.5627737,2.6142921,3.6676233,4.7191415,5.772473,6.825804,7.3479376,7.8700705,8.392203,8.914337,9.438283,8.080374,6.722465,5.3645563,4.00846,2.6505513,2.1501737,1.649796,1.1494182,0.6508536,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07977036,0.15954071,0.23931105,0.3208944,0.40066472,0.44780177,0.4949388,0.5420758,0.58921283,0.63816285,0.99531645,1.35247,1.7096237,2.0667772,2.4257438,2.467442,2.5091403,2.5526514,2.5943494,2.6378605,3.092914,3.5479677,4.0030212,4.458075,4.9131284,5.315606,5.718084,6.1205616,6.5230393,6.925517,7.208339,7.4893484,7.7721705,8.054993,8.337815,8.519112,8.70222,8.885329,9.066626,9.249735,9.817192,10.384649,10.952107,11.519565,12.087022,13.9507475,12.977186,12.005438,11.0318775,10.060129,9.088382,8.649645,8.212721,7.7757964,7.3370595,6.9001355,7.0524244,7.2047133,7.3570023,7.509291,7.66158,7.0433598,6.4233265,5.803293,5.18326,4.5632267,4.519716,4.478018,4.4345064,4.3928084,4.349297,4.537845,4.7245803,4.9131284,5.0998635,5.2865987,4.7771564,4.267714,3.7582715,3.247016,2.7375734,3.2198215,3.7020695,4.1843176,4.668379,5.1506267,5.475147,5.7996674,6.1241875,6.450521,6.775041,6.5592985,6.345369,6.1296263,5.915697,5.6999545,5.560356,5.4207582,5.279347,5.139749,5.0001507,4.8696175,4.740897,4.610364,4.4798307,4.349297,4.313038,4.274966,4.2368937,4.2006345,4.162562,4.227829,4.2930956,4.358362,4.421816,4.4870825,4.322103,4.157123,3.9921436,3.827164,3.6621845,3.83079,3.9975824,4.164375,4.3329806,4.499773,4.4743915,4.4508233,4.4254417,4.40006,4.3746786,4.2767787,4.1806917,4.082792,3.9848917,3.8869917,3.207131,2.5272698,1.8474089,1.167548,0.48768693,0.40429065,0.32270733,0.23931105,0.15772775,0.07433146,0.09064813,0.10515183,0.11965553,0.13415924,0.15047589,0.12690738,0.10515183,0.08339628,0.059827764,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.2991388,0.6000906,0.89922947,1.2001812,1.49932,1.6642996,1.8292793,1.9942589,2.1592383,2.324218,2.8953013,3.4645715,4.0356545,4.604925,5.1741953,4.439945,3.7056956,2.9696326,2.2353828,1.49932,1.5083848,1.5156367,1.5228885,1.5301404,1.5373923,1.2291887,0.922798,0.61459434,0.30820364,0.0,0.04169814,0.08520924,0.12690738,0.17041849,0.21211663,1.114972,2.0178273,2.9206827,3.8217251,4.7245803,4.360175,3.9957695,3.6295512,3.2651455,2.9007401,2.9369993,2.9750717,3.0131438,3.049403,3.0874753,3.4319382,3.778214,4.122677,4.4671397,4.8116026,4.610364,4.407312,4.2042603,4.0030212,3.7999697,3.5243993,3.2506418,2.9750717,2.6995013,2.4257438,1.9543737,1.4848163,1.015259,0.54570174,0.07433146,0.5728962,1.0696479,1.5682126,2.0649643,2.561716,2.817344,3.0729716,3.3267863,3.5824142,3.8380418,3.5443418,3.2524548,2.960568,2.666868,2.374981,2.269829,2.1646774,2.0595255,1.9543737,1.8492218,1.9797552,2.1102884,2.2408218,2.3695421,2.5000753,2.3441606,2.1900587,2.034144,1.8800422,1.7241274,2.3532255,2.9805105,3.6077955,4.2350807,4.8623657,4.439945,4.017525,3.5951047,3.1726844,2.7502642,2.8445382,2.9406252,3.0348995,3.1291735,3.2252605,3.150929,3.0747845,3.000453,2.9243085,2.8499773,2.4529383,2.0558996,1.6570477,1.260009,0.8629702,0.73424983,0.6073425,0.48043507,0.35171473,0.22480737,0.1794833,0.13415924,0.09064813,0.045324065,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.15772775,0.16497959,0.17223145,0.1794833,0.18673515,0.15772775,0.12690738,0.09789998,0.06707962,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.07977036,0.15954071,0.23931105,0.3208944,0.40066472,0.969935,1.5392052,2.1102884,2.6795588,3.2506418,2.7919624,2.335096,1.8782293,1.4195497,0.96268314,1.0406405,1.1167849,1.1947423,1.2726997,1.3506571,1.0950294,0.83940166,0.5855869,0.32995918,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.045324065,0.09064813,0.13415924,0.1794833,0.22480737,0.1794833,0.13415924,0.09064813,0.045324065,0.0,0.18492219,0.36984438,0.55476654,0.73968875,0.9246109,0.922798,0.91917205,0.91735905,0.9155461,0.9119202,1.5319533,2.1519866,2.7720199,3.392053,4.0120864,3.7347028,3.4573197,3.1799364,2.902553,2.6251698,3.966762,5.3101673,6.6517596,7.995165,9.336758,9.195346,9.052122,8.910711,8.767487,8.624263,7.909956,7.1956487,6.4795284,5.765221,5.050914,5.618371,6.185828,6.7532854,7.320743,7.8882003,7.507478,7.1267557,6.7478466,6.3671246,5.9882154,6.637256,7.28811,7.93715,8.588004,9.237044,10.594954,11.952863,13.310771,14.666867,16.024776,13.651608,11.280253,8.907085,6.53573,4.162562,3.7147603,3.2669585,2.819157,2.373168,1.9253663,2.032331,2.1392958,2.2480736,2.3550384,2.4620032,2.4420607,2.422118,2.4021754,2.382233,2.3622901,2.6922495,3.0222087,3.3521678,3.682127,4.0120864,3.6422417,3.2723975,2.902553,2.5327086,2.1628644,2.770207,3.3775494,3.9848917,4.592234,5.199577,4.7554007,4.309412,3.8652363,3.4192474,2.9750717,2.514579,2.0540867,1.5954071,1.1349145,0.6744221,0.7124943,0.7505665,0.7868258,0.824898,0.8629702,0.8448406,0.82671094,0.8103943,0.79226464,0.774135,0.7541924,0.73424983,0.71430725,0.69436467,0.6744221,0.55476654,0.43511102,0.3154555,0.19579996,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.6544795,1.310772,1.9652514,2.619731,3.2742105,3.0294604,2.7847104,2.5399606,2.2952106,2.0504606,3.247016,4.445384,5.6419396,6.8403077,8.036863,7.362441,6.688019,6.011784,5.337362,4.6629395,5.620184,6.5774283,7.5346723,8.491917,9.449161,8.696781,7.944402,7.192023,6.439643,5.6872635,5.384499,5.081734,4.780782,4.478018,4.175253,3.7147603,3.254268,2.7955883,2.335096,1.8746033,2.4257438,2.9750717,3.5243993,4.07554,4.6248674,4.2967215,3.9703882,3.6422417,3.3140955,2.9877625,3.4808881,3.972201,4.465327,4.95664,5.4497657,5.567608,5.6854506,5.803293,5.919323,6.037165,6.8983226,7.757667,8.617011,9.4781685,10.337513,12.07433,13.812962,15.54978,17.286598,19.025229,18.510347,17.995466,17.480585,16.965704,16.449009,15.906934,15.364858,14.8227825,14.280706,13.736817,14.964193,16.193382,17.420757,18.648132,19.87551,16.565039,13.254569,9.944099,6.635443,3.3249733,2.7194438,2.1157274,1.5101979,0.90466833,0.2991388,0.58921283,0.8792868,1.1693609,1.4594349,1.7495089,2.5671551,3.3848011,4.2024474,5.0200934,5.8377395,6.532104,7.228282,7.9226465,8.617011,9.313189,7.935337,6.5574856,5.179634,3.8017826,2.4257438,1.9616255,1.49932,1.0370146,0.5747091,0.11240368,0.09064813,0.06707962,0.045324065,0.02175555,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.059827764,0.11965553,0.1794833,0.23931105,0.2991388,0.3444629,0.38978696,0.43511102,0.48043507,0.52575916,0.7904517,1.0551442,1.3198367,1.5845293,1.8492218,2.0105755,2.1701162,2.3296568,2.4891977,2.6505513,3.247016,3.8452935,4.441758,5.040036,5.638314,5.8431783,6.0480433,6.2529078,6.4577727,6.6626377,6.9146395,7.166641,7.420456,7.6724577,7.9244595,8.339628,8.754796,9.169965,9.585134,10.000301,10.573197,11.144281,11.717177,12.290073,12.862969,14.05046,12.910107,11.769753,10.629399,9.490859,8.350506,8.036863,7.7250338,7.413204,7.0995617,6.787732,7.1847706,7.5818095,7.9806614,8.3777,8.774739,8.033237,7.2899227,6.546608,5.805106,5.0617914,4.893186,4.7227674,4.552349,4.3819304,4.213325,4.4127507,4.612177,4.8116026,5.0128417,5.2122674,4.7717175,4.3329806,3.8924308,3.4518807,3.0131438,3.3793623,3.7473936,4.115425,4.4816437,4.8496747,5.199577,5.5494785,5.89938,6.249282,6.599184,6.301858,6.004532,5.7072062,5.40988,5.1125546,4.9276323,4.74271,4.557788,4.3728657,4.1879435,3.930503,3.673062,3.4156215,3.1581807,2.9007401,2.8753586,2.8499773,2.8245957,2.7992141,2.7756457,2.8971143,3.0203958,3.141864,3.2651455,3.386614,3.2397642,3.092914,2.9442513,2.7974012,2.6505513,2.808279,2.9641938,3.1219215,3.2796493,3.437377,3.4627585,3.48814,3.5117085,3.53709,3.5624714,3.4482548,3.3322253,3.2180085,3.101979,2.9877625,2.4547513,1.9217403,1.3905423,0.8575313,0.3245203,0.27013144,0.21574254,0.15954071,0.10515183,0.05076295,0.059827764,0.07070554,0.07977036,0.09064813,0.099712946,0.08520924,0.07070554,0.054388877,0.03988518,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.41335547,0.824898,1.2382535,1.649796,2.0631514,2.1592383,2.2571385,2.3550384,2.4529383,2.5508385,2.7303216,2.909805,3.0892882,3.2705846,3.4500678,2.960568,2.469255,1.9797552,1.4902552,1.0007553,1.0043813,1.0098201,1.015259,1.020698,1.0243238,0.8194591,0.61459434,0.40972954,0.20486477,0.0,0.058014803,0.11421664,0.17223145,0.23024625,0.28826106,1.1222239,1.9579996,2.7919624,3.6277382,4.461701,4.164375,3.8670492,3.5697234,3.2723975,2.9750717,2.8372865,2.6995013,2.561716,2.4257438,2.2879589,2.7665808,3.247016,3.727451,4.207886,4.688321,4.552349,4.41819,4.2822175,4.1480584,4.0120864,3.7129474,3.4119956,3.1128569,2.811905,2.5127661,2.032331,1.551896,1.0732739,0.59283876,0.11240368,0.71430725,1.3180238,1.9199274,2.521831,3.1255474,3.4319382,3.7401419,4.0483456,4.3547363,4.6629395,4.41819,4.17344,3.926877,3.682127,3.437377,3.3050308,3.1726844,3.0403383,2.907992,2.7756457,2.9696326,3.1654327,3.3594196,3.5552197,3.7492065,3.4047437,3.0602808,2.715818,2.3695421,2.0250793,2.4348087,2.8445382,3.254268,3.6658103,4.07554,3.7220123,3.3702974,3.0167696,2.665055,2.3133402,2.280707,2.2480736,2.2154403,2.182807,2.1501737,2.0994108,2.0504606,1.9996977,1.9507477,1.8999848,1.6352923,1.3705997,1.1040943,0.83940166,0.5747091,0.4894999,0.40429065,0.3208944,0.23568514,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.10515183,0.11059072,0.11421664,0.11965553,0.12509441,0.10515183,0.08520924,0.065266654,0.045324065,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.058014803,0.11421664,0.17223145,0.23024625,0.28826106,0.6671702,1.0478923,1.4268016,1.8075237,2.1882458,1.8818551,1.5772774,1.2726997,0.968122,0.66173136,0.7106813,0.75781834,0.80495536,0.8520924,0.89922947,0.7306239,0.56020546,0.38978696,0.21936847,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06707962,0.13415924,0.2030518,0.27013144,0.33721104,0.27013144,0.2030518,0.13415924,0.06707962,0.0,0.27738327,0.55476654,0.8321498,1.1095331,1.3869164,1.3017071,1.2183108,1.1331016,1.0478923,0.96268314,1.6171626,2.2716422,2.9279346,3.5824142,4.2368937,4.0030212,3.7673361,3.531651,3.2977788,3.0620937,5.195951,7.327995,9.460039,11.592083,13.72594,12.792264,11.860401,10.926725,9.994863,9.063,7.951654,6.8421206,5.732588,4.6230545,3.5117085,4.9203806,6.3272395,7.7359114,9.142771,10.549629,9.579695,8.609759,7.6398244,6.6698895,5.6999545,6.9128265,8.125698,9.336758,10.549629,11.762501,11.9057255,12.047136,12.19036,12.331772,12.474996,10.734551,8.994107,7.2554765,5.5150323,3.774588,3.4482548,3.1201086,2.7919624,2.465629,2.137483,2.42937,2.72307,3.0149567,3.3068438,3.6005437,3.4192474,3.2397642,3.0602808,2.8807976,2.6995013,2.8826106,3.0657198,3.247016,3.4301252,3.6132345,3.2832751,2.953316,2.6233568,2.2915847,1.9616255,3.1309865,4.2967215,5.464269,6.6318173,7.799365,7.132195,6.4650245,5.7978544,5.130684,4.461701,3.6857529,2.907992,2.1302311,1.35247,0.5747091,0.5747091,0.5747091,0.5747091,0.5747091,0.5747091,0.61822027,0.65991837,0.7016165,0.7451276,0.7868258,0.7324369,0.678048,0.62184614,0.56745726,0.51306844,0.42060733,0.32814622,0.23568514,0.14322405,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.9826257,1.9652514,2.9478772,3.930503,4.9131284,4.5450974,4.177066,3.8108473,3.442816,3.0747845,3.7147603,4.3547363,4.994712,5.634688,6.2746634,5.8377395,5.4008155,4.9620786,4.5251546,4.0882306,5.4932766,6.8983226,8.303369,9.708415,11.111648,10.139899,9.168152,8.194591,7.2228427,6.249282,5.9519563,5.65463,5.3573046,5.0599785,4.762653,4.322103,3.8833659,3.442816,3.002266,2.561716,3.1744974,3.787279,4.40006,5.0128417,5.6256227,5.2032027,4.780782,4.358362,3.9341288,3.5117085,4.1317415,4.751775,5.371808,5.9918413,6.6118746,6.8203654,7.027043,7.2355337,7.4422116,7.650702,8.865387,10.080072,11.294757,12.509441,13.72594,15.662184,17.60024,19.538298,21.474543,23.4126,22.602205,21.791811,20.983229,20.172834,19.36244,18.417887,17.473333,16.526966,15.582414,14.63786,14.935185,15.2325115,15.529838,15.827164,16.124489,13.722314,11.320138,8.917963,6.5157876,4.1117992,3.3793623,2.6469254,1.9144884,1.1820517,0.44961473,0.7469406,1.0442665,1.3434052,1.6407311,1.938057,2.520018,3.101979,3.6857529,4.267714,4.8496747,5.718084,6.58468,7.453089,8.319685,9.188094,7.7903004,6.392506,4.994712,3.5969179,2.1991236,1.7748904,1.3506571,0.9246109,0.50037766,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03988518,0.07977036,0.11965553,0.15954071,0.19942589,0.24293698,0.28463513,0.32814622,0.36984438,0.41335547,0.5855869,0.75781834,0.9300498,1.1022812,1.2745126,1.551896,1.8292793,2.1066625,2.3858588,2.663242,3.4029307,4.1426196,4.882308,5.621997,6.3616858,6.3707504,6.378002,6.3852544,6.392506,6.399758,6.622752,6.8457465,7.066928,7.2899227,7.512917,8.160145,8.807372,9.4546,10.101828,10.750868,11.327391,11.9057255,12.482247,13.060582,13.637105,14.150173,12.843027,11.535881,10.226922,8.919776,7.61263,7.4258947,7.2373466,7.0506115,6.8620634,6.6753283,7.317117,7.9607186,8.602508,9.244296,9.8878975,9.023115,8.158332,7.2917356,6.4269524,5.562169,5.2648435,4.9675174,4.670192,4.3728657,4.07554,4.2876563,4.499773,4.7118897,4.9258194,5.137936,4.7680917,4.3982472,4.02659,3.6567454,3.2869012,3.540716,3.7927177,4.0447197,4.2967215,4.550536,4.9258194,5.2992897,5.674573,6.049856,6.4251394,6.0444174,5.6655083,5.2847857,4.9058766,4.5251546,4.2949085,4.064662,3.834416,3.6041696,3.3757362,2.9895754,2.6052272,2.2190661,1.8347181,1.4503701,1.4376793,1.4249886,1.4122978,1.3996071,1.3869164,1.5682126,1.7476959,1.9271792,2.1066625,2.2879589,2.1574254,2.0268922,1.8981718,1.7676386,1.6371052,1.7857682,1.9326181,2.079468,2.228131,2.374981,2.4493124,2.525457,2.5997884,2.6741197,2.7502642,2.617918,2.4855716,2.3532255,2.220879,2.08672,1.7023718,1.3180238,0.9318628,0.5475147,0.16316663,0.13415924,0.10696479,0.07977036,0.052575916,0.025381476,0.030820364,0.034446288,0.03988518,0.045324065,0.05076295,0.04169814,0.034446288,0.027194439,0.01994259,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.52575916,1.0497054,1.5754645,2.0994108,2.6251698,2.6541772,2.6849976,2.715818,2.7448254,2.7756457,2.565342,2.3550384,2.1447346,1.9344311,1.7241274,1.4793775,1.2346275,0.9898776,0.7451276,0.50037766,0.50219065,0.5058166,0.5076295,0.5094425,0.51306844,0.40972954,0.30820364,0.20486477,0.10333887,0.0,0.072518505,0.14503701,0.21755551,0.29007402,0.36259252,1.1294757,1.8981718,2.665055,3.4319382,4.2006345,3.9703882,3.7401419,3.5098956,3.2796493,3.049403,2.7375734,2.4257438,2.1121013,1.8002719,1.4866294,2.1030366,2.7176309,3.3322253,3.9468195,4.5632267,4.494334,4.4272547,4.360175,4.2930956,4.2242026,3.8996825,3.5751622,3.2506418,2.9243085,2.5997884,2.1102884,1.6207886,1.1294757,0.6399758,0.15047589,0.8575313,1.5645868,2.2716422,2.9805105,3.6875658,4.0483456,4.407312,4.7680917,5.127058,5.487838,5.290225,5.092612,4.894999,4.6973863,4.499773,4.3402324,4.1806917,4.019338,3.8597972,3.7002566,3.9595103,4.220577,4.4798307,4.740897,5.0001507,4.465327,3.930503,3.395679,2.8608549,2.324218,2.518205,2.7103791,2.902553,3.094727,3.2869012,3.005892,2.72307,2.4402475,2.1574254,1.8746033,1.7150626,1.5555218,1.3941683,1.2346275,1.0750868,1.0497054,1.0243238,1.0007553,0.97537386,0.9499924,0.81764615,0.6852999,0.5529536,0.42060733,0.28826106,0.24474995,0.2030518,0.15954071,0.11784257,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.052575916,0.054388877,0.058014803,0.059827764,0.06164073,0.052575916,0.04169814,0.032633327,0.02175555,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.034446288,0.07070554,0.10515183,0.13959812,0.17585737,0.36440548,0.55476654,0.7451276,0.9354887,1.1258497,0.97174793,0.8194591,0.6671702,0.5148814,0.36259252,0.38072214,0.39703882,0.41516843,0.43329805,0.44961473,0.36440548,0.27919623,0.19579996,0.11059072,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.09064813,0.1794833,0.27013144,0.36077955,0.44961473,0.36077955,0.27013144,0.1794833,0.09064813,0.0,0.36984438,0.73968875,1.1095331,1.4793775,1.8492218,1.6824293,1.5156367,1.3470312,1.1802386,1.0116332,1.7023718,2.3931105,3.0820365,3.7727752,4.461701,4.269527,4.077353,3.8851788,3.6930048,3.5008307,6.4233265,9.345822,12.268318,15.190813,18.11331,16.389181,14.666867,12.944552,11.222239,9.499924,7.995165,6.490406,4.985647,3.4790752,1.9743162,4.2223897,6.4704633,8.716724,10.964798,13.212872,11.651911,10.092763,8.531802,6.972654,5.411693,7.1883965,8.963287,10.738177,12.513068,14.287958,13.2146845,12.143224,11.069949,9.9966755,8.925215,7.817495,6.7097745,5.6020546,4.494334,3.386614,3.1799364,2.9732587,2.764768,2.5580902,2.3495996,2.8282216,3.3050308,3.7818398,4.2604623,4.7372713,4.3982472,4.0574102,3.7183862,3.3775494,3.0367124,3.0729716,3.1074178,3.141864,3.1781235,3.2125697,2.9224956,2.6324217,2.3423476,2.0522738,1.7621996,3.489953,5.217706,6.94546,8.673213,10.399154,9.510801,8.620637,7.7304726,6.8403077,5.9501433,4.855114,3.7600844,2.665055,1.5700256,0.4749962,0.43692398,0.40066472,0.36259252,0.3245203,0.28826106,0.38978696,0.49312583,0.5946517,0.6979906,0.7995165,0.7106813,0.6200332,0.5293851,0.4405499,0.34990177,0.28463513,0.21936847,0.15410182,0.09064813,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,1.310772,2.619731,3.930503,5.239462,6.550234,6.060734,5.569421,5.0799212,4.590421,4.100921,4.1825047,4.265901,4.347484,4.4308805,4.512464,4.313038,4.1117992,3.9123733,3.7129474,3.5117085,5.3645563,7.217404,9.070251,10.9230995,12.774135,11.583018,10.390089,9.197159,8.00423,6.813113,6.5194135,6.2275267,5.9356394,5.6419396,5.3500524,4.9294453,4.510651,4.0900435,3.6694362,3.2506418,3.925064,4.599486,5.275721,5.9501433,6.624565,6.107871,5.5893636,5.0726695,4.554162,4.0374675,4.784408,5.5331616,6.2801023,7.027043,7.7757964,8.073122,8.370448,8.667774,8.9651,9.262425,10.832452,12.402477,13.972503,15.542528,17.112555,19.250036,21.38752,23.525002,25.662485,27.799969,26.695873,25.589968,24.485872,23.379965,22.275871,20.927027,19.579996,18.232965,16.885933,15.537089,14.904366,14.271642,13.640731,13.008006,12.375282,10.879588,9.385707,7.890013,6.394319,4.900438,4.0392804,3.1799364,2.3205922,1.4594349,0.6000906,0.90466833,1.209246,1.5156367,1.8202144,2.124792,2.472881,2.819157,3.1672456,3.5153344,3.8616104,4.902251,5.942891,6.981719,8.02236,9.063,7.645263,6.2275267,4.8097897,3.392053,1.9743162,1.5881553,1.2001812,0.8122072,0.42423326,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.13959812,0.1794833,0.21936847,0.25925365,0.2991388,0.38072214,0.4604925,0.5402629,0.6200332,0.69980353,1.0950294,1.4902552,1.8854811,2.280707,2.6741197,3.5570326,4.439945,5.3228583,6.205771,7.0868707,6.8983226,6.7079616,6.5176005,6.3272395,6.1368785,6.3308654,6.5230393,6.7152133,6.9073873,7.0995617,7.9806614,8.859948,9.739235,10.620335,11.499621,12.083396,12.665357,13.247317,13.829279,14.413053,14.249886,12.774135,11.300196,9.824444,8.350506,6.874754,6.813113,6.7496595,6.688019,6.624565,6.5629244,7.4494634,8.337815,9.224354,10.112705,10.999244,10.012992,9.024928,8.036863,7.0506115,6.0625467,5.638314,5.2122674,4.788034,4.361988,3.9377546,4.162562,4.3873696,4.612177,4.836984,5.0617914,4.762653,4.461701,4.162562,3.8616104,3.5624714,3.7002566,3.8380418,3.975827,4.1117992,4.249584,4.650249,5.049101,5.4497657,5.8504305,6.249282,5.7869763,5.3246713,4.8623657,4.40006,3.9377546,3.6621845,3.386614,3.1128569,2.8372865,2.561716,2.0504606,1.5373923,1.0243238,0.51306844,0.0,0.0,0.0,0.0,0.0,0.0,0.2374981,0.4749962,0.7124943,0.9499924,1.1874905,1.0750868,0.96268314,0.85027945,0.73787576,0.62547207,0.76325727,0.89922947,1.0370146,1.1747998,1.3125849,1.4376793,1.5627737,1.6878681,1.8129625,1.938057,1.7875811,1.6371052,1.4866294,1.3379664,1.1874905,0.9499924,0.7124943,0.4749962,0.2374981,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.63816285,1.2745126,1.9126755,2.5508385,3.1871881,3.149116,3.1128569,3.0747845,3.0367124,3.000453,2.4003625,1.8002719,1.2001812,0.6000906,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0870222,0.17585737,0.26287958,0.34990177,0.43692398,1.1367276,1.8383441,2.5381477,3.2379513,3.9377546,3.774588,3.6132345,3.4500678,3.2869012,3.1255474,2.6378605,2.1501737,1.6624867,1.1747998,0.6871128,1.4376793,2.1882458,2.9369993,3.6875658,4.4381323,4.4381323,4.4381323,4.4381323,4.4381323,4.4381323,4.0882306,3.738329,3.386614,3.0367124,2.6868105,2.1882458,1.6878681,1.1874905,0.6871128,0.18673515,1.0007553,1.8129625,2.6251698,3.437377,4.249584,4.6629395,5.0744824,5.487838,5.89938,6.3127356,6.16226,6.011784,5.863121,5.712645,5.562169,5.375434,5.186886,5.0001507,4.8116026,4.6248674,4.949388,5.275721,5.600241,5.924762,6.249282,5.52591,4.800725,4.07554,3.350355,2.6251698,2.5997884,2.5744069,2.5508385,2.525457,2.5000753,2.2879589,2.0758421,1.8619126,1.649796,1.4376793,1.1494182,0.8629702,0.5747091,0.28826106,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.11240368,0.22480737,0.33721104,0.44961473,0.5620184,0.44961473,0.33721104,0.22480737,0.11240368,0.0,0.46230546,0.9246109,1.3869164,1.8492218,2.3133402,2.0631514,1.8129625,1.5627737,1.3125849,1.062396,1.7875811,2.5127661,3.2379513,3.9631362,4.688321,4.537845,4.3873696,4.2368937,4.0882306,3.9377546,7.650702,11.361836,15.074784,18.787731,22.500679,19.987913,17.475147,14.96238,12.449615,9.936848,8.036863,6.1368785,4.2368937,2.3369088,0.43692398,3.5243993,6.6118746,9.699349,12.786825,15.8743,13.724127,11.575767,9.425592,7.2754188,5.125245,7.462154,9.799063,12.137785,14.474693,16.811602,14.525456,12.237497,9.949538,7.66158,5.375434,4.900438,4.4254417,3.9504454,3.4754493,3.000453,2.911618,2.8245957,2.7375734,2.6505513,2.561716,3.2252605,3.8869917,4.550536,5.2122674,5.8758116,5.375434,4.8750563,4.3746786,3.874301,3.3757362,3.2633326,3.149116,3.0367124,2.9243085,2.811905,2.561716,2.3133402,2.0631514,1.8129625,1.5627737,3.8507326,6.1368785,8.424837,10.712796,13.000754,11.887595,10.774437,9.663091,8.549932,7.4367723,6.0244746,4.612177,3.199879,1.7875811,0.37528324,0.2991388,0.22480737,0.15047589,0.07433146,0.0,0.16316663,0.3245203,0.48768693,0.6508536,0.8122072,0.6871128,0.5620184,0.43692398,0.31182957,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.0,0.0,0.0,0.0,0.0,1.6371052,3.2742105,4.9131284,6.550234,8.187339,7.574558,6.9617763,6.350808,5.7380266,5.125245,4.650249,4.175253,3.7002566,3.2252605,2.7502642,2.7883365,2.8245957,2.8626678,2.9007401,2.9369993,5.237649,7.5382986,9.837135,12.137785,14.436621,13.024323,11.612025,10.199727,8.78743,7.3751316,7.0868707,6.8004227,6.5121617,6.2257137,5.9374523,5.5367875,5.137936,4.7372713,4.3366065,3.9377546,4.6756306,5.411693,6.149569,6.887445,7.6253204,7.0125394,6.399758,5.7869763,5.1741953,4.5632267,5.4370747,6.3127356,7.1883965,8.062244,8.937905,9.325879,9.712041,10.100015,10.487988,10.874149,12.799516,14.724882,16.650248,18.575615,20.499168,22.837889,25.174799,27.511707,29.85043,32.187336,30.787731,29.388123,27.986704,26.587097,25.187489,23.43798,21.686659,19.93715,18.187641,16.438131,14.875358,13.312584,11.74981,10.1870365,8.624263,8.036863,7.4494634,6.8620634,6.2746634,5.6872635,4.699199,3.7129474,2.7248828,1.7368182,0.7505665,1.062396,1.3742256,1.6878681,1.9996977,2.3133402,2.4257438,2.5381477,2.6505513,2.762955,2.8753586,4.0882306,5.2992897,6.5121617,7.7250338,8.937905,7.500226,6.0625467,4.6248674,3.1871881,1.7495089,1.3996071,1.0497054,0.69980353,0.34990177,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.17585737,0.16316663,0.15047589,0.13778515,0.12509441,0.63816285,1.1494182,1.6624867,2.175555,2.6868105,3.7129474,4.7372713,5.763408,6.787732,7.8120556,7.424082,7.037921,6.6499467,6.261973,5.8758116,6.037165,6.200332,6.3616858,6.5248523,6.688019,7.799365,8.912524,10.025683,11.137029,12.250188,12.837588,13.424988,14.012388,14.599788,15.187187,12.224807,11.057259,9.88971,8.722163,7.554615,6.3870673,6.3272395,6.2674117,6.207584,6.147756,6.0879283,6.9001355,7.7123427,8.52455,9.336758,10.150778,9.400211,8.649645,7.899078,7.1503243,6.399758,6.049856,5.6999545,5.3500524,5.0001507,4.650249,4.8297324,5.009216,5.1905117,5.369995,5.5494785,5.335549,5.1198063,4.9058766,4.690134,4.4743915,4.349297,4.2242026,4.099108,3.975827,3.8507326,4.0918565,4.3347936,4.5777307,4.8206677,5.0617914,4.6792564,4.2967215,3.9141862,3.531651,3.149116,2.9297476,2.7103791,2.4891977,2.269829,2.0504606,1.6407311,1.2291887,0.8194591,0.40972954,0.0,0.0,0.0,0.0,0.0,0.0,0.19036107,0.38072214,0.56927025,0.75963134,0.9499924,0.85934424,0.7705091,0.67986095,0.58921283,0.50037766,0.6091554,0.7197462,0.83033687,0.93911463,1.0497054,1.1494182,1.2491312,1.3506571,1.4503701,1.550083,1.4304274,1.310772,1.1893034,1.0696479,0.9499924,0.75963134,0.56927025,0.38072214,0.19036107,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.6544795,1.209246,1.7658255,2.3205922,2.8753586,2.7955883,2.715818,2.6342347,2.5544643,2.474694,1.9797552,1.4848163,0.9898776,0.4949388,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.17041849,0.34083697,0.5094425,0.67986095,0.85027945,1.5247015,2.1991236,2.8753586,3.5497808,4.2242026,4.0157123,3.8054085,3.5951047,3.3848011,3.1744974,2.7248828,2.275268,1.8256533,1.3742256,0.9246109,1.4956942,2.0649643,2.6342347,3.2053177,3.774588,3.8054085,3.834416,3.8652363,3.8942437,3.925064,3.7618973,3.6005437,3.437377,3.2742105,3.1128569,2.8282216,2.5417736,2.2571385,1.9725033,1.6878681,2.322405,2.956942,3.5932918,4.227829,4.8623657,5.105303,5.3482394,5.5893636,5.8323007,6.0752378,5.9882154,5.89938,5.812358,5.7253356,5.638314,5.368182,5.0980506,4.8279195,4.557788,4.2876563,4.465327,4.6429973,4.8206677,4.9983377,5.1741953,4.572292,3.9703882,3.3666716,2.764768,2.1628644,2.1302311,2.0975976,2.0649643,2.032331,1.9996977,1.8292793,1.6606737,1.4902552,1.3198367,1.1494182,0.91917205,0.69073874,0.4604925,0.23024625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.17041849,0.29007402,0.40972954,0.5293851,0.6508536,0.62547207,0.6000906,0.5747091,0.5493277,0.52575916,0.69255173,0.85934424,1.0279498,1.1947423,1.3633479,1.5301404,1.696933,1.8655385,2.032331,2.1991236,1.983381,1.7658255,1.54827,1.3307146,1.1131591,2.3133402,3.5117085,4.7118897,5.9120708,7.112252,6.794984,6.4777155,6.1604466,5.8431783,5.52591,8.415772,11.3056345,14.195497,17.08536,19.975222,17.937452,15.899682,13.861912,11.8241415,9.788185,8.455658,7.12313,5.7906027,4.458075,3.1255474,5.2104545,7.2953615,9.380268,11.465176,13.550082,12.329959,11.109835,9.88971,8.669587,7.4494634,9.576068,11.700861,13.825653,15.950445,18.075237,15.464571,12.855718,10.245051,7.6343856,5.0255322,5.0074024,4.989273,4.972956,4.954827,4.93851,4.8496747,4.762653,4.6756306,4.5867953,4.499773,4.5450974,4.590421,4.6357455,4.6792564,4.7245803,4.8116026,4.900438,4.98746,5.0744824,5.163317,4.974769,4.788034,4.599486,4.4127507,4.2242026,3.9141862,3.6059825,3.295966,2.9859493,2.675933,4.3855567,6.09518,7.804804,9.514427,11.224051,10.391902,9.5597515,8.727602,7.895452,7.063302,5.8794374,4.6973863,3.5153344,2.333283,1.1494182,1.0007553,0.85027945,0.69980353,0.5493277,0.40066472,0.55839247,0.71430725,0.872035,1.0297627,1.1874905,1.0569572,0.92823684,0.79770356,0.6671702,0.53663695,0.47318324,0.40791658,0.34264994,0.27738327,0.21211663,0.19942589,0.18673515,0.17585737,0.16316663,0.15047589,1.452183,2.7557032,4.0574102,5.3591175,6.6626377,6.2529078,5.8431783,5.431636,5.0219064,4.612177,4.1915693,3.7727752,3.3521678,2.9333735,2.5127661,2.5870976,2.663242,2.7375734,2.811905,2.8880494,4.8333583,6.776854,8.722163,10.667472,12.612781,11.42529,10.2378,9.050309,7.8628187,6.6753283,6.4795284,6.285541,6.089741,5.8957543,5.6999545,5.3500524,5.0001507,4.650249,4.3003473,3.9504454,4.572292,5.1941376,5.8177967,6.439643,7.063302,7.117691,7.17208,7.228282,7.2826705,7.3370595,7.7776093,8.21816,8.656897,9.097446,9.537996,9.731983,9.927783,10.12177,10.31757,10.51337,12.311829,14.112101,15.912373,17.712645,19.512917,21.329504,23.147905,24.964495,26.782896,28.599485,27.332224,26.064962,24.797703,23.530441,22.26318,20.77655,19.291735,17.80692,16.322102,14.837286,13.314397,11.793322,10.270433,8.747544,7.224656,6.7496595,6.2746634,5.7996674,5.3246713,4.8496747,4.137181,3.4246864,2.712192,1.9996977,1.2872034,1.6534219,2.0178273,2.382233,2.7466383,3.1128569,3.3304121,3.5479677,3.7655232,3.9830787,4.2006345,5.230397,6.26016,7.2899227,8.319685,9.349448,8.029612,6.7097745,5.389938,4.070101,2.7502642,2.2498865,1.7495089,1.2491312,0.7505665,0.25018883,0.20667773,0.16497959,0.12328146,0.07977036,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.032633327,0.065266654,0.09789998,0.13053331,0.16316663,0.15228885,0.14322405,0.13234627,0.12328146,0.11240368,0.53663695,0.96268314,1.3869164,1.8129625,2.2371957,3.0620937,3.8869917,4.7118897,5.5367875,6.3616858,6.2746634,6.187641,6.1006193,6.011784,5.924762,5.99728,6.069799,6.1423173,6.2148356,6.2873545,7.2427855,8.198216,9.151835,10.107266,11.062697,11.668227,12.271944,12.877473,13.483003,14.0867195,10.199727,9.340384,8.479226,7.6198816,6.7605376,5.89938,5.8431783,5.7851634,5.727149,5.669134,5.612932,6.350808,7.0868707,7.8247466,8.562622,9.300498,8.78743,8.274362,7.763106,7.250037,6.736969,6.4632115,6.187641,5.9120708,5.638314,5.3627434,5.4969025,5.632875,5.767034,5.903006,6.037165,5.906632,5.7779117,5.6473784,5.516845,5.388125,5.0001507,4.612177,4.2242026,3.8380418,3.4500678,3.5352771,3.6204863,3.7056956,3.7909048,3.874301,3.5733492,3.2705846,2.9678197,2.665055,2.3622901,2.1973107,2.032331,1.8673514,1.7023718,1.5373923,1.2291887,0.922798,0.61459434,0.30820364,0.0,0.0,0.0,0.0,0.0,0.0,0.14322405,0.28463513,0.42785916,0.56927025,0.7124943,0.64541465,0.57833505,0.5094425,0.44236287,0.37528324,0.45686656,0.5402629,0.62184614,0.70524246,0.7868258,0.8629702,0.93730164,1.0116332,1.0877775,1.162109,1.0732739,0.9826257,0.8919776,0.8031424,0.7124943,0.56927025,0.42785916,0.28463513,0.14322405,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03988518,0.07977036,0.11965553,0.15954071,0.19942589,0.6726091,1.1457924,1.6171626,2.0903459,2.561716,2.4402475,2.3169663,2.1954978,2.0722163,1.9507477,1.5591478,1.1693609,0.7795739,0.38978696,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.2520018,0.5058166,0.75781834,1.0098201,1.261822,1.9126755,2.561716,3.2125697,3.8616104,4.512464,4.255023,3.9975824,3.7401419,3.482701,3.2252605,2.811905,2.4003625,1.987007,1.5754645,1.162109,1.551896,1.9416829,2.333283,2.72307,3.1128569,3.1726844,3.2325122,3.29234,3.3521678,3.4119956,3.437377,3.4627585,3.48814,3.5117085,3.53709,3.4681973,3.397492,3.3267863,3.2578938,3.1871881,3.644055,4.102734,4.559601,5.0182805,5.475147,5.5476656,5.620184,5.6927023,5.765221,5.8377395,5.812358,5.7869763,5.7615952,5.7380266,5.712645,5.3591175,5.0074024,4.655688,4.3021603,3.9504454,3.9794528,4.0102735,4.0392804,4.070101,4.100921,3.6204863,3.1400511,2.659616,2.179181,1.7005589,1.6606737,1.6207886,1.5809034,1.5392052,1.49932,1.3724127,1.2455053,1.1167849,0.9898776,0.8629702,0.69073874,0.5166943,0.3444629,0.17223145,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.34083697,0.58014804,0.8194591,1.0605831,1.2998942,1.1367276,0.97537386,0.8122072,0.6508536,0.48768693,0.9354887,1.3832904,1.8292793,2.277081,2.7248828,2.5979755,2.469255,2.3423476,2.2154403,2.08672,1.9017978,1.7168756,1.5319533,1.3470312,1.162109,2.8372865,4.512464,6.187641,7.8628187,9.537996,9.052122,8.568061,8.082188,7.5981264,7.112252,9.180842,11.24762,13.314397,15.382988,17.449764,15.8869915,14.324218,12.763257,11.200482,9.637709,8.872639,8.107569,7.3424983,6.5774283,5.812358,6.8946967,7.9770355,9.059374,10.141713,11.225864,10.93579,10.645717,10.355642,10.065568,9.775495,11.6881695,13.599032,15.511708,17.424383,19.337059,16.405499,13.472125,10.540565,7.607191,4.6756306,5.1143675,5.5549173,5.995467,6.434204,6.874754,6.787732,6.70071,6.6118746,6.5248523,6.43783,5.864934,5.292038,4.7191415,4.1480584,3.5751622,4.249584,4.9258194,5.600241,6.2746634,6.9490857,6.688019,6.4251394,6.16226,5.89938,5.638314,5.2666564,4.896812,4.5269675,4.157123,3.787279,4.9203806,6.051669,7.1847706,8.317872,9.449161,8.898021,8.345067,7.7921133,7.2391596,6.688019,5.7344007,4.782595,3.83079,2.8771715,1.9253663,1.7005589,1.4757515,1.2491312,1.0243238,0.7995165,0.95180535,1.1040943,1.258196,1.4104849,1.5627737,1.4268016,1.2926424,1.1566701,1.0225109,0.8883517,0.79589057,0.7016165,0.6091554,0.5166943,0.42423326,0.40066472,0.37528324,0.34990177,0.3245203,0.2991388,1.2672608,2.2353828,3.2016919,4.169814,5.137936,4.9294453,4.7227674,4.514277,4.307599,4.100921,3.7347028,3.3702974,3.005892,2.6396735,2.275268,2.3876717,2.5000753,2.612479,2.7248828,2.8372865,4.4272547,6.017223,7.607191,9.197159,10.7871275,9.824444,8.861761,7.900891,6.9382076,5.975525,5.8721857,5.77066,5.667321,5.565795,5.462456,5.163317,4.8623657,4.5632267,4.262275,3.9631362,4.4707656,4.9783955,5.484212,5.9918413,6.4994707,7.2228427,7.944402,8.667774,9.389333,10.112705,10.118144,10.12177,10.127209,10.1326475,10.138086,10.139899,10.141713,10.145339,10.147152,10.150778,11.825955,13.499319,15.174497,16.849674,18.52485,19.822933,21.119202,22.417282,23.715364,25.013445,23.876717,22.741802,21.606888,20.471973,19.337059,18.116936,16.89681,15.676687,14.458377,13.238253,11.755249,10.272246,8.789243,7.308052,5.825049,5.462456,5.0998635,4.7372713,4.3746786,4.0120864,3.5751622,3.1382382,2.6995013,2.2625773,1.8256533,2.2426348,2.659616,3.0765975,3.4953918,3.9123733,4.2350807,4.557788,4.880495,5.2032027,5.524097,6.3725634,7.219217,8.067683,8.914337,9.762803,8.560809,7.3570023,6.155008,4.953014,3.7492065,3.100166,2.4493124,1.8002719,1.1494182,0.50037766,0.41516843,0.32995918,0.24474995,0.15954071,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.027194439,0.054388877,0.08339628,0.11059072,0.13778515,0.13053331,0.12328146,0.11421664,0.10696479,0.099712946,0.43692398,0.775948,1.1131591,1.4503701,1.7875811,2.4130533,3.0367124,3.6621845,4.2876563,4.9131284,5.125245,5.337362,5.5494785,5.7615952,5.975525,5.957395,5.9392653,5.922949,5.904819,5.8866897,6.684393,7.4820967,8.2798,9.077503,9.875207,10.497053,11.120712,11.7425585,12.364405,12.988064,8.174648,7.6216946,7.0705543,6.5176005,5.964647,5.411693,5.3573046,5.3029156,5.2467136,5.1923246,5.137936,5.7996674,6.4632115,7.124943,7.7866745,8.450218,8.174648,7.900891,7.6253204,7.3497505,7.07418,6.874754,6.6753283,6.4759026,6.2746634,6.0752378,6.165886,6.2547207,6.345369,6.434204,6.5248523,6.4795284,6.434204,6.390693,6.345369,6.300045,5.6491914,5.0001507,4.349297,3.7002566,3.049403,2.9768846,2.904366,2.8318477,2.759329,2.6868105,2.465629,2.2426348,2.0196402,1.7966459,1.5754645,1.4648738,1.3542831,1.2455053,1.1349145,1.0243238,0.8194591,0.61459434,0.40972954,0.20486477,0.0,0.0,0.0,0.0,0.0,0.0,0.09427405,0.19036107,0.28463513,0.38072214,0.4749962,0.42967212,0.38434806,0.34083697,0.2955129,0.25018883,0.3045777,0.36077955,0.41516843,0.46955732,0.52575916,0.5747091,0.62547207,0.6744221,0.72518504,0.774135,0.71430725,0.6544795,0.5946517,0.53482395,0.4749962,0.38072214,0.28463513,0.19036107,0.09427405,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.059827764,0.11965553,0.1794833,0.23931105,0.2991388,0.69073874,1.0805258,1.4703126,1.8600996,2.2498865,2.084907,1.9199274,1.7549478,1.5899682,1.4249886,1.1403534,0.8557183,0.56927025,0.28463513,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.33539808,0.67079616,1.0043813,1.3397794,1.6751775,2.3006494,2.9243085,3.5497808,4.175253,4.800725,4.494334,4.1897564,3.8851788,3.5806012,3.2742105,2.9007401,2.525457,2.1501737,1.7748904,1.3996071,1.6099107,1.8202144,2.030518,2.2408218,2.4493124,2.5399606,2.6306088,2.7194438,2.810092,2.9007401,3.1128569,3.3249733,3.53709,3.7492065,3.9631362,4.1081734,4.25321,4.3982472,4.5432844,4.688321,4.9675174,5.2467136,5.527723,5.806919,6.0879283,5.9900284,5.8921285,5.7942286,5.6981416,5.600241,5.638314,5.674573,5.712645,5.750717,5.7869763,5.351866,4.9167547,4.4816437,4.0483456,3.6132345,3.4953918,3.3775494,3.2597067,3.141864,3.0258346,2.666868,2.3097143,1.9525607,1.5954071,1.2382535,1.1893034,1.1421664,1.0950294,1.0478923,1.0007553,0.9155461,0.83033687,0.7451276,0.65991837,0.5747091,0.4604925,0.3444629,0.23024625,0.11421664,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.030820364,0.059827764,0.09064813,0.11965553,0.15047589,0.5094425,0.87022203,1.2291887,1.5899682,1.9507477,1.649796,1.3506571,1.0497054,0.7505665,0.44961473,1.1784257,1.9054236,2.6324217,3.3594196,4.0882306,3.6658103,3.24339,2.819157,2.3967366,1.9743162,1.8220274,1.6697385,1.5174497,1.3651608,1.2128719,3.3630457,5.5132194,7.663393,9.811753,11.961927,11.30926,10.658407,10.00574,9.353074,8.700407,9.945912,11.189605,12.43511,13.680615,14.924308,13.836531,12.750566,11.662788,10.57501,9.487233,9.28962,9.092008,8.894395,8.696781,8.500981,8.580752,8.660522,8.740293,8.820063,8.899834,9.539809,10.179785,10.81976,11.459737,12.099712,13.800271,15.50083,17.199575,18.900135,20.600695,17.344612,14.090345,10.834265,7.5799966,4.325729,5.223145,6.1205616,7.017978,7.915395,8.812811,8.725789,8.636953,8.549932,8.46291,8.375887,7.1847706,5.995467,4.804351,3.6150475,2.4257438,3.6875658,4.949388,6.2130227,7.474845,8.736667,8.399456,8.062244,7.7250338,7.3878226,7.0506115,6.6191263,6.189454,5.7597823,5.33011,4.900438,5.4552045,6.009971,6.5647373,7.119504,7.6742706,7.402326,7.130382,6.8566246,6.58468,6.3127356,5.5893636,4.8678045,4.1444325,3.4228733,2.6995013,2.4003625,2.0994108,1.8002719,1.49932,1.2001812,1.3470312,1.4956942,1.6425442,1.789394,1.938057,1.7966459,1.6570477,1.5174497,1.3778516,1.2382535,1.1167849,0.99712944,0.8774739,0.75781834,0.63816285,0.6000906,0.5620184,0.52575916,0.48768693,0.44961473,1.0823387,1.7150626,2.3477864,2.9805105,3.6132345,3.6077955,3.6023567,3.5969179,3.5932918,3.587853,3.2778363,2.9678197,2.657803,2.3477864,2.03777,2.1882458,2.3369088,2.4873846,2.6378605,2.7883365,4.022964,5.2575917,6.492219,7.7268467,8.963287,8.225411,7.4875355,6.7496595,6.011784,5.275721,5.2648435,5.2557783,5.2449007,5.235836,5.224958,4.974769,4.7245803,4.4743915,4.2242026,3.975827,4.367427,4.76084,5.1524396,5.5458527,5.9374523,7.327995,8.716724,10.107266,11.497808,12.888351,12.456866,12.027194,11.597522,11.16785,10.738177,10.547816,10.357455,10.167094,9.976733,9.788185,11.338268,12.8865385,14.436621,15.986704,17.536787,18.314548,19.092308,19.87007,20.647831,21.425592,20.423023,19.420456,18.417887,17.41532,16.41275,15.457319,14.501887,13.548269,12.592838,11.637406,10.194288,8.752983,7.309865,5.866747,4.4254417,4.175253,3.925064,3.6748753,3.4246864,3.1744974,3.0131438,2.8499773,2.6868105,2.525457,2.3622901,2.8318477,3.303218,3.7727752,4.2423325,4.7118897,5.139749,5.567608,5.995467,6.4233265,6.849373,7.51473,8.180087,8.845445,9.510801,10.174346,9.090195,8.00423,6.9200783,5.8359265,4.749962,3.9504454,3.150929,2.3495996,1.550083,0.7505665,0.62184614,0.4949388,0.3680314,0.23931105,0.11240368,0.09064813,0.06707962,0.045324065,0.02175555,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02175555,0.045324065,0.06707962,0.09064813,0.11240368,0.10696479,0.10333887,0.09789998,0.092461094,0.0870222,0.33721104,0.5873999,0.8375887,1.0877775,1.3379664,1.7621996,2.1882458,2.612479,3.0367124,3.4627585,3.975827,4.4870825,5.0001507,5.5132194,6.0244746,5.91751,5.810545,5.7017674,5.5948024,5.487838,6.1278133,6.7677894,7.407765,8.047741,8.6877165,9.327692,9.967669,10.607644,11.24762,11.887595,6.149569,5.904819,5.660069,5.4153194,5.1705694,4.9258194,4.8732433,4.8206677,4.7680917,4.7155156,4.6629395,5.2503395,5.8377395,6.4251394,7.0125394,7.5999393,7.5618668,7.5256076,7.4875355,7.4494634,7.413204,7.28811,7.1630154,7.037921,6.9128265,6.787732,6.833056,6.87838,6.921891,6.967215,7.0125394,7.0524244,7.0923095,7.132195,7.17208,7.211965,6.300045,5.388125,4.4743915,3.5624714,2.6505513,2.420305,2.1900587,1.9598125,1.7295663,1.49932,1.357909,1.214685,1.0732739,0.9300498,0.7868258,0.7324369,0.678048,0.62184614,0.56745726,0.51306844,0.40972954,0.30820364,0.20486477,0.10333887,0.0,0.0,0.0,0.0,0.0,0.0,0.047137026,0.09427405,0.14322405,0.19036107,0.2374981,0.21574254,0.19217403,0.17041849,0.14684997,0.12509441,0.15228885,0.1794833,0.20667773,0.23568514,0.26287958,0.28826106,0.31182957,0.33721104,0.36259252,0.387974,0.35715362,0.32814622,0.29732585,0.26831847,0.2374981,0.19036107,0.14322405,0.09427405,0.047137026,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07977036,0.15954071,0.23931105,0.3208944,0.40066472,0.7070554,1.015259,1.3216497,1.6298534,1.938057,1.7295663,1.5228885,1.3143979,1.1077201,0.89922947,0.7197462,0.5402629,0.36077955,0.1794833,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.4169814,0.83577573,1.2527572,1.6697385,2.08672,2.6868105,3.2869012,3.8869917,4.4870825,5.087173,4.7354584,4.3819304,4.0302157,3.6766882,3.3249733,2.9877625,2.6505513,2.3133402,1.9743162,1.6371052,1.6679256,1.696933,1.7277533,1.7567607,1.7875811,1.9072367,2.0268922,2.1483607,2.268016,2.3876717,2.7883365,3.1871881,3.587853,3.9867048,4.3873696,4.748149,5.1071157,5.467895,5.826862,6.187641,6.2891674,6.392506,6.495845,6.5973706,6.70071,6.432391,6.165886,5.8975673,5.6292486,5.3627434,5.462456,5.562169,5.661882,5.763408,5.863121,5.3446136,4.8279195,4.309412,3.7927177,3.2742105,3.009518,2.7448254,2.4801328,2.2154403,1.9507477,1.7150626,1.4793775,1.2455053,1.0098201,0.774135,0.7197462,0.6653573,0.6091554,0.55476654,0.50037766,0.45686656,0.41516843,0.37165734,0.32995918,0.28826106,0.23024625,0.17223145,0.11421664,0.058014803,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03988518,0.07977036,0.11965553,0.15954071,0.19942589,0.67986095,1.1602961,1.6407311,2.1193533,2.5997884,2.1628644,1.7241274,1.2872034,0.85027945,0.41335547,1.4195497,2.427557,3.435564,4.441758,5.4497657,4.7318325,4.0157123,3.2977788,2.5798457,1.8619126,1.742257,1.6226015,1.502946,1.3832904,1.261822,3.8869917,6.5121617,9.137331,11.762501,14.387671,13.568212,12.74694,11.927481,11.108022,10.28675,10.70917,11.13159,11.555823,11.978244,12.400664,11.787883,11.175101,10.56232,9.949538,9.336758,9.708415,10.078259,10.448103,10.817947,11.187792,10.264994,9.342196,8.419398,7.4966,6.5756154,8.145641,9.715667,11.285692,12.855718,14.425743,15.912373,17.400814,18.887444,20.375887,21.862516,18.285542,14.706753,11.129777,7.552802,3.975827,5.33011,6.684393,8.040489,9.394773,10.750868,10.662033,10.57501,10.487988,10.399154,10.312131,8.504607,6.697084,4.88956,3.0820365,1.2745126,3.1255474,4.974769,6.825804,8.675026,10.524248,10.112705,9.699349,9.287807,8.874452,8.46291,7.9715962,7.4820967,6.9925966,6.5030966,6.011784,5.9900284,5.9682727,5.9447045,5.922949,5.89938,5.906632,5.915697,5.922949,5.9302006,5.9374523,5.4443264,4.953014,4.459888,3.966762,3.4754493,3.100166,2.7248828,2.3495996,1.9743162,1.6008459,1.742257,1.8854811,2.0268922,2.1701162,2.3133402,2.1683033,2.0232663,1.8782293,1.7331922,1.5881553,1.4394923,1.2926424,1.1457924,0.99712944,0.85027945,0.7995165,0.7505665,0.69980353,0.6508536,0.6000906,0.8974165,1.1947423,1.4920682,1.789394,2.08672,2.2843328,2.4819458,2.6795588,2.8771715,3.0747845,2.819157,2.565342,2.3097143,2.0540867,1.8002719,1.987007,2.175555,2.3622901,2.5508385,2.7375734,3.6168604,4.49796,5.377247,6.258347,7.137634,6.624565,6.11331,5.600241,5.087173,4.574105,4.6575007,4.7390842,4.8224807,4.9058766,4.98746,4.788034,4.5867953,4.3873696,4.1879435,3.9867048,4.265901,4.5432844,4.8206677,5.0980506,5.375434,7.4331465,9.489046,11.546759,13.604471,15.662184,14.7974,13.932617,13.067834,12.203052,11.338268,10.955733,10.573197,10.190662,9.808127,9.425592,10.850581,12.27557,13.700559,15.125546,16.550535,16.807976,17.065416,17.322857,17.580297,17.837738,16.967516,16.097294,15.227073,14.356851,13.486629,12.797703,12.106964,11.418038,10.7273,10.038374,8.63514,7.231908,5.8304877,4.4272547,3.0258346,2.8880494,2.7502642,2.612479,2.474694,2.3369088,2.4493124,2.561716,2.6741197,2.7883365,2.9007401,3.4228733,3.9450066,4.4671397,4.989273,5.5132194,6.0444174,6.5774283,7.1104393,7.6416373,8.174648,8.656897,9.139144,9.623205,10.1054535,10.587702,9.619579,8.653271,7.6851482,6.717026,5.750717,4.800725,3.8507326,2.9007401,1.9507477,1.0007553,0.83033687,0.65991837,0.4894999,0.3208944,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.018129626,0.034446288,0.052575916,0.07070554,0.0870222,0.08520924,0.08339628,0.07977036,0.07795739,0.07433146,0.2374981,0.40066472,0.5620184,0.72518504,0.8883517,1.1131591,1.3379664,1.5627737,1.7875811,2.0123885,2.8245957,3.636803,4.4508233,5.2630305,6.0752378,5.8776245,5.6800117,5.482399,5.2847857,5.087173,5.569421,6.051669,6.53573,7.017978,7.500226,8.158332,8.814624,9.47273,10.130835,10.7871275,4.12449,4.1879435,4.249584,4.313038,4.3746786,4.4381323,4.3873696,4.3366065,4.2876563,4.2368937,4.1879435,4.699199,5.2122674,5.7253356,6.2384043,6.7496595,6.9508986,7.1503243,7.3497505,7.549176,7.750415,7.699652,7.650702,7.5999393,7.549176,7.500226,7.500226,7.500226,7.500226,7.500226,7.500226,7.6253204,7.750415,7.8755093,8.000604,8.125698,6.9508986,5.774286,4.599486,3.4246864,2.2498865,1.8619126,1.4757515,1.0877775,0.69980353,0.31182957,0.25018883,0.18673515,0.12509441,0.06164073,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.099712946,0.19942589,0.2991388,0.40066472,0.50037766,0.72518504,0.9499924,1.1747998,1.3996071,1.6244144,1.3742256,1.1258497,0.87566096,0.62547207,0.37528324,0.2991388,0.22480737,0.15047589,0.07433146,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.50037766,1.0007553,1.49932,1.9996977,2.5000753,3.0747845,3.6494937,4.2242026,4.800725,5.375434,4.974769,4.5759177,4.175253,3.774588,3.3757362,3.0747845,2.7756457,2.474694,2.175555,1.8746033,1.7241274,1.5754645,1.4249886,1.2745126,1.1258497,1.2745126,1.4249886,1.5754645,1.7241274,1.8746033,2.4620032,3.049403,3.636803,4.2242026,4.8116026,5.388125,5.962834,6.5375433,7.112252,7.686961,7.61263,7.5382986,7.462154,7.3878226,7.311678,6.874754,6.43783,5.999093,5.562169,5.125245,5.2865987,5.4497657,5.612932,5.774286,5.9374523,5.337362,4.7372713,4.137181,3.53709,2.9369993,2.525457,2.1121013,1.7005589,1.2872034,0.87566096,0.76325727,0.6508536,0.53663695,0.42423326,0.31182957,0.25018883,0.18673515,0.12509441,0.06164073,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,0.85027945,1.4503701,2.0504606,2.6505513,3.2506418,2.6741197,2.0994108,1.5247015,0.9499924,0.37528324,1.6624867,2.94969,4.2368937,5.52591,6.813113,5.7996674,4.788034,3.774588,2.762955,1.7495089,1.6624867,1.5754645,1.4866294,1.3996071,1.3125849,4.4127507,7.512917,10.613083,13.713249,16.811602,15.825351,14.837286,13.849221,12.862969,11.874905,11.47424,11.075388,10.674724,10.275872,9.875207,9.737422,9.599637,9.461852,9.325879,9.188094,10.125396,11.062697,11.999999,12.937301,13.874602,11.949236,10.025683,8.100317,6.1749506,4.249584,6.7496595,9.249735,11.74981,14.249886,16.749962,18.024473,19.3008,20.575312,21.849825,23.124338,19.224655,15.324973,11.42529,7.5256076,3.6241121,5.4370747,7.250037,9.063,10.874149,12.687112,12.60009,12.513068,12.4242325,12.337211,12.250188,9.824444,7.400513,4.974769,2.5508385,0.12509441,2.563529,5.0001507,7.4367723,9.875207,12.311829,11.8241415,11.338268,10.850581,10.362894,9.875207,9.324066,8.774739,8.225411,7.6742706,7.124943,6.5248523,5.924762,5.3246713,4.7245803,4.12449,4.4127507,4.699199,4.98746,5.275721,5.562169,5.2992897,5.038223,4.7753434,4.512464,4.249584,3.7999697,3.350355,2.9007401,2.4493124,1.9996977,2.137483,2.275268,2.4130533,2.5508385,2.6868105,2.5381477,2.3876717,2.2371957,2.08672,1.938057,1.7621996,1.5881553,1.4122978,1.2382535,1.062396,1.0007553,0.93730164,0.87566096,0.8122072,0.7505665,0.7124943,0.6744221,0.63816285,0.6000906,0.5620184,0.96268314,1.3633479,1.7621996,2.1628644,2.561716,2.3622901,2.1628644,1.9616255,1.7621996,1.5627737,1.7875811,2.0123885,2.2371957,2.4620032,2.6868105,3.2125697,3.738329,4.262275,4.788034,5.3119802,5.0255322,4.7372713,4.4508233,4.162562,3.874301,4.0501585,4.2242026,4.40006,4.574105,4.749962,4.599486,4.4508233,4.3003473,4.1498713,3.9993954,4.162562,4.325729,4.4870825,4.650249,4.8116026,7.5382986,10.263181,12.988064,15.712947,18.43783,17.137936,15.838041,14.538147,13.238253,11.938358,11.361836,10.7871275,10.212419,9.637709,9.063,10.362894,11.662788,12.962683,14.262577,15.56247,15.299591,15.036712,14.775645,14.512766,14.249886,13.512011,12.774135,12.038072,11.300196,10.56232,10.138086,9.712041,9.287807,8.861761,8.437528,7.07418,5.712645,4.349297,2.9877625,1.6244144,1.6008459,1.5754645,1.550083,1.5247015,1.49932,1.887294,2.275268,2.663242,3.049403,3.437377,4.0120864,4.5867953,5.163317,5.7380266,6.3127356,6.9508986,7.5872483,8.225411,8.861761,9.499924,9.800876,10.100015,10.399154,10.700105,10.999244,10.150778,9.300498,8.450218,7.5999393,6.7496595,5.6491914,4.550536,3.4500678,2.3495996,1.2491312,1.0370146,0.824898,0.61278135,0.40066472,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.13778515,0.21211663,0.28826106,0.36259252,0.43692398,0.46230546,0.48768693,0.51306844,0.53663695,0.5620184,1.6751775,2.7883365,3.8996825,5.0128417,6.1241875,5.8377395,5.5494785,5.2630305,4.974769,4.688321,5.0128417,5.337362,5.661882,5.9882154,6.3127356,6.987158,7.663393,8.337815,9.012237,9.686659,4.3746786,4.4526362,4.5305934,4.606738,4.6846952,4.762653,4.7372713,4.7118897,4.688321,4.6629395,4.6375585,5.029158,5.422571,5.814171,6.207584,6.599184,6.7297173,6.8602505,6.9907837,7.119504,7.250037,7.250037,7.250037,7.250037,7.250037,7.250037,7.1630154,7.07418,6.987158,6.9001355,6.813113,7.157576,7.502039,7.8483152,8.192778,8.537241,7.4820967,6.4269524,5.371808,4.3166637,3.2633326,2.6976883,2.132044,1.5682126,1.0025684,0.43692398,0.36984438,0.30276474,0.23568514,0.16679256,0.099712946,0.12690738,0.15591478,0.18310922,0.21030366,0.2374981,0.2574407,0.27738327,0.29732585,0.31726846,0.33721104,0.27013144,0.2030518,0.13415924,0.06707962,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.099712946,0.17585737,0.25018883,0.3245203,0.40066472,0.5982776,0.79589057,0.9916905,1.1893034,1.3869164,1.1693609,0.95180535,0.73424983,0.5166943,0.2991388,0.23931105,0.1794833,0.11965553,0.059827764,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.15772775,0.19036107,0.2229944,0.25562772,0.28826106,0.3245203,0.36259252,0.40066472,0.43692398,0.4749962,1.0243238,1.5754645,2.124792,2.675933,3.2252605,3.5606585,3.8942437,4.229642,4.5650396,4.900438,4.6593137,4.420003,4.1806917,3.9395678,3.7002566,3.489953,3.2796493,3.0693457,2.8608549,2.6505513,2.5381477,2.4257438,2.3133402,2.2009366,2.08672,2.280707,2.472881,2.665055,2.857229,3.049403,3.5534067,4.0555973,4.557788,5.0599785,5.562169,5.906632,6.2529078,6.5973706,6.9418335,7.28811,7.0705543,6.8529987,6.635443,6.4178877,6.200332,5.844991,5.4896507,5.1343102,4.780782,4.4254417,4.4925213,4.559601,4.6266804,4.695573,4.762653,4.2804046,3.7981565,3.3140955,2.8318477,2.3495996,2.0196402,1.6896812,1.3597219,1.0297627,0.69980353,0.6091554,0.52032024,0.42967212,0.34083697,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.11240368,0.19942589,0.28826106,0.37528324,0.46230546,1.015259,1.5682126,2.1193533,2.6723068,3.2252605,2.7466383,2.269829,1.79302,1.3143979,0.8375887,1.8673514,2.8971143,3.926877,4.95664,5.9882154,5.369995,4.751775,4.135368,3.5171473,2.9007401,2.7266958,2.5544643,2.382233,2.2100015,2.03777,4.539658,7.041547,9.545248,12.047136,14.549025,14.139296,13.729566,13.319836,12.910107,12.500377,11.894848,11.289318,10.685601,10.080072,9.474543,9.367578,9.2606125,9.151835,9.04487,8.937905,10.018432,11.097144,12.17767,13.258195,14.336908,12.843027,11.347333,9.853452,8.357758,6.8620634,8.410334,9.956791,11.50506,13.05333,14.599788,15.471823,16.34567,17.217705,18.08974,18.961775,15.848919,12.737875,9.625018,6.5121617,3.3993049,4.933071,6.4650245,7.996978,9.530745,11.062697,11.024626,10.986553,10.950294,10.912222,10.874149,9.164526,7.454902,5.7452784,4.0356545,2.326031,4.100921,5.8758116,7.650702,9.425592,11.200482,10.640278,10.080072,9.519867,8.9596615,8.399456,7.9752226,7.549176,7.124943,6.70071,6.2746634,6.115123,5.955582,5.7942286,5.634688,5.475147,5.4552045,5.4352617,5.4153194,5.3953767,5.375434,4.992899,4.610364,4.227829,3.8452935,3.4627585,3.1128569,2.762955,2.4130533,2.0631514,1.7132497,1.8093367,1.9072367,2.0051367,2.1030366,2.1991236,2.1066625,2.0142014,1.9217403,1.8292793,1.7368182,1.5917811,1.4467441,1.3017071,1.1566701,1.0116332,1.0424535,1.0732739,1.1022812,1.1331016,1.162109,1.1204109,1.0768998,1.0352017,0.9916905,0.9499924,1.3905423,1.8292793,2.269829,2.7103791,3.150929,3.0167696,2.8844235,2.752077,2.619731,2.4873846,2.6831846,2.8771715,3.0729716,3.2669585,3.4627585,3.8906176,4.3166637,4.744523,5.1723824,5.600241,5.239462,4.880495,4.519716,4.160749,3.7999697,3.9450066,4.0900435,4.2350807,4.3801174,4.5251546,4.3783045,4.229642,4.082792,3.9341288,3.787279,3.8471067,3.9069343,3.966762,4.02659,4.0882306,6.4106355,8.733041,11.055446,13.377851,15.700256,14.94425,14.190058,13.434052,12.67986,11.925668,11.254871,10.585889,9.915092,9.244296,8.575313,9.907841,11.240368,12.572895,13.905423,15.23795,14.839099,14.4420595,14.045021,13.647983,13.24913,12.654479,12.059827,11.465176,10.870523,10.275872,10.032935,9.789998,9.547061,9.305937,9.063,8.258044,7.453089,6.6481338,5.8431783,5.038223,5.1071157,5.177821,5.2485266,5.317419,5.388125,5.4207582,5.4533916,5.486025,5.516845,5.5494785,5.5929894,5.634688,5.678199,5.719897,5.7615952,6.285541,6.8076744,7.3298078,7.851941,8.374074,8.760235,9.144584,9.530745,9.915092,10.29944,9.487233,8.675026,7.8628187,7.0506115,6.2365913,5.2503395,4.262275,3.2742105,2.2879589,1.2998942,1.0696479,0.83940166,0.6091554,0.38072214,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.11240368,0.17585737,0.2374981,0.2991388,0.36259252,0.39159992,0.4224203,0.45324063,0.48224804,0.51306844,1.4431182,2.373168,3.303218,4.233268,5.163317,4.947575,4.7318325,4.517903,4.3021603,4.0882306,4.407312,4.7282066,5.047288,5.368182,5.6872635,6.8022356,7.9172077,9.03218,10.147152,11.262123,4.6248674,4.7173285,4.8097897,4.902251,4.994712,5.087173,5.087173,5.087173,5.087173,5.087173,5.087173,5.3591175,5.632875,5.904819,6.1767635,6.450521,6.510349,6.5701766,6.630004,6.6898317,6.7496595,6.8004227,6.849373,6.9001355,6.9508986,6.9998484,6.825804,6.6499467,6.4759026,6.300045,6.1241875,6.6898317,7.2554765,7.819308,8.384952,8.950596,8.015107,7.079619,6.14413,5.2104545,4.274966,3.531651,2.7901495,2.0468347,1.305333,0.5620184,0.4894999,0.4169814,0.3444629,0.27194437,0.19942589,0.25562772,0.3100166,0.36440548,0.42060733,0.4749962,0.5148814,0.55476654,0.5946517,0.6345369,0.6744221,0.5402629,0.40429065,0.27013144,0.13415924,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,0.2991388,0.46955732,0.6399758,0.8103943,0.9808127,1.1494182,0.9644961,0.7795739,0.5946517,0.40972954,0.22480737,0.1794833,0.13415924,0.09064813,0.045324065,0.0,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,0.3154555,0.38072214,0.44417584,0.5094425,0.5747091,0.6508536,0.72518504,0.7995165,0.87566096,0.9499924,1.550083,2.1501737,2.7502642,3.350355,3.9504454,4.0447197,4.1408067,4.2350807,4.329355,4.4254417,4.345671,4.265901,4.1843176,4.1045475,4.024777,3.9051213,3.785466,3.6658103,3.5443418,3.4246864,3.350355,3.2742105,3.199879,3.1255474,3.049403,3.2850883,3.5207734,3.7546456,3.9903307,4.2242026,4.6429973,5.0599785,5.47696,5.8957543,6.3127356,6.4269524,6.542982,6.6571984,6.773228,6.887445,6.526665,6.167699,5.806919,5.4479527,5.087173,4.8152285,4.5432844,4.269527,3.9975824,3.7256382,3.6966307,3.6694362,3.6422417,3.6150475,3.587853,3.2216346,2.857229,2.4928236,2.128418,1.7621996,1.5156367,1.2672608,1.020698,0.77232206,0.52575916,0.45686656,0.38978696,0.32270733,0.25562772,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.17585737,0.2991388,0.42423326,0.5493277,0.6744221,1.1802386,1.6842422,2.1900587,2.6958754,3.199879,2.819157,2.4402475,2.0595255,1.6806163,1.2998942,2.0722163,2.8445382,3.6168604,4.3891826,5.163317,4.940323,4.7173285,4.494334,4.273153,4.0501585,3.7927177,3.5352771,3.2778363,3.0203958,2.762955,4.668379,6.5719895,8.477413,10.382836,12.28826,12.455053,12.621845,12.790451,12.957244,13.125849,12.3154545,11.50506,10.694666,9.884272,9.07569,8.997733,8.919776,8.841819,8.765674,8.6877165,9.909654,11.13159,12.35534,13.577277,14.799213,13.735004,12.670795,11.6047735,10.540565,9.474543,10.069194,10.665659,11.26031,11.854962,12.449615,12.920984,13.390542,13.860099,14.329657,14.801026,12.474996,10.150778,7.8247466,5.5005283,3.1744974,4.4272547,5.6800117,6.932769,8.185526,9.438283,9.449161,9.461852,9.474543,9.487233,9.499924,8.504607,7.509291,6.5157876,5.520471,4.5251546,5.638314,6.7496595,7.8628187,8.974165,10.087324,9.4546,8.821876,8.189152,7.558241,6.925517,6.624565,6.3254266,6.0244746,5.7253356,5.424384,5.7053933,5.9845896,6.265599,6.544795,6.825804,6.497658,6.169512,5.8431783,5.5150323,5.186886,4.6846952,4.1825047,3.680314,3.1781235,2.6741197,2.4257438,2.175555,1.9253663,1.6751775,1.4249886,1.4830034,1.5392052,1.5972201,1.6552348,1.7132497,1.6769904,1.6425442,1.6080978,1.5718386,1.5373923,1.4231756,1.3071461,1.1929294,1.0768998,0.96268314,1.0841516,1.2074331,1.3307146,1.452183,1.5754645,1.5283275,1.4793775,1.4322405,1.3851035,1.3379664,1.8184015,2.2970235,2.7774587,3.2578938,3.738329,3.673062,3.6077955,3.5425289,3.4772623,3.4119956,3.576975,3.7419548,3.9069343,4.071914,4.2368937,4.5668526,4.896812,5.2267714,5.5567303,5.8866897,5.4552045,5.0219064,4.590421,4.157123,3.7256382,3.8398547,3.9558845,4.070101,4.1843176,4.3003473,4.15531,4.0102735,3.8652363,3.720199,3.5751622,3.531651,3.489953,3.4482548,3.4047437,3.3630457,5.282973,7.2029004,9.122828,11.042755,12.962683,12.752378,12.542075,12.331772,12.123281,11.912977,11.147907,10.382836,9.617766,8.852696,8.087626,9.452786,10.817947,12.183108,13.548269,14.911617,14.380419,13.847408,13.314397,12.783199,12.250188,11.7969475,11.34552,10.89228,10.440851,9.987611,9.927783,9.867955,9.808127,9.7483,9.686659,9.440096,9.19172,8.945157,8.696781,8.450218,8.615198,8.780178,8.945157,9.110137,9.275117,8.952409,8.629702,8.306994,7.9842873,7.66158,7.17208,6.68258,6.19308,5.7017674,5.2122674,5.620184,6.0281005,6.434204,6.8421206,7.250037,7.7195945,8.189152,8.660522,9.130079,9.599637,8.825501,8.049554,7.2754188,6.4994707,5.7253356,4.8496747,3.975827,3.100166,2.2245052,1.3506571,1.1022812,0.8557183,0.6073425,0.36077955,0.11240368,0.09064813,0.06707962,0.045324065,0.02175555,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.0870222,0.13778515,0.18673515,0.2374981,0.28826106,0.32270733,0.35715362,0.39159992,0.42785916,0.46230546,1.209246,1.9579996,2.70494,3.4518807,4.2006345,4.0574102,3.9141862,3.7727752,3.6295512,3.48814,3.8017826,4.117238,4.4326935,4.748149,5.0617914,6.6173134,8.172835,9.728357,11.282066,12.837588,4.8750563,4.9820213,5.090799,5.197764,5.3047285,5.411693,5.4370747,5.462456,5.487838,5.5132194,5.5367875,5.6908894,5.8431783,5.995467,6.147756,6.300045,6.2891674,6.2801023,6.2692246,6.26016,6.249282,6.350808,6.450521,6.550234,6.6499467,6.7496595,6.48678,6.2257137,5.962834,5.6999545,5.4370747,6.2220874,7.0071006,7.7921133,8.577126,9.362139,8.548119,7.7322855,6.9182653,6.1024323,5.2884116,4.367427,3.4482548,2.5272698,1.6080978,0.6871128,0.6091554,0.533011,0.4550536,0.3770962,0.2991388,0.3825351,0.46411842,0.5475147,0.630911,0.7124943,0.77232206,0.8321498,0.8919776,0.95180535,1.0116332,0.8103943,0.6073425,0.40429065,0.2030518,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.099712946,0.12509441,0.15047589,0.17585737,0.19942589,0.34264994,0.48587397,0.62728506,0.7705091,0.9119202,0.75963134,0.6073425,0.4550536,0.30276474,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.07433146,0.15047589,0.22480737,0.2991388,0.37528324,0.47318324,0.56927025,0.6671702,0.7650702,0.8629702,0.97537386,1.0877775,1.2001812,1.3125849,1.4249886,2.0758421,2.7248828,3.3757362,4.024777,4.6756306,4.5305934,4.3855567,4.2405195,4.0954823,3.9504454,4.0302157,4.1099863,4.1897564,4.269527,4.349297,4.3202896,4.2894692,4.2604623,4.229642,4.2006345,4.162562,4.12449,4.0882306,4.0501585,4.0120864,4.2894692,4.5668526,4.844236,5.123432,5.4008155,5.732588,6.0643597,6.397945,6.7297173,7.063302,6.947273,6.833056,6.717026,6.60281,6.48678,5.9845896,5.482399,4.9802084,4.478018,3.975827,3.785466,3.5951047,3.4047437,3.2143826,3.0258346,2.902553,2.7792716,2.657803,2.5345216,2.4130533,2.1646774,1.9181144,1.6697385,1.4231756,1.1747998,1.0098201,0.8448406,0.67986095,0.5148814,0.34990177,0.3045777,0.25925365,0.21574254,0.17041849,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.2374981,0.40066472,0.5620184,0.72518504,0.8883517,1.3452182,1.8020848,2.2607644,2.7176309,3.1744974,2.8916752,2.610666,2.327844,2.0450218,1.7621996,2.277081,2.7919624,3.3068438,3.8217251,4.3366065,4.510651,4.6828823,4.855114,5.027345,5.199577,4.856927,4.514277,4.171627,3.83079,3.48814,4.795286,6.1024323,7.409578,8.716724,10.025683,10.770811,11.514126,12.259253,13.00438,13.749508,12.734249,11.720803,10.705544,9.690285,8.675026,8.627889,8.580752,8.531802,8.484665,8.437528,9.802689,11.16785,12.5330105,13.898171,15.263332,14.626982,13.992445,13.357908,12.7233715,12.087022,11.729868,11.372714,11.015561,10.656594,10.29944,10.36652,10.435412,10.502492,10.5695715,10.636651,9.099259,7.5618668,6.0244746,4.4870825,2.94969,3.923251,4.894999,5.866747,6.8403077,7.8120556,7.8755093,7.93715,8.000604,8.062244,8.125698,7.844689,7.5654926,7.2844834,7.0052876,6.7242785,7.175706,7.6253204,8.074935,8.52455,8.974165,8.270736,7.5654926,6.8602505,6.155008,5.4497657,5.275721,5.0998635,4.9258194,4.749962,4.574105,5.295664,6.01541,6.735156,7.454902,8.174648,7.5401115,6.9055743,6.2692246,5.634688,5.0001507,4.3783045,3.7546456,3.1327994,2.5091403,1.887294,1.7368182,1.5881553,1.4376793,1.2872034,1.1367276,1.1548572,1.1729867,1.1893034,1.2074331,1.2255627,1.2473183,1.2708868,1.2926424,1.3143979,1.3379664,1.2527572,1.167548,1.0823387,0.99712944,0.9119202,1.1276628,1.3415923,1.5573349,1.7730774,1.987007,1.9344311,1.8818551,1.8292793,1.7767034,1.7241274,2.2444477,2.764768,3.2850883,3.8054085,4.325729,4.327542,4.329355,4.3329806,4.3347936,4.3384194,4.4725785,4.606738,4.74271,4.876869,5.0128417,5.2449007,5.47696,5.710832,5.942891,6.1749506,5.669134,5.1651306,4.6593137,4.15531,3.6494937,3.7347028,3.8199122,3.9051213,3.9903307,4.07554,3.9323158,3.7890918,3.6476808,3.5044568,3.3630457,3.2180085,3.0729716,2.9279346,2.7828975,2.6378605,4.15531,5.67276,7.1902094,8.70766,10.225109,10.560507,10.894093,11.22949,11.564888,11.900287,11.039129,10.179785,9.32044,8.459284,7.5999393,8.997733,10.395528,11.793322,13.189302,14.587097,13.919927,13.252756,12.585587,11.916603,11.249433,10.939416,10.629399,10.319383,10.009366,9.699349,9.822631,9.944099,10.067381,10.190662,10.312131,10.622148,10.932164,11.242181,11.552197,11.862214,12.123281,12.382534,12.6417885,12.902855,13.162108,12.485873,11.807825,11.129777,10.451729,9.775495,8.752983,7.7304726,6.7079616,5.6854506,4.6629395,4.954827,5.2467136,5.540414,5.8323007,6.1241875,6.680767,7.2355337,7.7903004,8.345067,8.899834,8.161958,7.4258947,6.688019,5.9501433,5.2122674,4.4508233,3.6875658,2.9243085,2.1628644,1.3996071,1.1349145,0.87022203,0.6055295,0.34083697,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.06164073,0.099712946,0.13778515,0.17585737,0.21211663,0.2520018,0.291887,0.33177215,0.37165734,0.41335547,0.97718686,1.5428312,2.1066625,2.6723068,3.2379513,3.1672456,3.0983531,3.0276475,2.956942,2.8880494,3.198066,3.5080826,3.8180993,4.1281157,4.4381323,6.432391,8.428463,10.422722,12.416981,14.413053,5.125245,5.2467136,5.369995,5.4932766,5.614745,5.7380266,5.7869763,5.8377395,5.8866897,5.9374523,5.9882154,6.0208488,6.051669,6.0843024,6.1169357,6.149569,6.069799,5.9900284,5.910258,5.8304877,5.750717,5.89938,6.049856,6.200332,6.350808,6.4994707,6.149569,5.7996674,5.4497657,5.0998635,4.749962,5.754343,6.7605376,7.764919,8.7693,9.775495,9.079316,8.384952,7.690587,6.9944096,6.300045,5.2032027,4.1045475,3.007705,1.9108626,0.8122072,0.7306239,0.64722764,0.5656443,0.48224804,0.40066472,0.5094425,0.6200332,0.7306239,0.83940166,0.9499924,1.0297627,1.1095331,1.1893034,1.2708868,1.3506571,1.0805258,0.8103943,0.5402629,0.27013144,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.099712946,0.099712946,0.099712946,0.099712946,0.099712946,0.21574254,0.32995918,0.44417584,0.56020546,0.6744221,0.55476654,0.43511102,0.3154555,0.19579996,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.099712946,0.19942589,0.2991388,0.40066472,0.50037766,0.629098,0.75963134,0.8901646,1.020698,1.1494182,1.2998942,1.4503701,1.6008459,1.7495089,1.8999848,2.5997884,3.299592,3.9993954,4.699199,5.4008155,5.0146546,4.6303062,4.2441454,3.8597972,3.4754493,3.7147603,3.9558845,4.195195,4.4345064,4.6756306,4.7354584,4.795286,4.855114,4.914942,4.974769,4.974769,4.974769,4.974769,4.974769,4.974769,5.295664,5.614745,5.9356394,6.2547207,6.5756154,6.8221784,7.0705543,7.317117,7.5654926,7.8120556,7.4675927,7.12313,6.776854,6.432391,6.0879283,5.4425135,4.797099,4.1516843,3.5080826,2.8626678,2.7557032,2.6469254,2.5399606,2.4329958,2.324218,2.1066625,1.889107,1.6733645,1.455809,1.2382535,1.1077201,0.97718686,0.8466535,0.7179332,0.5873999,0.5058166,0.4224203,0.34083697,0.2574407,0.17585737,0.15228885,0.13053331,0.10696479,0.08520924,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.2991388,0.50037766,0.69980353,0.89922947,1.1004683,1.5101979,1.9199274,2.3296568,2.7393866,3.149116,2.9641938,2.7792716,2.5943494,2.4094272,2.2245052,2.4819458,2.7393866,2.9968271,3.254268,3.5117085,4.079166,4.646623,5.2158933,5.7833505,6.350808,5.922949,5.4950895,5.06723,4.6393714,4.213325,4.9221935,5.632875,6.341743,7.0524244,7.763106,9.084756,10.408218,11.729868,13.05333,14.37498,13.154857,11.934732,10.714609,9.494485,8.274362,8.258044,8.239915,8.221786,8.205468,8.187339,9.695724,11.202296,12.710681,14.217253,15.725637,15.520773,15.3159075,15.10923,14.904366,14.699501,13.390542,12.07977,10.770811,9.460039,8.149267,7.8156815,7.4802837,7.1448855,6.8094873,6.474089,5.7253356,4.974769,4.2242026,3.4754493,2.7248828,3.4174345,4.1099863,4.802538,5.4950895,6.187641,6.300045,6.412449,6.5248523,6.637256,6.7496595,7.1847706,7.6198816,8.054993,8.490104,8.925215,8.713099,8.499168,8.287052,8.074935,7.8628187,7.0850577,6.3072968,5.529536,4.751775,3.975827,3.925064,3.874301,3.825351,3.774588,3.7256382,4.8859344,6.0444174,7.2047133,8.365009,9.525306,8.582565,7.6398244,6.697084,5.754343,4.8116026,4.070101,3.3267863,2.5852847,1.84197,1.1004683,1.0497054,1.0007553,0.9499924,0.89922947,0.85027945,0.82671094,0.80495536,0.78319985,0.75963134,0.73787576,0.81764615,0.8974165,0.97718686,1.0569572,1.1367276,1.0823387,1.0279498,0.97174793,0.91735905,0.8629702,1.1693609,1.4775645,1.7857682,2.0921588,2.4003625,2.3423476,2.2843328,2.228131,2.1701162,2.1121013,2.6723068,3.2325122,3.7927177,4.3529234,4.9131284,4.9820213,5.0527267,5.121619,5.1923246,5.2630305,5.368182,5.473334,5.576673,5.6818247,5.7869763,5.922949,6.057108,6.19308,6.3272395,6.4632115,5.8848767,5.3083544,4.7300196,4.1516843,3.5751622,3.6295512,3.6857529,3.7401419,3.7945306,3.8507326,3.7093215,3.5697234,3.4301252,3.290527,3.149116,2.902553,2.6541772,2.4076142,2.1592383,1.9126755,3.0276475,4.1426196,5.2575917,6.3725634,7.4875355,8.366822,9.247922,10.127209,11.008308,11.887595,10.932164,9.976733,9.023115,8.067683,7.112252,8.54268,9.973107,11.401722,12.8321495,14.262577,13.4594345,12.658105,11.854962,11.05182,10.25049,10.081885,9.915092,9.7483,9.579695,9.412902,9.71748,10.022058,10.326634,10.633025,10.937603,11.804199,12.672608,13.539205,14.407614,15.27421,15.62955,15.984891,16.34023,16.695572,17.050913,16.017525,14.985949,13.95256,12.920984,11.887595,10.332074,8.778365,7.2228427,5.667321,4.1117992,4.2894692,4.4671397,4.64481,4.8224807,5.0001507,5.6401267,6.2801023,6.9200783,7.560054,8.200029,7.500226,6.8004227,6.1006193,5.4008155,4.699199,4.0501585,3.3993049,2.7502642,2.0994108,1.4503701,1.167548,0.88472575,0.60190356,0.3208944,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.038072214,0.06164073,0.0870222,0.11240368,0.13778515,0.18310922,0.22662032,0.27194437,0.31726846,0.36259252,0.7451276,1.1276628,1.5101979,1.892733,2.275268,2.277081,2.280707,2.2825198,2.2843328,2.2879589,2.5925364,2.8971143,3.2016919,3.5080826,3.8126602,6.247469,8.682278,11.117086,13.551895,15.986704,5.375434,5.5132194,5.6491914,5.7869763,5.924762,6.0625467,6.1368785,6.2130227,6.2873545,6.3616858,6.43783,6.350808,6.261973,6.1749506,6.0879283,6.000906,5.8504305,5.6999545,5.5494785,5.4008155,5.2503395,5.4497657,5.6491914,5.8504305,6.049856,6.249282,5.812358,5.375434,4.936697,4.499773,4.062849,5.2865987,6.5121617,7.7377243,8.963287,10.1870365,9.612328,9.037619,8.46291,7.8882003,7.311678,6.037165,4.762653,3.48814,2.2118144,0.93730164,0.85027945,0.76325727,0.6744221,0.5873999,0.50037766,0.63816285,0.774135,0.9119202,1.0497054,1.1874905,1.2872034,1.3869164,1.4866294,1.5881553,1.6878681,1.3506571,1.0116332,0.6744221,0.33721104,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0870222,0.17585737,0.26287958,0.34990177,0.43692398,0.34990177,0.26287958,0.17585737,0.0870222,0.0,0.0,0.0,0.0,0.0,0.0,0.12509441,0.25018883,0.37528324,0.50037766,0.62547207,0.7868258,0.9499924,1.1131591,1.2745126,1.4376793,1.6244144,1.8129625,1.9996977,2.1882458,2.374981,3.1255474,3.874301,4.6248674,5.375434,6.1241875,5.5005283,4.8750563,4.249584,3.6241121,3.000453,3.3993049,3.7999697,4.2006345,4.599486,5.0001507,5.1506267,5.2992897,5.4497657,5.600241,5.750717,5.7869763,5.825049,5.863121,5.89938,5.9374523,6.300045,6.6626377,7.02523,7.3878226,7.750415,7.911769,8.074935,8.238102,8.399456,8.562622,7.987913,7.413204,6.836682,6.261973,5.6872635,4.900438,4.1117992,3.3249733,2.5381477,1.7495089,1.7241274,1.7005589,1.6751775,1.649796,1.6244144,1.3125849,1.0007553,0.6871128,0.37528324,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.36259252,0.6000906,0.8375887,1.0750868,1.3125849,1.6751775,2.03777,2.4003625,2.762955,3.1255474,3.0367124,2.94969,2.8626678,2.7756457,2.6868105,2.6868105,2.6868105,2.6868105,2.6868105,2.6868105,3.6494937,4.612177,5.57486,6.5375433,7.500226,6.987158,6.4759026,5.962834,5.4497657,4.936697,5.049101,5.163317,5.275721,5.388125,5.5005283,7.400513,9.300498,11.200482,13.100468,15.000452,13.575464,12.1504755,10.725487,9.300498,7.8755093,7.8882003,7.900891,7.911769,7.9244595,7.93715,9.5869465,11.236742,12.888351,14.538147,16.187943,16.41275,16.637558,16.862366,17.087172,17.31198,15.049402,12.786825,10.524248,8.26167,6.000906,5.2630305,4.5251546,3.787279,3.049403,2.3133402,2.3495996,2.3876717,2.4257438,2.4620032,2.5000753,2.913431,3.3249733,3.738329,4.1498713,4.5632267,4.7245803,4.8877473,5.049101,5.2122674,5.375434,6.5248523,7.6742706,8.825501,9.97492,11.124338,10.25049,9.374829,8.499168,7.6253204,6.7496595,5.89938,5.050914,4.2006345,3.350355,2.5000753,2.5744069,2.6505513,2.7248828,2.7992141,2.8753586,4.4743915,6.0752378,7.6742706,9.275117,10.874149,9.625018,8.375887,7.124943,5.8758116,4.6248674,3.7618973,2.9007401,2.03777,1.1747998,0.31182957,0.36259252,0.41335547,0.46230546,0.51306844,0.5620184,0.50037766,0.43692398,0.37528324,0.31182957,0.25018883,0.387974,0.52575916,0.66173136,0.7995165,0.93730164,0.9119202,0.8883517,0.8629702,0.8375887,0.8122072,1.2128719,1.6117238,2.0123885,2.4130533,2.811905,2.7502642,2.6868105,2.6251698,2.561716,2.5000753,3.100166,3.7002566,4.3003473,4.900438,5.5005283,5.638314,5.774286,5.9120708,6.049856,6.187641,6.261973,6.338117,6.412449,6.48678,6.5629244,6.599184,6.637256,6.6753283,6.7134004,6.7496595,6.1006193,5.4497657,4.800725,4.1498713,3.5008307,3.5243993,3.5497808,3.5751622,3.6005437,3.6241121,3.48814,3.350355,3.2125697,3.0747845,2.9369993,2.5870976,2.2371957,1.887294,1.5373923,1.1874905,1.8999848,2.612479,3.3249733,4.0374675,4.749962,6.1749506,7.5999393,9.024928,10.449916,11.874905,10.825199,9.775495,8.725789,7.6742706,6.624565,8.087626,9.550687,11.011934,12.474996,13.938056,13.000754,12.06164,11.124338,10.1870365,9.249735,9.224354,9.200785,9.175404,9.1500225,9.12464,9.612328,10.100015,10.587702,11.075388,11.563075,12.988064,14.413053,15.838041,17.26303,18.688019,19.137632,19.587248,20.036863,20.48829,20.937904,19.549175,18.16226,16.775343,15.388427,13.999697,11.912977,9.824444,7.7377243,5.6510043,3.5624714,3.6241121,3.6875658,3.7492065,3.8126602,3.874301,4.599486,5.3246713,6.049856,6.775041,7.500226,6.836682,6.1749506,5.5132194,4.8496747,4.1879435,3.6494937,3.1128569,2.5744069,2.03777,1.49932,1.2001812,0.89922947,0.6000906,0.2991388,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.11240368,0.16316663,0.21211663,0.26287958,0.31182957,0.51306844,0.7124943,0.9119202,1.1131591,1.3125849,1.3869164,1.4630609,1.5373923,1.6117238,1.6878681,1.987007,2.2879589,2.5870976,2.8880494,3.1871881,6.0625467,8.937905,11.813264,14.68681,17.562168,7.112252,7.1466985,7.1829576,7.217404,7.25185,7.28811,7.217404,7.1466985,7.077806,7.0071006,6.9382076,6.7605376,6.582867,6.4051967,6.2275267,6.049856,5.915697,5.7797246,5.6455655,5.5095935,5.375434,5.562169,5.750717,5.9374523,6.1241875,6.3127356,5.9392653,5.567608,5.1941376,4.8224807,4.4508233,5.371808,6.294606,7.217404,8.140202,9.063,8.564435,8.067683,7.569119,7.072367,6.5756154,5.524097,4.4743915,3.4246864,2.374981,1.3252757,1.2491312,1.1747998,1.1004683,1.0243238,0.9499924,1.0406405,1.1294757,1.2201238,1.310772,1.3996071,1.3977941,1.3941683,1.3923552,1.3905423,1.3869164,1.1294757,0.872035,0.61459434,0.35715362,0.099712946,0.17767033,0.25562772,0.33177215,0.40972954,0.48768693,0.4169814,0.3480888,0.27738327,0.20667773,0.13778515,0.12328146,0.10696479,0.092461094,0.07795739,0.06164073,0.21755551,0.37165734,0.5275721,0.68167394,0.8375887,0.67079616,0.50219065,0.33539808,0.16679256,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.36440548,0.7306239,1.0950294,1.4594349,1.8256533,1.6298534,1.4358664,1.2400664,1.0442665,0.85027945,0.67986095,0.5094425,0.34083697,0.17041849,0.0,0.045324065,0.09064813,0.13415924,0.1794833,0.22480737,0.2229944,0.21936847,0.21755551,0.21574254,0.21211663,0.28463513,0.35715362,0.42967212,0.50219065,0.5747091,0.46774435,0.36077955,0.2520018,0.14503701,0.038072214,0.059827764,0.08339628,0.10515183,0.12690738,0.15047589,0.33539808,0.52032024,0.70524246,0.8901646,1.0750868,1.2708868,1.4648738,1.6606737,1.8546607,2.0504606,2.1392958,2.229944,2.3205922,2.4094272,2.5000753,3.0421512,3.584227,4.1281157,4.670192,5.2122674,4.800725,4.3873696,3.975827,3.5624714,3.149116,3.7727752,4.3946214,5.0182805,5.6401267,6.261973,6.414262,6.5683637,6.720652,6.872941,7.02523,6.8620634,6.70071,6.5375433,6.3743763,6.2130227,6.4650245,6.717026,6.970841,7.2228427,7.474845,7.5419245,7.610817,7.6778965,7.744976,7.8120556,7.262728,6.7115874,6.16226,5.612932,5.0617914,4.3420453,3.6222992,2.902553,2.182807,1.4630609,1.4304274,1.3977941,1.3651608,1.3325275,1.2998942,1.0497054,0.7995165,0.5493277,0.2991388,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.11240368,0.12509441,0.13778515,0.15047589,0.16316663,0.13053331,0.09789998,0.065266654,0.032633327,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.047137026,0.09427405,0.14322405,0.19036107,0.2374981,0.43692398,0.63816285,0.8375887,1.0370146,1.2382535,1.5355793,1.8329052,2.1302311,2.427557,2.7248828,2.6995013,2.6741197,2.6505513,2.6251698,2.5997884,2.5907235,2.5798457,2.570781,2.5599031,2.5508385,3.3848011,4.220577,5.0545397,5.8903155,6.7242785,6.2746634,5.825049,5.375434,4.9258194,4.4743915,4.6194286,4.764466,4.9095025,5.0545397,5.199577,6.8004227,8.399456,10.000301,11.599335,13.200181,12.06164,10.924912,9.788185,8.649645,7.512917,7.5056653,7.4966,7.4893484,7.4820967,7.474845,8.939718,10.4045925,11.869466,13.33434,14.799213,15.734702,16.67019,17.60568,18.539356,19.474844,16.982021,14.49101,11.998186,9.5053625,7.0125394,6.4831543,5.9519563,5.422571,4.893186,4.361988,4.2949085,4.227829,4.160749,4.0918565,4.024777,4.1408067,4.255023,4.36924,4.4852695,4.599486,4.8678045,5.1343102,5.4026284,5.669134,5.9374523,6.796797,7.6579537,8.517298,9.376642,10.2378,9.271491,8.306994,7.3424983,6.378002,5.411693,4.7300196,4.0483456,3.3648586,2.6831846,1.9996977,2.1429217,2.2843328,2.427557,2.570781,2.712192,3.9576974,5.2032027,6.446895,7.6924005,8.937905,7.938963,6.9418335,5.9447045,4.947575,3.9504454,3.2306993,2.5091403,1.789394,1.0696479,0.34990177,0.42967212,0.5094425,0.58921283,0.67079616,0.7505665,0.69073874,0.630911,0.56927025,0.5094425,0.44961473,0.5293851,0.6091554,0.69073874,0.7705091,0.85027945,0.87566096,0.89922947,0.9246109,0.9499924,0.97537386,1.3923552,1.8093367,2.228131,2.6451125,3.0620937,3.007705,2.953316,2.8971143,2.8427253,2.7883365,3.5080826,4.227829,4.947575,5.667321,6.3870673,6.392506,6.397945,6.4033837,6.4070096,6.412449,6.6155005,6.816739,7.019791,7.2228427,7.4258947,7.230095,7.0342946,6.8403077,6.644508,6.450521,5.77066,5.090799,4.409125,3.729264,3.049403,3.1454902,3.2397642,3.3358512,3.4301252,3.5243993,3.5534067,3.5806012,3.6077955,3.63499,3.6621845,3.350355,3.0367124,2.7248828,2.4130533,2.0994108,2.810092,3.5207734,4.229642,4.940323,5.6491914,6.742408,7.835624,8.927028,10.020245,11.111648,10.41547,9.71748,9.019489,8.323311,7.6253204,9.11195,10.600392,12.087022,13.575464,15.062093,14.356851,13.653421,12.948178,12.242936,11.537694,11.019187,10.502492,9.985798,9.467291,8.950596,9.077503,9.2044115,9.333132,9.460039,9.5869465,10.839704,12.092461,13.345218,14.597975,15.850732,16.4617,17.074482,17.687263,18.300045,18.912827,18.575615,18.238403,17.89938,17.562168,17.224958,15.263332,13.299893,11.338268,9.374829,7.413204,6.880193,6.347182,5.815984,5.282973,4.749962,5.1923246,5.634688,6.0770507,6.5194135,6.9617763,6.300045,5.638314,4.974769,4.313038,3.6494937,3.1690586,2.6904364,2.2100015,1.7295663,1.2491312,1.0442665,0.83940166,0.6345369,0.42967212,0.22480737,0.18310922,0.13959812,0.09789998,0.054388877,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.02175555,0.032633327,0.04169814,0.052575916,0.06164073,0.11240368,0.16316663,0.21211663,0.26287958,0.31182957,0.52575916,0.73787576,0.9499924,1.162109,1.3742256,1.4268016,1.4793775,1.5319533,1.5845293,1.6371052,2.034144,2.4329958,2.8300345,3.2270734,3.625925,6.0226617,8.419398,10.817947,13.2146845,15.613234,8.849071,8.781991,8.714911,8.647832,8.580752,8.511859,8.29793,8.082188,7.8682575,7.652515,7.4367723,7.170267,6.9019485,6.635443,6.3671246,6.1006193,5.979151,5.859495,5.7398396,5.620184,5.5005283,5.674573,5.8504305,6.0244746,6.200332,6.3743763,6.0679855,5.7597823,5.4515786,5.145188,4.836984,5.4570174,6.0770507,6.697084,7.317117,7.93715,7.518356,7.0977483,6.677141,6.258347,5.8377395,5.0128417,4.1879435,3.3630457,2.5381477,1.7132497,1.649796,1.5881553,1.5247015,1.4630609,1.3996071,1.4431182,1.4848163,1.5283275,1.5700256,1.6117238,1.5083848,1.403233,1.2980812,1.1929294,1.0877775,0.9101072,0.7324369,0.55476654,0.3770962,0.19942589,0.35534066,0.5094425,0.6653573,0.8194591,0.97537386,0.83577573,0.69436467,0.55476654,0.41516843,0.2755703,0.24474995,0.21574254,0.18492219,0.15410182,0.12509441,0.43511102,0.7451276,1.0551442,1.3651608,1.6751775,1.3397794,1.0043813,0.67079616,0.33539808,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.7306239,1.4594349,2.1900587,2.9206827,3.6494937,3.2597067,2.8699198,2.4801328,2.0903459,1.7005589,1.3597219,1.020698,0.67986095,0.34083697,0.0,0.065266654,0.13053331,0.19579996,0.25925365,0.3245203,0.3444629,0.36440548,0.38434806,0.40429065,0.42423326,0.48224804,0.5402629,0.5982776,0.6544795,0.7124943,0.5855869,0.45686656,0.32995918,0.2030518,0.07433146,0.11965553,0.16497959,0.21030366,0.25562772,0.2991388,0.54570174,0.7904517,1.0352017,1.2799516,1.5247015,1.7531348,1.9797552,2.2081885,2.4348087,2.663242,2.6541772,2.6469254,2.6396735,2.6324217,2.6251698,2.960568,3.294153,3.6295512,3.9649491,4.3003473,4.100921,3.8996825,3.7002566,3.5008307,3.299592,4.1444325,4.989273,5.8341136,6.680767,7.5256076,7.6797094,7.835624,7.989726,8.145641,8.299743,7.93715,7.574558,7.211965,6.849373,6.48678,6.630004,6.773228,6.9146395,7.057863,7.1992745,7.17208,7.1448855,7.117691,7.0904965,7.063302,6.5375433,6.011784,5.487838,4.9620786,4.4381323,3.785466,3.1327994,2.4801328,1.8274662,1.1747998,1.1349145,1.0950294,1.0551442,1.015259,0.97537386,0.7868258,0.6000906,0.41335547,0.22480737,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03988518,0.07977036,0.11965553,0.15954071,0.19942589,0.22480737,0.25018883,0.2755703,0.2991388,0.3245203,0.25925365,0.19579996,0.13053331,0.065266654,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07070554,0.13959812,0.21030366,0.27919623,0.34990177,0.51306844,0.6744221,0.8375887,1.0007553,1.162109,1.3941683,1.6280404,1.8600996,2.0921588,2.324218,2.3622901,2.4003625,2.4366217,2.474694,2.5127661,2.4928236,2.472881,2.4529383,2.4329958,2.4130533,3.1201086,3.827164,4.5342193,5.243088,5.9501433,5.562169,5.1741953,4.788034,4.40006,4.0120864,4.1897564,4.367427,4.5450974,4.7227674,4.900438,6.200332,7.500226,8.80012,10.100015,11.399909,10.549629,9.699349,8.8508835,8.000604,7.1503243,7.12313,7.0941224,7.066928,7.039734,7.0125394,8.292491,9.572442,10.852394,12.132345,13.412297,15.058467,16.702824,18.347181,19.993351,21.637709,18.914639,16.193382,13.470312,10.747242,8.024173,7.703278,7.380571,7.057863,6.735156,6.412449,6.240217,6.0679855,5.8957543,5.7217097,5.5494785,5.368182,5.185073,5.0019636,4.8206677,4.6375585,5.009216,5.382686,5.754343,6.1278133,6.4994707,7.0705543,7.6398244,8.210908,8.780178,9.349448,8.294304,7.2391596,6.185828,5.130684,4.07554,3.5606585,3.045777,2.5308957,2.0142014,1.49932,1.7096237,1.9199274,2.1302311,2.3405347,2.5508385,3.43919,4.329355,5.219519,6.109684,6.9998484,6.2547207,5.5095935,4.764466,4.019338,3.2742105,2.6976883,2.1193533,1.5428312,0.9644961,0.387974,0.49675176,0.6073425,0.7179332,0.82671094,0.93730164,0.8792868,0.823085,0.7650702,0.7070554,0.6508536,0.6726091,0.69436467,0.7179332,0.73968875,0.76325727,0.8375887,0.9119202,0.9880646,1.062396,1.1367276,1.5718386,2.0069497,2.4420607,2.8771715,3.3122826,3.2651455,3.2180085,3.1708715,3.1219215,3.0747845,3.9141862,4.7554007,5.5948024,6.434204,7.2754188,7.1466985,7.019791,6.892884,6.7641635,6.637256,6.967215,7.2971745,7.6271334,7.957093,8.287052,7.859193,7.4331465,7.0052876,6.5774283,6.149569,5.4407005,4.7300196,4.019338,3.3104696,2.5997884,2.764768,2.9297476,3.094727,3.2597067,3.4246864,3.6168604,3.8108473,4.0030212,4.195195,4.3873696,4.1117992,3.8380418,3.5624714,3.2869012,3.0131438,3.720199,4.4272547,5.1343102,5.8431783,6.550234,7.309865,8.069496,8.829127,9.590572,10.3502035,10.00574,9.659465,9.3150015,8.970539,8.624263,10.138086,11.650098,13.162108,14.674119,16.187943,15.71476,15.241576,14.770206,14.297023,13.825653,12.814019,11.804199,10.794379,9.784559,8.774739,8.54268,8.31062,8.076748,7.844689,7.61263,8.693155,9.771869,10.852394,11.9329195,13.013446,13.7875805,14.561715,15.337664,16.1118,16.887747,17.60024,18.312735,19.025229,19.737724,20.450218,18.611874,16.775343,14.936998,13.100468,11.262123,10.13446,9.006798,7.8791356,6.7532854,5.6256227,5.7851634,5.9447045,6.104245,6.265599,6.4251394,5.7615952,5.0998635,4.4381323,3.774588,3.1128569,2.6904364,2.268016,1.845596,1.4231756,1.0007553,0.8901646,0.7795739,0.67079616,0.56020546,0.44961473,0.36440548,0.27919623,0.19579996,0.11059072,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.032633327,0.03988518,0.047137026,0.054388877,0.06164073,0.11240368,0.16316663,0.21211663,0.26287958,0.31182957,0.53663695,0.76325727,0.9880646,1.2128719,1.4376793,1.4666867,1.4975071,1.5283275,1.5573349,1.5881553,2.0830941,2.5780327,3.0729716,3.5679104,4.062849,5.9827766,7.902704,9.822631,11.7425585,13.662486,10.587702,10.417283,10.246864,10.078259,9.907841,9.737422,9.376642,9.017676,8.656897,8.29793,7.93715,7.5799966,7.2228427,6.8656893,6.506723,6.149569,6.0444174,5.9392653,5.8341136,5.730775,5.6256227,5.7869763,5.9501433,6.11331,6.2746634,6.43783,6.1948934,5.9519563,5.710832,5.467895,5.224958,5.542227,5.859495,6.1767635,6.495845,6.813113,6.4704633,6.1278133,5.7851634,5.4425135,5.0998635,4.499773,3.8996825,3.299592,2.6995013,2.0994108,2.0504606,1.9996977,1.9507477,1.8999848,1.8492218,1.845596,1.840157,1.8347181,1.8292793,1.8256533,1.6171626,1.4104849,1.2019942,0.99531645,0.7868258,0.69073874,0.59283876,0.4949388,0.39703882,0.2991388,0.533011,0.7650702,0.99712944,1.2291887,1.4630609,1.2527572,1.0424535,0.8321498,0.62184614,0.41335547,0.3680314,0.32270733,0.27738327,0.23205921,0.18673515,0.6526665,1.1167849,1.5827163,2.0468347,2.5127661,2.0105755,1.5083848,1.0043813,0.50219065,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.0950294,2.1900587,3.2850883,4.3801174,5.475147,4.88956,4.305786,3.720199,3.1346123,2.5508385,2.039583,1.5301404,1.020698,0.5094425,0.0,0.08520924,0.17041849,0.25562772,0.34083697,0.42423326,0.46774435,0.5094425,0.5529536,0.5946517,0.63816285,0.67986095,0.72337204,0.7650702,0.80676836,0.85027945,0.7016165,0.55476654,0.40791658,0.25925365,0.11240368,0.1794833,0.24837588,0.3154555,0.3825351,0.44961473,0.7541924,1.0605831,1.3651608,1.6697385,1.9743162,2.2353828,2.4946365,2.7557032,3.0149567,3.2742105,3.1708715,3.0657198,2.960568,2.855416,2.7502642,2.8771715,3.005892,3.1327994,3.2597067,3.386614,3.3993049,3.4119956,3.4246864,3.437377,3.4500678,4.517903,5.5857377,6.6517596,7.7195945,8.78743,8.945157,9.102885,9.2606125,9.418341,9.574255,9.012237,8.450218,7.8882003,7.324369,6.7623506,6.794984,6.827617,6.8602505,6.892884,6.925517,6.8022356,6.680767,6.5574856,6.434204,6.3127356,5.812358,5.3119802,4.8116026,4.313038,3.8126602,3.2270734,2.6432993,2.0577126,1.4721256,0.8883517,0.83940166,0.79226464,0.7451276,0.6979906,0.6508536,0.52575916,0.40066472,0.2755703,0.15047589,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.059827764,0.11965553,0.1794833,0.23931105,0.2991388,0.33721104,0.37528324,0.41335547,0.44961473,0.48768693,0.38978696,0.291887,0.19579996,0.09789998,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.092461094,0.18492219,0.27738327,0.36984438,0.46230546,0.5873999,0.7124943,0.8375887,0.96268314,1.0877775,1.2545701,1.4231756,1.5899682,1.7567607,1.9253663,2.0250793,2.124792,2.2245052,2.324218,2.4257438,2.3949237,2.3641033,2.335096,2.3042755,2.275268,2.855416,3.435564,4.0157123,4.59586,5.1741953,4.8496747,4.5251546,4.2006345,3.874301,3.5497808,3.7600844,3.9703882,4.1806917,4.3891826,4.599486,5.600241,6.599184,7.5999393,8.600695,9.599637,9.037619,8.4756,7.911769,7.3497505,6.787732,6.740595,6.6916447,6.644508,6.5973706,6.550234,7.645263,8.740293,9.835322,10.930351,12.025381,14.380419,16.735458,19.090496,21.445534,23.800573,20.847258,17.895754,14.942437,11.989121,9.037619,8.923402,8.807372,8.693155,8.577126,8.46291,8.185526,7.9081426,7.6307597,7.3533764,7.07418,6.5955577,6.115123,5.634688,5.1542525,4.6756306,5.1524396,5.6292486,6.107871,6.58468,7.063302,7.3424983,7.6216946,7.902704,8.1819,8.46291,7.317117,6.1731377,5.027345,3.881553,2.7375734,2.3894846,2.0432088,1.69512,1.3470312,1.0007553,1.2781386,1.5555218,1.8329052,2.1102884,2.3876717,2.9224956,3.4573197,3.9921436,4.5269675,5.0617914,4.5704784,4.077353,3.584227,3.092914,2.5997884,2.1646774,1.7295663,1.2944553,0.85934424,0.42423326,0.5656443,0.70524246,0.8448406,0.98443866,1.1258497,1.0696479,1.015259,0.96087015,0.90466833,0.85027945,0.81583315,0.7795739,0.7451276,0.7106813,0.6744221,0.7995165,0.9246109,1.0497054,1.1747998,1.2998942,1.7531348,2.2045624,2.657803,3.1092308,3.5624714,3.5225863,3.482701,3.442816,3.4029307,3.3630457,4.322103,5.282973,6.24203,7.2029004,8.161958,7.902704,7.6416373,7.382384,7.12313,6.8620634,7.320743,7.7776093,8.234476,8.693155,9.1500225,8.490104,7.8301854,7.170267,6.510349,5.8504305,5.1107416,4.36924,3.6295512,2.8898623,2.1501737,2.3858588,2.619731,2.855416,3.0892882,3.3249733,3.682127,4.0392804,4.3982472,4.7554007,5.1125546,4.8750563,4.6375585,4.40006,4.162562,3.925064,4.6303062,5.335549,6.0407915,6.7442207,7.4494634,7.877322,8.3051815,8.733041,9.1609,9.5869465,9.594198,9.603263,9.610515,9.617766,9.625018,11.162411,12.699803,14.237195,15.774588,17.31198,17.072668,16.833357,16.592234,16.352922,16.1118,14.610665,13.107719,11.6047735,10.101828,8.600695,8.007855,7.415017,6.8221784,6.2293396,5.638314,6.544795,7.453089,8.3595705,9.267865,10.174346,11.111648,12.050762,12.988064,13.925365,14.862667,16.624866,18.387066,20.149265,21.913279,23.675478,21.962229,20.250792,18.537542,16.826105,15.112856,13.390542,11.668227,9.945912,8.221786,6.4994707,6.378002,6.2547207,6.1332526,6.009971,5.8866897,5.224958,4.5632267,3.8996825,3.2379513,2.5744069,2.2100015,1.845596,1.4793775,1.114972,0.7505665,0.73424983,0.7197462,0.70524246,0.69073874,0.6744221,0.5475147,0.42060733,0.291887,0.16497959,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.04169814,0.047137026,0.052575916,0.058014803,0.06164073,0.11240368,0.16316663,0.21211663,0.26287958,0.31182957,0.5493277,0.7868258,1.0243238,1.261822,1.49932,1.5083848,1.5156367,1.5228885,1.5301404,1.5373923,2.1302311,2.72307,3.3159087,3.9069343,4.499773,5.942891,7.3860097,8.827314,10.270433,11.711739,12.32452,12.052575,11.780631,11.506873,11.234929,10.962985,10.457169,9.953164,9.447348,8.943344,8.437528,7.989726,7.5419245,7.0941224,6.6481338,6.200332,6.109684,6.0208488,5.9302006,5.8395524,5.750717,5.89938,6.049856,6.200332,6.350808,6.4994707,6.3218007,6.14413,5.9682727,5.7906027,5.612932,5.6274357,5.6419396,5.658256,5.67276,5.6872635,5.422571,5.1578784,4.893186,4.6266804,4.361988,3.9867048,3.6132345,3.2379513,2.8626678,2.4873846,2.4493124,2.4130533,2.374981,2.3369088,2.3006494,2.2480736,2.1954978,2.1429217,2.0903459,2.03777,1.7277533,1.4177368,1.1077201,0.79770356,0.48768693,0.46955732,0.45324063,0.43511102,0.4169814,0.40066472,0.7106813,1.020698,1.3307146,1.6407311,1.9507477,1.6697385,1.3905423,1.1095331,0.83033687,0.5493277,0.4894999,0.42967212,0.36984438,0.3100166,0.25018883,0.87022203,1.4902552,2.1102884,2.7303216,3.350355,2.6795588,2.0105755,1.3397794,0.67079616,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.4594349,2.9206827,4.3801174,5.8395524,7.3008003,6.5194135,5.7398396,4.9602656,4.1806917,3.3993049,2.7194438,2.039583,1.3597219,0.67986095,0.0,0.10515183,0.21030366,0.3154555,0.42060733,0.52575916,0.58921283,0.6544795,0.7197462,0.7850128,0.85027945,0.8774739,0.90466833,0.9318628,0.96087015,0.9880646,0.8194591,0.6526665,0.48587397,0.31726846,0.15047589,0.23931105,0.32995918,0.42060733,0.5094425,0.6000906,0.9644961,1.3307146,1.69512,2.0595255,2.4257438,2.7176309,3.009518,3.303218,3.5951047,3.8869917,3.6857529,3.482701,3.2796493,3.0765975,2.8753586,2.7955883,2.715818,2.6342347,2.5544643,2.474694,2.6995013,2.9243085,3.149116,3.3757362,3.6005437,4.88956,6.1803894,7.4694057,8.760235,10.049252,10.210606,10.370146,10.529687,10.689227,10.850581,10.087324,9.325879,8.562622,7.799365,7.037921,6.9599633,6.882006,6.8058615,6.7279043,6.6499467,6.432391,6.2148356,5.99728,5.7797246,5.562169,5.087173,4.612177,4.137181,3.6621845,3.1871881,2.6704938,2.1519866,1.6352923,1.1167849,0.6000906,0.54570174,0.4894999,0.43511102,0.38072214,0.3245203,0.26287958,0.19942589,0.13778515,0.07433146,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07977036,0.15954071,0.23931105,0.3208944,0.40066472,0.44961473,0.50037766,0.5493277,0.6000906,0.6508536,0.52032024,0.38978696,0.25925365,0.13053331,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.11421664,0.23024625,0.3444629,0.4604925,0.5747091,0.66173136,0.7505665,0.8375887,0.9246109,1.0116332,1.114972,1.2183108,1.3198367,1.4231756,1.5247015,1.6878681,1.8492218,2.0123885,2.175555,2.3369088,2.2970235,2.2571385,2.2172532,2.1773682,2.137483,2.5907235,3.0421512,3.4953918,3.9468195,4.40006,4.137181,3.874301,3.6132345,3.350355,3.0874753,3.3304121,3.5733492,3.8144734,4.0574102,4.3003473,5.0001507,5.6999545,6.399758,7.0995617,7.799365,7.5256076,7.250037,6.9744673,6.70071,6.4251394,6.35806,6.2891674,6.2220874,6.155008,6.0879283,6.9980354,7.9081426,8.81825,9.728357,10.636651,13.702372,16.768091,19.831997,22.897717,25.963438,22.779875,19.598125,16.414564,13.232814,10.049252,10.141713,10.234174,10.326634,10.420909,10.51337,10.130835,9.7483,9.365765,8.98323,8.600695,7.8229337,7.0451727,6.2674117,5.4896507,4.7118897,5.295664,5.8776245,6.4595857,7.0433598,7.6253204,7.614443,7.605378,7.5945,7.5854354,7.574558,6.33993,5.105303,3.870675,2.6342347,1.3996071,1.2201238,1.0406405,0.85934424,0.67986095,0.50037766,0.8448406,1.1893034,1.5355793,1.8800422,2.2245052,2.4058013,2.5852847,2.764768,2.9442513,3.1255474,2.8844235,2.6451125,2.4058013,2.1646774,1.9253663,1.6316663,1.3397794,1.0478923,0.7541924,0.46230546,0.6327239,0.8031424,0.97174793,1.1421664,1.3125849,1.260009,1.2074331,1.1548572,1.1022812,1.0497054,0.9572442,0.86478317,0.77232206,0.67986095,0.5873999,0.76325727,0.93730164,1.1131591,1.2872034,1.4630609,1.9326181,2.4021754,2.8717327,3.343103,3.8126602,3.780027,3.7473936,3.7147603,3.682127,3.6494937,4.7300196,5.810545,6.889258,7.9697833,9.050309,8.656897,8.265296,7.8718834,7.4802837,7.0868707,7.6724577,8.258044,8.841819,9.427405,10.012992,9.119202,8.227224,7.3352466,6.4432693,5.5494785,4.780782,4.0102735,3.2397642,2.469255,1.7005589,2.0051367,2.3097143,2.6142921,2.9206827,3.2252605,3.7473936,4.269527,4.7916603,5.315606,5.8377395,5.638314,5.4370747,5.237649,5.038223,4.836984,5.540414,6.24203,6.94546,7.647076,8.350506,8.444779,8.540867,8.63514,8.729415,8.825501,9.184468,9.545248,9.904215,10.264994,10.625773,12.186734,13.749508,15.312282,16.875055,18.43783,18.430578,18.423326,18.41426,18.40701,18.399757,16.405499,14.409427,12.415168,10.420909,8.424837,7.473032,6.5194135,5.567608,4.615803,3.6621845,4.3982472,5.132497,5.866747,6.60281,7.3370595,8.437528,9.537996,10.636651,11.73712,12.837588,15.649493,18.463211,21.275116,24.08702,26.90074,25.312584,23.724428,22.138086,20.54993,18.961775,16.64481,14.327844,12.009064,9.692098,7.3751316,6.970841,6.5647373,6.1604466,5.754343,5.3500524,4.688321,4.024777,3.3630457,2.6995013,2.03777,1.7295663,1.4231756,1.114972,0.80676836,0.50037766,0.58014804,0.65991837,0.73968875,0.8194591,0.89922947,0.7306239,0.56020546,0.38978696,0.21936847,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.052575916,0.054388877,0.058014803,0.059827764,0.06164073,0.11240368,0.16316663,0.21211663,0.26287958,0.31182957,0.5620184,0.8122072,1.062396,1.3125849,1.5627737,1.54827,1.5319533,1.5174497,1.502946,1.4866294,2.1773682,2.8681068,3.5570326,4.2477713,4.936697,5.903006,6.867502,7.8319983,8.798307,9.762803,14.06315,13.687867,13.312584,12.937301,12.562017,12.186734,11.537694,10.88684,10.2378,9.5869465,8.937905,8.399456,7.8628187,7.324369,6.787732,6.249282,6.1749506,6.1006193,6.0244746,5.9501433,5.8758116,6.011784,6.149569,6.2873545,6.4251394,6.5629244,6.450521,6.338117,6.2257137,6.11331,6.000906,5.712645,5.424384,5.137936,4.8496747,4.5632267,4.3746786,4.1879435,3.9993954,3.8126602,3.6241121,3.4754493,3.3249733,3.1744974,3.0258346,2.8753586,2.8499773,2.8245957,2.7992141,2.7756457,2.7502642,2.6505513,2.5508385,2.4493124,2.3495996,2.2498865,1.8383441,1.4249886,1.0116332,0.6000906,0.18673515,0.25018883,0.31182957,0.37528324,0.43692398,0.50037766,0.8883517,1.2745126,1.6624867,2.0504606,2.4366217,2.08672,1.7368182,1.3869164,1.0370146,0.6871128,0.61278135,0.53663695,0.46230546,0.387974,0.31182957,1.0877775,1.8619126,2.6378605,3.4119956,4.1879435,3.350355,2.5127661,1.6751775,0.8375887,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.8256533,3.6494937,5.475147,7.3008003,9.12464,8.149267,7.175706,6.200332,5.224958,4.249584,3.3993049,2.5508385,1.7005589,0.85027945,0.0,0.12509441,0.25018883,0.37528324,0.50037766,0.62547207,0.7124943,0.7995165,0.8883517,0.97537386,1.062396,1.0750868,1.0877775,1.1004683,1.1131591,1.1258497,0.93730164,0.7505665,0.5620184,0.37528324,0.18673515,0.2991388,0.41335547,0.52575916,0.63816285,0.7505665,1.1747998,1.6008459,2.0250793,2.4493124,2.8753586,3.199879,3.5243993,3.8507326,4.175253,4.499773,4.2006345,3.8996825,3.6005437,3.299592,3.000453,2.712192,2.4257438,2.137483,1.8492218,1.5627737,1.9996977,2.4366217,2.8753586,3.3122826,3.7492065,5.2630305,6.775041,8.287052,9.800876,11.312886,11.47424,11.637406,11.800573,11.961927,12.125093,11.162411,10.199727,9.237044,8.274362,7.311678,7.124943,6.9382076,6.7496595,6.5629244,6.3743763,6.0625467,5.750717,5.4370747,5.125245,4.8116026,4.361988,3.9123733,3.4627585,3.0131438,2.561716,2.1121013,1.6624867,1.2128719,0.76325727,0.31182957,0.25018883,0.18673515,0.12509441,0.06164073,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.099712946,0.19942589,0.2991388,0.40066472,0.50037766,0.5620184,0.62547207,0.6871128,0.7505665,0.8122072,0.6508536,0.48768693,0.3245203,0.16316663,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13778515,0.2755703,0.41335547,0.5493277,0.6871128,0.73787576,0.7868258,0.8375887,0.8883517,0.93730164,0.97537386,1.0116332,1.0497054,1.0877775,1.1258497,1.3506571,1.5754645,1.8002719,2.0250793,2.2498865,2.1991236,2.1501737,2.0994108,2.0504606,1.9996977,2.324218,2.6505513,2.9750717,3.299592,3.6241121,3.4246864,3.2252605,3.0258346,2.8245957,2.6251698,2.9007401,3.1744974,3.4500678,3.7256382,3.9993954,4.40006,4.800725,5.199577,5.600241,6.000906,6.011784,6.0244746,6.037165,6.049856,6.0625467,5.975525,5.8866897,5.7996674,5.712645,5.6256227,6.350808,7.07418,7.799365,8.52455,9.249735,13.026136,16.800724,20.575312,24.349901,28.124489,24.712494,21.300497,17.886688,14.474693,11.062697,11.361836,11.662788,11.961927,12.262879,12.562017,12.07433,11.586644,11.10077,10.613083,10.125396,9.050309,7.9752226,6.9001355,5.825049,4.749962,5.4370747,6.1241875,6.813113,7.500226,8.187339,7.8882003,7.5872483,7.28811,6.987158,6.688019,5.3627434,4.0374675,2.712192,1.3869164,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.41335547,0.824898,1.2382535,1.649796,2.0631514,1.887294,1.7132497,1.5373923,1.3633479,1.1874905,1.2001812,1.2128719,1.2255627,1.2382535,1.2491312,1.1004683,0.9499924,0.7995165,0.6508536,0.50037766,0.69980353,0.89922947,1.1004683,1.2998942,1.49932,1.4503701,1.3996071,1.3506571,1.2998942,1.2491312,1.1004683,0.9499924,0.7995165,0.6508536,0.50037766,0.72518504,0.9499924,1.1747998,1.3996071,1.6244144,2.1121013,2.5997884,3.0874753,3.5751622,4.062849,4.0374675,4.0120864,3.9867048,3.9631362,3.9377546,5.137936,6.338117,7.5382986,8.736667,9.936848,9.412902,8.887142,8.363196,7.837437,7.311678,8.024173,8.736667,9.449161,10.161655,10.874149,9.750113,8.624263,7.500226,6.3743763,5.2503395,4.4508233,3.6494937,2.8499773,2.0504606,1.2491312,1.6244144,1.9996977,2.374981,2.7502642,3.1255474,3.8126602,4.499773,5.186886,5.8758116,6.5629244,6.399758,6.2384043,6.0752378,5.9120708,5.750717,6.450521,7.1503243,7.850128,8.549932,9.249735,9.012237,8.774739,8.537241,8.299743,8.062244,8.774739,9.487233,10.199727,10.912222,11.624716,13.212872,14.799213,16.38737,17.975525,19.561867,19.786674,20.013294,20.238102,20.462908,20.687716,18.20033,15.712947,13.225562,10.738177,8.2507925,6.9382076,5.6256227,4.313038,3.000453,1.6878681,2.2498865,2.811905,3.3757362,3.9377546,4.499773,5.763408,7.02523,8.287052,9.550687,10.812509,14.675932,18.537542,22.400965,26.262575,30.124186,28.66294,27.199877,25.736816,24.27557,22.812508,19.899076,16.98746,14.074029,11.162411,8.2507925,7.5618668,6.874754,6.187641,5.5005283,4.8116026,4.1498713,3.48814,2.8245957,2.1628644,1.49932,1.2491312,1.0007553,0.7505665,0.50037766,0.25018883,0.42423326,0.6000906,0.774135,0.9499924,1.1258497,0.9119202,0.69980353,0.48768693,0.2755703,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.11240368,0.16316663,0.21211663,0.26287958,0.31182957,0.5747091,0.8375887,1.1004683,1.3633479,1.6244144,1.5881553,1.550083,1.5120108,1.4757515,1.4376793,2.2245052,3.0131438,3.7999697,4.5867953,5.375434,5.863121,6.350808,6.836682,7.324369,7.8120556,15.263332,14.777458,14.293397,13.807523,13.321649,12.837588,12.077957,11.318325,10.556881,9.79725,9.037619,8.42665,7.817495,7.208339,6.5973706,5.9882154,5.903006,5.8177967,5.732588,5.6473784,5.562169,5.7072062,5.8522434,5.99728,6.1423173,6.2873545,6.240217,6.19308,6.14413,6.096993,6.049856,6.000906,5.9501433,5.89938,5.8504305,5.7996674,5.542227,5.2847857,5.027345,4.7699046,4.512464,4.2368937,3.9631362,3.6875658,3.4119956,3.1382382,3.1708715,3.2016919,3.2343252,3.2669585,3.299592,3.2216346,3.1454902,3.0675328,2.9895754,2.913431,2.5907235,2.268016,1.9453088,1.6226015,1.2998942,1.3742256,1.4503701,1.5247015,1.6008459,1.6751775,2.079468,2.4855716,2.8898623,3.295966,3.7002566,3.3630457,3.0258346,2.6868105,2.3495996,2.0123885,1.9181144,1.8220274,1.7277533,1.6334792,1.5373923,2.0432088,2.5472124,3.053029,3.5570326,4.062849,3.6531196,3.24339,2.8318477,2.422118,2.0123885,1.8075237,1.6026589,1.3977941,1.1929294,0.9880646,0.79589057,0.60190356,0.40972954,0.21755551,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,1.5917811,3.159994,4.7282066,6.294606,7.8628187,7.0016613,6.1423173,5.282973,4.421816,3.5624714,2.8517902,2.1429217,1.4322405,0.72337204,0.012690738,0.11059072,0.20667773,0.3045777,0.40247768,0.50037766,0.56927025,0.6399758,0.7106813,0.7795739,0.85027945,0.86478317,0.8792868,0.89560354,0.9101072,0.9246109,0.8466535,0.7705091,0.69255173,0.61459434,0.53663695,0.6852999,0.8321498,0.9808127,1.1276628,1.2745126,2.039583,2.8046532,3.5697234,4.3347936,5.0998635,5.0744824,5.050914,5.0255322,5.0001507,4.974769,4.59586,4.215138,3.834416,3.4555066,3.0747845,2.8844235,2.6958754,2.5055144,2.3151531,2.124792,2.6723068,3.2198215,3.7673361,4.314851,4.8623657,5.9356394,7.0071006,8.080374,9.151835,10.225109,10.324821,10.424535,10.524248,10.625773,10.725487,9.935035,9.144584,8.354132,7.5654926,6.775041,6.439643,6.104245,5.77066,5.4352617,5.0998635,4.8496747,4.599486,4.349297,4.099108,3.8507326,3.489953,3.1291735,2.770207,2.4094272,2.0504606,1.6896812,1.3307146,0.969935,0.6091554,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07977036,0.15954071,0.23931105,0.3208944,0.40066472,0.44961473,0.50037766,0.5493277,0.6000906,0.6508536,0.52032024,0.38978696,0.25925365,0.13053331,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.018129626,0.034446288,0.052575916,0.07070554,0.0870222,0.14503701,0.2030518,0.25925365,0.31726846,0.37528324,0.51306844,0.6508536,0.7868258,0.9246109,1.062396,1.1095331,1.1566701,1.2056202,1.2527572,1.2998942,1.452183,1.6044719,1.7567607,1.9108626,2.0631514,2.1102884,2.1574254,2.2045624,2.2516994,2.3006494,2.2172532,2.13567,2.0522738,1.9706904,1.887294,2.1683033,2.4474995,2.7266958,3.007705,3.2869012,3.2216346,3.1581807,3.092914,3.0276475,2.962381,3.3757362,3.787279,4.2006345,4.612177,5.0255322,5.230397,5.4352617,5.6401267,5.844991,6.049856,5.9483304,5.844991,5.7416525,5.6401267,5.5367875,5.3573046,5.177821,4.9983377,4.8170414,4.6375585,5.732588,6.827617,7.9226465,9.017676,10.112705,13.185677,16.256836,19.329807,22.402779,25.473938,22.562319,19.650702,16.73727,13.825653,10.912222,11.156972,11.401722,11.648285,11.893035,12.137785,11.592083,11.048194,10.502492,9.956791,9.412902,8.756609,8.10213,7.4476504,6.793171,6.1368785,6.7097745,7.2826705,7.855567,8.428463,8.999546,8.531802,8.06587,7.5981264,7.130382,6.6626377,5.3645563,4.068288,2.770207,1.4721256,0.17585737,0.14684997,0.11965553,0.092461094,0.065266654,0.038072214,0.3680314,0.6979906,1.0279498,1.357909,1.6878681,1.5555218,1.4231756,1.2908293,1.1566701,1.0243238,1.0370146,1.0497054,1.062396,1.0750868,1.0877775,0.9572442,0.82671094,0.6979906,0.56745726,0.43692398,0.6091554,0.78319985,0.9554313,1.1276628,1.2998942,1.3397794,1.3796645,1.4195497,1.4594349,1.49932,1.4576219,1.4159238,1.3724127,1.3307146,1.2872034,1.504759,1.7223145,1.93987,2.1574254,2.374981,2.8245957,3.2742105,3.7256382,4.175253,4.6248674,4.6593137,4.695573,4.7300196,4.764466,4.800725,5.7869763,6.775041,7.763106,8.749357,9.737422,9.340384,8.943344,8.544493,8.147454,7.750415,8.557183,9.365765,10.172533,10.979301,11.787883,10.830639,9.873394,8.914337,7.957093,6.9998484,5.922949,4.844236,3.7673361,2.6904364,1.6117238,2.0232663,2.4329958,2.8427253,3.2524548,3.6621845,4.4852695,5.3083544,6.1296263,6.9527116,7.7757964,7.752228,7.7304726,7.706904,7.6851482,7.663393,8.025986,8.386765,8.749357,9.11195,9.474543,9.382081,9.28962,9.197159,9.104698,9.012237,9.947725,10.883214,11.81689,12.752378,13.687867,14.639673,15.593291,16.545097,17.496902,18.45052,18.671701,18.894695,19.117691,19.340685,19.561867,17.513218,15.462758,13.412297,11.361836,9.313189,8.174648,7.037921,5.89938,4.762653,3.625925,3.9848917,4.345671,4.704638,5.0654173,5.424384,6.510349,7.5945,8.680465,9.764616,10.850581,14.003323,17.154251,20.306993,23.459736,26.612478,25.163921,23.717176,22.270432,20.821875,19.375132,16.956638,14.53996,12.121468,9.704789,7.28811,6.6499467,6.011784,5.375434,4.7372713,4.099108,3.5225863,2.9442513,2.3677292,1.789394,1.2128719,1.0279498,0.8430276,0.65810543,0.47318324,0.28826106,0.5275721,0.7668832,1.0080072,1.2473183,1.4866294,1.2418793,0.99712944,0.7523795,0.5076295,0.26287958,0.25925365,0.2574407,0.25562772,0.2520018,0.25018883,0.21211663,0.17585737,0.13778515,0.099712946,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.06707962,0.072518505,0.07795739,0.08339628,0.0870222,0.12509441,0.16316663,0.19942589,0.2374981,0.2755703,0.49675176,0.7197462,0.94274056,1.1657349,1.3869164,1.4449311,1.502946,1.5591478,1.6171626,1.6751775,2.2843328,2.8953013,3.5044568,4.115425,4.7245803,5.658256,6.590119,7.5219817,8.455658,9.38752,16.4617,15.867048,15.272397,14.677745,14.083094,13.486629,12.618219,11.747997,10.877775,10.007553,9.137331,8.455658,7.7721705,7.0904965,6.4070096,5.7253356,5.6292486,5.5349746,5.4407005,5.3446136,5.2503395,5.4026284,5.5549173,5.7072062,5.859495,6.011784,6.0299134,6.0480433,6.0643597,6.0824895,6.1006193,6.2873545,6.474089,6.6626377,6.849373,7.037921,6.7097745,6.3816285,6.055295,5.727149,5.4008155,5.0001507,4.599486,4.2006345,3.7999697,3.3993049,3.489953,3.5806012,3.6694362,3.7600844,3.8507326,3.7945306,3.7401419,3.6857529,3.6295512,3.5751622,3.343103,3.1092308,2.8771715,2.6451125,2.4130533,2.5000753,2.5870976,2.6741197,2.762955,2.8499773,3.2723975,3.6948178,4.117238,4.539658,4.9620786,4.6375585,4.313038,3.9867048,3.6621845,3.3376641,3.2216346,3.1074178,2.9932013,2.8771715,2.762955,2.9968271,3.2325122,3.4681973,3.7020695,3.9377546,3.9558845,3.972201,3.9903307,4.006647,4.024777,3.6150475,3.2053177,2.7955883,2.3858588,1.9743162,1.5899682,1.2056202,0.8194591,0.43511102,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,1.3597219,2.6704938,3.9794528,5.290225,6.599184,5.8558693,5.1107416,4.365614,3.6204863,2.8753586,2.3042755,1.7350051,1.1657349,0.5946517,0.025381476,0.09427405,0.16497959,0.23568514,0.3045777,0.37528324,0.42785916,0.48043507,0.533011,0.5855869,0.63816285,0.6544795,0.6726091,0.69073874,0.7070554,0.72518504,0.75781834,0.7904517,0.823085,0.8557183,0.8883517,1.0696479,1.2527572,1.4358664,1.6171626,1.8002719,2.904366,4.0102735,5.1143675,6.2202744,7.324369,6.9490857,6.5756154,6.200332,5.825049,5.4497657,4.989273,4.5305934,4.070101,3.6096084,3.149116,3.056655,2.9641938,2.8717327,2.7792716,2.6868105,3.3449159,4.0030212,4.6593137,5.317419,5.975525,6.6082487,7.2391596,7.8718834,8.504607,9.137331,9.175404,9.211663,9.249735,9.287807,9.325879,8.70766,8.089439,7.473032,6.8548117,6.2384043,5.754343,5.272095,4.7898474,4.307599,3.825351,3.636803,3.4500678,3.2633326,3.0747845,2.8880494,2.617918,2.3477864,2.077655,1.8075237,1.5373923,1.2672608,0.99712944,0.726998,0.45686656,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.059827764,0.11965553,0.1794833,0.23931105,0.2991388,0.33721104,0.37528324,0.41335547,0.44961473,0.48768693,0.38978696,0.291887,0.19579996,0.09789998,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.034446288,0.07070554,0.10515183,0.13959812,0.17585737,0.29007402,0.40429065,0.52032024,0.6345369,0.7505665,0.8883517,1.0243238,1.162109,1.2998942,1.4376793,1.4830034,1.5283275,1.5718386,1.6171626,1.6624867,1.9308052,2.1973107,2.465629,2.7321346,3.000453,2.8699198,2.7393866,2.610666,2.4801328,2.3495996,2.2353828,2.1193533,2.0051367,1.889107,1.7748904,2.0105755,2.2444477,2.4801328,2.715818,2.94969,3.0203958,3.0892882,3.159994,3.2306993,3.299592,3.8507326,4.40006,4.949388,5.5005283,6.049856,6.060734,6.069799,6.0806766,6.089741,6.1006193,5.883064,5.6655083,5.4479527,5.230397,5.0128417,4.740897,4.4671397,4.195195,3.923251,3.6494937,5.1143675,6.5792413,8.045928,9.510801,10.975676,13.345218,15.71476,18.084301,20.455656,22.8252,20.412146,18.000906,15.5878525,13.174799,10.761745,10.952107,11.142468,11.332829,11.5231905,11.711739,11.109835,10.507931,9.904215,9.302311,8.700407,8.464723,8.23085,7.995165,7.75948,7.5256076,7.9824743,8.439341,8.898021,9.354887,9.811753,9.177217,8.54268,7.9081426,7.271793,6.637256,5.368182,4.0972953,2.8282216,1.5573349,0.28826106,0.24474995,0.2030518,0.15954071,0.11784257,0.07433146,0.32270733,0.56927025,0.81764615,1.064209,1.3125849,1.2219368,1.1331016,1.0424535,0.95180535,0.8629702,0.87566096,0.8883517,0.89922947,0.9119202,0.9246109,0.81583315,0.70524246,0.5946517,0.48587397,0.37528324,0.52032024,0.6653573,0.8103943,0.9554313,1.1004683,1.2291887,1.3597219,1.4902552,1.6207886,1.7495089,1.8147756,1.8800422,1.9453088,2.0105755,2.0758421,2.2843328,2.4946365,2.70494,2.9152439,3.1255474,3.53709,3.9504454,4.361988,4.7753434,5.186886,5.282973,5.377247,5.473334,5.567608,5.661882,6.43783,7.211965,7.987913,8.762048,9.537996,9.267865,8.997733,8.727602,8.457471,8.187339,9.090195,9.99305,10.8959055,11.7969475,12.699803,11.909351,11.120712,10.330261,9.539809,8.749357,7.3950744,6.0407915,4.6846952,3.3304121,1.9743162,2.420305,2.864481,3.3104696,3.7546456,4.2006345,5.1578784,6.115123,7.072367,8.029612,8.9868555,9.104698,9.222541,9.340384,9.458226,9.574255,9.599637,9.625018,9.6504,9.675781,9.699349,9.751925,9.804502,9.857078,9.909654,9.96223,11.120712,12.277383,13.435865,14.592536,15.749206,16.068287,16.385555,16.702824,17.020092,17.33736,17.55673,17.77791,17.99728,18.216648,18.43783,16.824293,15.212569,13.600845,11.9873085,10.375585,9.412902,8.450218,7.4875355,6.5248523,5.562169,5.719897,5.8776245,6.035352,6.19308,6.350808,7.2572894,8.165584,9.072064,9.980359,10.88684,13.330714,15.772775,18.214834,20.656897,23.100769,21.666716,20.234476,18.802235,17.369995,15.937754,14.014201,12.092461,10.17072,8.247167,6.3254266,5.7380266,5.1506267,4.5632267,3.975827,3.388427,2.8953013,2.4021754,1.9108626,1.4177368,0.9246109,0.80495536,0.6852999,0.5656443,0.44417584,0.3245203,0.630911,0.9354887,1.2400664,1.5446441,1.8492218,1.5718386,1.2944553,1.017072,0.73968875,0.46230546,0.46955732,0.47680917,0.48587397,0.49312583,0.50037766,0.42423326,0.34990177,0.2755703,0.19942589,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.072518505,0.08339628,0.092461094,0.10333887,0.11240368,0.13778515,0.16316663,0.18673515,0.21211663,0.2374981,0.42060733,0.60190356,0.7850128,0.968122,1.1494182,1.3017071,1.455809,1.6080978,1.7603867,1.9126755,2.3441606,2.7774587,3.2107568,3.6422417,4.07554,5.4533916,6.82943,8.207282,9.585134,10.962985,17.661882,16.956638,16.25321,15.547967,14.842725,14.137483,13.15667,12.17767,11.1968565,10.217857,9.237044,8.482852,7.7268467,6.972654,6.2166486,5.462456,5.3573046,5.2521524,5.147001,5.041849,4.936697,5.0980506,5.2575917,5.4171324,5.576673,5.7380266,5.81961,5.903006,5.9845896,6.0679855,6.149569,6.5756154,6.9998484,7.4258947,7.850128,8.274362,7.877322,7.4802837,7.083245,6.684393,6.2873545,5.763408,5.237649,4.7118897,4.1879435,3.6621845,3.8108473,3.9576974,4.1045475,4.25321,4.40006,4.367427,4.3347936,4.3021603,4.269527,4.2368937,4.0954823,3.9522583,3.8108473,3.6676233,3.5243993,3.625925,3.7256382,3.825351,3.925064,4.024777,4.465327,4.9058766,5.3446136,5.7851634,6.2257137,5.9120708,5.600241,5.2884116,4.974769,4.6629395,4.5269675,4.3928084,4.256836,4.122677,3.9867048,3.9522583,3.917812,3.8833659,3.8471067,3.8126602,4.256836,4.702825,5.147001,5.5929894,6.037165,5.422571,4.8079767,4.1933823,3.576975,2.962381,2.3858588,1.8075237,1.2291887,0.6526665,0.07433146,0.07433146,0.07433146,0.07433146,0.07433146,0.07433146,1.1276628,2.179181,3.2325122,4.2858434,5.337362,4.708264,4.077353,3.4482548,2.817344,2.1882458,1.7567607,1.3270886,0.8974165,0.46774435,0.038072214,0.07977036,0.12328146,0.16497959,0.20667773,0.25018883,0.28463513,0.3208944,0.35534066,0.38978696,0.42423326,0.44417584,0.46411842,0.48587397,0.5058166,0.52575916,0.6671702,0.8103943,0.95180535,1.0950294,1.2382535,1.455809,1.6733645,1.8909199,2.1066625,2.324218,3.7691493,5.2158933,6.6608243,8.105756,9.550687,8.825501,8.100317,7.3751316,6.6499467,5.924762,5.384499,4.844236,4.305786,3.7655232,3.2252605,3.2306993,3.2343252,3.2397642,3.245203,3.2506418,4.017525,4.784408,5.5531044,6.319988,7.0868707,7.2808576,7.473032,7.665206,7.85738,8.049554,8.024173,8.000604,7.9752226,7.949841,7.9244595,7.4802837,7.0342946,6.590119,6.14413,5.6999545,5.0708566,4.439945,3.8108473,3.1799364,2.5508385,2.4257438,2.3006494,2.175555,2.0504606,1.9253663,1.74407,1.5645868,1.3851035,1.2056202,1.0243238,0.8448406,0.6653573,0.48587397,0.3045777,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03988518,0.07977036,0.11965553,0.15954071,0.19942589,0.22480737,0.25018883,0.2755703,0.2991388,0.3245203,0.25925365,0.19579996,0.13053331,0.065266654,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.052575916,0.10515183,0.15772775,0.21030366,0.26287958,0.43511102,0.6073425,0.7795739,0.95180535,1.1258497,1.261822,1.3996071,1.5373923,1.6751775,1.8129625,1.8546607,1.8981718,1.93987,1.983381,2.0250793,2.4076142,2.7901495,3.1726844,3.5552197,3.9377546,3.6295512,3.3231604,3.0149567,2.7067533,2.4003625,2.2516994,2.1048496,1.9579996,1.8093367,1.6624867,1.8528478,2.0432088,2.231757,2.422118,2.612479,2.817344,3.0222087,3.2270734,3.4319382,3.636803,4.325729,5.0128417,5.6999545,6.3870673,7.07418,6.889258,6.7043357,6.5194135,6.3344913,6.149569,5.8177967,5.484212,5.1524396,4.8206677,4.4870825,4.122677,3.7582715,3.392053,3.0276475,2.663242,4.49796,6.3326783,8.167397,10.002114,11.836833,13.504758,15.172684,16.840609,18.506721,20.174648,18.261972,16.349297,14.436621,12.525759,10.613083,10.747242,10.883214,11.017374,11.153346,11.287505,10.627586,9.967669,9.30775,8.647832,7.987913,8.172835,8.357758,8.54268,8.727602,8.912524,9.255174,9.597824,9.940474,10.283124,10.625773,9.822631,9.019489,8.21816,7.415017,6.6118746,5.369995,4.1281157,2.8844235,1.6425442,0.40066472,0.34264994,0.28463513,0.22662032,0.17041849,0.11240368,0.27738327,0.44236287,0.6073425,0.77232206,0.93730164,0.8901646,0.8430276,0.79589057,0.7469406,0.69980353,0.7124943,0.72518504,0.73787576,0.7505665,0.76325727,0.6726091,0.581961,0.49312583,0.40247768,0.31182957,0.42967212,0.5475147,0.6653573,0.78319985,0.89922947,1.1204109,1.3397794,1.5591478,1.7803292,1.9996977,2.1719291,2.3441606,2.518205,2.6904364,2.8626678,3.0657198,3.2669585,3.4700103,3.673062,3.874301,4.249584,4.6248674,5.0001507,5.375434,5.750717,5.904819,6.060734,6.2148356,6.3707504,6.5248523,7.0868707,7.650702,8.212721,8.774739,9.336758,9.195346,9.052122,8.910711,8.767487,8.624263,9.623205,10.620335,11.617464,12.6145935,13.611723,12.989877,12.368031,11.744371,11.122525,10.500679,8.8672,7.2355337,5.6020546,3.9703882,2.3369088,2.817344,3.2977788,3.778214,4.256836,4.7372713,5.8304877,6.921891,8.015107,9.108324,10.199727,10.457169,10.714609,10.97205,11.22949,11.486931,11.175101,10.863272,10.549629,10.2378,9.924157,10.12177,10.319383,10.516996,10.714609,10.912222,12.291886,13.673364,15.053028,16.432693,17.812357,17.495089,17.17782,16.860552,16.543283,16.224201,16.441757,16.659313,16.87687,17.094423,17.31198,16.13718,14.96238,13.7875805,12.612781,11.437981,10.649343,9.862516,9.07569,8.287052,7.500226,7.454902,7.409578,7.364254,7.320743,7.2754188,8.00423,8.734854,9.465478,10.194288,10.924912,12.658105,14.389484,16.122677,17.854055,19.587248,18.169512,16.751774,15.334038,13.918114,12.500377,11.071762,9.644961,8.21816,6.789545,5.3627434,4.8242936,4.2876563,3.7492065,3.2125697,2.6741197,2.268016,1.8600996,1.452183,1.0442665,0.63816285,0.581961,0.5275721,0.47318324,0.4169814,0.36259252,0.7324369,1.1022812,1.4721256,1.84197,2.2118144,1.9017978,1.5917811,1.2817645,0.97174793,0.66173136,0.67986095,0.6979906,0.71430725,0.7324369,0.7505665,0.63816285,0.52575916,0.41335547,0.2991388,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.07795739,0.092461094,0.10696479,0.12328146,0.13778515,0.15047589,0.16316663,0.17585737,0.18673515,0.19942589,0.34264994,0.48587397,0.62728506,0.7705091,0.9119202,1.1602961,1.4068589,1.6552348,1.9017978,2.1501737,2.4058013,2.659616,2.9152439,3.1708715,3.4246864,5.2467136,7.0705543,8.892582,10.714609,12.538449,18.862062,18.048042,17.23221,16.41819,15.602356,14.788336,13.696932,12.607342,11.517752,10.428161,9.336758,8.510046,7.6833353,6.8548117,6.0281005,5.199577,5.08536,4.9693303,4.855114,4.740897,4.6248674,4.7916603,4.9602656,5.127058,5.295664,5.462456,5.6093063,5.7579694,5.904819,6.051669,6.200332,6.8620634,7.5256076,8.187339,8.8508835,9.512614,9.04487,8.577126,8.109382,7.6416373,7.175706,6.5248523,5.8758116,5.224958,4.574105,3.925064,4.1299286,4.3347936,4.539658,4.744523,4.949388,4.940323,4.9294453,4.9203806,4.9095025,4.900438,4.847862,4.795286,4.74271,4.690134,4.6375585,4.749962,4.8623657,4.974769,5.087173,5.199577,5.658256,6.115123,6.5719895,7.0306687,7.4875355,7.1883965,6.887445,6.588306,6.2873545,5.9882154,5.8323007,5.678199,5.522284,5.368182,5.2122674,4.9076896,4.603112,4.2967215,3.9921436,3.6875658,4.559601,5.431636,6.305484,7.177519,8.049554,7.230095,6.4106355,5.5893636,4.7699046,3.9504454,3.1799364,2.4094272,1.6407311,0.87022203,0.099712946,0.099712946,0.099712946,0.099712946,0.099712946,0.099712946,0.89560354,1.6896812,2.4855716,3.2796493,4.07554,3.5606585,3.045777,2.5290828,2.0142014,1.49932,1.209246,0.91917205,0.629098,0.34083697,0.05076295,0.065266654,0.07977036,0.09427405,0.11059072,0.12509441,0.14322405,0.15954071,0.17767033,0.19579996,0.21211663,0.23568514,0.2574407,0.27919623,0.30276474,0.3245203,0.57833505,0.83033687,1.0823387,1.3343405,1.5881553,1.840157,2.0921588,2.3441606,2.5979755,2.8499773,4.6357455,6.4197006,8.205468,9.989424,11.775192,10.700105,9.625018,8.549932,7.474845,6.399758,5.7797246,5.1596913,4.539658,3.919625,3.299592,3.4029307,3.5044568,3.6077955,3.7093215,3.8126602,4.690134,5.567608,6.445082,7.322556,8.200029,7.951654,7.705091,7.456715,7.210152,6.9617763,6.874754,6.787732,6.70071,6.6118746,6.5248523,6.2529078,5.979151,5.7072062,5.4352617,5.163317,4.3855567,3.6077955,2.8300345,2.0522738,1.2745126,1.2128719,1.1494182,1.0877775,1.0243238,0.96268314,0.872035,0.78319985,0.69255173,0.60190356,0.51306844,0.4224203,0.33177215,0.24293698,0.15228885,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.11240368,0.12509441,0.13778515,0.15047589,0.16316663,0.13053331,0.09789998,0.065266654,0.032633327,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07070554,0.13959812,0.21030366,0.27919623,0.34990177,0.58014804,0.8103943,1.0406405,1.2708868,1.49932,1.6371052,1.7748904,1.9126755,2.0504606,2.1882458,2.228131,2.268016,2.3079014,2.3477864,2.3876717,2.8844235,3.3829882,3.87974,4.3783045,4.8750563,4.3891826,3.9051213,3.4192474,2.9351864,2.4493124,2.269829,2.0903459,1.9108626,1.7295663,1.550083,1.69512,1.840157,1.9851941,2.1302311,2.275268,2.6142921,2.955129,3.294153,3.63499,3.975827,4.800725,5.6256227,6.450521,7.2754188,8.100317,7.7195945,7.3406854,6.9599633,6.5792413,6.200332,5.75253,5.3047285,4.856927,4.409125,3.9631362,3.5044568,3.04759,2.5907235,2.132044,1.6751775,3.87974,6.0843024,8.290678,10.49524,12.699803,13.664299,14.630608,15.595104,16.5596,17.524096,16.1118,14.699501,13.287203,11.874905,10.462607,10.542377,10.622148,10.701918,10.781689,10.863272,10.145339,9.427405,8.709473,7.993352,7.2754188,7.8791356,8.484665,9.090195,9.695724,10.29944,10.527874,10.754494,10.982927,11.209548,11.437981,10.468046,9.498111,8.528176,7.558241,6.588306,5.371808,4.157123,2.9424384,1.7277533,0.51306844,0.4405499,0.3680314,0.2955129,0.2229944,0.15047589,0.23205921,0.3154555,0.39703882,0.48043507,0.5620184,0.55839247,0.5529536,0.5475147,0.5420758,0.53663695,0.5493277,0.5620184,0.5747091,0.5873999,0.6000906,0.5293851,0.4604925,0.38978696,0.3208944,0.25018883,0.34083697,0.42967212,0.52032024,0.6091554,0.69980353,1.0098201,1.3198367,1.6298534,1.93987,2.2498865,2.5308957,2.810092,3.0892882,3.3702974,3.6494937,3.8452935,4.0392804,4.2350807,4.4308805,4.6248674,4.9620786,5.2992897,5.638314,5.975525,6.3127356,6.526665,6.742408,6.9581504,7.17208,7.3878226,7.7377243,8.087626,8.437528,8.78743,9.137331,9.122828,9.108324,9.092008,9.077503,9.063,10.154404,11.24762,12.340837,13.43224,14.525456,14.070402,13.615349,13.1602955,12.705242,12.250188,10.339326,8.430276,6.5194135,4.610364,2.6995013,3.2143826,3.729264,4.2441454,4.76084,5.275721,6.5030966,7.7304726,8.957849,10.185224,11.4126,11.809638,12.206677,12.605529,13.002567,13.399607,12.750566,12.099712,11.450671,10.799818,10.150778,10.493427,10.834265,11.176914,11.519565,11.862214,13.464873,15.067532,16.67019,18.27285,19.87551,18.92189,17.970085,17.01828,16.064661,15.112856,15.326786,15.542528,15.758271,15.9722,16.187943,15.4500675,14.712192,13.974316,13.238253,12.500377,11.887595,11.274815,10.662033,10.049252,9.438283,9.189907,8.943344,8.694968,8.448405,8.200029,8.752983,9.304124,9.857078,10.410031,10.962985,11.985496,13.008006,14.030518,15.053028,16.075539,14.672306,13.270886,11.867653,10.46442,9.063,8.129324,7.1974616,6.265599,5.331923,4.40006,3.9123733,3.4246864,2.9369993,2.4493124,1.9616255,1.6407311,1.3180238,0.99531645,0.6726091,0.34990177,0.36077955,0.36984438,0.38072214,0.38978696,0.40066472,0.83577573,1.2708868,1.7041848,2.1392958,2.5744069,2.231757,1.8909199,1.54827,1.2056202,0.8629702,0.8901646,0.91735905,0.9445535,0.97174793,1.0007553,0.85027945,0.69980353,0.5493277,0.40066472,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.08339628,0.10333887,0.12328146,0.14322405,0.16316663,0.16316663,0.16316663,0.16316663,0.16316663,0.16316663,0.26469254,0.3680314,0.46955732,0.5728962,0.6744221,1.017072,1.3597219,1.7023718,2.0450218,2.3876717,2.465629,2.5417736,2.619731,2.6976883,2.7756457,5.041849,7.309865,9.577881,11.844085,14.112101,20.062244,19.137632,18.213022,17.286598,16.361988,15.437376,14.237195,13.037014,11.836833,10.636651,9.438283,8.537241,7.6380115,6.736969,5.8377395,4.936697,4.8116026,4.688321,4.5632267,4.4381323,4.313038,4.4870825,4.6629395,4.836984,5.0128417,5.186886,5.4008155,5.612932,5.825049,6.037165,6.249282,7.1503243,8.049554,8.950596,9.849826,10.750868,10.212419,9.675781,9.137331,8.600695,8.062244,7.28811,6.5121617,5.7380266,4.9620786,4.1879435,4.4508233,4.7118897,4.974769,5.237649,5.5005283,5.5132194,5.524097,5.5367875,5.5494785,5.562169,5.600241,5.638314,5.674573,5.712645,5.750717,5.8758116,5.999093,6.1241875,6.249282,6.3743763,6.849373,7.324369,7.799365,8.274362,8.749357,8.46291,8.174648,7.8882003,7.5999393,7.311678,7.137634,6.9617763,6.787732,6.6118746,6.43783,5.863121,5.2884116,4.7118897,4.137181,3.5624714,4.8623657,6.16226,7.462154,8.762048,10.061942,9.037619,8.013294,6.987158,5.962834,4.936697,3.975827,3.0131438,2.0504606,1.0877775,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.12509441,0.66173136,1.2001812,1.7368182,2.275268,2.811905,2.4130533,2.0123885,1.6117238,1.2128719,0.8122072,0.66173136,0.51306844,0.36259252,0.21211663,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.48768693,0.85027945,1.2128719,1.5754645,1.938057,2.2245052,2.5127661,2.7992141,3.0874753,3.3757362,5.5005283,7.6253204,9.750113,11.874905,13.999697,12.574709,11.14972,9.724731,8.299743,6.874754,6.1749506,5.475147,4.7753434,4.07554,3.3757362,3.5751622,3.774588,3.975827,4.175253,4.3746786,5.3627434,6.350808,7.3370595,8.325124,9.313189,8.624263,7.93715,7.250037,6.5629244,5.8758116,5.7253356,5.57486,5.424384,5.275721,5.125245,5.0255322,4.9258194,4.8242936,4.7245803,4.6248674,3.7002566,2.7756457,1.8492218,0.9246109,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0870222,0.17585737,0.26287958,0.34990177,0.43692398,0.72518504,1.0116332,1.2998942,1.5881553,1.8746033,2.0123885,2.1501737,2.2879589,2.4257438,2.561716,2.5997884,2.6378605,2.6741197,2.712192,2.7502642,3.3630457,3.975827,4.5867953,5.199577,5.812358,5.1506267,4.4870825,3.825351,3.1618068,2.5000753,2.2879589,2.0758421,1.8619126,1.649796,1.4376793,1.5373923,1.6371052,1.7368182,1.8383441,1.938057,2.4130533,2.8880494,3.3630457,3.8380418,4.313038,5.275721,6.2365913,7.1992745,8.161958,9.12464,8.549932,7.9752226,7.400513,6.825804,6.249282,5.6872635,5.125245,4.5632267,3.9993954,3.437377,2.8880494,2.3369088,1.7875811,1.2382535,0.6871128,3.2633326,5.8377395,8.412147,10.988366,13.562773,13.825653,14.0867195,14.349599,14.612478,14.875358,13.961625,13.049705,12.137785,11.225864,10.312131,10.337513,10.362894,10.388275,10.411844,10.437225,9.663091,8.887142,8.113008,7.3370595,6.5629244,7.5872483,8.611572,9.637709,10.662033,11.6881695,11.800573,11.912977,12.025381,12.137785,12.250188,11.111648,9.97492,8.838193,7.699652,6.5629244,5.375434,4.1879435,3.000453,1.8129625,0.62547207,0.53663695,0.44961473,0.36259252,0.2755703,0.18673515,0.18673515,0.18673515,0.18673515,0.18673515,0.18673515,0.22480737,0.26287958,0.2991388,0.33721104,0.37528324,0.387974,0.40066472,0.41335547,0.42423326,0.43692398,0.387974,0.33721104,0.28826106,0.2374981,0.18673515,0.25018883,0.31182957,0.37528324,0.43692398,0.50037766,0.89922947,1.2998942,1.7005589,2.0994108,2.5000753,2.8880494,3.2742105,3.6621845,4.0501585,4.4381323,4.6248674,4.8116026,5.0001507,5.186886,5.375434,5.674573,5.975525,6.2746634,6.5756154,6.874754,7.1503243,7.4258947,7.699652,7.9752226,8.2507925,8.386765,8.52455,8.662335,8.80012,8.937905,9.050309,9.162713,9.275117,9.38752,9.499924,10.687414,11.874905,13.062395,14.249886,15.437376,15.149116,14.862667,14.574407,14.287958,13.999697,11.813264,9.625018,7.4367723,5.2503395,3.0620937,3.6132345,4.162562,4.7118897,5.2630305,5.812358,7.175706,8.537241,9.900589,11.262123,12.625471,13.162108,13.700559,14.237195,14.775645,15.312282,14.324218,13.337966,12.349901,11.361836,10.375585,10.863272,11.349146,11.836833,12.32452,12.812206,14.63786,16.4617,18.287354,20.113007,21.936848,20.350506,18.76235,17.174194,15.5878525,13.999697,14.211814,14.425743,14.63786,14.849977,15.062093,14.762955,14.462003,14.162864,13.861912,13.562773,13.125849,12.687112,12.250188,11.813264,11.374527,10.924912,10.475298,10.025683,9.574255,9.12464,9.499924,9.875207,10.25049,10.625773,10.999244,11.312886,11.624716,11.938358,12.250188,12.562017,11.175101,9.788185,8.399456,7.0125394,5.6256227,5.186886,4.749962,4.313038,3.874301,3.437377,3.000453,2.561716,2.124792,1.6878681,1.2491312,1.0116332,0.774135,0.53663695,0.2991388,0.06164073,0.13778515,0.21211663,0.28826106,0.36259252,0.43692398,0.93730164,1.4376793,1.938057,2.4366217,2.9369993,2.561716,2.1882458,1.8129625,1.4376793,1.062396,1.1004683,1.1367276,1.1747998,1.2128719,1.2491312,1.062396,0.87566096,0.6871128,0.50037766,0.31182957,0.25018883,0.18673515,0.12509441,0.06164073,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.0870222,0.11240368,0.13778515,0.16316663,0.18673515,0.17585737,0.16316663,0.15047589,0.13778515,0.12509441,0.18673515,0.25018883,0.31182957,0.37528324,0.43692398,0.87566096,1.3125849,1.7495089,2.1882458,2.6251698,2.525457,2.4257438,2.324218,2.2245052,2.124792,4.836984,7.550989,10.263181,12.975373,15.687565,18.425138,18.729717,19.034294,19.340685,19.645262,19.94984,19.744976,19.540112,19.335245,19.13038,18.925516,17.698141,16.470764,15.243389,14.016014,12.788638,12.11059,11.432542,10.754494,10.078259,9.400211,8.963287,8.52455,8.087626,7.650702,7.211965,7.1068134,7.003474,6.8983226,6.793171,6.688019,7.3316207,7.9770355,8.62245,9.267865,9.91328,9.510801,9.108324,8.705847,8.303369,7.900891,7.1974616,6.495845,5.7924156,5.090799,4.3873696,4.597673,4.8079767,5.0182805,5.2267714,5.4370747,5.411693,5.388125,5.3627434,5.337362,5.3119802,5.328297,5.3428006,5.3573046,5.371808,5.388125,5.4515786,5.516845,5.582112,5.6473784,5.712645,6.049856,6.3870673,6.7242785,7.063302,7.400513,7.217404,7.0342946,6.8529987,6.6698895,6.48678,6.4650245,6.4432693,6.4197006,6.397945,6.3743763,5.7978544,5.219519,4.6429973,4.064662,3.48814,4.505212,5.522284,6.539356,7.558241,8.575313,7.783048,6.9907837,6.1967063,5.4044414,4.612177,3.8398547,3.0675328,2.2952106,1.5228885,0.7505665,0.7777609,0.80495536,0.8321498,0.85934424,0.8883517,1.310772,1.7331922,2.1556125,2.5780327,3.000453,2.665055,2.3296568,1.9942589,1.6606737,1.3252757,1.1367276,0.9499924,0.76325727,0.5747091,0.387974,0.36984438,0.35171473,0.33539808,0.31726846,0.2991388,0.3480888,0.39522585,0.44236287,0.4894999,0.53663695,0.6508536,0.76325727,0.87566096,0.9880646,1.1004683,1.3542831,1.6099107,1.8655385,2.1193533,2.374981,2.6777458,2.9805105,3.2832751,3.584227,3.8869917,5.5349746,7.1829576,8.829127,10.477111,12.125093,11.019187,9.915092,8.809185,7.705091,6.599184,5.977338,5.3554916,4.7318325,4.1099863,3.48814,3.489953,3.491766,3.4953918,3.4972048,3.5008307,4.2949085,5.090799,5.8848767,6.680767,7.474845,6.967215,6.4595857,5.9519563,5.4443264,4.936697,4.7771564,4.6176157,4.458075,4.2967215,4.137181,4.0501585,3.9631362,3.874301,3.787279,3.7002566,2.960568,2.220879,1.4793775,0.73968875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.13053331,0.25925365,0.38978696,0.52032024,0.6508536,0.97537386,1.2998942,1.6244144,1.9507477,2.275268,2.2408218,2.2045624,2.1701162,2.13567,2.0994108,2.126605,2.1556125,2.182807,2.2100015,2.2371957,2.8354735,3.4319382,4.0302157,4.6266804,5.224958,4.6774435,4.1299286,3.5824142,3.0348995,2.4873846,2.7847104,3.0820365,3.3793623,3.6785011,3.975827,3.9848917,3.9957695,4.004834,4.0157123,4.024777,4.227829,4.4308805,4.632119,4.835171,5.038223,5.658256,6.2782893,6.8983226,7.518356,8.136576,7.558241,6.978093,6.397945,5.8177967,5.237649,4.8841214,4.5324063,4.1806917,3.827164,3.4754493,3.5606585,3.6458678,3.729264,3.8144734,3.8996825,6.198519,8.495543,10.792566,13.08959,15.388427,15.174497,14.96238,14.750263,14.538147,14.324218,13.305332,12.284635,11.26575,10.245051,9.224354,9.264238,9.304124,9.345822,9.385707,9.425592,8.762048,8.100317,7.4367723,6.775041,6.11331,7.02523,7.93715,8.8508835,9.762803,10.674724,10.705544,10.734551,10.765372,10.794379,10.825199,9.824444,8.825501,7.8247466,6.825804,5.825049,4.8279195,3.83079,2.8318477,1.8347181,0.8375887,0.72337204,0.6073425,0.49312583,0.3770962,0.26287958,0.24293698,0.2229944,0.2030518,0.18310922,0.16316663,0.19761293,0.23205921,0.26831847,0.30276474,0.33721104,0.3480888,0.35715362,0.3680314,0.3770962,0.387974,0.37165734,0.35715362,0.34264994,0.32814622,0.31182957,0.4224203,0.533011,0.6417888,0.7523795,0.8629702,1.1856775,1.5083848,1.8292793,2.1519866,2.474694,2.762955,3.049403,3.3376641,3.6241121,3.9123733,4.327542,4.74271,5.1578784,5.573047,5.9882154,6.4251394,6.8620634,7.3008003,7.7377243,8.174648,8.283426,8.39039,8.497355,8.604321,8.713099,9.171778,9.63227,10.092763,10.553255,11.011934,11.202296,11.392657,11.583018,11.773379,11.961927,13.035201,14.108475,15.179935,16.25321,17.32467,17.288412,17.25034,17.212267,17.176008,17.137936,15.125546,13.113158,11.10077,9.088382,7.075993,6.963589,6.849373,6.736969,6.624565,6.5121617,7.478471,8.442966,9.407463,10.371959,11.338268,11.934732,12.5330105,13.129475,13.727753,14.324218,13.729566,13.134913,12.540262,11.94561,11.350959,11.735307,12.119655,12.5058155,12.890164,13.274512,14.851789,16.429068,18.008158,19.585434,21.162712,20.229036,19.297174,18.36531,17.433449,16.499773,16.57773,16.655687,16.731833,16.80979,16.887747,16.450823,16.012085,15.575162,15.138238,14.699501,14.010575,13.319836,12.629097,11.940171,11.249433,10.701918,10.154404,9.606889,9.059374,8.511859,8.629702,8.747544,8.865387,8.98323,9.099259,9.309563,9.519867,9.73017,9.940474,10.148965,9.023115,7.895452,6.7677894,5.6401267,4.512464,4.160749,3.8072214,3.4555066,3.101979,2.7502642,2.4003625,2.0504606,1.7005589,1.3506571,1.0007553,0.8103943,0.6200332,0.42967212,0.23931105,0.05076295,0.11059072,0.17041849,0.23024625,0.29007402,0.34990177,0.7505665,1.1494182,1.550083,1.9507477,2.3495996,2.0504606,1.7495089,1.4503701,1.1494182,0.85027945,0.88291276,0.9155461,0.9481794,0.9808127,1.0116332,0.85934424,0.7070554,0.55476654,0.40247768,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.02175555,0.01994259,0.018129626,0.014503701,0.012690738,0.01994259,0.027194439,0.034446288,0.04169814,0.05076295,0.07977036,0.11059072,0.13959812,0.17041849,0.19942589,0.22662032,0.25562772,0.28282216,0.3100166,0.33721104,0.37165734,0.40791658,0.44236287,0.47680917,0.51306844,0.88472575,1.258196,1.6298534,2.0033236,2.374981,2.3006494,2.2245052,2.1501737,2.0758421,1.9996977,4.4671397,6.9345818,9.402024,11.869466,14.336908,16.788034,18.3218,19.85738,21.392958,22.926725,24.462305,25.252756,26.041395,26.831846,27.622297,28.41275,26.857227,25.301706,23.747997,22.192474,20.636953,19.407764,18.176764,16.947575,15.716573,14.487384,13.437678,12.387974,11.338268,10.28675,9.237044,8.814624,8.392203,7.9697833,7.5473633,7.124943,7.51473,7.9045167,8.294304,8.685904,9.07569,8.807372,8.540867,8.272549,8.00423,7.7377243,7.1068134,6.4777155,5.846804,5.217706,4.5867953,4.744523,4.902251,5.0599785,5.217706,5.375434,5.3119802,5.2503395,5.186886,5.125245,5.0617914,5.0545397,5.047288,5.040036,5.032784,5.0255322,5.029158,5.034597,5.040036,5.045475,5.050914,5.2503395,5.4497657,5.6491914,5.8504305,6.049856,5.9718986,5.8957543,5.8177967,5.7398396,5.661882,5.7924156,5.922949,6.051669,6.1822023,6.3127356,5.732588,5.1524396,4.572292,3.9921436,3.4119956,4.1480584,4.882308,5.618371,6.352621,7.0868707,6.526665,5.9682727,5.408067,4.847862,4.2876563,3.7056956,3.1219215,2.5399606,1.9579996,1.3742256,1.4304274,1.4848163,1.5392052,1.5954071,1.649796,1.9579996,2.2643902,2.572594,2.8807976,3.1871881,2.9170568,2.6469254,2.3767939,2.1066625,1.8383441,1.6117238,1.3869164,1.162109,0.93730164,0.7124943,0.69073874,0.6671702,0.64541465,0.62184614,0.6000906,0.69436467,0.7904517,0.88472575,0.9808127,1.0750868,1.2745126,1.4757515,1.6751775,1.8746033,2.0758421,2.222692,2.3695421,2.518205,2.665055,2.811905,3.1291735,3.4482548,3.7655232,4.082792,4.40006,5.569421,6.740595,7.909956,9.079316,10.25049,9.465478,8.680465,7.895452,7.1104393,6.3254266,5.7797246,5.235836,4.690134,4.1444325,3.6005437,3.4047437,3.2107568,3.0149567,2.819157,2.6251698,3.2270734,3.83079,4.4326935,5.034597,5.638314,5.3101673,4.9820213,4.655688,4.327542,3.9993954,3.83079,3.6603715,3.489953,3.3195345,3.150929,3.0747845,3.000453,2.9243085,2.8499773,2.7756457,2.220879,1.6642996,1.1095331,0.55476654,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.17223145,0.3444629,0.5166943,0.69073874,0.8629702,1.2255627,1.5881553,1.9507477,2.3133402,2.6741197,2.467442,2.2607644,2.0522738,1.845596,1.6371052,1.6552348,1.6733645,1.6896812,1.7078108,1.7241274,2.3079014,2.8898623,3.4718235,4.0555973,4.6375585,4.2042603,3.7727752,3.339477,2.907992,2.474694,3.2832751,4.0900435,4.896812,5.7053933,6.5121617,6.432391,6.352621,6.2728505,6.19308,6.11331,6.0426044,5.9718986,5.903006,5.8323007,5.7615952,6.0407915,6.3181744,6.5955577,6.872941,7.1503243,6.5647373,5.979151,5.3953767,4.8097897,4.2242026,4.082792,3.9395678,3.7981565,3.6549325,3.5117085,4.233268,4.953014,5.67276,6.392506,7.112252,9.131892,11.151533,13.172986,15.192626,17.212267,16.525154,15.838041,15.149116,14.462003,13.77489,12.647227,11.519565,10.391902,9.264238,8.138389,8.192778,8.247167,8.303369,8.357758,8.412147,7.8628187,7.311678,6.7623506,6.2130227,5.661882,6.4632115,7.262728,8.062244,8.861761,9.663091,9.610515,9.557939,9.5053625,9.452786,9.400211,8.537241,7.6742706,6.813113,5.9501433,5.087173,4.2804046,3.4718235,2.665055,1.8582866,1.0497054,0.90829426,0.7650702,0.62184614,0.48043507,0.33721104,0.29732585,0.2574407,0.21755551,0.17767033,0.13778515,0.17041849,0.2030518,0.23568514,0.26831847,0.2991388,0.30820364,0.3154555,0.32270733,0.32995918,0.33721104,0.35715362,0.3770962,0.39703882,0.4169814,0.43692398,0.5946517,0.7523795,0.9101072,1.067835,1.2255627,1.4703126,1.7150626,1.9598125,2.2045624,2.4493124,2.6378605,2.8245957,3.0131438,3.199879,3.386614,4.0302157,4.6720047,5.315606,5.957395,6.599184,7.175706,7.750415,8.325124,8.899834,9.474543,9.414715,9.354887,9.295059,9.235231,9.175404,9.956791,10.73999,11.5231905,12.304577,13.087777,13.354282,13.622601,13.889107,14.157425,14.425743,15.382988,16.34023,17.297476,18.25472,19.211964,19.424082,19.63801,19.850128,20.062244,20.27436,18.43783,16.599485,14.762955,12.92461,11.088079,10.312131,9.537996,8.762048,7.987913,7.211965,7.7794223,8.34688,8.914337,9.481794,10.049252,10.707357,11.365462,12.021755,12.67986,13.337966,13.134913,12.931862,12.730623,12.527572,12.32452,12.607342,12.890164,13.172986,13.455809,13.736817,15.067532,16.398247,17.727148,19.057863,20.386765,20.10938,19.831997,19.554615,19.277231,18.999847,18.941833,18.885632,18.827616,18.769602,18.711586,18.136877,17.562168,16.98746,16.41275,15.838041,14.895301,13.95256,13.009819,12.067079,11.124338,10.480737,9.835322,9.189907,8.544493,7.900891,7.75948,7.6198816,7.4802837,7.3406854,7.1992745,7.308052,7.415017,7.5219817,7.6307597,7.7377243,6.869315,6.002719,5.1343102,4.267714,3.3993049,3.1327994,2.864481,2.5979755,2.3296568,2.0631514,1.8002719,1.5373923,1.2745126,1.0116332,0.7505665,0.6073425,0.46411842,0.32270733,0.1794833,0.038072214,0.08339628,0.12690738,0.17223145,0.21755551,0.26287958,0.5620184,0.8629702,1.162109,1.4630609,1.7621996,1.5373923,1.3125849,1.0877775,0.8629702,0.63816285,0.6653573,0.69255173,0.7197462,0.7469406,0.774135,0.65810543,0.5402629,0.4224203,0.3045777,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.045324065,0.03988518,0.034446288,0.030820364,0.025381476,0.027194439,0.030820364,0.032633327,0.034446288,0.038072214,0.072518505,0.10696479,0.14322405,0.17767033,0.21211663,0.27919623,0.3480888,0.41516843,0.48224804,0.5493277,0.55839247,0.5656443,0.5728962,0.58014804,0.5873999,0.89560354,1.2019942,1.5101979,1.8165885,2.124792,2.0758421,2.0250793,1.9743162,1.9253663,1.8746033,4.0972953,6.319988,8.54268,10.765372,12.988064,15.149116,17.915697,20.680464,23.445232,26.210001,28.974768,30.760536,32.54449,34.33026,36.116028,37.899982,36.018127,34.13446,32.252605,30.370749,28.487082,26.704939,24.922796,23.140654,21.358513,19.574556,17.912071,16.249584,14.587097,12.92461,11.262123,10.522435,9.782746,9.043057,8.303369,7.5618668,7.6978393,7.8319983,7.9679704,8.10213,8.238102,8.105756,7.9715962,7.83925,7.706904,7.574558,7.017978,6.4595857,5.903006,5.3446136,4.788034,4.893186,4.9983377,5.101677,5.2068286,5.3119802,5.2122674,5.1125546,5.0128417,4.9131284,4.8116026,4.782595,4.751775,4.7227674,4.691947,4.6629395,4.606738,4.552349,4.49796,4.441758,4.3873696,4.4508233,4.512464,4.574105,4.6375585,4.699199,4.7282066,4.7554007,4.782595,4.8097897,4.836984,5.1198063,5.4026284,5.6854506,5.9682727,6.249282,5.667321,5.08536,4.501586,3.919625,3.3376641,3.7890918,4.2423325,4.695573,5.147001,5.600241,5.272095,4.945762,4.6176157,4.2894692,3.9631362,3.5697234,3.1781235,2.7847104,2.3931105,1.9996977,2.0830941,2.1646774,2.2480736,2.3296568,2.4130533,2.6052272,2.7974012,2.9895754,3.1817493,3.3757362,3.1708715,2.9641938,2.759329,2.5544643,2.3495996,2.08672,1.8256533,1.5627737,1.2998942,1.0370146,1.0098201,0.9826257,0.9554313,0.92823684,0.89922947,1.0424535,1.1856775,1.3270886,1.4703126,1.6117238,1.8999848,2.1882458,2.474694,2.762955,3.049403,3.0892882,3.1291735,3.1708715,3.2107568,3.2506418,3.5824142,3.9141862,4.2477713,4.5795436,4.9131284,5.6056805,6.298232,6.9907837,7.6833353,8.374074,7.909956,7.4458375,6.979906,6.5157876,6.049856,5.582112,5.1143675,4.646623,4.1806917,3.7129474,3.3195345,2.9279346,2.5345216,2.1429217,1.7495089,2.1592383,2.570781,2.9805105,3.39024,3.7999697,3.6531196,3.5044568,3.3576066,3.2107568,3.0620937,2.8826106,2.7031271,2.521831,2.3423476,2.1628644,2.0994108,2.03777,1.9743162,1.9126755,1.8492218,1.4793775,1.1095331,0.73968875,0.36984438,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.21574254,0.42967212,0.64541465,0.85934424,1.0750868,1.4757515,1.8746033,2.275268,2.6741197,3.0747845,2.6958754,2.3151531,1.9344311,1.5555218,1.1747998,1.1820517,1.1893034,1.1983683,1.2056202,1.2128719,1.7803292,2.3477864,2.9152439,3.482701,4.0501585,3.73289,3.4156215,3.0983531,2.7792716,2.4620032,3.780027,5.0980506,6.414262,7.7322855,9.050309,8.87989,8.709473,8.540867,8.370448,8.200029,7.85738,7.51473,7.17208,6.82943,6.48678,6.4233265,6.35806,6.2927933,6.2275267,6.16226,5.573047,4.9820213,4.3928084,3.8017826,3.2125697,3.2796493,3.346729,3.4156215,3.482701,3.5497808,4.9058766,6.26016,7.614443,8.970539,10.324821,12.067079,13.809336,15.553406,17.295664,19.03792,17.87581,16.71189,15.54978,14.387671,13.225562,11.989121,10.754494,9.519867,8.285239,7.0506115,7.119504,7.1902094,7.2591023,7.3298078,7.400513,6.9617763,6.5248523,6.0879283,5.6491914,5.2122674,5.89938,6.588306,7.2754188,7.9625316,8.649645,8.515485,8.379513,8.245354,8.109382,7.9752226,7.250037,6.5248523,5.7996674,5.0744824,4.349297,3.73289,3.1146698,2.4982624,1.8800422,1.261822,1.0932164,0.922798,0.7523795,0.581961,0.41335547,0.35171473,0.291887,0.23205921,0.17223145,0.11240368,0.14322405,0.17223145,0.2030518,0.23205921,0.26287958,0.26831847,0.27194437,0.27738327,0.28282216,0.28826106,0.34264994,0.39703882,0.45324063,0.5076295,0.5620184,0.7668832,0.97174793,1.1766127,1.3832904,1.5881553,1.7549478,1.9217403,2.0903459,2.2571385,2.4257438,2.5127661,2.5997884,2.6868105,2.7756457,2.8626678,3.73289,4.603112,5.473334,6.341743,7.211965,7.9244595,8.636953,9.349448,10.061942,10.774437,10.547816,10.319383,10.092763,9.864329,9.637709,10.741803,11.847711,12.951805,14.057712,15.161806,15.508082,15.852545,16.197008,16.543283,16.887747,17.730774,18.57199,19.415016,20.258043,21.099258,21.563377,22.025682,22.487988,22.950293,23.4126,21.750113,20.087626,18.425138,16.762651,15.100165,13.662486,12.224807,10.7871275,9.349448,7.911769,8.082188,8.252605,8.423024,8.59163,8.762048,9.479981,10.197914,10.915848,11.631968,12.349901,12.540262,12.730623,12.919171,13.109532,13.299893,13.479377,13.660673,13.840157,14.01964,14.199123,15.283275,16.365614,17.447952,18.53029,19.612629,19.989725,20.366821,20.745731,21.122828,21.499924,21.307749,21.115576,20.9234,20.729414,20.537241,19.824745,19.112251,18.399757,17.687263,16.97477,15.780026,14.585284,13.390542,12.195799,10.999244,10.257742,9.514427,8.772926,8.029612,7.28811,6.889258,6.492219,6.09518,5.6981416,5.2992897,5.3047285,5.3101673,5.315606,5.319232,5.3246713,4.7173285,4.1099863,3.5026438,2.8953013,2.2879589,2.1048496,1.9217403,1.7404441,1.5573349,1.3742256,1.2001812,1.0243238,0.85027945,0.6744221,0.50037766,0.40429065,0.3100166,0.21574254,0.11965553,0.025381476,0.054388877,0.08520924,0.11421664,0.14503701,0.17585737,0.37528324,0.5747091,0.774135,0.97537386,1.1747998,1.0243238,0.87566096,0.72518504,0.5747091,0.42423326,0.44780177,0.46955732,0.49312583,0.5148814,0.53663695,0.4550536,0.37165734,0.29007402,0.20667773,0.12509441,0.099712946,0.07433146,0.05076295,0.025381476,0.0,0.014503701,0.030820364,0.045324065,0.059827764,0.07433146,0.06707962,0.059827764,0.052575916,0.045324065,0.038072214,0.034446288,0.032633327,0.030820364,0.027194439,0.025381476,0.065266654,0.10515183,0.14503701,0.18492219,0.22480737,0.33177215,0.4405499,0.5475147,0.6544795,0.76325727,0.7433147,0.72337204,0.7016165,0.68167394,0.66173136,0.90466833,1.1476053,1.3905423,1.6316663,1.8746033,1.8492218,1.8256533,1.8002719,1.7748904,1.7495089,3.727451,5.7053933,7.6833353,9.659465,11.637406,13.512011,17.50778,21.501736,25.497505,29.493275,33.487232,36.26832,39.04759,41.82686,44.607944,47.387215,45.177216,42.967213,40.757214,38.54721,36.337208,34.002113,31.667017,29.331923,26.996826,24.66173,22.388275,20.113007,17.837738,15.56247,13.287203,12.230246,11.173288,10.114518,9.057561,8.000604,7.8791356,7.75948,7.6398244,7.520169,7.400513,7.402326,7.404139,7.407765,7.409578,7.413204,6.92733,6.4432693,5.957395,5.473334,4.98746,5.040036,5.092612,5.145188,5.197764,5.2503395,5.1125546,4.974769,4.836984,4.699199,4.5632267,4.510651,4.458075,4.405499,4.3529234,4.3003473,4.1843176,4.070101,3.9558845,3.8398547,3.7256382,3.6494937,3.5751622,3.5008307,3.4246864,3.350355,3.482701,3.6150475,3.7473936,3.87974,4.0120864,4.4471974,4.882308,5.317419,5.75253,6.187641,5.6020546,5.0182805,4.4326935,3.8471067,3.2633326,3.4319382,3.6023567,3.7727752,3.9431937,4.1117992,4.017525,3.923251,3.827164,3.73289,3.636803,3.435564,3.2325122,3.0294604,2.8282216,2.6251698,2.7357605,2.8445382,2.955129,3.0657198,3.1744974,3.2524548,3.3304121,3.4083695,3.484514,3.5624714,3.4228733,3.2832751,3.141864,3.002266,2.8626678,2.561716,2.2625773,1.9616255,1.6624867,1.3633479,1.3307146,1.2980812,1.2654479,1.2328146,1.2001812,1.3905423,1.5809034,1.7694515,1.9598125,2.1501737,2.525457,2.9007401,3.2742105,3.6494937,4.024777,3.9576974,3.8906176,3.8217251,3.7546456,3.6875658,4.0356545,4.3819304,4.7300196,5.0781083,5.424384,5.6401267,5.8558693,6.069799,6.285541,6.4994707,6.354434,6.209397,6.0643597,5.919323,5.774286,5.384499,4.994712,4.604925,4.215138,3.825351,3.2343252,2.6451125,2.0540867,1.4648738,0.87566096,1.0932164,1.310772,1.5283275,1.745883,1.9616255,1.9942589,2.0268922,2.0595255,2.0921588,2.124792,1.9344311,1.745883,1.5555218,1.3651608,1.1747998,1.1258497,1.0750868,1.0243238,0.97537386,0.9246109,0.73968875,0.55476654,0.36984438,0.18492219,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.2574407,0.5148814,0.77232206,1.0297627,1.2872034,1.7241274,2.1628644,2.5997884,3.0367124,3.4754493,2.9224956,2.3695421,1.8165885,1.2654479,0.7124943,0.7106813,0.7070554,0.70524246,0.7016165,0.69980353,1.2527572,1.8057107,2.3568513,2.909805,3.4627585,3.2597067,3.056655,2.855416,2.6523643,2.4493124,4.2767787,6.104245,7.931711,9.759177,11.586644,11.327391,11.068136,10.80707,10.547816,10.28675,9.672155,9.057561,8.442966,7.8283725,7.211965,6.8058615,6.397945,5.9900284,5.582112,5.1741953,4.5795436,3.9848917,3.39024,2.7955883,2.1991236,2.47832,2.7557032,3.0330863,3.3104696,3.587853,5.578486,7.567306,9.557939,11.546759,13.537392,15.002265,16.467138,17.932013,19.396887,20.861761,19.224655,17.58755,15.950445,14.313339,12.674421,11.332829,9.989424,8.647832,7.304426,5.962834,6.0480433,6.1332526,6.2166486,6.301858,6.3870673,6.0625467,5.7380266,5.411693,5.087173,4.762653,5.337362,5.9120708,6.48678,7.063302,7.6380115,7.420456,7.2029004,6.985345,6.7677894,6.550234,5.962834,5.375434,4.788034,4.2006345,3.6132345,3.1853752,2.7575161,2.3296568,1.9017978,1.4757515,1.2781386,1.0805258,0.88291276,0.6852999,0.48768693,0.40791658,0.32814622,0.24837588,0.16679256,0.0870222,0.11421664,0.14322405,0.17041849,0.19761293,0.22480737,0.22662032,0.23024625,0.23205921,0.23568514,0.2374981,0.32814622,0.4169814,0.5076295,0.5982776,0.6871128,0.93911463,1.1929294,1.4449311,1.696933,1.9507477,2.039583,2.1302311,2.220879,2.3097143,2.4003625,2.3876717,2.374981,2.3622901,2.3495996,2.3369088,3.435564,4.5324063,5.6292486,6.7279043,7.8247466,8.675026,9.525306,10.375585,11.225864,12.07433,11.679105,11.285692,10.890467,10.49524,10.100015,11.526816,12.955431,14.382232,15.810846,17.237648,17.660069,18.082489,18.50491,18.92733,19.34975,20.076748,20.80556,21.532557,22.259554,22.988365,23.70086,24.413355,25.125849,25.838343,26.550837,25.062395,23.575766,22.087322,20.600695,19.112251,17.01284,14.91343,12.812206,10.712796,8.613385,8.384952,8.158332,7.9298983,7.703278,7.474845,8.252605,9.030367,9.808127,10.585889,11.361836,11.94561,12.527572,13.109532,13.693306,14.275268,14.353225,14.429369,14.507326,14.585284,14.663241,15.497204,16.33298,17.166943,18.002718,18.836681,19.87007,20.901646,21.935034,22.968424,23.999998,23.671852,23.34552,23.017372,22.689226,22.362894,21.512613,20.662334,19.812056,18.961775,18.11331,16.664753,15.218008,13.769451,12.322706,10.874149,10.034748,9.195346,8.354132,7.51473,6.6753283,6.0208488,5.3645563,4.710077,4.0555973,3.3993049,3.303218,3.2053177,3.1074178,3.009518,2.911618,2.565342,2.2172532,1.8691645,1.5228885,1.1747998,1.0768998,0.9808127,0.88291276,0.7850128,0.6871128,0.6000906,0.51306844,0.42423326,0.33721104,0.25018883,0.2030518,0.15410182,0.10696479,0.059827764,0.012690738,0.027194439,0.04169814,0.058014803,0.072518505,0.0870222,0.18673515,0.28826106,0.387974,0.48768693,0.5873999,0.51306844,0.43692398,0.36259252,0.28826106,0.21211663,0.23024625,0.24837588,0.26469254,0.28282216,0.2991388,0.2520018,0.20486477,0.15772775,0.11059072,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.01994259,0.03988518,0.059827764,0.07977036,0.099712946,0.09064813,0.07977036,0.07070554,0.059827764,0.05076295,0.04169814,0.034446288,0.027194439,0.01994259,0.012690738,0.058014803,0.10333887,0.14684997,0.19217403,0.2374981,0.38434806,0.533011,0.67986095,0.82671094,0.97537386,0.92823684,0.8792868,0.8321498,0.7850128,0.73787576,0.9155461,1.0932164,1.2708868,1.4467441,1.6244144,1.6244144,1.6244144,1.6244144,1.6244144,1.6244144,3.3576066,5.090799,6.8221784,8.55537,10.28675,11.874905,17.099863,22.324821,27.54978,32.77474,37.999695,41.774284,45.550686,49.32527,53.09986,56.87445,54.338116,51.79997,49.261818,46.725483,44.187336,41.299286,38.41305,35.525,32.63695,29.750715,26.862667,23.974617,21.086567,18.20033,15.312282,13.938056,12.562017,11.187792,9.811753,8.437528,8.062244,7.686961,7.311678,6.9382076,6.5629244,6.70071,6.836682,6.9744673,7.112252,7.250037,6.836682,6.4251394,6.011784,5.600241,5.186886,5.186886,5.186886,5.186886,5.186886,5.186886,5.0128417,4.836984,4.6629395,4.4870825,4.313038,4.2368937,4.162562,4.0882306,4.0120864,3.9377546,3.7618973,3.587853,3.4119956,3.2379513,3.0620937,2.8499773,2.6378605,2.4257438,2.2118144,1.9996977,2.2371957,2.474694,2.712192,2.94969,3.1871881,3.774588,4.361988,4.949388,5.5367875,6.1241875,5.5367875,4.949388,4.361988,3.774588,3.1871881,3.0747845,2.962381,2.8499773,2.7375734,2.6251698,2.762955,2.9007401,3.0367124,3.1744974,3.3122826,3.299592,3.2869012,3.2742105,3.2633326,3.2506418,3.386614,3.5243993,3.6621845,3.7999697,3.9377546,3.8996825,3.8616104,3.825351,3.787279,3.7492065,3.6748753,3.6005437,3.5243993,3.4500678,3.3757362,3.0367124,2.6995013,2.3622901,2.0250793,1.6878681,1.649796,1.6117238,1.5754645,1.5373923,1.49932,1.7368182,1.9743162,2.2118144,2.4493124,2.6868105,3.149116,3.6132345,4.07554,4.537845,5.0001507,4.8242936,4.650249,4.4743915,4.3003473,4.12449,4.4870825,4.8496747,5.2122674,5.57486,5.9374523,5.674573,5.411693,5.1506267,4.8877473,4.6248674,4.800725,4.974769,5.1506267,5.3246713,5.5005283,5.186886,4.8750563,4.5632267,4.249584,3.9377546,3.149116,2.3622901,1.5754645,0.7868258,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.33721104,0.5493277,0.76325727,0.97537386,1.1874905,0.9880646,0.7868258,0.5873999,0.387974,0.18673515,0.15047589,0.11240368,0.07433146,0.038072214,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.2991388,0.6000906,0.89922947,1.2001812,1.49932,1.9743162,2.4493124,2.9243085,3.3993049,3.874301,3.149116,2.4257438,1.7005589,0.97537386,0.25018883,0.2374981,0.22480737,0.21211663,0.19942589,0.18673515,0.72518504,1.261822,1.8002719,2.3369088,2.8753586,2.7883365,2.6995013,2.612479,2.525457,2.4366217,4.7753434,7.112252,9.4509735,11.787883,14.124791,13.77489,13.424988,13.075087,12.725184,12.375282,11.486931,10.600392,9.712041,8.825501,7.93715,7.1865835,6.43783,5.6872635,4.936697,4.1879435,3.587853,2.9877625,2.3876717,1.7875811,1.1874905,1.6751775,2.1628644,2.6505513,3.1382382,3.6241121,6.249282,8.874452,11.499621,14.124791,16.749962,17.937452,19.124943,20.312433,21.499924,22.687414,20.575312,18.463211,16.349297,14.237195,12.125093,10.674724,9.224354,7.7757964,6.3254266,4.8750563,4.974769,5.0744824,5.1741953,5.275721,5.375434,5.163317,4.949388,4.7372713,4.5251546,4.313038,4.7753434,5.237649,5.6999545,6.16226,6.624565,6.3254266,6.0244746,5.7253356,5.424384,5.125245,4.6756306,4.2242026,3.774588,3.3249733,2.8753586,2.6378605,2.4003625,2.1628644,1.9253663,1.6878681,1.4630609,1.2382535,1.0116332,0.7868258,0.5620184,0.46230546,0.36259252,0.26287958,0.16316663,0.06164073,0.0870222,0.11240368,0.13778515,0.16316663,0.18673515,0.18673515,0.18673515,0.18673515,0.18673515,0.18673515,0.31182957,0.43692398,0.5620184,0.6871128,0.8122072,1.1131591,1.4122978,1.7132497,2.0123885,2.3133402,2.324218,2.3369088,2.3495996,2.3622901,2.374981,2.2625773,2.1501737,2.03777,1.9253663,1.8129625,3.1382382,4.461701,5.7869763,7.112252,8.437528,9.425592,10.411844,11.399909,12.387974,13.374225,12.812206,12.250188,11.6881695,11.124338,10.56232,12.311829,14.06315,15.812659,17.562168,19.311678,19.812056,20.312433,20.81281,21.313189,21.811752,22.424534,23.037315,23.650097,24.262878,24.87566,25.838343,26.799213,27.761896,28.724579,29.687262,28.374678,27.062092,25.749508,24.436922,23.124338,20.363195,17.60024,14.837286,12.07433,9.313189,8.6877165,8.062244,7.4367723,6.813113,6.187641,7.02523,7.8628187,8.700407,9.537996,10.375585,11.350959,12.32452,13.299893,14.275268,15.250641,15.22526,15.199879,15.174497,15.149116,15.125546,15.712947,16.300346,16.887747,17.475147,18.062546,19.750414,21.438282,23.124338,24.812206,26.500074,26.03777,25.575462,25.113157,24.650852,24.186733,23.200481,22.212418,21.224354,20.238102,19.250036,17.549479,15.850732,14.150173,12.449615,10.750868,9.811753,8.874452,7.93715,6.9998484,6.0625467,5.1506267,4.2368937,3.3249733,2.4130533,1.49932,1.2998942,1.1004683,0.89922947,0.69980353,0.50037766,0.41335547,0.3245203,0.2374981,0.15047589,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.0,0.0,0.0,0.0,0.0,0.025381476,0.05076295,0.07433146,0.099712946,0.12509441,0.11240368,0.099712946,0.0870222,0.07433146,0.06164073,0.05076295,0.038072214,0.025381476,0.012690738,0.0,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,0.43692398,0.62547207,0.8122072,1.0007553,1.1874905,1.1131591,1.0370146,0.96268314,0.8883517,0.8122072,0.9246109,1.0370146,1.1494182,1.261822,1.3742256,1.3996071,1.4249886,1.4503701,1.4757515,1.49932,2.9877625,4.4743915,5.962834,7.4494634,8.937905,10.312131,14.529082,18.747847,22.964798,27.181747,31.398699,34.471672,37.544643,40.617615,43.688774,46.761745,44.736664,42.711586,40.68651,38.661427,36.63635,35.18054,33.722916,32.265297,30.807673,29.350052,27.47726,25.604471,23.733494,21.860703,19.987913,18.372562,16.757214,15.141864,13.528327,11.912977,11.650098,11.3872175,11.124338,10.863272,10.600392,11.722616,12.84484,13.967064,15.091101,16.213324,16.200634,16.187943,16.175253,16.162561,16.14987,15.54978,14.951503,14.351412,13.751321,13.151231,13.410484,13.669738,13.930804,14.190058,14.451125,14.757515,15.065719,15.373922,15.680313,15.988517,14.568967,13.147605,11.728055,10.308505,8.887142,7.763106,6.637256,5.5132194,4.3873696,3.2633326,3.2306993,3.198066,3.1654327,3.1327994,3.100166,3.5352771,3.9703882,4.405499,4.84061,5.275721,4.751775,4.229642,3.7075086,3.1853752,2.663242,2.5870976,2.5127661,2.4366217,2.3622901,2.2879589,2.42937,2.572594,2.715818,2.857229,3.000453,3.1327994,3.2651455,3.397492,3.529838,3.6621845,4.0392804,4.41819,4.795286,5.1723824,5.5494785,5.522284,5.4950895,5.467895,5.4407005,5.4135065,5.0545397,4.6973863,4.3402324,3.9830787,3.6241121,3.2705846,2.9152439,2.5599031,2.2045624,1.8492218,1.7694515,1.6896812,1.6099107,1.5301404,1.4503701,1.6425442,1.8347181,2.0268922,2.220879,2.4130533,2.8626678,3.3122826,3.7618973,4.213325,4.6629395,4.505212,4.347484,4.1897564,4.0320287,3.874301,4.1045475,4.3347936,4.5650396,4.795286,5.0255322,4.7699046,4.514277,4.2604623,4.004834,3.7492065,3.9522583,4.15531,4.358362,4.559601,4.762653,4.458075,4.1516843,3.8471067,3.5425289,3.2379513,2.5925364,1.9471219,1.3017071,0.65810543,0.012690738,0.04169814,0.072518505,0.10333887,0.13234627,0.16316663,0.3208944,0.47680917,0.6345369,0.79226464,0.9499924,0.7904517,0.629098,0.46955732,0.3100166,0.15047589,0.11965553,0.09064813,0.059827764,0.030820364,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.058014803,0.065266654,0.072518505,0.07977036,0.0870222,0.11784257,0.14684997,0.17767033,0.20667773,0.2374981,0.2574407,0.27738327,0.29732585,0.31726846,0.33721104,0.70524246,1.0732739,1.4394923,1.8075237,2.175555,2.4384346,2.6995013,2.962381,3.2252605,3.48814,2.8372865,2.1882458,1.5373923,0.8883517,0.2374981,0.25018883,0.26287958,0.2755703,0.28826106,0.2991388,0.80676836,1.3143979,1.8220274,2.3296568,2.8372865,2.6995013,2.561716,2.4257438,2.2879589,2.1501737,4.4834566,6.814926,9.14821,11.479679,13.812962,13.325275,12.837588,12.349901,11.862214,11.374527,10.455356,9.53437,8.615198,7.6942134,6.775041,6.19308,5.6093063,5.027345,4.445384,3.8616104,3.3775494,2.8916752,2.4076142,1.9217403,1.4376793,2.228131,3.0167696,3.8072214,4.597673,5.388125,7.993352,10.596766,13.201994,15.80722,18.412449,18.767788,19.123129,19.476658,19.831997,20.187338,18.307297,16.427254,14.547212,12.66717,10.7871275,9.759177,8.733041,7.705091,6.677141,5.6491914,5.6981416,5.7452784,5.7924156,5.8395524,5.8866897,5.540414,5.1923246,4.844236,4.49796,4.1498713,4.554162,4.9602656,5.3645563,5.77066,6.1749506,5.979151,5.7851634,5.5893636,5.3953767,5.199577,4.782595,4.365614,3.9468195,3.529838,3.1128569,2.7828975,2.4529383,2.1229792,1.79302,1.4630609,1.2690738,1.0768998,0.88472575,0.69255173,0.50037766,0.40972954,0.3208944,0.23024625,0.13959812,0.05076295,0.07977036,0.11059072,0.13959812,0.17041849,0.19942589,0.2755703,0.34990177,0.42423326,0.50037766,0.5747091,0.67986095,0.7850128,0.8901646,0.99531645,1.1004683,1.2781386,1.455809,1.6316663,1.8093367,1.987007,2.0250793,2.0631514,2.0994108,2.137483,2.175555,2.0975976,2.0196402,1.9416829,1.8655385,1.7875811,3.0421512,4.2967215,5.5531044,6.8076744,8.062244,8.930654,9.79725,10.665659,11.532255,12.400664,12.077957,11.755249,11.432542,11.109835,10.7871275,12.183108,13.577277,14.973258,16.367426,17.761595,18.102432,18.443268,18.782291,19.123129,19.462152,20.093063,20.722162,21.353073,21.982172,22.613083,23.606586,24.601902,25.59722,26.592535,27.587852,26.670492,25.753134,24.835773,23.916603,22.999243,20.736666,18.475903,16.213324,13.9507475,11.6881695,10.810696,9.933222,9.055748,8.178274,7.3008003,7.895452,8.490104,9.084756,9.679407,10.275872,11.050007,11.8241415,12.60009,13.374225,14.150173,14.249886,14.349599,14.449312,14.5508375,14.650551,15.23795,15.825351,16.41275,17.00015,17.58755,18.992596,20.397642,21.802689,23.207733,24.61278,24.07433,23.537693,22.999243,22.462606,21.924156,20.914337,19.904516,18.894695,17.884876,16.875055,15.509895,14.144734,12.779573,11.4144125,10.049252,9.023115,7.995165,6.967215,5.9392653,4.9131284,4.169814,3.4283123,2.6849976,1.9416829,1.2001812,1.0406405,0.8792868,0.7197462,0.56020546,0.40066472,0.32995918,0.25925365,0.19036107,0.11965553,0.05076295,0.03988518,0.030820364,0.01994259,0.010877775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.18673515,0.36259252,0.53663695,0.7124943,0.8883517,0.7106813,0.533011,0.35534066,0.17767033,0.0,0.058014803,0.11421664,0.17223145,0.23024625,0.28826106,0.27738327,0.26831847,0.2574407,0.24837588,0.2374981,0.20486477,0.17223145,0.13959812,0.10696479,0.07433146,0.10333887,0.13053331,0.15772775,0.18492219,0.21211663,0.21936847,0.22662032,0.23568514,0.24293698,0.25018883,0.42967212,0.6091554,0.7904517,0.969935,1.1494182,1.0805258,1.0098201,0.93911463,0.87022203,0.7995165,0.9880646,1.1747998,1.3633479,1.550083,1.7368182,1.7368182,1.7368182,1.7368182,1.7368182,1.7368182,3.0367124,4.3384194,5.638314,6.9382076,8.238102,8.749357,11.9601145,15.170871,18.379814,21.59057,24.799515,27.17087,29.540413,31.909954,34.279495,36.650852,35.137028,33.625015,32.113007,30.600996,29.087172,29.059977,29.032784,29.005589,28.978394,28.949387,28.091856,27.234324,26.376793,25.51926,24.66173,22.80707,20.952408,19.097748,17.243088,15.386614,15.23795,15.087475,14.936998,14.786523,14.63786,16.744522,18.852999,20.95966,23.068136,25.174799,25.562773,25.948933,26.336908,26.724882,27.112856,25.912674,24.712494,23.512312,22.31213,21.11195,21.808126,22.502491,23.196856,23.893034,24.587399,25.276325,25.967064,26.657803,27.346727,28.037466,25.372412,22.707355,20.042301,17.377247,14.712192,12.674421,10.636651,8.600695,6.5629244,4.5251546,4.2223897,3.919625,3.6168604,3.3140955,3.0131438,3.294153,3.576975,3.8597972,4.1426196,4.4254417,3.966762,3.5098956,3.053029,2.5943494,2.137483,2.0994108,2.0631514,2.0250793,1.987007,1.9507477,2.0975976,2.2444477,2.3931105,2.5399606,2.6868105,2.9641938,3.24339,3.5207734,3.7981565,4.07554,4.691947,5.3101673,5.9283876,6.544795,7.1630154,7.1448855,7.1267557,7.1104393,7.0923095,7.07418,6.434204,5.7942286,5.1542525,4.514277,3.874301,3.5026438,3.1291735,2.7575161,2.3858588,2.0123885,1.889107,1.7676386,1.6443571,1.5228885,1.3996071,1.54827,1.69512,1.84197,1.9906329,2.137483,2.5744069,3.0131438,3.4500678,3.8869917,4.325729,4.1843176,4.0447197,3.9051213,3.7655232,3.6241121,3.7220123,3.8199122,3.917812,4.0157123,4.1117992,3.8652363,3.6168604,3.3702974,3.1219215,2.8753586,3.105605,3.3358512,3.5642843,3.7945306,4.024777,3.727451,3.4301252,3.1327994,2.8354735,2.5381477,2.034144,1.5319533,1.0297627,0.5275721,0.025381476,0.059827764,0.09427405,0.13053331,0.16497959,0.19942589,0.30276474,0.40429065,0.5076295,0.6091554,0.7124943,0.59283876,0.47318324,0.35171473,0.23205921,0.11240368,0.09064813,0.06707962,0.045324065,0.02175555,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.052575916,0.06707962,0.08339628,0.09789998,0.11240368,0.18492219,0.2574407,0.32995918,0.40247768,0.4749962,0.5148814,0.55476654,0.5946517,0.6345369,0.6744221,1.1095331,1.5446441,1.9797552,2.4148662,2.8499773,2.9007401,2.94969,3.000453,3.049403,3.100166,2.525457,1.9507477,1.3742256,0.7995165,0.22480737,0.26287958,0.2991388,0.33721104,0.37528324,0.41335547,0.8901646,1.3669738,1.845596,2.322405,2.7992141,2.612479,2.4257438,2.2371957,2.0504606,1.8619126,4.1897564,6.5176005,8.845445,11.173288,13.499319,12.87566,12.250188,11.624716,10.999244,10.375585,9.421967,8.470161,7.518356,6.5647373,5.612932,5.197764,4.782595,4.367427,3.9522583,3.53709,3.1672456,2.7974012,2.427557,2.0577126,1.6878681,2.7792716,3.872488,4.9657044,6.057108,7.1503243,9.735609,12.31908,14.904366,17.48965,20.074934,19.598125,19.119503,18.642694,18.165886,17.687263,16.03928,14.39311,12.745127,11.097144,9.449161,8.845445,8.239915,7.6343856,7.0306687,6.4251394,6.4197006,6.414262,6.4106355,6.4051967,6.399758,5.91751,5.4352617,4.953014,4.4707656,3.9867048,4.3347936,4.6828823,5.029158,5.377247,5.7253356,5.634688,5.5458527,5.4552045,5.3645563,5.275721,4.88956,4.505212,4.120864,3.7347028,3.350355,2.9279346,2.5055144,2.0830941,1.6606737,1.2382535,1.0768998,0.91735905,0.75781834,0.5982776,0.43692398,0.35715362,0.27738327,0.19761293,0.11784257,0.038072214,0.072518505,0.10696479,0.14322405,0.17767033,0.21211663,0.36259252,0.51306844,0.66173136,0.8122072,0.96268314,1.0478923,1.1331016,1.2183108,1.3017071,1.3869164,1.4431182,1.4975071,1.551896,1.6080978,1.6624867,1.7241274,1.7875811,1.8492218,1.9126755,1.9743162,1.9326181,1.889107,1.8474089,1.8057107,1.7621996,2.9478772,4.1317415,5.317419,6.5030966,7.686961,8.435715,9.182655,9.929596,10.6783495,11.42529,11.341894,11.26031,11.176914,11.095331,11.011934,12.052575,13.093216,14.132043,15.172684,16.213324,16.392807,16.57229,16.751774,16.933071,17.112555,17.75978,18.40701,19.054237,19.703278,20.350506,21.378454,22.404593,23.43254,24.460491,25.488441,24.964495,24.442362,23.920229,23.398094,22.87415,21.11195,19.34975,17.58755,15.825351,14.06315,12.931862,11.802386,10.672911,9.541622,8.412147,8.765674,9.117389,9.469104,9.822631,10.174346,10.750868,11.325577,11.900287,12.474996,13.049705,13.274512,13.499319,13.724127,13.9507475,14.175554,14.762955,15.350354,15.937754,16.525154,17.112555,18.234777,19.357002,20.479225,21.603262,22.725487,22.112705,21.499924,20.887142,20.27436,19.663393,18.630003,17.598429,16.565039,15.5334635,14.500074,13.470312,12.440549,11.410787,10.37921,9.349448,8.232663,7.115878,5.99728,4.880495,3.7618973,3.1908143,2.617918,2.0450218,1.4721256,0.89922947,0.7795739,0.65991837,0.5402629,0.42060733,0.2991388,0.24837588,0.19579996,0.14322405,0.09064813,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.36259252,0.69980353,1.0370146,1.3742256,1.7132497,1.3705997,1.0279498,0.6852999,0.34264994,0.0,0.11421664,0.23024625,0.3444629,0.4604925,0.5747091,0.5293851,0.48587397,0.4405499,0.39522585,0.34990177,0.29732585,0.24474995,0.19217403,0.13959812,0.0870222,0.15410182,0.2229944,0.29007402,0.35715362,0.42423326,0.38978696,0.35534066,0.3208944,0.28463513,0.25018883,0.4224203,0.5946517,0.7668832,0.93911463,1.1131591,1.0478923,0.9826257,0.91735905,0.8520924,0.7868258,1.0497054,1.3125849,1.5754645,1.8383441,2.0994108,2.0758421,2.0504606,2.0250793,1.9996977,1.9743162,3.0874753,4.2006345,5.3119802,6.4251394,7.5382986,7.1865835,9.389333,11.592083,13.794832,15.9975815,18.20033,19.866444,21.53437,23.202295,24.87022,26.536333,25.537392,24.536636,23.537693,22.536938,21.537996,22.939415,24.34265,25.744068,27.147303,28.550535,28.708263,28.864178,29.021906,29.179632,29.33736,27.24339,25.147604,23.051819,20.957848,18.862062,18.825804,18.787731,18.749659,18.7134,18.675327,21.768242,24.859343,27.952257,31.045172,34.138084,34.92491,35.71355,36.500374,37.2872,38.07584,36.27557,34.475296,32.675026,30.874752,29.07448,30.20577,31.335245,32.46472,33.59601,34.725487,35.796947,36.87022,37.943493,39.014954,40.08823,36.17767,32.26711,28.35836,24.4478,20.537241,17.58755,14.63786,11.6881695,8.736667,5.7869763,5.2158933,4.6429973,4.070101,3.4972048,2.9243085,3.054842,3.1853752,3.3140955,3.444629,3.5751622,3.1817493,2.7901495,2.3967366,2.0051367,1.6117238,1.6117238,1.6117238,1.6117238,1.6117238,1.6117238,1.7658255,1.9181144,2.0704033,2.222692,2.374981,2.7974012,3.2198215,3.6422417,4.064662,4.4870825,5.3446136,6.202145,7.059676,7.9172077,8.774739,8.767487,8.760235,8.752983,8.745731,8.736667,7.8156815,6.892884,5.9700856,5.047288,4.12449,3.7347028,3.3449159,2.955129,2.565342,2.175555,2.0105755,1.845596,1.6806163,1.5156367,1.3506571,1.452183,1.5555218,1.6570477,1.7603867,1.8619126,2.2879589,2.712192,3.1382382,3.5624714,3.9867048,3.8652363,3.7419548,3.6204863,3.4972048,3.3757362,3.339477,3.3050308,3.2705846,3.2343252,3.199879,2.960568,2.7194438,2.4801328,2.2408218,1.9996977,2.2571385,2.514579,2.7720199,3.0294604,3.2869012,2.9968271,2.7067533,2.4166791,2.126605,1.8383441,1.4775645,1.1167849,0.75781834,0.39703882,0.038072214,0.07795739,0.11784257,0.15772775,0.19761293,0.2374981,0.28463513,0.33177215,0.38072214,0.42785916,0.4749962,0.39522585,0.3154555,0.23568514,0.15410182,0.07433146,0.059827764,0.045324065,0.030820364,0.014503701,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0054388875,0.010877775,0.014503701,0.01994259,0.025381476,0.047137026,0.07070554,0.092461094,0.11421664,0.13778515,0.2520018,0.3680314,0.48224804,0.5982776,0.7124943,0.77232206,0.8321498,0.8919776,0.95180535,1.0116332,1.5156367,2.0178273,2.520018,3.0222087,3.5243993,3.3630457,3.199879,3.0367124,2.8753586,2.712192,2.2118144,1.7132497,1.2128719,0.7124943,0.21211663,0.2755703,0.33721104,0.40066472,0.46230546,0.52575916,0.97174793,1.4195497,1.8673514,2.3151531,2.762955,2.525457,2.2879589,2.0504606,1.8129625,1.5754645,3.8978696,6.2202744,8.54268,10.865085,13.1874895,12.4242325,11.662788,10.899531,10.138086,9.374829,8.39039,7.404139,6.4197006,5.4352617,4.4508233,4.2024474,3.9558845,3.7075086,3.4591327,3.2125697,2.956942,2.7031271,2.4474995,2.1918716,1.938057,3.3322253,4.7282066,6.1223745,7.518356,8.912524,11.477866,14.043208,16.606737,19.17208,21.737421,20.42665,19.117691,17.80692,16.49796,15.187187,13.773077,12.357153,10.943042,9.527119,8.113008,7.9298983,7.746789,7.5654926,7.382384,7.1992745,7.1430726,7.0850577,7.027043,6.970841,6.9128265,6.294606,5.678199,5.0599785,4.441758,3.825351,4.115425,4.405499,4.695573,4.985647,5.275721,5.290225,5.3047285,5.319232,5.335549,5.3500524,4.9983377,4.64481,4.2930956,3.9395678,3.587853,3.0729716,2.5580902,2.0432088,1.5283275,1.0116332,0.88472575,0.75781834,0.629098,0.50219065,0.37528324,0.3045777,0.23568514,0.16497959,0.09427405,0.025381476,0.065266654,0.10515183,0.14503701,0.18492219,0.22480737,0.44961473,0.6744221,0.89922947,1.1258497,1.3506571,1.4141108,1.4793775,1.5446441,1.6099107,1.6751775,1.6080978,1.5392052,1.4721256,1.405046,1.3379664,1.4249886,1.5120108,1.6008459,1.6878681,1.7748904,1.7676386,1.7603867,1.7531348,1.745883,1.7368182,2.8517902,3.966762,5.081734,6.1967063,7.311678,7.9407763,8.568061,9.195346,9.822631,10.449916,10.607644,10.765372,10.9230995,11.080828,11.236742,11.922042,12.607342,13.292642,13.9779415,14.663241,14.683184,14.703127,14.723069,14.743011,14.762955,15.428311,16.091856,16.757214,17.422571,18.087927,19.146698,20.207281,21.267864,22.326633,23.387217,23.26031,23.13159,23.004683,22.877775,22.750868,21.487232,20.22541,18.961775,17.699953,16.438131,15.054841,13.673364,12.290073,10.906783,9.525306,9.635896,9.744674,9.855265,9.965856,10.074633,10.449916,10.825199,11.200482,11.575767,11.949236,12.299138,12.650853,13.000754,13.3506565,13.700559,14.287958,14.875358,15.462758,16.050158,16.637558,17.47696,18.318174,19.157576,19.996977,20.838192,20.149265,19.462152,18.77504,18.087927,17.400814,16.34567,15.290526,14.235382,13.180238,12.125093,11.430729,10.734551,10.040187,9.345822,8.649645,7.4422116,6.2347784,5.027345,3.8199122,2.612479,2.2100015,1.8075237,1.405046,1.0025684,0.6000906,0.52032024,0.4405499,0.36077955,0.27919623,0.19942589,0.16497959,0.13053331,0.09427405,0.059827764,0.025381476,0.01994259,0.014503701,0.010877775,0.0054388875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0072518503,0.014503701,0.02175555,0.030820364,0.038072214,0.53663695,1.0370146,1.5373923,2.03777,2.5381477,2.030518,1.5228885,1.015259,0.5076295,0.0,0.17223145,0.3444629,0.5166943,0.69073874,0.8629702,0.78319985,0.7016165,0.62184614,0.5420758,0.46230546,0.38978696,0.31726846,0.24474995,0.17223145,0.099712946,0.20667773,0.3154555,0.4224203,0.5293851,0.63816285,0.56020546,0.48224804,0.40429065,0.32814622,0.25018883,0.41516843,0.58014804,0.7451276,0.9101072,1.0750868,1.015259,0.9554313,0.89560354,0.83577573,0.774135,1.1131591,1.4503701,1.7875811,2.124792,2.4620032,2.4130533,2.3622901,2.3133402,2.2625773,2.2118144,3.1382382,4.062849,4.98746,5.9120708,6.836682,5.6256227,6.8203654,8.015107,9.20985,10.4045925,11.599335,12.565643,13.53014,14.494636,15.459132,16.425442,15.937754,15.4500675,14.96238,14.474693,13.987006,16.820667,19.652514,22.484362,25.318022,28.14987,29.322857,30.495844,31.667017,32.840004,34.012993,31.677895,29.3428,27.007704,24.672607,22.337511,22.411844,22.487988,22.562319,22.638464,22.712795,26.790148,30.8675,34.944855,39.022205,43.09956,44.28705,45.47454,46.66203,47.84952,49.03701,46.638462,44.2381,41.837738,39.437374,37.037014,38.603413,40.168,41.732586,43.297173,44.86176,46.31757,47.773376,49.22737,50.68318,52.137177,46.982925,41.828674,36.672607,31.518354,26.36229,22.500679,18.637255,14.775645,10.912222,7.0506115,6.207584,5.3645563,4.5233417,3.680314,2.8372865,2.8155308,2.7919624,2.770207,2.7466383,2.7248828,2.3967366,2.0704033,1.742257,1.4141108,1.0877775,1.1258497,1.162109,1.2001812,1.2382535,1.2745126,1.4322405,1.5899682,1.7476959,1.9054236,2.0631514,2.6306088,3.198066,3.7655232,4.3329806,4.900438,5.99728,7.0941224,8.192778,9.28962,10.388275,10.390089,10.391902,10.395528,10.397341,10.399154,9.195346,7.989726,6.784106,5.580299,4.3746786,3.966762,3.5606585,3.152742,2.7448254,2.3369088,2.1302311,1.9217403,1.7150626,1.5083848,1.2998942,1.357909,1.4141108,1.4721256,1.5301404,1.5881553,1.9996977,2.4130533,2.8245957,3.2379513,3.6494937,3.5443418,3.43919,3.3358512,3.2306993,3.1255474,2.956942,2.7901495,2.6233568,2.4547513,2.2879589,2.0540867,1.8220274,1.5899682,1.357909,1.1258497,1.4104849,1.69512,1.9797552,2.2643902,2.5508385,2.268016,1.9851941,1.7023718,1.4195497,1.1367276,0.91917205,0.7016165,0.48587397,0.26831847,0.05076295,0.09427405,0.13959812,0.18492219,0.23024625,0.2755703,0.26831847,0.25925365,0.2520018,0.24474995,0.2374981,0.19761293,0.15772775,0.11784257,0.07795739,0.038072214,0.030820364,0.02175555,0.014503701,0.0072518503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0018129626,0.0054388875,0.0072518503,0.010877775,0.012690738,0.04169814,0.072518505,0.10333887,0.13234627,0.16316663,0.3208944,0.47680917,0.6345369,0.79226464,0.9499924,1.0297627,1.1095331,1.1893034,1.2708868,1.3506571,1.9199274,2.4891977,3.0602808,3.6295512,4.2006345,3.825351,3.4500678,3.0747845,2.6995013,2.324218,1.8999848,1.4757515,1.0497054,0.62547207,0.19942589,0.28826106,0.37528324,0.46230546,0.5493277,0.63816285,1.0551442,1.4721256,1.889107,2.3079014,2.7248828,2.4366217,2.1501737,1.8619126,1.5754645,1.2872034,3.6059825,5.922949,8.239915,10.556881,12.87566,11.974618,11.075388,10.174346,9.275117,8.375887,7.3570023,6.33993,5.3228583,4.305786,3.2869012,3.207131,3.1273603,3.04759,2.9678197,2.8880494,2.7466383,2.6070402,2.467442,2.327844,2.1882458,3.8851788,5.582112,7.2808576,8.977791,10.674724,13.220123,15.765523,18.310923,20.85451,23.399908,21.256987,19.115877,16.972956,14.830034,12.687112,11.50506,10.323009,9.139144,7.957093,6.775041,7.0143523,7.2554765,7.494787,7.7359114,7.9752226,7.8646317,7.755854,7.645263,7.5346723,7.4258947,6.6717024,5.919323,5.1669436,4.4145637,3.6621845,3.8942437,4.1281157,4.360175,4.592234,4.8242936,4.945762,5.0654173,5.185073,5.3047285,5.424384,5.105303,4.784408,4.465327,4.1444325,3.825351,3.2180085,2.610666,2.0033236,1.3941683,0.7868258,0.69255173,0.5982776,0.50219065,0.40791658,0.31182957,0.2520018,0.19217403,0.13234627,0.072518505,0.012690738,0.058014803,0.10333887,0.14684997,0.19217403,0.2374981,0.53663695,0.8375887,1.1367276,1.4376793,1.7368182,1.7821422,1.8274662,1.8727903,1.9181144,1.9616255,1.7730774,1.5827163,1.3923552,1.2019942,1.0116332,1.1258497,1.2382535,1.3506571,1.4630609,1.5754645,1.6026589,1.6298534,1.6570477,1.6842422,1.7132497,2.7575161,3.8017826,4.847862,5.8921285,6.9382076,7.4458375,7.951654,8.459284,8.966913,9.474543,9.873394,10.270433,10.667472,11.06451,11.463363,11.793322,12.123281,12.45324,12.783199,13.113158,12.971747,12.8321495,12.692551,12.552953,12.413355,13.095029,13.776703,14.46019,15.141864,15.825351,16.916754,18.00997,19.103188,20.19459,21.287807,21.554312,21.82263,22.089136,22.357454,22.625772,21.862516,21.099258,20.337814,19.574556,18.813112,17.17782,15.542528,13.907236,12.271944,10.636651,10.504305,10.371959,10.239613,10.107266,9.97492,10.150778,10.324821,10.500679,10.674724,10.850581,11.325577,11.800573,12.27557,12.750566,13.225562,13.812962,14.400362,14.9877615,15.575162,16.162561,16.719141,17.277533,17.834112,18.392506,18.949085,18.187641,17.424383,16.66294,15.899682,15.138238,14.059525,12.982625,11.9057255,10.827013,9.750113,9.389333,9.030367,8.669587,8.31062,7.949841,6.6517596,5.3554916,4.0574102,2.759329,1.4630609,1.2291887,0.99712944,0.7650702,0.533011,0.2991388,0.25925365,0.21936847,0.1794833,0.13959812,0.099712946,0.08339628,0.065266654,0.047137026,0.030820364,0.012690738,0.010877775,0.0072518503,0.0054388875,0.0018129626,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.010877775,0.01994259,0.030820364,0.03988518,0.05076295,0.7124943,1.3742256,2.03777,2.6995013,3.3630457,2.6904364,2.0178273,1.3452182,0.6726091,0.0,0.23024625,0.4604925,0.69073874,0.91917205,1.1494182,1.0352017,0.91917205,0.80495536,0.69073874,0.5747091,0.48224804,0.38978696,0.29732585,0.20486477,0.11240368,0.25925365,0.40791658,0.55476654,0.7016165,0.85027945,0.7306239,0.6091554,0.4894999,0.36984438,0.25018883,0.40791658,0.5656443,0.72337204,0.8792868,1.0370146,0.9826257,0.92823684,0.872035,0.81764615,0.76325727,1.1747998,1.5881553,1.9996977,2.4130533,2.8245957,2.7502642,2.6741197,2.5997884,2.525457,2.4493124,3.1871881,3.925064,4.6629395,5.4008155,6.1368785,4.062849,4.249584,4.4381323,4.6248674,4.8116026,5.0001507,5.2630305,5.524097,5.7869763,6.049856,6.3127356,6.338117,6.3616858,6.3870673,6.412449,6.43783,10.700105,14.96238,19.224655,23.48693,27.749205,29.93745,32.125698,34.31213,36.500374,38.68681,36.1124,33.537994,30.961775,28.387367,25.812962,25.999697,26.188244,26.374979,26.561714,26.750263,31.812054,36.87566,41.93745,46.99924,52.062847,53.64919,55.237343,56.8255,58.411842,59.999996,56.999542,54.000904,51.00045,47.999996,44.999546,46.99924,49.00075,51.00045,53.00015,54.999847,56.83819,58.67472,60.513065,62.349598,64.18794,57.78818,51.388424,44.986855,38.587097,32.187336,27.411995,22.638464,17.863121,13.087777,8.312433,7.1992745,6.0879283,4.974769,3.8616104,2.7502642,2.5744069,2.4003625,2.2245052,2.0504606,1.8746033,1.6117238,1.3506571,1.0877775,0.824898,0.5620184,0.63816285,0.7124943,0.7868258,0.8629702,0.93730164,1.1004683,1.261822,1.4249886,1.5881553,1.7495089,2.4620032,3.1744974,3.8869917,4.599486,5.3119802,6.6499467,7.987913,9.325879,10.662033,11.999999,12.012691,12.025381,12.038072,12.050762,12.06164,10.57501,9.088382,7.5999393,6.11331,4.6248674,4.2006345,3.774588,3.350355,2.9243085,2.5000753,2.2498865,1.9996977,1.7495089,1.49932,1.2491312,1.261822,1.2745126,1.2872034,1.2998942,1.3125849,1.7132497,2.1121013,2.5127661,2.911618,3.3122826,3.2252605,3.1382382,3.049403,2.962381,2.8753586,2.5744069,2.275268,1.9743162,1.6751775,1.3742256,1.1494182,0.9246109,0.69980353,0.4749962,0.25018883,0.5620184,0.87566096,1.1874905,1.49932,1.8129625,1.5373923,1.261822,0.9880646,0.7124943,0.43692398,0.36259252,0.28826106,0.21211663,0.13778515,0.06164073,0.11240368,0.16316663,0.21211663,0.26287958,0.31182957,0.25018883,0.18673515,0.12509441,0.06164073,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.038072214,0.07433146,0.11240368,0.15047589,0.18673515,0.387974,0.5873999,0.7868258,0.9880646,1.1874905,1.2872034,1.3869164,1.4866294,1.5881553,1.6878681,2.324218,2.962381,3.6005437,4.2368937,4.8750563,4.2876563,3.7002566,3.1128569,2.525457,1.938057,1.5881553,1.2382535,0.8883517,0.53663695,0.18673515,0.2991388,0.41335547,0.52575916,0.63816285,0.7505665,1.1367276,1.5247015,1.9126755,2.3006494,2.6868105,2.3495996,2.0123885,1.6751775,1.3379664,1.0007553,3.3122826,5.6256227,7.93715,10.25049,12.562017,11.525003,10.487988,9.449161,8.412147,7.3751316,6.3254266,5.275721,4.2242026,3.1744974,2.124792,2.2118144,2.3006494,2.3876717,2.474694,2.561716,2.5381477,2.5127661,2.4873846,2.4620032,2.4366217,4.4381323,6.43783,8.437528,10.437225,12.436923,14.96238,17.487837,20.013294,22.536938,25.062395,22.087322,19.112251,16.13718,13.162108,10.1870365,9.237044,8.287052,7.3370595,6.3870673,5.4370747,6.1006193,6.7623506,7.4258947,8.087626,8.749357,8.588004,8.424837,8.26167,8.100317,7.93715,7.0506115,6.16226,5.275721,4.3873696,3.5008307,3.6748753,3.8507326,4.024777,4.2006345,4.3746786,4.599486,4.8242936,5.049101,5.275721,5.5005283,5.2122674,4.9258194,4.6375585,4.349297,4.062849,3.3630457,2.663242,1.9616255,1.261822,0.5620184,0.50037766,0.43692398,0.37528324,0.31182957,0.25018883,0.19942589,0.15047589,0.099712946,0.05076295,0.0,0.05076295,0.099712946,0.15047589,0.19942589,0.25018883,0.62547207,1.0007553,1.3742256,1.7495089,2.124792,2.1501737,2.175555,2.1991236,2.2245052,2.2498865,1.938057,1.6244144,1.3125849,1.0007553,0.6871128,0.824898,0.96268314,1.1004683,1.2382535,1.3742256,1.4376793,1.49932,1.5627737,1.6244144,1.6878681,2.663242,3.636803,4.612177,5.5875506,6.5629244,6.9508986,7.3370595,7.7250338,8.113008,8.499168,9.137331,9.775495,10.411844,11.050007,11.6881695,11.662788,11.637406,11.612025,11.586644,11.563075,11.262123,10.962985,10.662033,10.362894,10.061942,10.761745,11.463363,12.163166,12.862969,13.562773,14.68681,15.812659,16.936697,18.062546,19.188396,19.850128,20.511858,21.175404,21.837133,22.500679,22.237799,21.97492,21.71204,21.44916,21.188093,19.298986,17.411694,15.524399,13.637105,11.74981,11.374527,10.999244,10.625773,10.25049,9.875207,9.849826,9.824444,9.800876,9.775495,9.750113,10.3502035,10.950294,11.5503845,12.1504755,12.750566,13.337966,13.925365,14.512766,15.100165,15.687565,15.963136,16.236893,16.512463,16.788034,17.06179,16.224201,15.388427,14.5508375,13.713249,12.87566,11.775192,10.674724,9.574255,8.4756,7.3751316,7.3497505,7.324369,7.3008003,7.2754188,7.250037,5.863121,4.4743915,3.0874753,1.7005589,0.31182957,0.25018883,0.18673515,0.12509441,0.06164073,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.012690738,0.025381476,0.038072214,0.05076295,0.06164073,0.8883517,1.7132497,2.5381477,3.3630457,4.1879435,3.350355,2.5127661,1.6751775,0.8375887,0.0,0.28826106,0.5747091,0.8629702,1.1494182,1.4376793,1.2872034,1.1367276,0.9880646,0.8375887,0.6871128,0.5747091,0.46230546,0.34990177,0.2374981,0.12509441,0.31182957,0.50037766,0.6871128,0.87566096,1.062396,0.89922947,0.73787576,0.5747091,0.41335547,0.25018883,0.40066472,0.5493277,0.69980353,0.85027945,1.0007553,0.9499924,0.89922947,0.85027945,0.7995165,0.7505665,1.2382535,1.7259403,2.2118144,2.6995013,3.1871881,3.0874753,2.9877625,2.8880494,2.7883365,2.6868105,3.2379513,3.787279,4.3384194,4.8877473,5.4370747;
 } 
