netcdf QPE_CPC_CMORPH.2018062700{
dimensions: 
 lat = 180; 
 lon = 281; 
variables:  
float lat(lat) ; 
   lat:long_name = "latitude" ;
   lat:units = "degrees_north" ;
   lat:standard_name = "latitude" ;
float lon(lon) ;
   lon:long_name = "longitude" ;
   lon:units = "degrees_east" ;
   lon:standard_name = "longitude" ;
float APCP_24(lat, lon) ;
   APCP_24:name = "APCP_24" ;
   APCP_24:long_name = "Total Precipitation" ;
   APCP_24:level = "A24" ;
   APCP_24:units = "kg/m^2" ;
   APCP_24:_FillValue = -9999.f ;
   APCP_24:init_time = "20180626_000000" ;
   APCP_24:init_time_ut = "1529971200.0" ;
   APCP_24:valid_time = "20180627_000000" ;
   APCP_24:valid_time_ut = "1530057600.0" ;
   APCP_24:accum_time = "240000" ;
   APCP_24:_FillValue = -9.99e8 ;
   APCP_24:accum_time_sec = 86400 ;
 // global attributes: 
 :_NCProperties = "version=1|netcdflibversion=4.4.1.1|hdf5libversion=1.8.12" ;
	:FileOrigins = "CPC_CMORPH_DAILY_PRCP" ; 
	:MET_version = "V7.0" ;
	:Projection = "LatLon" ;
	:lat_ll = "15.125 degrees_north" ; 
	:lon_ll = "70.125 degrees_east" ; 
	:delta_lat = "0.250000 degrees" ;
	:delta_lon = "0.250000 degrees" ;
	:Nlat = "180 grid_points" ; 
	:Nlon = "281 grid_points" ; 
data:
lat = 15.125,15.375,15.625,15.875,16.125,16.375,16.625,16.875,17.125,17.375,17.625,17.875,18.125,18.375,18.625,18.875,19.125,19.375,19.625,19.875,20.125,20.375,20.625,20.875,21.125,21.375,21.625,21.875,22.125,22.375,22.625,22.875,23.125,23.375,23.625,23.875,24.125,24.375,24.625,24.875,25.125,25.375,25.625,25.875,26.125,26.375,26.625,26.875,27.125,27.375,27.625,27.875,28.125,28.375,28.625,28.875,29.125,29.375,29.625,29.875,30.125,30.375,30.625,30.875,31.125,31.375,31.625,31.875,32.125,32.375,32.625,32.875,33.125,33.375,33.625,33.875,34.125,34.375,34.625,34.875,35.125,35.375,35.625,35.875,36.125,36.375,36.625,36.875,37.125,37.375,37.625,37.875,38.125,38.375,38.625,38.875,39.125,39.375,39.625,39.875,40.125,40.375,40.625,40.875,41.125,41.375,41.625,41.875,42.125,42.375,42.625,42.875,43.125,43.375,43.625,43.875,44.125,44.375,44.625,44.875,45.125,45.375,45.625,45.875,46.125,46.375,46.625,46.875,47.125,47.375,47.625,47.875,48.125,48.375,48.625,48.875,49.125,49.375,49.625,49.875,50.125,50.375,50.625,50.875,51.125,51.375,51.625,51.875,52.125,52.375,52.625,52.875,53.125,53.375,53.625,53.875,54.125,54.375,54.625,54.875,55.125,55.375,55.625,55.875,56.125,56.375,56.625,56.875,57.125,57.375,57.625,57.875,58.125,58.375,58.625,58.875,59.125,59.375,59.625,59.875;
lon = 70.125,70.375,70.625,70.875,71.125,71.375,71.625,71.875,72.125,72.375,72.625,72.875,73.125,73.375,73.625,73.875,74.125,74.375,74.625,74.875,75.125,75.375,75.625,75.875,76.125,76.375,76.625,76.875,77.125,77.375,77.625,77.875,78.125,78.375,78.625,78.875,79.125,79.375,79.625,79.875,80.125,80.375,80.625,80.875,81.125,81.375,81.625,81.875,82.125,82.375,82.625,82.875,83.125,83.375,83.625,83.875,84.125,84.375,84.625,84.875,85.125,85.375,85.625,85.875,86.125,86.375,86.625,86.875,87.125,87.375,87.625,87.875,88.125,88.375,88.625,88.875,89.125,89.375,89.625,89.875,90.125,90.375,90.625,90.875,91.125,91.375,91.625,91.875,92.125,92.375,92.625,92.875,93.125,93.375,93.625,93.875,94.125,94.375,94.625,94.875,95.125,95.375,95.625,95.875,96.125,96.375,96.625,96.875,97.125,97.375,97.625,97.875,98.125,98.375,98.625,98.875,99.125,99.375,99.625,99.875,100.125,100.375,100.625,100.875,101.125,101.375,101.625,101.875,102.125,102.375,102.625,102.875,103.125,103.375,103.625,103.875,104.125,104.375,104.625,104.875,105.125,105.375,105.625,105.875,106.125,106.375,106.625,106.875,107.125,107.375,107.625,107.875,108.125,108.375,108.625,108.875,109.125,109.375,109.625,109.875,110.125,110.375,110.625,110.875,111.125,111.375,111.625,111.875,112.125,112.375,112.625,112.875,113.125,113.375,113.625,113.875,114.125,114.375,114.625,114.875,115.125,115.375,115.625,115.875,116.125,116.375,116.625,116.875,117.125,117.375,117.625,117.875,118.125,118.375,118.625,118.875,119.125,119.375,119.625,119.875,120.125,120.375,120.625,120.875,121.125,121.375,121.625,121.875,122.125,122.375,122.625,122.875,123.125,123.375,123.625,123.875,124.125,124.375,124.625,124.875,125.125,125.375,125.625,125.875,126.125,126.375,126.625,126.875,127.125,127.375,127.625,127.875,128.125,128.375,128.625,128.875,129.125,129.375,129.625,129.875,130.125,130.375,130.625,130.875,131.125,131.375,131.625,131.875,132.125,132.375,132.625,132.875,133.125,133.375,133.625,133.875,134.125,134.375,134.625,134.875,135.125,135.375,135.625,135.875,136.125,136.375,136.625,136.875,137.125,137.375,137.625,137.875,138.125,138.375,138.625,138.875,139.125,139.375,139.625,139.875,140.125;
APCP_24 = 0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.041666668,0.9777778,2.0833335,5.0444446,3.8416667,1.5777779,0.3,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06666667,0.44444445,2.677778,4.1333337,2.4777777,0.68333334,0.5222223,1.2750001,1.0888889,0.32222223,0.0,0.0,0.175,2.688889,9.5,15.288889,18.955557,24.541668,29.622225,28.000004,27.288887,24.941666,24.644445,11.891666,3.488889,5.633334,11.241666,13.9,18.941668,22.677778,17.525,14.044445,12.733334,7.2000003,6.455556,6.816666,9.366667,15.733334,30.277779,40.19167,41.755554,81.82222,62.033333,55.68889,51.300003,52.91111,46.625,46.877777,49.511112,51.566673,57.577778,55.825005,45.67778,34.841667,25.466667,25.366667,29.616667,30.988888,20.941668,14.211112,13.816667,16.57778,22.350002,21.333334,21.3,23.65,28.9,33.983334,39.177776,38.000004,26.722223,19.466667,18.016666,18.266668,19.191668,28.266666,33.46667,22.188889,7.7,4.7000003,6.477778,6.658334,5.3555555,6.191667,4.5111113,3.9250002,2.4444442,3.0555556,1.7749999,3.5111113,10.0,22.155556,12.058334,11.677778,26.144445,31.008335,20.188887,10.874999,10.155557,9.633334,7.111111,7.675,10.455556,12.411111,15.391667,10.622223,1.5333334,1.5111113,6.8250003,25.51111,44.344448,48.274998,18.51111,8.675,4.966667,0.8833334,3.777778,9.183333,14.277778,10.077778,28.041668,44.27778,7.566666,2.0222223,0.45833334,0.07777778,0.011111111,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.3,2.4250002,7.188889,14.591665,16.2,11.325001,8.477777,10.144444,10.641666,13.688889,11.816668,15.577778,19.891666,27.955555,30.308334,33.733334,31.811113,27.541666,35.711113,50.425003,54.444443,51.108334,50.444443,41.955555,27.6,19.522223,12.541668,5.8444448,0.6750001,0.3333333,0.78333336,1.4444445,5.366667,10.583334,11.088889,15.358334,8.688889,1.9583334,0.988889,1.0222223,0.33333337,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.26666668,1.5,4.8444443,11.116666,12.944445,3.2333336,1.075,2.5444443,2.9333334,0.8666667,0.19166669,0.0,0.0,0.0,0.022222223,0.23333333,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.075,0.7777778,1.0666668,0.5083334,0.50000006,0.8666667,0.74444443,0.60833335,0.97777784,3.1333337,10.466667,16.41111,17.866667,19.466667,21.433334,23.288889,21.755556,20.416668,12.533333,6.6000004,2.6444445,0.84999996,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.033333335,0.033333335,0.9444445,2.5,6.777778,7.966666,4.8,2.3555558,0.85833335,0.5222222,0.40833333,0.34444445,0.21666667,0.1,0.044444446,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.033333335,0.9000001,3.85,6.1333337,2.7,0.35555556,0.45833334,1.2777778,1.7,0.8833334,1.2333332,4.05,5.833334,8.316667,12.522222,19.477777,26.016668,33.144447,37.85,40.544445,47.383335,62.98889,28.691668,10.955557,8.777779,7.533334,8.911112,10.258334,13.055555,10.858333,8.077778,6.777778,7.0583344,7.822222,8.633333,10.233334,14.966667,27.7,50.13333,70.7,97.16667,97.37501,79.21111,62.000004,45.18889,44.100006,42.211113,44.677776,44.833336,46.58889,41.725002,30.255558,24.833334,27.811111,29.844444,32.3,35.944447,33.258335,24.055555,21.991669,24.0,25.533333,21.966667,20.344444,22.125,24.866665,30.941666,37.52222,37.800003,28.47778,21.944445,18.749998,19.28889,26.483334,30.866673,29.741669,25.444445,10.191667,5.566667,7.2777777,8.2,7.822222,7.175,6.0555553,3.2333333,1.8111112,1.4444445,1.1666666,1.4222223,4.525,20.044445,25.766665,16.433334,22.955559,35.483334,34.36667,14.800001,7.4000006,8.233334,8.077778,5.3,8.111111,14.388888,21.383333,9.277778,1.6333333,0.94444454,5.683333,22.955559,39.01111,45.55,11.900001,10.6,7.6888885,3.8250003,5.5000005,13.775,27.833334,34.4,30.833332,28.011112,12.266666,1.8444446,0.5666666,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.4222222,2.5083337,5.3,13.683333,13.511111,9.258333,7.955556,8.5222225,12.599999,22.38889,20.566668,23.344444,25.116669,37.988888,50.75833,59.81111,58.566666,41.575,34.52222,34.850002,31.944447,33.55,40.622227,43.72222,39.608334,42.844448,49.591663,16.866667,4.4583335,0.7111112,0.87499994,1.4666667,9.4777775,13.424999,18.422222,20.24167,13.755555,4.491667,0.72222227,0.96666676,0.7916666,0.055555556,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06666667,0.21666667,1.4444445,12.216666,10.344444,2.9444447,0.9333334,0.48888892,1.4,0.4333333,0.025000002,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.116666675,0.57777774,1.9555556,2.3333335,1.7666668,1.7583331,2.0555556,1.3833333,0.96666664,2.1444447,8.491667,20.8,30.916666,35.86667,35.733334,31.533333,32.755558,35.041664,24.766666,14.25,8.3,3.9166667,0.08125,0.10833335,0.0,0.08125,0.7666667,0.19375,0.0,0.0,0.0,0.0,0.05,0.083333336,0.23750001,2.025,6.1375,14.633333,17.675001,13.625,7.891667,2.8625,0.85833335,0.33125,0.17500001,0.15,0.083333336,0.033333335,0.0,0.0,0.00625,0.0,0.0,0.0,0.0,0.1,0.19999999,0.83125,1.5333333,1.2125,1.0166667,0.20625,0.40833336,1.7250001,2.3625,2.075,4.30625,8.241667,13.03125,16.7,20.008333,25.66875,32.71667,37.068752,43.11667,45.75625,42.9,32.60625,19.25,10.45,5.2875,4.7750006,6.33125,6.55,6.625,6.641667,7.4000006,8.23125,9.933333,11.806251,14.666666,16.824999,23.15,40.93125,80.96667,110.05833,124.8375,117.125,95.256256,60.408337,53.91875,45.308334,42.641666,44.387505,47.7,41.2,33.508335,24.025002,25.566666,23.716667,25.35625,26.0,31.10625,36.691666,38.675,36.64167,34.212505,20.416668,16.758335,15.2875,15.391667,18.1375,22.275,21.33125,24.508333,26.191668,20.593752,14.799999,16.0375,16.116667,18.70625,19.000002,13.8625,11.991668,9.058333,9.34375,14.316667,22.7125,26.8,18.65625,8.166666,2.675,2.6312501,1.2333335,3.6062503,13.283334,16.10625,12.891668,12.575001,15.825,23.483335,23.78125,12.233334,11.981251,15.691667,3.54375,4.6749997,12.441667,17.475,11.941666,5.09375,1.8083335,2.8062499,7.4333334,13.783334,20.9375,8.191667,6.1562505,5.7666674,4.825,6.1,21.574999,34.93333,43.933334,23.8625,6.241667,10.31875,3.4666667,0.21875001,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.6666667,7.0812507,7.158334,6.45,9.841666,12.841666,15.250001,32.508335,34.7625,24.491667,24.90625,29.39167,30.012499,29.491665,28.500002,29.35,33.183334,37.4375,41.324997,39.04375,34.4,38.574997,40.906246,42.908337,52.962505,36.716667,12.91875,5.5750003,3.1687498,4.008333,12.283333,13.00625,12.716668,8.43125,7.6916666,8.30625,3.0583334,1.1833333,1.2,0.23333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.275,2.2666667,6.1187506,11.425,12.13125,7.975,10.737501,9.283334,3.4333332,1.5500001,0.09166667,0.0125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.24166667,1.1250001,3.525,4.55,3.5875003,2.1166668,2.28125,1.85,2.8583333,6.5,13.1,25.281252,34.65,42.287502,43.85833,42.091667,43.425003,35.800003,23.00625,14.650002,11.106252,0.0,0.0,0.0,0.108333334,0.46666667,0.35833335,0.0,0.0,0.07777778,0.22222224,0.4916667,1.111111,1.2666667,1.6222223,3.4083333,5.1888895,9.541666,7.211111,4.277778,1.9416666,0.78888893,0.275,0.1,0.0,0.0,0.0,0.0,0.0,0.058333337,0.25555557,0.18333334,0.022222223,1.2750001,0.62222224,0.9555557,3.3583336,1.4888889,0.016666668,0.32222223,0.9666667,0.5777778,0.7222222,1.1333332,1.6777776,4.0916667,6.0000005,9.591667,12.511111,14.944445,17.85,21.733334,28.341667,33.888885,36.24167,28.633335,24.883335,25.66667,17.633333,7.25,5.633333,6.5250006,7.411111,6.925,7.111111,9.2,10.333334,11.933334,14.700001,18.555555,23.24167,29.266666,35.43334,52.255558,65.57778,81.50833,88.0,89.674995,81.03333,69.833336,70.6,77.27779,75.416664,65.66667,57.775005,49.755558,37.566666,25.47778,23.377777,21.791666,21.2,29.291666,45.077778,53.208336,43.444443,38.608334,30.177776,15.300001,6.6750007,3.6777775,3.2416668,7.8333335,12.983334,19.677776,23.677776,25.458334,25.311111,21.866667,18.1,15.15,14.866667,9.35,14.6,24.044445,14.049999,8.633334,25.933334,45.06667,50.90833,37.633335,17.600002,4.6333337,4.211111,4.091667,6.9555554,14.891666,17.733334,17.033335,16.008335,16.533333,26.466667,25.022223,9.116667,14.755556,10.008333,1.8111112,3.8222225,7.2666664,7.9555554,5.525,2.3777778,3.3083334,3.8000004,3.3555555,4.858333,3.1777782,2.716667,2.4222224,3.4166667,4.677778,21.566668,42.555557,46.26667,26.2,5.1555557,1.5083333,3.1333337,0.11666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.022222223,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.42222226,2.325,3.7111113,8.408334,10.411112,10.022222,14.608334,25.933332,21.608334,17.811111,21.416668,22.755556,11.316667,3.6333334,5.3888893,14.491667,26.099998,38.375,46.91111,48.10833,49.15556,53.67778,52.016663,42.488888,49.90833,56.000004,32.46667,22.633333,20.916666,16.722223,16.288887,17.16667,12.133334,10.025001,5.133333,5.6916666,4.9,2.5333335,1.2416668,0.56666666,0.1,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.7222222,3.4833336,9.244444,18.033335,24.211111,20.658333,12.51111,3.388889,0.5833333,0.022222223,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011111111,3.477778,6.7916665,10.688889,13.575,14.2,10.775,6.2222223,3.4,2.0249999,5.3111115,11.05,15.866667,19.291668,21.01111,20.677778,19.891666,17.844444,15.166665,12.0,12.666667,0.13749999,0.2,0.17500001,0.2875,0.21666665,0.30625,0.5416667,0.6625,0.775,1.0833334,1.6250001,3.5749998,6.2749996,6.633333,10.61875,12.758334,10.10625,7.05,5.2833333,3.7125,2.3250003,1.1375,0.40000004,0.0375,0.0,0.0,0.0,0.0,0.0,0.0,0.06875,0.0,0.51875,0.93333334,0.67499995,1.9562501,3.0333333,1.6187502,0.7333334,0.20625001,0.24166667,0.4583333,1.075,1.7583334,3.2124999,4.35,4.0687504,5.3500004,6.9750004,8.8375,10.033335,14.356251,18.941668,21.368752,21.7,19.95625,17.258335,14.483333,8.500001,5.325,5.925,7.983333,7.8375006,6.8500004,8.708334,11.85,13.291668,19.556248,27.783335,34.193752,39.766666,43.925003,51.174995,60.658333,64.793755,66.091675,62.468754,64.4,61.387497,73.274994,79.433334,82.43751,71.691666,63.9375,67.541664,63.687504,45.008335,32.658333,24.300001,23.916668,33.93125,54.0,71.0625,75.7,57.59375,50.316666,40.850002,19.337502,6.3583336,1.3750001,0.40833336,2.90625,6.616667,9.033333,11.93125,14.216667,14.950001,18.341667,14.675,8.966667,4.70625,9.45,19.283335,20.012499,9.391667,8.581249,15.75,26.000002,33.808334,32.625,14.487499,3.0333333,4.0062504,6.0333333,6.7875,14.458333,21.691666,20.99375,17.408333,19.44375,25.59167,9.1125,2.1083333,8.862501,3.4333334,0.30833334,1.7125,3.741667,2.68125,3.3916667,2.3624997,3.1833334,3.1416667,3.10625,2.4916668,4.36875,2.7833333,2.3937502,2.6166666,8.70625,23.366669,42.13334,19.525,3.5333335,0.30625,0.24166667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.050000004,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.24166667,2.1499999,4.491667,6.8999996,7.1083336,8.683332,11.650001,8.741667,7.6999993,12.133333,24.1875,25.833334,15.493751,4.333333,1.6999999,3.66875,9.874999,19.08125,31.266666,39.1625,43.14167,40.808334,31.443748,26.849998,30.918753,58.56667,45.34375,23.699999,14.13125,7.6333337,3.6916668,4.1125,4.333333,6.2374997,3.7499998,1.01875,1.6083335,0.9833333,0.51875,0.5416667,0.29375002,0.041666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.18125,0.8166667,2.15625,3.5333335,3.9499998,3.0,2.166667,1.08125,0.60833335,0.10000001,0.0,0.0,0.05,0.0625,0.06666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05,0.54375005,2.6250002,5.6,7.3250003,11.7125,16.658335,15.724999,12.299999,12.1,13.706251,15.133333,13.4875,8.799999,4.9166665,2.8437498,2.891667,4.50625,4.908334,6.4875,8.85,11.35,13.25,14.141667,14.8875,15.316665,15.51875,0.275,0.07777778,0.22222222,0.25,0.022222223,0.38333333,1.8222222,1.9666667,2.3555558,3.7,6.4500003,10.677776,15.608334,13.266666,9.433333,10.388888,11.333334,7.7333336,6.255556,4.425,2.7777777,1.7666668,0.62222224,0.116666675,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011111111,0.05555556,0.18333334,0.3,0.19166666,0.13333333,0.07500001,0.0,0.45555556,1.8583333,3.3111115,2.4916668,3.3666668,2.4416668,2.488889,3.5444446,4.9833336,5.311111,6.908334,8.722222,9.616667,10.788889,12.025,9.122222,5.777778,3.6583333,2.8777778,4.266667,7.2777777,8.608334,7.8444448,9.011111,12.116666,14.1,18.458334,28.266666,41.516666,49.77778,55.408333,58.47778,62.61111,60.350002,63.177773,57.041664,54.499996,55.891666,62.933334,72.12222,77.3,75.511116,68.00833,67.9,71.05,66.600006,48.5,35.841667,32.377777,45.583336,73.9,82.39167,75.333336,76.89166,72.91112,68.94445,49.75833,26.588892,8.424999,1.3222222,2.1166666,2.1555555,0.9,2.3166666,2.7888892,5.758333,11.4777775,10.25,4.877778,3.8416667,3.5333335,5.0666666,9.216667,10.788889,9.366667,11.1,13.008333,13.588888,17.044445,13.300002,5.1000004,1.9583334,4.855556,9.816668,12.122222,18.655556,30.1,29.433334,26.816668,26.98889,14.891668,0.8111111,4.383333,5.0444446,1.4666667,0.6166667,0.8111111,1.6833334,2.3666666,1.3000001,1.9777778,1.6222224,2.0,2.488889,2.2833335,3.2111113,2.0333333,0.6222222,3.091667,7.5888886,11.855556,11.950001,3.688889,0.36666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.43333334,2.1916666,5.3888893,4.633333,5.211111,8.244445,7.5083337,4.8888893,6.8916674,11.766667,20.866667,25.78889,23.224998,12.177778,5.088889,1.1000001,0.055555556,0.041666668,1.0222223,6.033334,23.033333,32.122223,31.683334,34.122223,29.84167,30.055557,26.75,24.077778,13.358334,5.0,2.4666667,0.675,0.61111116,1.075,3.8111115,0.475,0.011111111,0.011111111,0.15,0.13333334,0.20833336,0.0,0.0,0.0,0.0,0.0,0.0,0.3,0.73333335,1.15,1.4666667,0.20000002,0.0,0.0,0.0,0.0,0.0,0.0,0.050000004,0.0,0.0,0.033333335,2.0666666,1.1999999,0.0,0.008333334,0.24444444,0.46666667,1.7333333,2.7222223,2.475,1.4777777,0.38333333,0.0,0.0,0.0,0.0,0.0,0.055555556,1.25,4.022222,7.2833333,11.044445,14.075,18.011112,17.111113,12.541667,10.300001,9.991667,11.355556,12.316668,10.555555,8.422222,6.4500003,4.8222227,4.0916667,3.3000002,3.7083335,4.677778,6.61111,9.400002,11.833334,13.416668,12.533334,13.041667,0.29999998,0.8666667,0.8666666,0.98749995,0.7416666,1.1437501,1.6583333,1.6125,0.775,1.3333334,2.28125,4.6083336,4.95625,5.008333,3.2812502,4.0499997,3.53125,1.4416666,1.2416667,0.9250001,0.8000001,0.66875005,0.57500005,0.23750001,0.075,0.19166668,0.043750003,0.0,0.0,0.13333334,0.2875,0.24166666,0.2875,0.20833334,0.15,0.081250004,0.09166667,0.35625,0.45833337,0.056250002,0.0,0.29166666,1.625,2.3666668,2.1687498,2.05,1.7125,0.7416667,0.6333333,0.8125,1.6666667,4.5875006,5.5249996,4.1125,3.9666667,4.18125,4.008333,2.9166665,2.03125,2.0916667,2.93125,5.691667,8.475,10.208334,11.691667,14.44375,17.075,20.200003,26.174997,35.625,48.016666,60.3,67.21667,68.575005,64.799995,62.266666,60.337494,55.19167,56.537502,69.13334,70.200005,77.3875,86.524994,81.98125,68.8,57.962498,58.575,62.233334,52.693752,39.041668,44.725002,70.291664,73.05626,56.716667,53.406254,53.783333,67.425,53.5125,28.041662,10.8125,4.1,4.86875,7.891667,14.266668,20.83125,18.541666,6.9437504,8.691668,9.93125,3.2416668,1.40625,1.025,0.9583333,1.1374999,3.9000006,6.9312496,12.175,13.800001,13.25,15.674999,13.825,7.5750003,3.40625,2.6666665,7.58125,14.883333,20.175001,28.518753,33.3,28.45,28.183332,15.63125,3.6333332,1.6249999,2.5500002,2.2333333,2.15,1.4916668,1.25625,1.7583332,1.0,0.5333333,0.40833336,3.1500003,1.4333334,1.00625,2.2500002,1.3874999,0.7916667,2.1000001,2.8500001,2.1000001,3.2624998,2.35,0.23750003,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.16666667,1.9750003,3.1333332,3.50625,5.7833333,6.833333,5.05625,5.758333,8.525001,11.625,15.21875,16.391666,15.4375,8.741667,3.75,1.11875,0.28333336,0.26875,0.44166672,4.09375,13.15,18.491667,21.206251,22.533333,25.181252,33.649998,33.48125,26.416668,16.737501,7.4833336,6.408334,3.25,1.4583334,0.35625002,2.2250001,0.65625,0.0,0.0,0.0,0.0,0.00625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016666668,0.2,0.28125,0.008333334,0.0,0.0,0.0,0.0,0.0,0.0,0.31666666,0.25,0.083333336,0.05625,0.24166667,0.56875,2.0750003,3.2583334,1.95,1.1,0.38125,0.0,0.0,0.0,0.0,0.0,0.008333334,0.075,0.48333335,2.05,4.758333,8.08125,10.8,11.641666,12.30625,10.983334,12.53125,15.166668,15.975,15.5,14.399999,14.21875,12.908334,10.65,9.408334,8.36875,9.675,11.933333,15.387502,18.908335,19.925,16.425001,12.24375,0.041666668,0.23333335,0.5555556,1.8583335,2.011111,1.775,0.8777778,0.98333335,0.47777775,0.6888889,0.97499996,2.2444444,2.9250002,5.322222,7.1833334,6.422222,4.208333,1.4000001,1.0111111,0.33333337,0.4,0.275,0.011111111,0.09166667,0.10000001,0.25555557,0.24166667,0.033333335,0.0,0.0,0.0,0.0,0.0,0.011111111,0.022222223,0.0,0.0,0.0,0.25555557,0.4666667,0.044444446,0.0,0.21666668,0.25555557,0.06666667,0.12222223,0.14166668,0.07777778,0.044444446,0.09166667,0.21111111,2.5500002,5.1444445,4.2250004,2.788889,1.5333333,1.0666667,0.77777785,0.8000001,1.5333333,2.875,5.322222,8.208334,12.344444,15.033333,18.199999,21.844446,25.9,29.01111,34.44167,44.300003,59.508335,72.355545,75.08889,77.61667,68.81112,68.04167,64.23334,64.35833,76.76666,88.01111,80.84167,87.50001,103.12501,84.83334,58.51667,47.399998,52.84445,55.708332,46.47778,37.7,42.244442,52.233334,42.88889,42.55,30.266666,42.27778,56.858337,30.577782,12.266667,4.9777775,3.8083336,10.1888895,18.555555,35.333336,22.744444,10.908334,8.811111,13.475001,3.0555556,0.6333334,0.16666667,0.5666667,0.29166672,1.1777778,4.008333,8.644445,13.783333,12.022222,9.377778,10.55,11.122222,8.008333,4.322222,6.341667,14.988888,24.58889,32.6,35.244442,36.933334,29.788887,18.841667,6.833333,3.7083333,1.2333335,2.3333333,2.5750003,5.6111107,0.3666667,4.7333336,1.3833334,1.2222223,2.288889,5.008334,2.2000003,1.925,1.1222223,1.3916669,1.8555555,2.6916666,2.2555556,1.0333333,0.05,0.16666667,0.05,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.008333334,0.43333334,0.69166666,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.35555553,1.9166666,3.411111,6.7750006,9.888889,11.877779,9.633333,9.233334,12.575001,20.622223,24.641666,21.588888,16.8,12.388889,9.000001,7.083333,5.1222224,2.8166666,1.1555556,1.6583334,3.5111113,4.211111,6.0750003,9.588888,15.85,25.855555,30.341667,35.922222,38.158333,26.044445,9.4777775,2.15,0.23333332,0.0,0.08888889,1.9833335,0.21111111,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06666667,0.39999998,0.0,0.0,0.19166666,1.3666667,1.2222223,0.13333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06666667,0.975,3.5888891,3.4,0.7416666,0.07777777,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.15000002,0.6666666,1.5333334,3.1555555,5.9833336,9.911112,13.055555,14.775001,15.51111,16.216667,16.933332,17.391666,16.511112,15.800001,14.841666,14.3,15.15,15.933333,15.775,15.688889,16.033333,16.508333,16.544443,14.3,12.977779,12.591666,0.075,0.041666668,0.033333335,0.5187501,1.5666668,2.1937501,1.4333334,0.9625,1.175,2.1166666,2.3375,1.9749999,1.21875,1.9166666,2.2187502,2.483333,1.24375,0.075,0.058333337,0.10000001,0.116666675,0.10625,0.008333334,0.0,0.025000002,0.033333335,0.0375,0.225,0.1375,0.0,0.0,0.0,0.0125,0.008333334,0.050000004,0.20625001,0.40000004,0.16250001,0.0,0.0,0.016666668,0.19166666,6.668751,13.041668,9.3,5.4833336,3.175,1.0916666,1.4166667,2.5937502,2.8083334,1.8812501,3.7916665,4.81875,5.491667,2.7250001,0.35833338,0.33333334,0.45000005,1.0,2.225,4.3416667,8.00625,12.525,17.05,21.750002,26.716667,31.737501,36.841663,39.587505,44.23333,58.018753,70.48334,74.925,81.806244,84.233345,77.2125,76.958336,87.256256,90.975,104.12501,101.043755,93.23334,97.31251,97.09167,73.95625,52.483334,46.275,47.45,53.76667,48.781254,41.44166,37.99375,42.550003,31.3375,24.808334,24.508335,38.56875,29.083334,11.625,4.191667,1.425,2.3250003,5.125,8.343749,5.258333,3.7625,7.0166674,12.1875,4.2,1.2375,0.5,0.5500001,0.1,0.28333333,2.2625003,5.566667,11.9125,13.083333,13.416666,9.94375,10.641666,10.125,8.333333,6.9437504,9.391667,18.650002,29.868748,40.14167,39.45625,28.275,11.531249,5.316667,7.8062496,2.325,1.4583335,1.525,9.058334,15.7625,21.416668,8.13125,2.3916664,1.5833333,2.4562502,3.4416668,1.98125,1.075,3.6687503,4.366667,4.9,2.75,1.0583334,0.0,0.0,0.0,0.0,0.0125,0.016666668,0.0,0.0,0.0,0.0,0.0,0.00625,2.0083334,1.6500001,1.4333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.30833334,1.5750002,3.1750002,5.0937505,8.833334,11.508333,14.175,17.75,21.400002,32.850002,45.5125,42.625,30.35625,23.566666,18.258333,13.75,11.941668,5.75,2.5833335,1.7249999,2.2333336,2.65,3.5875,6.75,17.987501,22.125,19.33125,27.175,59.39375,57.43333,33.25,11.731251,1.5166669,0.0625,0.0,0.80625004,0.8083333,0.24166667,0.80625,0.975,0.57500005,0.20000002,0.0125,0.0,0.36666667,2.3687499,1.4833335,0.45,1.3333334,0.68125,0.0,0.0125,0.4916667,0.8416667,0.26875,0.008333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.056250002,0.2916667,0.2125,0.31666666,0.90625,1.6500002,0.75,0.48125002,0.33333334,0.0375,0.0,0.0,0.016666668,0.050000004,0.16875002,0.30833334,1.0812501,3.0833333,5.19375,6.3416667,8.69375,12.950001,19.3,24.84375,24.516668,19.862501,16.083334,11.062499,8.7,7.3666673,5.70625,6.4083343,9.05,12.558333,14.368751,12.675,9.449999,7.2937503,5.7250004,4.3,3.4583333,5.825,0.35,0.29999998,0.5222223,1.2916666,1.3333336,2.0,2.6222224,2.8833332,4.4888887,6.4,11.125001,9.755557,6.2333336,2.3777778,4.408334,1.9111112,0.9333334,0.9222222,0.6444444,0.55833334,0.36666667,0.14166668,0.055555556,0.0,0.0,0.0,0.0,0.0,0.008333334,0.0,0.016666668,0.0,0.13333334,0.5555556,0.85555553,0.6666667,0.47777778,1.0083334,0.8333334,0.225,0.1777778,1.5555557,4.5249996,6.2222223,9.633333,17.11111,18.408333,15.577778,11.177778,7.4916673,6.7666664,2.55,2.4333334,2.766667,3.3333333,2.516667,0.7777778,0.48888892,0.6500001,1.1444446,2.1833336,3.733333,7.925,13.0222225,18.388887,24.925001,30.666662,40.641666,44.922222,47.866665,51.46667,58.808334,66.38889,72.68889,75.67501,81.78888,80.983345,74.35555,78.425,89.32223,96.288895,100.98333,101.55555,109.91667,115.0,104.625,67.744446,51.43333,42.09167,49.422222,57.016666,42.81111,32.383335,31.944447,31.241663,20.022223,24.9,33.775,18.28889,9.366668,4.8666673,1.3833333,1.1333336,2.7222223,7.4083333,11.144444,7.85,1.4111111,1.8666666,2.4333334,1.7333333,0.9777778,0.6888889,0.16666667,0.21111111,3.9333334,7.833333,10.825001,12.466667,14.588888,17.683334,11.3,9.041667,9.088889,8.483334,7.1222224,12.955557,22.333334,28.97778,30.041666,25.611113,11.208333,2.6555557,10.208334,13.055556,7.166667,1.4833333,6.9777775,21.45,20.633335,14.35,16.4,1.7888889,0.5,1.0666667,1.5666667,2.1555555,5.6333337,7.4000006,5.766667,3.4111109,1.5222223,0.0,0.0,0.0,0.022222223,0.8166667,1.0555555,0.0,0.0,0.0,0.0,0.0,0.0,0.055555556,4.4583335,1.388889,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.3416667,0.8555556,1.9916668,6.2555556,7.911112,8.066668,12.644445,23.091665,31.7,25.55,25.033335,20.433332,19.2,16.566668,9.691667,4.2444444,2.075,0.82222223,0.5166667,1.4666667,3.0333333,6.275,10.88889,23.824999,42.67778,39.858337,33.86667,38.841663,28.911112,15.455556,4.7000003,0.28888887,0.0,0.0,0.26666665,0.7222222,0.15555556,0.6583333,0.7555555,0.53333336,0.1,0.5416666,1.5222223,4.4888887,11.35,6.466667,1.9083334,1.1777779,0.37500003,0.0,0.033333335,0.07777778,0.24444446,0.025,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.22500001,1.1777779,1.45,0.48888886,0.4666667,0.8555556,0.011111111,0.28333336,0.1888889,0.0,0.0,0.008333334,0.13333334,0.37777779,0.8000001,1.7111112,3.3333335,6.588889,9.55,10.900001,12.466667,16.11111,22.3,35.350002,45.27778,38.941666,31.500002,24.325,17.1,11.366668,6.1166673,4.455556,3.8750005,3.9111109,5.366667,5.8666663,3.8,2.65,2.5222223,2.6000001,2.6555557,4.258333,0.06666667,0.25555554,0.34444442,1.1583333,1.5555557,1.475,1.3555555,2.1833336,3.9222224,5.644445,9.708333,10.422222,7.5916667,2.1777775,6.3,5.388889,1.1333334,0.54444444,0.4555556,0.4,0.15555556,0.016666668,0.0,0.0,0.0,0.0,0.0,0.0,0.033333335,0.7333333,0.55,0.3888889,0.20000002,0.10000001,0.25555557,0.9083333,0.35555556,0.42499998,1.488889,0.93333334,0.88888884,1.1777778,3.141667,6.2777777,12.516668,20.48889,26.541668,28.522224,26.577778,21.900002,18.844444,11.916666,5.7222223,2.6916668,2.4333334,3.475,5.6555552,5.211111,3.2250001,2.2777777,2.9083333,4.377778,7.1249995,12.733334,19.344444,29.575,40.555553,58.149994,61.666664,63.0,66.37778,74.78333,74.922226,72.87778,73.26666,76.899994,78.575,74.022224,70.166664,73.62222,86.700005,97.049995,104.27778,111.69167,119.08889,118.924995,88.55556,71.922226,61.750004,55.27778,63.508335,59.166668,44.166668,39.233337,37.541664,31.9,30.522224,33.608334,28.1,13.508334,5.1000004,1.8166667,0.8,1.2777779,2.275,4.1555557,3.875,0.65555555,0.3166667,1.6333333,1.8166665,1.8333334,1.4,1.0166667,0.8333334,3.3083334,9.88889,14.033335,12.411111,11.622223,16.983334,16.677778,13.058333,12.0,10.449999,8.922222,9.322222,14.616666,21.544445,24.558334,24.2,9.416667,4.033334,5.3333335,20.38889,23.166668,9.225,7.2000003,19.116669,18.2,11.366668,15.600001,1.4666667,0.083333336,0.6,0.7166667,2.277778,5.2416663,6.1555552,4.516667,2.211111,0.5,0.0,0.0,0.083333336,0.36666667,8.908333,5.2777777,0.33333334,0.0,0.0,0.0,0.0,0.0,0.0,0.875,0.6666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.2,0.8,2.341667,5.3444448,7.6777782,6.275,5.7444444,8.633334,12.433332,10.441667,8.400001,7.9416666,13.922224,15.577778,11.666667,5.1777782,3.8500001,0.95555556,0.0,0.044444446,0.8444444,3.85,9.133334,25.608334,56.733337,51.616665,35.155556,24.908333,6.6444445,1.3555558,0.35000002,0.0,0.0,0.0,0.0,0.22222222,0.5222222,0.48333335,1.2444445,1.7249999,2.1111112,2.9,4.9555554,6.788889,9.225,8.255556,4.825,2.0333335,0.31666666,0.06666667,0.116666675,0.0,0.0,0.23333335,0.5222222,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.19166668,1.2111111,1.225,0.06666667,0.4166667,0.21111113,0.0,0.0,0.0,0.0,0.0,0.0,0.06666667,0.41111112,2.016667,4.5,8.5,9.433333,10.975,13.611111,17.649998,26.344444,37.08889,52.016666,60.77778,59.733334,53.366665,41.83333,34.57778,27.01111,14.2,6.377778,3.9333334,2.066667,1.3166667,1.2333333,1.2777778,1.5833334,2.0555556,3.775,7.944444,10.483334,0.0,0.0,0.075,0.01875,0.19166666,0.7625,0.8416667,1.1,2.6166666,2.591667,2.2,1.3750001,1.09375,0.6333333,1.9999999,2.425,0.40625003,0.15833333,0.108333334,0.0,0.025000002,0.00625,0.0,0.0,0.0,0.0,0.0,0.0,0.025,2.3666668,3.3125,2.7833335,2.1375003,1.3000001,0.87500006,1.175,1.6500001,1.1,1.0416667,1.53125,2.3416667,2.4333334,1.73125,2.5833335,3.325,5.741667,10.19375,15.241667,19.241667,23.875,24.3,23.556252,17.316668,11.975,5.425,4.9312496,7.683334,9.325,7.18125,4.375,9.175,17.366667,23.6375,38.76667,50.291668,66.83125,91.125,92.29375,82.18334,84.68125,81.41667,77.15626,75.791664,74.975006,74.9875,72.75835,70.737495,66.84167,63.112507,61.09167,61.525,61.55,60.466667,59.999996,58.325,69.91875,72.75001,70.26667,66.675,57.56667,51.818752,52.408333,48.575,43.383335,36.4125,33.75,32.958336,36.025005,36.658333,23.812502,18.8,11.293751,3.9250002,1.5083333,0.48125005,2.0666668,2.6999998,0.75000006,0.375,1.5583334,3.16875,4.016667,3.5333333,2.29375,2.5083334,2.99375,8.066667,13.18125,15.141668,13.783333,11.44375,11.625,12.387501,11.116667,11.699999,12.966667,11.950001,11.162499,11.433333,11.5,16.841667,14.481249,9.158332,5.26875,12.683334,29.841667,28.093752,13.883333,14.5625,15.75,9.6,8.916666,0.45000005,0.0125,0.09166667,0.67499995,0.8333334,2.0375,3.525,4.2875,3.0916665,0.35,0.05,0.075,0.375,1.4,26.41875,22.325,4.5249996,0.50624996,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.35625002,0.70000005,1.425,3.483333,5.0666666,5.36875,3.7750003,3.59375,3.766667,3.575,3.7083335,3.7375,9.083334,15.183332,13.7125,7.191667,4.05,1.725,1.4312501,1.0500001,0.5833334,0.55625004,1.9583333,10.9,19.375,24.906248,19.075,18.906248,6.5166664,1.4416666,0.33125,0.0,0.0625,0.15,0.112500004,0.083333336,0.14166668,0.17500001,0.27500004,0.51875,0.8166667,1.1125,2.1,3.1833334,4.5062504,4.4166665,3.3000002,1.6,0.35000002,0.058333337,0.05625,0.025,0.09166667,0.64375,2.3083334,2.125,0.425,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.008333334,0.275,0.025,0.0,0.0,0.0,0.0,0.0,0.0,0.033333335,0.33333334,1.5562501,3.8333333,6.1062503,8.858334,11.1625,14.341667,18.387499,24.183332,31.683334,37.71875,42.541664,45.2,43.891666,45.218746,46.316666,43.40834,32.325,22.275,16.868752,11.816668,6.4062505,3.5333335,3.016667,3.6312501,6.316667,10.075001,13.766667,17.0625,0.0,0.0,0.0,0.008333334,0.05555556,0.13333334,0.21111111,0.22500001,2.1444445,2.3444445,2.4583333,1.3111111,1.5083333,1.8222222,2.8833332,2.5555556,1.9666667,1.3444445,0.8222223,0.108333334,0.0,0.0,0.0,0.0,0.0,0.0,0.008333334,0.26666668,0.30833337,1.3111111,4.558334,5.644445,5.6,4.6111116,3.4555557,2.5416667,2.4555557,2.6333332,2.1222222,0.77500004,0.6666666,1.4444445,2.425,2.0555556,1.9416667,0.46666667,0.5583333,1.4555557,1.9,2.575,4.4888887,9.950001,13.444445,13.666668,13.211111,12.633333,11.066667,14.144445,12.991667,13.422222,20.966665,57.06667,91.46666,124.64445,141.13333,144.44167,154.75555,165.93333,158.82224,132.18333,98.922226,71.90834,66.477776,64.18889,63.791668,58.944447,54.51667,50.255554,49.391666,50.000004,52.822224,57.8,57.011112,54.56667,47.8,41.70833,33.71111,30.07778,31.4,30.877777,30.991665,35.966667,34.55834,38.711113,39.333332,37.68889,34.555557,36.425003,29.933334,20.966667,13.222221,7.25,3.188889,0.3333333,0.06666667,0.26666668,0.9166666,0.78888893,1.175,1.3111112,1.5833333,2.9222224,2.511111,3.5749998,3.1555557,3.716666,5.2999997,6.333333,9.122222,10.333334,8.108334,7.7888894,8.75,5.9777784,8.075,12.733333,17.933332,16.808334,13.633333,11.308333,11.211111,14.175001,14.066668,8.883333,6.488889,18.58889,29.125002,26.744446,16.291668,8.588889,6.4916673,1.4777778,0.0,0.008333334,0.011111111,0.15,1.3777778,2.8000002,4.166667,3.225,2.2333333,0.9666666,0.5,1.3666668,2.15,2.6777778,32.233334,39.73333,18.344444,4.7333336,0.08888889,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.16666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.26666665,0.8333334,1.2666667,1.8222222,2.3333333,2.4222221,0.9250001,0.18888889,0.33333334,0.9833334,2.9555557,3.0166667,2.688889,2.8833334,3.3,1.8444445,1.2916666,1.3444444,3.5916667,8.911112,9.583334,9.355556,4.6666665,8.755555,3.4666667,0.375,0.0,0.008333334,0.044444446,0.033333335,0.033333335,0.1,0.2,0.21111111,0.55833334,0.61111116,0.2916667,0.37777776,0.4666667,0.8000001,0.92222226,0.80833334,0.5555556,0.050000004,0.022222223,0.15,0.6,1.4555557,2.4583335,1.7444446,4.008333,0.7444445,0.64166665,1.5222223,1.5999999,0.62499994,0.27777776,0.025,0.06666667,0.3416667,0.49999997,0.06666667,0.0,0.0,0.0,0.0,0.0,0.0,0.008333334,0.11111111,0.35555556,0.9250001,2.1333334,4.3583336,9.377778,14.550001,17.188889,17.016666,20.688889,25.822222,20.925001,19.966667,20.775,22.955557,24.183334,26.122225,28.155558,25.258333,24.566664,25.71667,23.5,18.0,13.122223,8.777778,9.691667,14.388889,17.116669,18.711113,22.475002,0.0,0.05,0.20833331,0.5375001,0.3083333,0.53125,0.5583334,0.80625004,2.7166667,3.1833332,1.925,1.3416667,0.825,0.65833336,0.925,0.7833333,0.525,0.36666664,0.19999999,0.0,0.23333333,0.53749996,0.40833336,0.325,0.45833334,0.058333334,0.00625,0.5166667,1.225,1.1666667,2.5625002,6.2166667,9.800001,9.891667,8.566667,6.89375,5.533334,4.5312505,3.4916666,3.21875,1.4416667,1.6583333,1.8375002,2.1916666,2.05625,1.1583334,0.91875005,0.6333334,0.45833337,0.5,0.38333333,0.60625005,1.2833334,3.4375,4.8250003,5.6375,6.8500004,9.233334,14.756249,16.466667,19.556252,41.6,90.625,156.725,148.43333,126.08751,129.90001,154.4,148.94168,126.562515,90.84166,72.21875,70.4,65.99167,58.149998,48.583336,46.90625,45.5,45.53125,46.983334,52.783333,61.975002,65.89168,65.44375,58.2,47.5,32.25,23.491667,21.987501,21.083334,23.33125,27.525,29.3375,34.033337,36.525,35.983334,29.108332,19.712502,12.391668,10.20625,7.5166664,5.1500006,2.2749999,0.3416667,0.20625003,0.9916667,1.7187499,1.8500001,2.2687502,2.3083334,2.7937498,4.408334,4.2333336,4.925,5.8,3.6937497,3.016667,3.35625,4.225,6.708333,5.5875006,5.55,10.1625,9.533335,8.7375,10.683334,14.833334,17.106253,17.616667,15.943749,13.491668,13.418751,15.075001,10.518751,7.450001,15.2,27.8125,23.225002,15.412501,7.5000005,4.09375,0.4416667,0.0,0.0125,0.008333334,0.0,0.083333336,0.050000004,0.041666668,0.125,0.9,4.4083333,3.5812502,4.383333,5.7,7.5916667,16.525002,20.5,28.275,10.168749,0.48333335,0.0,0.025000002,0.0125,0.0,0.0,0.0,0.0,0.65625,0.22500001,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03125,0.27500004,0.7062501,2.2583332,2.375,0.6583334,1.425,1.675,0.725,0.5125,0.55,2.3375,5.016667,5.5916667,3.2312503,2.7250001,1.70625,2.3583333,4.5187497,3.3249998,0.84375,0.65,2.5500002,0.6875,0.0,0.01875,0.008333334,0.0,0.016666668,0.17500001,0.37500006,0.40833336,1.0625,1.9416667,1.3499999,0.26666668,0.32500002,1.0375001,1.375,1.5375001,1.5333333,1.6125,1.425,1.1875001,1.6916666,2.6166666,4.975,5.4166665,3.3125,2.2833333,4.3375,9.1,6.833333,4.33125,4.366667,4.425,2.8000002,2.35,2.2083335,0.112500004,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.125,0.73333335,2.1375003,5.4083333,10.375,13.75,12.51875,11.900001,12.283335,12.793751,15.325,19.256248,23.491667,24.34375,25.391668,24.483334,20.9125,20.883333,24.050003,28.96667,32.46875,31.866669,26.90833,22.525,17.908333,16.7125,18.199999,19.837502,0.0,0.033333335,0.23333332,0.29999998,0.43333328,1.3916668,0.73333335,0.625,1.488889,2.5222225,0.70000005,0.45555556,0.3166667,0.20000002,0.008333334,0.0,0.0,0.0,0.0,0.0,0.08888889,0.36666667,0.54444444,1.6083333,1.9000001,1.488889,0.23333335,0.12222223,0.5916667,1.1555554,2.425,2.7333336,8.025,14.544444,15.422223,15.041666,14.066667,10.816668,8.1888895,6.1249995,4.177778,2.777778,1.8916667,2.4,1.7500001,0.84444445,1.1416669,2.7555556,2.8555558,1.7083333,0.36666667,0.25833336,0.20000002,0.4,0.6777778,1.6,3.377778,5.8888884,10.116667,13.444445,22.725002,34.91111,57.88333,99.100006,117.14444,116.46666,114.67778,127.72502,106.466675,99.61667,83.422226,84.041664,75.01111,71.44444,69.43334,71.5,74.89167,80.06667,80.05,81.68889,75.94444,66.31667,63.35556,68.575,69.58889,60.60833,45.46667,35.4,27.633335,21.244446,19.091667,20.166666,21.941668,23.344444,27.391665,32.633335,24.044445,13.241668,9.944445,14.825001,9.833334,3.95,1.1444445,0.022222223,0.0,0.0,0.050000004,0.08888889,0.7666667,2.9333334,3.7250001,4.133333,3.7444446,2.9250002,3.6888885,5.933334,2.9222224,3.1666665,4.7777777,4.7888894,3.8583333,4.3888893,8.441667,9.955555,7.75,9.222221,9.055555,10.641666,13.555557,16.591667,15.900001,14.849999,13.8111105,11.941667,6.911111,8.322223,15.6,22.255554,11.374999,6.9333334,3.691667,0.90000004,0.06666667,0.016666668,0.15555556,0.18333334,0.022222223,0.025,0.0,0.0,0.3111111,11.933334,8.300001,6.5444436,6.0583334,9.5222225,12.716666,9.0222225,7.311111,3.5333338,0.16666669,0.0,1.7111111,0.7583333,0.022222223,0.0,0.0,0.0,0.09166667,0.011111111,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011111111,0.23333333,0.26666668,0.18888888,0.083333336,0.0,0.0,0.0,0.25,2.7444446,5.391667,4.0666666,4.7222223,4.625,2.577778,1.1000001,0.2777778,1.6666667,5.1222224,7.1444445,8.183333,9.933333,7.408333,0.82222223,1.075,1.5444446,0.30833334,0.0,0.07777778,0.18333334,0.4,0.4166667,0.099999994,0.0,0.033333335,0.033333335,0.116666675,0.56666666,1.2083334,1.9888889,3.3833334,1.9000001,1.1111112,1.6750001,2.477778,2.5583336,3.0333333,3.3333335,3.5777779,3.5666668,3.7555554,4.577778,7.833333,6.7333336,4.225,3.566667,7.6500006,15.266666,10.511111,4.525,6.7777777,4.908334,2.4444447,1.0916667,0.48888886,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.45555556,1.1916667,3.0333333,5.1583333,7.5444446,6.883333,4.366667,4.0111113,7.133333,13.388889,21.624998,29.08889,33.624996,35.344444,33.844444,30.516666,29.8,29.858334,32.288895,36.100002,40.711113,36.0,32.383335,23.533333,20.149998,22.4,23.008331,0.51875,1.025,0.375,0.16250001,0.30833334,0.45,0.19166669,0.68125,1.675,2.8583333,0.24375,0.058333337,1.2125001,0.55833334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025,0.8416667,4.05,6.175,3.6583335,2.0125,1.2083333,1.4812499,3.3416667,3.0625,4.1583333,5.25,9.341667,13.733333,15.06875,18.808332,23.212502,26.308332,24.606255,14.549999,8.325001,3.19375,1.8166667,2.3999999,1.9833333,1.69375,1.8416667,1.85,0.6499999,0.05,0.0375,0.108333334,0.36875004,0.86666673,1.925,3.8,6.4500003,10.90625,16.866667,26.618752,38.916668,52.443756,74.441666,103.95,125.056244,113.325,95.36875,78.65833,71.83126,64.941666,59.4,66.78334,75.63333,92.4625,117.816666,127.39375,109.950005,97.9875,72.14167,59.850002,54.15625,55.491665,62.075005,61.71667,53.374996,45.808334,40.291668,32.46875,22.150002,13.84375,10.958335,10.05,6.5583334,3.78125,3.9,2.6916666,4.0,13.116667,20.3625,10.2,3.96875,1.3499999,0.25,0.0125,0.0,0.112500004,0.4666667,1.39375,1.975,4.25,8.258333,9.550001,6.96875,5.5250006,3.925,2.016667,3.8250003,6.7416673,6.491667,4.53125,3.9333334,3.15625,3.4,2.7312503,2.625,6.166667,10.231251,10.6,12.112501,12.900001,12.975001,14.908333,12.387501,7.6833344,5.316667,5.8062496,14.975,12.30625,4.041667,2.1749997,0.8000001,0.13333334,0.05,0.39999998,0.3125,0.0,0.0,0.0,0.0,0.041666668,4.9000006,5.99375,4.233333,4.7562504,6.1083336,12.36875,11.658334,3.7583334,0.9437501,0.3666667,0.0,2.4166667,2.53125,0.4416667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06666667,0.65625,0.7416667,0.52500004,0.23750001,0.008333334,0.0,0.0,0.025,1.8166667,6.7125,7.925,4.8916664,4.3562503,2.4083335,0.7625,0.15,0.26875,2.8500004,8.475,16.85625,18.358334,13.88125,5.858333,1.1375,0.39999998,0.1875,0.2,0.4166667,0.83125,1.4,0.975,0.0,0.0625,0.51666665,1.3833332,0.44999996,0.675,1.6812501,2.6750002,4.0,4.9249997,4.058333,4.6375003,5.7,5.99375,6.3916664,7.26875,7.8166666,8.43125,9.541667,8.866667,8.66875,10.391666,9.96875,4.3750005,6.63125,13.275,9.516666,3.98125,2.9583335,2.1000001,1.1,0.125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.008333334,0.14375001,0.4166667,1.1062502,2.2,3.4375002,4.3583336,5.18125,4.4666667,4.191666,6.05,10.299999,17.2125,25.924997,33.443752,38.358334,40.1,37.64375,32.116665,24.212498,20.224998,17.90625,20.575,25.541668,26.925003,27.733335,27.175001,26.441666,25.868752,0.55833334,1.2777779,0.9000001,0.95000017,0.8333334,0.45,0.11111112,0.27500004,1.0111111,1.1444443,0.44166666,0.022222223,0.008333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.4499998,5.388889,8.655556,10.425,6.633333,6.9833336,5.2222223,5.0083337,4.0444446,5.9416666,6.988889,11.211111,16.366669,19.644445,24.758337,35.8,39.533337,33.08889,22.077778,9.666667,2.8555558,1.3750002,1.7666669,1.1,0.97777784,1.0777779,0.90833336,1.0333333,1.1666666,0.70000005,0.4666667,1.3444445,2.625,5.0333333,9.033333,15.958334,23.11111,38.308334,58.577778,77.808334,94.76667,110.26667,131.46667,133.06668,112.20833,89.36666,77.03334,56.344444,47.600006,57.766663,73.77778,87.22499,125.566666,140.20834,147.22223,109.25834,71.48889,62.855553,56.991665,49.644444,44.966667,38.455555,34.21667,27.055553,24.822222,19.291666,16.066668,10.341666,5.766667,4.8333335,3.2111113,1.5000002,0.21111111,0.044444446,1.1749998,6.2444444,7.541667,6.4888887,4.5166664,1.9000002,0.93333334,0.29999998,0.022222223,0.075,0.4111111,1.125,2.8444448,6.25,10.411111,11.688889,8.591666,6.6,4.6,3.3111112,4.2333336,6.411111,5.988889,5.175,4.9444447,4.791667,2.6333334,2.2083335,1.3333334,0.82222223,2.8999999,5.466667,4.533334,4.3777776,4.8249993,7.8888893,9.883332,6.4666667,2.7666667,1.4333334,3.6222222,10.175,4.1555557,1.0166668,0.10000001,0.022222223,0.008333334,0.26666668,0.05,0.0,0.0,0.0,0.0,0.0,0.14444444,1.2333332,1.8555555,3.3083332,5.955556,12.033333,23.844444,26.266668,8.058332,0.22222221,0.008333334,0.26666665,3.25,1.0999999,0.20000002,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011111111,0.28333336,0.888889,0.988889,0.625,0.24444446,0.025000002,0.0,0.05,2.3444448,7.416667,9.011111,5.577778,2.6166668,0.7000001,0.10000001,0.0,0.0,0.08888889,2.5111113,5.158334,7.0111113,6.741667,5.922222,2.3333333,0.9777777,0.8666668,1.4222223,1.5555555,2.4166667,1.7777777,0.60833335,0.6111111,0.13333334,1.5777779,2.311111,0.4166667,0.13333334,0.49166667,1.3111111,2.3500001,3.888889,5.7,7.125,9.144444,11.025001,11.566666,11.641666,10.122222,10.341667,10.566668,7.288889,4.625,5.077778,2.8166666,2.5111113,2.4083333,3.5333338,2.4777777,1.7583334,1.3999999,1.0833335,0.6444445,0.075,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.044444446,0.44166666,1.2555556,2.775,4.2444444,5.3583336,5.544444,5.2,3.7444446,2.5111113,5.1083336,9.144444,14.724999,19.01111,22.108335,26.155556,29.500002,31.091667,30.755558,24.741665,21.2,20.366669,22.922222,25.588892,25.991667,25.0,25.0,25.455557,24.958334,0.058333337,0.8777778,0.8777778,1.0416667,0.8333333,0.75,0.2888889,0.30833334,0.20000002,0.044444446,0.0,0.10000001,0.39166668,0.79999995,1.1500001,0.51111114,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.43333334,3.4333332,7.111111,16.408333,18.333334,14.249999,15.822223,17.891666,13.922222,11.475,11.288888,9.544444,9.208334,14.8,19.891666,25.211111,33.416668,35.011112,26.5,14.55,5.6444445,3.1249995,2.3444448,2.1,1.8555557,1.5777779,1.6583333,2.2222223,2.775,2.677778,1.5916667,1.6222224,4.308333,6.533334,9.866666,17.066666,28.82222,43.7,67.344444,93.71667,113.14444,121.46666,134.36667,137.07779,125.674995,102.37778,82.43334,57.7,46.050003,52.644444,64.81112,69.34999,85.85555,101.433334,118.355545,108.35,81.111115,77.58889,70.683334,52.844444,45.26667,32.51111,25.558332,20.022223,18.444447,14.608334,13.488889,9.500001,5.722222,3.983333,2.2333336,0.725,0.055555556,0.0,0.016666668,0.5777778,1.3499999,1.8333333,2.983333,1.8555555,1.2444444,0.43333334,0.011111111,0.125,0.53333336,1.3,2.266667,4.166667,9.333334,15.077777,15.525001,9.755556,6.533333,6.9888887,4.7166667,3.5444446,4.6222224,6.266667,7.866667,8.275,4.377778,1.025,0.7111111,0.23333332,0.20000002,1.8000001,1.45,1.2888889,1.1416667,1.922222,2.7916665,2.9333334,0.90000015,0.43333334,2.1222222,4.591667,6.4333334,1.4583333,0.23333335,0.0,0.0,0.24444446,0.21666667,0.0,0.0,0.0,0.0,0.0,0.0,0.16666667,2.7555556,4.858333,11.566668,21.800001,35.377777,35.255554,26.641666,7.177778,0.40000004,0.08888889,1.6083333,2.0555556,0.52500004,0.022222223,0.0,0.0,0.0,0.0,0.044444446,0.06666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.11111112,0.3111111,0.2166667,0.13333334,0.033333335,0.0,0.0,1.1111112,2.5833335,2.7111115,2.5222223,2.0,1.1111112,0.25,0.0,0.0,0.0,0.35555556,0.8000001,1.1777778,1.3916667,1.888889,1.2083333,0.6333333,1.3166666,1.8666668,1.1666667,1.1916667,0.39999998,0.0,1.2888889,1.6500001,2.4444444,1.211111,0.21666667,0.055555556,0.16666667,0.34444445,0.89166665,2.5,3.0555556,3.9666667,4.7666664,4.825,5.6222224,5.3333335,4.9111114,5.3583336,6.0222225,5.3333335,3.8999999,4.7888894,1.4750001,0.3888889,1.4583333,2.2444446,2.7444444,2.2916667,1.8333333,1.4500002,0.8000001,0.15000002,0.0,0.125,0.31111112,0.12222222,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.008333334,0.05555556,0.083333336,0.3,0.26666665,0.53333336,1.1,2.688889,6.222222,10.933333,13.866667,16.083334,17.566668,19.925001,22.311111,24.488888,29.341663,31.677778,27.708336,24.855556,26.541668,29.499998,30.866669,32.433334,32.76667,33.266666,36.233334,35.433334,0.28125,0.46666667,0.5416667,1.03125,1.2166666,0.91875005,0.7416667,0.2875,0.625,0.38333333,0.0,0.0,0.01875,0.033333335,0.056250002,0.083333336,0.0,0.0,0.0,0.0,0.05,0.25,0.275,0.5375,1.575,4.491667,10.54375,12.008333,9.700001,8.508333,9.10625,8.616668,7.51875,6.700001,5.3166666,3.0687501,3.1666665,7.9625006,13.166668,16.59375,22.433332,27.658335,19.35,9.466667,4.56875,3.65,2.6562498,2.4499998,2.2250001,2.35625,2.8416667,3.6000001,5.5249996,5.35625,5.775,7.39375,11.608334,12.291666,16.90625,23.6,33.74375,50.2,73.23125,90.341675,101.075,107.19999,108.35834,98.46875,82.16667,66.4375,53.733334,44.975,49.166668,56.86667,56.456257,59.575,61.981255,70.38334,68.4,63.80833,51.116665,43.0875,35.86667,33.8,32.058334,25.0125,24.166666,21.825,21.131252,20.400002,21.2125,19.475,17.343752,11.183334,5.0125,1.5833334,0.25000003,0.0,0.0,0.0,0.050000004,0.18750001,0.19166668,0.13333334,0.056250002,0.0,0.0,0.0,0.18124998,0.5333333,1.55625,4.725,9.758334,15.806251,19.0,19.66875,18.383333,12.206249,7.975,6.1083336,5.7062507,7.25,9.55,8.575001,3.7437499,1.6166666,1.2416667,0.16250001,0.975,1.575,1.075,1.69375,3.2416668,1.7625,1.2333335,1.6166666,0.76875,1.2583334,3.30625,4.6,2.9125001,0.44166672,0.06666667,0.0,0.16666667,0.22500001,0.0,0.0,0.0,0.0,0.2916667,0.33333334,0.0,0.55833334,5.45,21.183334,43.6125,65.916664,64.11667,32.475,11.175,0.6,0.0,0.13125001,1.4166667,0.49375004,0.025,0.0,0.0,0.0,0.081250004,0.16666669,0.087500006,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.28333333,1.6000001,1.9000001,3.6,6.89375,6.041667,3.61875,1.4333333,0.76875,0.3916667,0.17500001,0.13125001,0.28333333,0.37500003,0.20000002,0.10000001,0.06666667,0.7875001,2.8583336,3.9,1.6875,0.325,0.89375,1.4333333,3.5937502,3.8666668,0.775,0.25,0.083333336,0.1,0.083333336,0.0625,0.23333335,0.26666668,0.23125,0.31666666,0.17500001,0.23333335,0.65625,2.0166667,3.725,6.108333,8.416666,11.512501,11.3,3.7999997,0.30833334,0.46875,0.0,0.15,0.13125,0.108333334,0.087500006,0.058333337,0.01875,0.041666668,0.45625004,0.43333337,0.2,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.033333335,0.34375,1.0083333,1.95,2.8083336,4.1125,7.55,11.300001,14.031251,15.233334,15.30625,15.674999,17.1375,18.816666,20.7,21.56875,22.466667,24.2,25.408333,25.743752,24.35,24.308334,26.06875,26.641668,27.8,32.600002,31.900002,0.4166667,0.44444445,0.011111111,1.1666666,1.4666667,0.8833333,0.7,0.65,1.0444444,0.022222223,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.008333334,0.044444446,0.0,0.022222223,0.0,0.055555556,3.288889,13.183335,21.38889,11.491667,9.333333,7.275,4.4,2.4583333,1.2777778,1.4444445,1.4000001,2.0111113,3.8583336,7.0222225,14.525,16.622225,16.48889,17.758333,11.266666,6.0583334,3.7,2.3166668,1.6333334,1.488889,1.325,2.477778,5.2333326,7.5000005,9.083334,10.411112,14.316666,16.088888,19.633333,21.108334,24.833336,30.116665,36.500004,51.491673,67.63334,73.08889,70.450005,64.32223,56.166668,49.311108,44.750004,37.7,33.091667,31.944445,34.600002,35.63333,37.999996,37.9,41.244446,37.416664,29.0,20.377777,17.675001,23.233334,23.083336,19.888891,20.008333,20.511112,20.67778,24.775,23.688889,20.316666,19.533335,16.491667,10.111111,5.0499997,1.6444445,0.42222226,0.70000005,2.2222223,1.7416666,0.79999995,1.8583333,3.8777778,2.0444446,0.78333336,0.3666667,0.475,0.3888889,0.14166667,0.08888889,0.44166672,2.5,4.955556,10.616667,21.47778,34.308334,43.644444,33.075,22.811111,15.766666,8.083334,6.622222,8.275002,10.3,9.633333,3.5444443,2.6555555,2.1833334,3.6000001,4.375,3.8222222,3.691667,9.900001,6.5916667,2.4777777,2.0444443,1.9000001,1.488889,5.1500006,9.000001,7.633333,0.97777784,0.1777778,0.016666668,0.0,0.10000001,0.0,0.0,0.0,0.0,0.28888887,0.25555557,0.0,0.0,1.4833332,15.966668,43.975002,73.08889,82.57778,49.258335,20.777779,7.316667,0.0,1.325,4.8,0.5666667,0.022222223,0.0,0.0,0.0,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.6166666,1.9555554,3.3555555,7.291667,7.1555557,4.7833333,1.5444446,0.39166668,0.14444445,0.0,0.0,0.011111111,0.033333335,0.022222223,0.0,0.022222223,0.058333337,1.6444445,3.011111,2.55,1.9222221,3.516667,2.4444447,2.641667,1.5666666,0.22222222,0.0,0.0,0.016666668,0.044444446,0.016666668,0.0,0.0,0.0,0.0,0.0,0.0,0.05,0.15555556,0.25833336,0.37777779,0.42222223,0.82500005,0.6666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.033333335,0.5083334,0.22222224,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.16666669,0.5111111,1.2166667,2.0777779,3.225,5.022222,5.9,6.65,6.977778,7.008333,7.4777784,10.558334,15.266667,16.577778,17.725,17.122223,18.291668,18.477777,16.183334,14.577779,15.277778,16.541668,19.077778,25.316666,30.122223,30.85,0.0,0.0,0.0,0.24374999,0.6166667,0.48124996,0.7,0.70000005,0.275,0.033333335,0.0,0.0,0.0,0.39166665,1.2625,0.7916667,0.0,0.675,0.075,0.16250002,1.1083332,1.5187501,1.6583333,3.775,3.7916667,3.4333332,4.8250003,2.8833334,3.1499999,6.4333334,5.3187504,5.5,4.475,5.1749997,4.5083337,3.71875,2.4333332,0.8125,1.1666666,2.275,6.7666664,7.0,5.5875,3.0833335,1.5187501,0.5416667,0.21875,0.35833335,0.49166667,0.61875,1.3333333,3.8687499,7.1750007,12.2875,13.283333,13.6,14.291669,16.133335,22.55625,27.616669,32.19375,34.899998,43.125,53.69167,52.550007,47.156254,42.641666,37.15625,35.93334,35.84375,35.175,34.58125,35.858334,38.125,37.774998,33.783333,29.65,26.225002,23.225002,19.341665,16.308334,13.762501,15.208334,23.4875,21.758335,20.6,22.291668,24.599998,22.66875,20.408335,15.925,10.599999,8.275001,5.616667,4.16875,3.5833335,3.4916668,3.9000003,3.783333,2.6187499,1.3,1.41875,2.4166667,2.4583337,2.1875,1.6500001,1.4999999,1.075,0.35625002,0.05,0.2375,0.25000003,1.075,4.425,10.858334,14.875,15.941666,13.6625,12.625001,9.175,4.4375,2.6750002,3.3125,3.9500005,6.043751,5.9083333,5.15,7.8,11.191667,13.2375,13.366667,12.21875,11.425,12.012501,9.266666,5.8333335,5.9437504,8.333333,10.987498,25.86667,24.4,12.300001,3.0500002,0.375,0.0,0.0,0.033333335,0.025,0.0,0.0,0.016666668,0.0,0.3625,0.48333335,0.38125,5.233333,20.387503,38.899998,43.341667,39.9375,31.025002,22.618752,0.033333335,0.225,5.2416663,0.71875006,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.4125,1.7416668,2.125,4.7,5.116667,4.71875,3.6416667,0.25,0.0,0.0,0.0,0.0,0.0,0.0,0.03125,0.425,0.71250004,0.7166667,1.8583335,1.7749999,1.6416667,2.9250004,4.166667,5.96875,2.6333334,1.6500001,0.28125,0.0,0.0,0.0,0.09375,0.083333336,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025,0.06666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0125,0.15833336,0.21249999,0.008333334,0.0,0.0,0.0,0.0,0.0,0.0,0.025,0.19166666,0.025,0.0,0.0,0.0,0.0125,0.10000001,1.2062501,4.0083337,7.0416665,9.05,8.333334,7.3125,7.391667,6.84375,8.883333,9.166667,10.293751,12.241667,16.087502,16.983334,13.4875,13.433333,14.958334,21.84375,30.25,39.862503,40.675003,41.6375,0.008333334,0.033333335,0.22222224,1.125,0.08888889,0.0,0.37777776,0.70833325,0.48888886,0.73333335,0.041666668,0.0,0.075,4.0,11.5,11.677777,4.7833333,1.8,1.9333335,1.0333333,0.6222222,2.0249999,4.5333333,8.3,11.344445,11.522222,9.041666,3.6555557,1.1333333,1.2111112,2.9333334,5.2222223,5.8500004,6.044444,7.188889,6.0166674,5.611111,2.7166665,1.7333336,0.8666667,0.7555556,0.78888893,1.0666667,1.8555555,1.675,1.988889,2.2333333,1.8444445,0.5111111,0.14166668,0.53333336,2.35,4.877778,8.125001,9.877779,11.674999,12.78889,13.177778,13.775002,15.9,20.183334,24.3,42.65,68.52222,52.888893,33.008335,28.233335,30.891666,37.42222,43.725002,48.699997,47.44167,50.21111,48.511112,44.658337,37.68889,28.366667,20.333334,16.741667,12.955556,11.233334,10.6,9.755555,15.474998,24.866667,27.216667,25.8,22.666668,17.241665,14.744445,11.191666,6.0111113,3.6583333,3.6111112,3.0,3.088889,3.8444445,5.125,5.5333333,4.358333,3.1111112,2.1749997,1.6111112,1.6666669,1.3083334,1.2333332,1.9416667,2.222222,1.625,1.2555556,1.2583334,2.2111108,1.9666667,1.6916667,1.9444444,3.3333335,7.7222223,10.091667,10.966667,9.3555565,5.008333,1.3777778,0.9583335,0.8333333,1.1999998,2.0555556,1.7666668,3.5916667,10.866667,17.641666,18.644444,17.666666,14.144444,10.633333,9.766666,8.655556,10.108334,12.988889,12.516667,14.144445,12.416668,7.9777784,5.1444445,0.8166667,0.022222223,0.11666667,0.45555553,0.7916666,1.3444445,1.5750002,0.5222222,0.07777778,0.9000001,1.4000001,1.3750001,0.6333334,3.0166664,10.411112,22.444445,20.458332,10.766667,7.1083336,0.2,0.0,0.26666668,0.24166666,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05,0.92222226,1.2666667,3.6250005,4.677778,8.283334,11.28889,1.05,0.033333335,0.0,0.0,0.0,0.0,0.0,0.22500001,1.9000001,3.1916666,2.1333334,2.1888888,3.3083332,2.5666668,2.125,2.9555557,6.025,3.811111,3.0777776,1.5166668,0.0,0.033333335,0.06666667,0.28333336,1.6555557,1.7222223,1.1583334,0.45555553,0.075,0.12222223,0.16666667,0.21111111,0.19166666,0.35555556,0.44444448,0.34166667,0.29999998,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.4416667,2.3666666,2.788889,6.883333,8.755555,8.0,5.8444448,3.8833337,5.277777,7.5777783,14.466667,14.433333,8.591667,13.688889,16.216665,20.755554,22.266666,29.05,35.17778,43.01667,54.122223,54.166668,0.3375,0.48333335,0.0,0.2625,0.033333335,0.112500004,0.25833333,0.73125,1.15,2.175,0.2625,0.0,0.28750002,3.9250002,9.900001,12.641667,14.4125,15.508334,7.441666,1.9625,0.7416668,0.8125,6.133333,10.31875,17.625004,19.433334,19.65,14.6,10.21875,7.9750004,7.1125,6.958333,9.7875,11.458334,10.433333,5.9625006,2.6750002,1.3812499,1.6666665,3.11875,3.9583335,3.9833333,3.2250001,2.3666668,1.9,0.32500002,1.2812501,2.075,2.9500003,3.9562502,2.2083333,3.31875,2.8666666,2.1750002,4.5083337,5.0937505,7.758333,9.541667,15.18125,17.866667,24.7875,33.39167,41.274998,46.8,44.725002,40.187504,36.466667,37.30625,43.7,46.187496,49.741665,57.05,55.391663,53.350002,52.912506,42.60833,27.800001,16.650002,12.55625,11.858334,10.541668,9.231251,9.616667,13.793751,18.183334,19.99375,19.241665,15.124999,12.331249,9.025001,6.3,3.766667,1.8687499,1.9666667,2.66875,3.4916668,4.8750005,8.01875,7.6583333,6.0812497,4.2583337,2.7875001,1.4916667,1.7999998,0.975,0.28333336,0.4625,0.6583333,1.34375,2.2833333,2.25,2.141667,2.4416666,2.425,1.5,1.40625,3.1083333,7.856251,8.158334,7.8583336,7.3250003,3.491667,0.71875006,0.28333333,0.25625,0.5,0.7749999,1.5562501,4.3916664,10.300001,14.075,20.38125,24.608332,23.150002,14.416668,8.674999,11.981251,16.841667,18.306252,15.775,8.612499,8.566667,5.3083334,2.3999996,1.1,2.3187501,5.4583335,13.26875,23.975,21.5,5.125,2.3166668,1.9687502,2.1833334,3.025,5.5249996,9.562499,14.291665,22.9,22.062502,23.149998,4.3812504,0.125,0.00625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.8833334,2.1333334,2.75,3.425,8.868751,12.558333,2.1375,0.06666667,0.0,0.0,0.0,0.0,0.0,0.0,1.1666667,3.4937503,4.1666665,2.5916667,1.45,1.9583336,1.4437501,0.9,1.0500001,0.7666667,1.4166666,2.0874999,1.0916666,0.7624999,0.35833338,0.25,0.70000005,1.3416666,1.0625,0.6166667,0.40000004,0.4916667,0.71875,0.4416667,0.52500004,1.5500001,2.0833335,1.0125,0.25833333,0.01875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06666667,0.4,0.8333334,1.68125,2.15,4.141667,10.362501,13.875,11.53125,9.266667,10.75625,11.825001,13.358334,17.11875,21.699999,28.45625,28.808334,19.86875,20.166666,24.833336,32.3125,37.8,48.1375,63.14167,58.2375,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.5083333,1.1555555,2.2555559,0.2,0.011111111,0.23333332,3.2333336,9.891666,12.8555565,13.174999,9.733334,6.1999993,1.1750002,0.76666665,3.0500002,1.5111113,7.2000003,5.333333,5.222222,3.1999998,2.777778,3.8500001,4.1333337,4.508333,5.2777777,5.5499997,6.788889,7.7111115,8.591666,6.6333337,5.375,4.766667,5.491667,6.4888887,9.033334,11.008332,12.955557,15.508334,18.311111,5.233333,2.0777779,1.5444444,3.0083334,4.6444445,7.466667,7.755556,6.3166666,5.6111116,4.6916666,6.5444446,8.466666,9.966667,12.466666,18.858332,25.733334,31.258337,34.18889,36.72222,38.608334,38.111115,35.2,41.244446,45.241673,42.800003,38.5,35.266666,36.255554,34.325,28.777779,18.875,12.9,8.575001,7.6777782,6.5222225,5.341667,4.966667,4.608333,5.633333,8.291667,9.022222,7.6777773,5.3666663,2.911111,2.1333334,1.1222223,0.525,0.12222223,0.42500004,0.9777779,1.3777778,1.9333333,1.7777778,0.7916667,0.6444445,0.6333333,0.78888893,1.3,0.9916666,0.47777778,0.5083334,0.72222227,2.6916666,4.266667,5.0916667,4.1444445,4.711111,3.7416668,2.622222,1.9999999,5.1444445,12.241667,16.944445,18.91111,17.133335,10.411111,2.8333335,0.57777774,0.33333334,0.6111111,0.5444445,1.2333333,2.0555556,4.783334,6.666667,13.925,18.266666,22.95,22.055557,16.511108,15.075001,25.077778,32.691666,36.08889,28.891666,12.133334,5.3222227,2.5000002,1.2555556,5.9583335,24.555557,51.533337,65.566666,67.933334,59.97778,15.166666,10.75,7.422222,5.025,6.8,7.366667,12.8555565,22.277777,32.091667,57.022224,26.591667,2.4888892,0.041666668,1.6666667,0.9833334,0.9888889,0.6,0.3,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.4,3.9333336,3.4833333,2.9444447,7.65,9.3111105,1.75,0.05555556,0.0,0.0,0.0,0.0,0.0,0.108333334,0.22222224,0.275,1.0333334,1.8222224,1.2833334,0.4,0.55833334,0.53333336,0.3916667,0.46666664,0.6111111,0.97499996,2.6555557,1.6750002,0.2777778,0.16666669,0.05555556,0.11111112,0.28333333,1.1777778,3.15,5.3555555,5.4750004,3.5333338,3.8583333,6.1000004,4.0222225,1.8249999,0.41111112,0.025,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011111111,0.24166666,0.53333336,0.8916667,0.7555556,0.47777778,1.1416667,2.9333334,5.05,8.933333,10.933332,14.544445,20.97778,30.85,46.833336,57.949997,51.788887,36.725002,30.322226,32.444443,33.225,28.41111,28.508335,34.377777,30.999998,0.0625,0.016666668,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.008333334,0.00625,0.008333334,0.025,0.69166666,5.6562495,11.633333,9.300001,3.125,1.5666666,0.7125,0.64166665,0.025,0.05,0.91875005,1.5,0.95000005,0.35000002,0.17500001,0.18750001,0.24166669,0.15,0.225,0.8,1.25,1.7750001,2.9812498,4.1,4.6312504,6.291666,8.21875,10.041666,13.583334,16.7875,21.158335,30.0125,27.058334,31.393751,25.35,14.508333,7.7000003,6.950001,8.174999,5.6000004,3.38125,2.4750001,2.9125,4.158334,5.8499994,8.0,11.891665,14.9625,17.791666,20.506248,22.333332,25.18333,26.5375,28.825,36.899998,48.41667,52.012505,48.533337,37.625,33.441666,28.350002,20.775,17.425,15.21875,11.783334,7.8375,5.833334,5.0333333,4.2125006,3.3416667,3.01875,2.975,3.16875,3.3583336,2.2333333,1.36875,0.80833334,0.63125,0.30833337,0.15,0.108333334,0.25625002,0.85833335,1.1416667,1.50625,1.2666667,0.36874998,0.016666668,0.0,0.0,0.13333336,0.33749992,0.25833336,0.36875,1.2916667,3.625,4.95,7.0874996,7.4000006,6.8833337,7.2437496,5.941666,4.66875,4.6916676,7.75625,11.25,12.625001,12.675,11.216666,3.875,1.525,1.5375,0.6916667,1.0500001,2.225,3.45,5.1687503,4.883333,5.125,6.5,7.2937493,15.174999,15.958334,12.243751,15.516667,22.75625,24.074999,26.731249,27.891666,13.233334,16.3625,20.125,8.85625,40.558334,87.41875,106.8,117.90625,88.38334,45.716667,24.668749,17.241667,12.900001,4.375,4.05,9.816666,22.800001,29.175,57.425003,62.96875,17.825,3.4125001,4.5166674,5.3125,11.966667,13.083334,1.8312501,0.51666665,0.2125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05,2.15,4.616667,2.1374998,1.2833333,3.96875,3.5166667,1.0374999,0.0,0.0,0.0,0.016666668,0.06875,0.5833333,0.50625,0.47500002,0.38750002,0.31666666,0.33333334,0.5500001,0.32500005,0.06875,0.89166677,2.45,3.7416666,3.666667,1.40625,0.7083333,0.15000002,0.016666668,0.4375,1.6916668,2.95,4.9749994,7.4666667,9.5375,11.208334,13.231251,9.508332,5.21875,1.8750001,0.21666667,0.0125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016666668,0.47499996,1.4166666,2.7562504,3.8750002,3.2250001,2.75,2.141667,2.1,3.3500001,5.1500006,7.4500003,12.975,16.91875,22.291668,25.29375,21.858332,18.73125,17.4,17.066668,19.762499,25.800003,25.893751,25.708334,25.21875,0.06666667,0.044444446,0.06666667,0.06666667,0.055555556,0.06666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.033333335,1.0666667,3.3111112,2.8083334,0.82222223,0.4666667,2.0083334,2.6000001,0.6583333,0.022222223,1.9416668,2.9666667,1.7444446,2.0333333,1.9444444,0.41666666,0.41111112,0.9083334,1.3444445,1.3916667,1.1555556,2.0666666,2.983333,4.7333336,6.9416666,6.2333336,6.5166674,10.044445,12.900001,19.375,25.488888,31.683332,37.28889,44.758327,45.56667,41.54444,25.400002,16.699999,16.458334,5.111111,1.3416667,0.42222223,1.0916667,2.2444444,3.966667,4.6583333,6.5,8.141666,10.422222,13.758335,18.066668,22.1,24.183332,26.277779,31.433334,48.255558,57.141666,53.81111,42.125,34.433334,28.7,24.416666,21.333332,18.041666,15.322222,11.216667,8.1,5.8444448,4.2000003,3.0555556,3.1,2.7111113,3.7166667,2.8333335,2.2,2.05,2.3222222,1.85,1.4666667,0.15833335,0.0,0.0,0.022222223,0.06666667,0.12500001,0.18888889,0.3,0.3222222,0.37500003,0.51111114,0.6,0.7416667,0.6,0.8083334,1.4000001,1.9083333,2.7777777,3.1833334,5.711111,6.1555557,4.5583334,5.955556,6.875,7.4444447,7.8500004,8.344444,8.3,6.1000004,6.244445,6.083333,4.2333336,2.1916668,1.2222223,1.111111,1.6416667,5.211111,7.691667,8.355556,6.6,5.6444445,6.133333,5.744444,9.133333,9.366668,11.3,14.800001,17.51111,15.849999,24.68889,20.31111,22.741667,30.93333,18.575,16.244446,35.083336,55.255558,68.73334,59.65556,50.388885,46.550003,32.0,21.550001,9.944446,10.075,7.9222226,18.100002,34.366665,59.877777,51.125004,21.366665,16.458332,7.9111104,10.466666,10.666667,16.722221,8.508334,3.377778,0.84166664,0.022222223,0.06666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.70000005,1.8999999,0.8833334,0.44444448,1.4333334,0.97777784,0.18333334,0.022222223,0.0,0.0,0.08888889,0.54166675,1.0888889,1.9583335,1.0888889,0.7333334,1.0,0.8333333,0.2916667,0.033333335,0.22500001,1.1555555,2.4,2.9222224,1.9666667,0.46666667,0.16666669,0.033333335,0.0,0.125,0.6777778,1.6888889,2.8833332,4.1444445,5.666667,6.777778,7.5166674,7.8666663,4.0499997,1.3777778,0.18888889,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.008333334,0.23333335,1.0666666,2.3999999,3.6666665,3.9333336,2.4555554,1.2666668,1.1333334,1.4416667,2.677778,5.9444447,6.7166667,6.555556,5.508333,5.133333,5.8333335,7.1888895,8.9,16.583334,28.055555,29.466665,26.588892,19.483334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.25,0.40000004,0.45000005,0.22222224,0.9111111,1.6,1.0777779,3.1416664,8.588888,7.1166673,5.477778,6.433334,2.4333334,2.4222221,1.2083334,0.23333335,1.225,3.2666667,4.641667,4.133333,4.288889,5.1416664,3.6555557,3.825,5.411111,10.7,13.744444,15.144444,20.05,27.366667,31.025,33.644444,44.116665,50.722225,52.02223,42.733337,26.133331,16.625,5.2666664,2.6833332,1.1555556,1.4333334,2.4333334,4.077778,7.4333334,11.1,13.575001,13.855556,17.116667,20.244446,22.144445,21.625,20.52222,22.791666,31.655558,44.76667,44.18889,39.766663,42.522224,44.95556,43.63333,37.266663,30.316668,25.288889,20.316666,15.211111,11.777779,7.766667,5.0111113,3.2333336,2.7444446,3.208333,1.6555556,1.3333334,0.85,0.48888892,0.28333336,0.91111124,0.7333334,0.7444445,0.59166664,0.3888889,0.39999998,0.9166666,1.1,1.1916666,1.3333334,1.4833333,1.9333332,2.3222222,3.1333334,3.5,3.666667,3.8222222,2.5583332,2.233333,2.2,2.6111112,3.9333334,3.7583332,5.7777786,8.3,7.877778,6.5583334,8.777779,11.177778,11.833332,8.3,9.35,14.577778,12.275,6.4,4.866667,5.0666666,8.166667,10.041666,9.933332,8.316667,5.0333333,7.825,8.877777,10.544444,11.441667,10.122222,8.975,7.0333333,10.333333,33.7,47.511112,29.425,19.777779,14.533333,11.655556,19.191668,32.166668,37.950005,40.61111,34.611107,25.533333,34.644444,26.483334,7.633333,4.775,7.533333,15.3,31.866667,50.2,21.808336,11.444444,15.175,17.766666,23.741667,37.31111,16.2,8.558333,3.177778,0.65833336,1.1666667,0.93333334,0.13333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.033333335,0.47777778,1.5083333,0.58888894,0.37500003,0.10000001,0.0,0.0,0.0,0.0,0.011111111,0.32500002,1.1777779,5.6333337,5.4666667,2.4499998,0.8,0.23333333,0.075,0.0,0.23333333,0.9333333,1.1083333,0.9111111,0.48888886,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.24444443,1.0583335,2.1000001,3.2333333,2.9583335,1.6111112,0.6916666,0.3888889,0.14166668,0.12222222,0.42222223,0.5,0.42222223,0.5083333,1.9222223,4.4,6.7666674,11.155556,21.775,32.51111,32.325,23.677778,12.700001,0.0375,0.008333334,0.008333334,0.01875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.15,0.24166667,1.4125,0.49166667,0.09166668,0.80625,4.083334,7.325,6.1583333,5.7125,4.758333,7.2083335,5.95625,1.35,0.28125,0.17500001,1.0437502,2.3666668,3.69375,3.0583334,3.4500003,4.1062503,4.016667,4.36875,5.208333,4.90625,5.8083334,7.7750006,11.50625,22.0,31.956247,36.158337,31.85,34.025,37.65,44.162502,40.333336,20.29375,6.166667,3.7687502,2.725,2.83125,4.95,9.483334,15.26875,20.416668,20.66875,19.816666,20.65625,20.483332,19.358334,18.675001,17.991665,19.55,24.566666,27.175,26.616669,28.84375,31.758333,30.116669,28.893751,23.966667,18.706251,13.775,10.3,7.608333,4.533334,2.85625,1.85,1.61875,1.7250001,2.725,1.9166667,1.2166667,0.74375,0.40833333,0.225,0.20833334,0.15625,0.041666668,0.41250002,0.48333335,0.6916667,0.725,1.2083334,2.1937501,2.6916666,2.9375,4.366667,5.5666666,8.28125,13.025001,15.543749,13.933333,10.118751,6.7083335,5.175,5.3500004,4.3583336,4.15,5.216667,7.2,8.875001,8.5875,11.683333,14.724999,16.900002,15.283332,13.525001,15.691668,17.531252,13.683334,7.6833344,3.55625,5.591667,10.21875,10.066667,7.2687497,4.05,4.325,5.416667,7.8,11.76875,14.658334,16.712502,14.658334,13.681251,19.033333,34.858337,31.29375,22.400002,14.21875,9.55,12.66875,15.35,16.14375,18.608334,25.199999,21.381252,29.583334,21.068748,14.608333,17.625,16.408333,11.041667,16.775,44.233334,15.831249,14.433333,6.5375,7.3083334,8.637501,28.75,14.408335,8.181251,4.8500004,1.03125,1.0666667,1.4749999,0.099999994,0.016666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.074999996,2.4375,3.2083335,1.00625,0.008333334,0.0,0.0,0.0,0.0,0.0,0.0,0.008333334,0.9375,1.85,2.69375,1.8416666,0.8333333,0.28750002,0.09166667,0.043750003,0.25,0.77500004,0.75,0.40833336,0.0625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.11250001,0.33333334,0.075,0.025,0.01875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01875,0.28333336,1.04375,2.1999998,3.1333332,2.8124998,1.5999999,1.5312501,1.5916667,0.8375001,0.25,0.0,0.0,0.0,0.13125,0.925,3.1187499,5.641666,7.933334,11.462501,13.191667,10.762501,6.6166673,3.2187502,0.058333337,0.044444446,0.011111111,0.025000002,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.0,0.0,0.0,0.0,0.0,0.51666677,2.711111,4.2583327,5.111111,2.2333336,0.45555556,3.1000001,2.325,1.1444445,0.45833334,0.8555556,1.3166667,1.2111111,2.25,3.1777778,3.377778,2.7250001,2.6222222,3.7166667,5.3222227,7.5,9.422222,9.166667,12.991667,16.144444,22.983335,24.0,15.991668,11.177778,12.8,15.783336,18.01111,9.408332,2.5555553,0.79999995,0.7444445,2.075,4.8,7.622222,10.299999,13.688889,17.258335,20.233335,22.458332,23.511114,21.1,19.733332,21.444447,21.050003,21.48889,16.724998,13.266668,12.516667,11.9777775,10.677778,7.933334,5.4666667,4.5250006,3.4333336,2.3500001,1.1222222,0.6888889,0.45833334,0.3,0.3166667,0.18888889,0.016666668,0.044444446,0.0,0.0,0.0,0.05,0.12222223,0.12500001,0.16666667,0.15833335,0.13333334,0.08888889,0.31666666,0.96666664,1.8333335,2.7444446,4.833334,7.711111,10.400001,13.758333,18.255552,22.59167,24.022223,20.958334,14.744445,10.483335,7.144445,7.122223,6.5083337,5.6444445,5.4750004,7.8222227,9.95,12.444445,15.111113,17.5,17.666668,15.566666,10.611112,6.533334,4.633333,3.2888892,2.1166668,1.3222222,4.5583334,9.377778,4.875,3.0,5.925,7.866667,9.688889,14.908334,17.666666,22.45,18.411112,14.966667,8.033334,4.8444448,5.7750006,7.6444445,7.2333336,4.966667,7.1333337,10.722221,8.975,7.611111,9.733334,12.641667,17.833334,10.35,19.066666,34.45,43.022224,30.455555,15.1,20.555557,22.449999,4.5888886,1.3583335,0.9111111,0.2,2.5444446,2.9666667,2.35,2.0,0.65000004,0.6555556,1.4666666,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.325,4.6111107,4.133333,0.5222222,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011111111,0.15555556,0.36666667,0.2888889,0.2916667,0.2888889,0.5166667,1.1555556,1.7111111,1.2833334,0.3555556,0.29166666,0.16666667,0.13333334,0.044444446,0.0,0.0,0.0,0.025,0.15555556,0.058333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011111111,0.075,0.25555557,0.45555556,0.46666667,0.97777784,3.8,4.622222,3.208333,1.3000001,0.41111112,0.041666668,0.011111111,0.43333337,1.4444445,2.6833334,2.9555554,1.6666667,2.575,4.0111113,4.491667,2.788889,2.1333334,0.0375,0.008333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.225,0.77500004,2.08125,0.0,0.0,0.0,0.0,3.30625,5.4000006,10.9875,14.724999,13.525,1.7583334,0.9333333,0.26875,0.36666664,0.087500006,0.15000002,0.65625,0.9583334,2.0500002,3.375,4.45,6.025,6.058333,7.05625,8.391667,10.987501,12.566667,16.725,21.324999,18.041666,20.85625,25.216667,28.593748,19.425,17.591667,18.962498,22.541668,13.018751,3.516667,1.1,0.44166666,3.2125,7.775,13.091668,18.850002,21.933334,21.0625,20.791668,22.75,20.25,14.974999,13.53125,15.35,15.68125,11.95,11.437499,10.616667,9.25,7.8666663,5.8333335,4.59375,3.5333335,0.8625,0.3416667,0.23750003,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00625,0.050000004,0.056250006,0.050000004,0.016666668,0.0,0.125,0.4375,0.875,1.8437501,3.4333336,4.583333,7.6687503,11.0,13.793751,14.958334,14.993751,13.9416685,11.70625,10.250001,9.775001,9.043751,10.975,13.20625,14.55,14.45,14.549999,15.058332,16.08125,18.133331,18.8375,17.95,10.34375,4.0916667,1.6666666,2.18125,5.5666666,6.3625,8.383333,7.3374996,5.1916666,4.5625,7.4,8.641666,6.625,11.066667,15.218751,14.133333,7.1250005,4.25,3.5916667,4.0,4.175,5.8999996,6.2083335,4.86875,8.825,5.1437507,5.2166667,6.4,7.71875,8.666668,4.7437506,3.741667,5.8125,8.716666,9.291667,6.15,2.4,7.0250006,1.1916667,0.1625,0.15,1.10625,0.81666666,0.925,0.20625001,1.4083333,0.28125,1.1666667,0.57500005,0.0,0.0,0.0,0.0,0.0,0.0,0.00625,0.05,0.05,0.01875,0.0,0.00625,0.0,0.0,0.0,0.0,0.0,0.0,0.025,0.7083334,1.4875,0.5500001,0.125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.008333334,0.19375,0.25,0.30625,0.56666666,0.9666665,0.90625,0.54999995,0.4375,0.23333335,0.13125001,0.05,0.0,0.0,0.008333334,0.04375,0.083333336,0.09375,0.025,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05625,0.025000002,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.075,0.525,1.0916666,1.7833334,1.5999999,0.9166666,1.31875,2.3666668,3.1562495,2.4083333,2.766667,1.09375,0.0,0.0,0.0,0.0,0.016666668,0.108333334,0.6312501,1.1333333,2.1750002,2.6916668,1.95,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.45833334,0.12222223,0.0,0.033333335,0.12500001,0.0,0.0,0.0,0.0,0.475,14.444445,29.133335,21.088888,21.166668,9.333333,4.3777776,1.6166666,0.42222226,0.15,0.08888889,0.48333335,0.67777777,0.7416667,0.8555556,1.4111112,2.8833332,3.5444446,10.200001,15.388889,20.591667,25.055557,27.644445,27.85,26.277779,28.366667,32.4,35.824997,38.422222,39.97778,42.241665,38.85556,25.591667,8.666667,4.216667,1.7555556,2.675,4.8444443,7.955555,9.075001,8.722222,8.483335,9.633333,13.208334,13.9777775,11.366668,9.383333,10.555555,11.025,10.622222,8.208334,6.088889,3.7916667,2.8555555,2.8222222,2.8166666,2.6222224,1.4499999,0.73333335,0.3,0.07777778,0.011111111,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13333334,0.3111111,0.60833335,0.6333333,0.425,0.08888889,0.0,0.0,0.0,0.0,0.0,0.0,0.0888889,0.10000002,0.13333334,0.2777778,0.86666673,1.9888891,4.8083334,8.4777775,11.175,13.98889,15.916667,18.144445,20.022224,16.233334,13.277778,16.341667,20.38889,21.708334,21.51111,20.744444,18.058332,15.966666,18.083336,20.255556,15.500001,8.88889,5.755555,5.458334,5.911112,5.2250004,7.5444446,9.541667,7.111111,5.125,4.111111,4.455556,3.6083336,6.322222,9.733334,9.3555565,6.0166664,3.511111,4.2666664,4.075,6.288889,10.049999,3.4333334,1.2833333,3.388889,6.4249997,8.955556,10.100002,5.983334,5.8,4.566667,5.2222223,2.4333332,0.96666676,1.1222222,0.9250001,0.9333334,1.8666667,1.4777777,0.30833337,0.4555556,2.6000001,3.8999999,2.7222223,1.5833334,1.1333333,1.9666666,1.3666668,1.35,1.1555556,0.9888889,0.11666667,0.0,0.0,0.0,0.0,0.011111111,0.06666667,0.108333334,0.022222223,0.008333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.033333335,0.0,0.0,0.0,0.0,0.0,0.39166665,1.1888889,0.82500005,0.26666665,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011111111,0.022222223,0.025000002,0.033333335,0.06666667,0.011111111,0.0,0.0,0.0,0.0,0.0,0.06666667,0.22222224,0.36666667,0.044444446,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.2,0.17777778,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.17777778,0.23333335,0.42222223,1.1500001,2.4111114,6.411111,6.275,0.3111111,0.0,0.0,0.008333334,0.2777778,1.8888891,5.7416673,4.411111,6.25,6.566667,6.875001,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.17500001,0.17500001,0.48125,1.375,0.1375,0.0,0.0,0.0,0.0,0.0,0.0,0.08125,4.2583337,12.212501,4.8166666,7.00625,10.308332,11.358334,8.275,3.9333334,0.74375004,0.041666668,0.0125,0.325,1.825,1.6000001,1.85,1.625,1.9666667,7.2375,11.400001,14.40625,17.933332,24.483332,26.500002,25.266668,27.1625,26.274998,23.78125,21.958334,18.891666,16.075,14.083333,7.7125006,3.6583333,1.6312501,0.83333325,0.47500002,0.43333334,0.39166668,0.6125,0.8666667,2.4187503,7.6166663,11.6875,12.541667,10.425001,10.400001,11.391666,10.7125,8.733334,6.96875,6.508333,5.53125,5.9583335,5.416667,4.44375,3.3916667,2.5812502,1.8833334,1.225,0.6666667,0.32500002,0.10625001,0.1,0.087500006,0.19166666,0.4125,0.48333335,0.59999996,0.8187501,1.3583333,2.0125,2.6999998,3.4374998,3.6499999,2.9562502,1.8083334,1.2833334,0.74375004,0.5,0.3125,0.10000001,0.19375,0.4166667,0.4666667,0.58124995,1.0,1.225,1.4166667,2.90625,5.133333,8.11875,11.208334,12.933332,16.487501,16.566668,14.512499,13.691668,15.650001,16.858334,20.066668,18.84375,18.808334,15.568748,15.108333,12.8,9.358334,8.275,8.543751,7.116667,5.0687504,2.675,3.09375,1.325,0.13125,0.083333336,0.0,0.12500001,0.65833336,1.96875,1.8,0.79999995,0.98333335,1.6333334,3.05625,6.2833333,10.250001,4.8500004,0.7875,0.4916667,1.7749999,3.025,4.0416665,2.3125,2.2666664,1.5062499,1.1916667,3.1124997,2.3999999,0.925,1.09375,0.25,0.043750003,0.025000002,0.1125,1.1833334,5.14375,9.708334,7.7916665,4.1499996,2.4750001,1.3,0.9916667,0.82500005,0.9083333,0.8,0.075,0.0,0.0,0.0,0.0,0.0,0.0,0.01875,0.058333337,0.0125,0.008333334,0.0125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.39375,2.0749998,1.6375,1.0166667,0.087500006,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.18333334,0.36666664,0.21875,0.008333334,0.00625,0.025000002,0.025,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.96875,0.22500001,0.0,0.0,0.0,0.0,0.0,0.1,1.5333333,3.91875,1.7,0.73333335,0.59375,0.025,0.0,0.13333334,0.69375,0.40833333,1.9333334,10.362499,12.708334,5.325,4.775,9.256249,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.9333334,4.6777782,2.15,3.9222226,8.05,12.311111,13.766667,12.05,7.244444,3.6083333,1.6333333,0.64166665,0.67777777,1.8416667,0.47777778,0.32222223,0.33333334,0.97777784,5.7750006,9.144444,13.4,12.3555565,11.711111,10.958334,10.644444,11.341666,10.655556,10.45,8.088889,4.366667,2.841667,2.2111113,1.5833334,1.4777778,0.90833336,1.0444443,0.675,0.8111111,0.76666665,0.6333334,1.0111111,8.166667,16.211111,19.408333,16.844444,17.233334,17.041666,16.266666,15.716667,13.366666,11.549999,8.855556,8.650001,9.8,8.4,6.183334,4.366667,2.9666667,2.0777779,0.8,0.24444443,0.022222223,0.05,0.17777778,0.26666665,0.45555556,1.0666666,1.8222224,2.3222225,2.4,1.8888888,1.0166668,0.48888892,0.32500002,0.58888894,1.4666667,3.0777779,3.3111112,3.3833334,2.6333332,1.7499999,0.73333335,0.23333335,0.31111112,0.5555556,1.0250001,1.888889,2.4250002,2.4777777,2.7166667,3.5,5.433334,6.877778,7.077778,7.5166664,9.522223,12.283333,11.944445,12.158335,10.800001,12.677778,12.658334,11.400001,8.866667,7.244445,7.025,5.8555555,3.4444447,2.725,2.9222221,3.1083333,2.3333333,2.0916667,1.3777778,0.33333334,0.055555556,0.35555556,0.033333335,0.0,0.0,0.0,0.13333334,0.2888889,0.022222223,0.51666665,2.011111,1.1999999,1.1444445,0.40833336,0.37777779,1.15,1.3888888,1.6777776,0.98333335,0.33333337,0.25000003,0.033333335,0.53333336,1.2111112,3.766667,7.4083333,9.355556,8.733334,4.8888893,2.4833338,2.3888888,12.666667,33.211113,35.755558,21.958332,12.400002,3.216667,1.1222224,1.8833333,2.766667,2.377778,0.8916667,0.5777778,0.16666667,0.0,0.0,0.0,0.0,0.0,0.0,0.008333334,0.0,0.0,0.011111111,0.008333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06666667,0.0,0.1777778,0.34444445,0.20000003,0.06666667,0.008333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.033333335,0.7000001,1.9833333,1.8555557,0.9666667,0.3888889,0.4,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.2333332,3.0888886,3.6583333,2.0666666,3.1,3.3333335,2.3,4.0000005,12.1,14.716667,9.166668,8.883334,12.91111,15.811112,20.233335,15.6,7.5583334,1.388889,0.41666672,0.22222222,0.22500001,0.16666667,0.42222226,0.7833333,1.4444444,7.016667,15.177779,18.95,17.0,15.511112,12.725001,10.911112,11.266666,12.755556,11.799998,7.511111,4.0333333,2.4250002,1.5555555,1.2666667,1.7333333,1.3833334,1.3111111,1.3833334,1.3888888,1.2444445,1.358333,1.5111111,1.3416667,3.255556,4.4333334,4.511111,4.2666664,4.116667,4.377778,5.766667,6.3444448,6.133333,6.0555553,5.225,6.077778,6.188889,4.8166666,1.8888891,0.48333335,0.29999998,0.475,0.9111111,1.2222223,1.45,1.7555556,1.9250001,2.7666667,4.15,4.933333,6.1666665,6.45,6.3444443,4.8916664,2.0888891,0.8666667,0.5222222,1.1833334,1.7555555,1.6,0.82500005,0.21111111,0.116666675,0.08888889,0.43333334,0.21111111,0.16666667,0.4166667,0.56666666,0.95000005,1.3222221,2.8,4.666667,6.633334,8.222222,7.200001,5.7916675,6.566667,7.0583334,8.388889,8.175001,8.522223,8.577779,7.8250003,5.577778,4.0750003,2.6555557,1.8499999,2.0222223,2.0666668,1.6500001,0.5888889,0.8,0.6111111,0.17500001,0.61111116,0.116666675,0.28888887,0.033333335,0.1,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.12222222,0.33333334,0.23333335,0.21666667,0.8666667,1.2583334,1.4000001,1.7444445,1.825,1.1111112,0.33333337,0.15555558,0.275,2.6444445,13.0,26.183334,30.233334,26.175001,14.455555,7.6250005,2.8111112,4.6083336,17.544445,29.088888,23.441668,15.177777,8.191668,3.8333335,5.2166667,5.0777774,3.733333,1.4416667,0.58888894,0.025000002,0.0,0.0,0.0,0.044444446,0.27500004,0.07777778,0.0,0.0,0.0,0.0,0.0,0.011111111,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.21111111,0.46666664,0.46666667,0.28333336,0.011111111,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.8875,8.35,11.387501,19.5,24.775,22.074999,24.349998,26.841667,27.0,19.01875,7.7166667,1.7625,1.925,4.54375,10.358333,22.524998,31.243752,22.816668,10.224999,4.875,3.84375,2.8000002,2.5062504,2.6666667,5.491667,7.75,10.141666,10.731251,11.85,12.931252,8.791666,9.216667,8.59375,7.9333334,10.01875,14.633333,16.175001,13.466667,11.8,10.48125,9.400001,11.83125,12.441667,6.84375,1.7916667,0.9875,1.1333332,1.25,1.29375,2.025,2.4,2.5500002,2.325,3.3000004,3.3083334,2.1187499,1.8833333,2.2374997,2.0,1.4437501,0.7833333,0.49375004,0.3,0.13333334,0.39374998,1.025,1.2562499,1.475,2.125,2.8916664,3.7583334,4.80625,6.1500006,6.7562504,8.666666,11.18125,15.883334,22.491667,27.431252,24.641666,16.124998,8.983333,4.05,1.6166667,0.91875005,1.05,1.0416666,0.74375,0.3916667,0.31875002,0.26666668,0.2875,0.25,0.06666667,0.25625,1.5666667,2.65,4.05,3.925,5.391667,8.1,11.391667,11.225001,9.456249,7.191667,7.0000005,8.633332,9.468751,7.1333337,5.2,3.875,3.266667,2.125,1.4583334,0.4375,0.22500001,0.35833338,0.66875005,0.6,0.5375,0.39166668,0.0375,0.26666665,0.425,0.0,0.0,0.01875,0.0,0.0,0.0,0.0,0.0,0.425,0.39375,0.4583333,0.41875005,0.26666668,0.17500001,0.5500001,0.6,0.85833335,1.3833334,1.5124999,0.40000004,0.112500004,0.09166667,0.0375,0.89166665,6.650001,21.90625,27.175,23.75625,22.691666,26.95,16.916668,11.881249,9.041667,3.9333339,1.23125,0.90000004,1.25625,1.7249999,1.7312497,0.5083333,0.0,0.0,0.0,0.0125,0.49166667,1.2937499,3.0000002,0.38333336,0.63125,0.44166666,0.17500001,0.05,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,9.822222,44.516663,67.31111,68.76667,63.444443,59.633335,64.422226,49.544445,33.908333,8.633333,1.45,1.0222222,4.25,20.977776,32.18889,31.699999,24.233334,12.991667,7.8555555,5.25,2.8444443,1.9416666,2.1222222,3.4444447,4.3666663,4.2444444,4.2083335,3.3666668,4.516667,5.766667,5.5666666,4.6083336,4.4,7.008333,12.333334,16.933332,16.88889,17.311111,19.4,21.900002,26.441666,21.344444,12.058334,6.1444445,1.9333334,0.4555556,0.6555556,0.87500006,0.8777778,0.6500001,0.8555556,0.7916667,1.9777777,2.588889,1.8416667,0.9666667,0.7750001,0.82222223,1.4583334,1.9444444,2.1083336,2.3555558,2.4777777,3.7916667,3.877778,5.75,6.455556,5.825,5.711111,6.0,6.908334,10.622223,14.816667,19.955557,26.133335,31.233334,36.555553,43.11667,43.755554,31.125,18.533333,8.3,4.0222225,2.0333335,1.1888889,1.2222223,0.7416666,0.3,0.108333334,0.06666667,0.25833333,0.9,0.7777778,0.7916667,1.8555555,2.3999999,2.6222224,4.308333,6.1777782,8.358334,10.044445,9.166666,9.091667,7.4888887,5.3833337,4.9111114,6.466667,7.0000005,6.4333334,4.4583335,3.0222223,1.9916666,1.2888889,0.71666664,0.1,0.033333335,0.18333334,0.2,0.21666667,0.08888889,0.10000001,0.022222223,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.044444446,2.0444443,4.1499996,0.26666668,0.52500004,0.33333334,0.33333334,0.33333334,0.28333336,1.1888889,1.7444444,2.0500002,0.88888884,0.016666668,0.0,0.0,0.07777778,1.1222223,4.8250003,5.466667,6.466667,15.766667,28.983332,22.144444,13.350001,9.266667,11.6,10.05,2.2555556,0.14166667,0.1,0.35833338,0.044444446,0.0,0.0,0.0,0.008333334,0.31111112,1.8333333,4.366667,1.8222221,0.17500001,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,4.083333,29.750002,64.89166,83.21875,74.59167,71.79375,74.70833,68.77501,38.343754,15.183334,5.725,4.158334,19.650002,34.491665,25.691668,22.425,15.866666,4.51875,2.2250001,1.2437499,0.7416667,0.65000004,0.89166665,2.9666665,6.59375,10.525001,15.350001,15.6,12.637501,10.233335,6.4583335,4.63125,3.3416672,3.34375,3.6333332,5.5062494,6.9000006,8.775,9.88125,10.658333,11.643751,13.433333,16.512499,12.466666,4.0,0.34166667,0.42499998,0.5625,0.5833333,0.48125002,0.4833334,0.89375,1.2083334,1.0416667,1.0125,1.3083335,2.9750001,5.1333337,8.412499,10.808333,12.5125,14.016668,14.016666,15.5,18.708332,20.256248,21.40833,19.00625,14.108334,13.6833315,14.625,15.591666,14.94375,12.683333,10.450001,10.658333,13.183332,16.725,23.066666,26.568748,17.258335,7.9125004,2.5833335,2.2187502,2.7583332,2.2416666,1.4062501,0.62500006,0.15625,0.075,0.6312501,0.85833335,0.84999996,0.875,2.0,2.1375003,2.075,2.40625,3.05,3.0,3.141667,3.2333333,3.30625,3.275,2.16875,1.9416668,2.78125,3.525,3.5083332,3.0812502,2.2083335,1.3437501,0.8833333,0.47500005,0.18333334,0.058333337,0.0,0.0,0.00625,0.15833335,0.27499998,0.13333334,1.15625,2.1,2.575,1.8,0.7,0.225,0.075,0.0,0.116666675,0.8583334,1.15625,0.35,0.10000001,0.0,0.20000002,0.5500001,0.6875001,1.1166667,0.8083334,0.69375,0.5,0.13750002,0.033333335,0.04375,0.6416667,1.375,1.64375,2.2166667,4.3625,8.833333,11.325,7.8583336,3.59375,1.8583333,7.6000004,22.431252,10.624999,0.65000004,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05625,0.4416667,0.3333333,0.06875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.9166667,4.088889,20.141666,46.15556,54.29167,47.68889,40.658333,42.522224,33.4,18.466667,8.077778,3.3416667,8.888889,12.666669,14.077778,9.611111,9.125,3.8111112,3.0583334,1.7000002,0.6,0.1888889,0.083333336,0.022222223,2.3888888,6.6833334,12.633334,21.558332,28.266666,17.608334,14.444446,9.677777,6.4083333,4.722222,3.4,2.4333334,1.9750001,2.7555556,4.9555554,6.083333,3.5555558,4.6499996,10.088888,22.716667,36.100002,29.76667,7.5333343,2.211111,1.8416667,1.111111,0.5,0.44444448,0.39166668,0.2,0.41111112,1.4333334,3.5555556,5.8083334,8.288889,10.483334,11.1888895,12.441666,12.788889,11.733334,10.525,10.055555,10.591666,10.077778,7.0333333,3.566667,2.2555554,2.9333332,3.6777778,3.6916666,2.511111,1.5333333,1.4,1.2555554,1.9250001,2.5555553,4.616667,5.022222,5.3750005,5.4111114,4.8500004,4.1,3.5555558,3.225,1.8444446,1.25,0.34444445,0.0,0.033333335,0.32222223,1.5583334,3.266667,4.7333336,4.7222223,3.6000001,2.9888887,2.6333332,2.1777778,1.3111111,0.9583334,0.9888889,1.3416667,1.3333334,1.8,4.9222226,7.0555553,4.6083336,3.4444447,2.5749998,1.6555556,1.5333333,0.8222223,0.17777778,0.14166668,0.11111111,0.13333333,0.08888889,0.675,1.3666668,10.566666,18.7,21.400002,23.450003,12.455555,2.9916668,0.6888889,0.14166668,0.022222223,0.13333334,0.84166664,0.50000006,0.016666668,0.0,0.0,0.22222222,0.4833334,1.0333333,0.7777778,0.016666668,0.0,0.0,0.0,0.0,0.0,0.10000001,1.0250001,2.677778,2.9250004,4.466667,13.641666,26.066666,19.083336,5.0444446,1.4,0.28333336,0.15555555,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.4666667,1.3555555,0.4666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0375,1.5083333,10.162499,27.391668,37.09375,25.416668,18.09375,12.474999,10.075,7.462501,2.5749998,3.4562497,7.266667,7.2999997,5.3083334,7.3083334,8.712501,10.766667,7.693751,5.283333,5.1625004,6.5333333,7.0375,6.825001,3.95,4.25625,5.1833334,9.43125,13.266666,6.7562504,4.758333,4.6250005,4.33125,5.0833335,5.45,4.008333,3.2749999,4.0833335,6.825,6.3624997,4.983333,5.93125,12.991666,29.393751,34.0,30.625,12.449999,4.066667,3.3125005,1.8833333,0.81875,0.18333334,0.10625,0.375,0.9999999,2.6437502,3.9916663,5.10625,4.708333,4.6375,4.25,4.075,3.6666667,2.9583333,2.1187499,1.8333333,1.475,1.4666667,1.3687501,1.2500001,1.2333333,1.24375,1.475,1.275,0.94166666,0.4375,0.26666668,0.108333334,0.5187501,0.89166677,1.58125,2.275,3.28125,4.6750007,5.26875,5.2750006,3.966667,3.1687498,2.2083335,1.6125,0.7166667,0.43124998,0.14166668,0.06666667,0.09375001,0.38333336,1.1812501,3.1499996,3.0562503,1.2666668,1.20625,1.3416667,2.0083332,2.0375,1.2583333,1.3875,1.9916667,1.83125,2.3333333,4.4583335,4.9312506,3.6416667,2.7687502,1.9916666,1.4562501,0.8083334,0.43333334,0.13749999,0.058333337,0.0,0.0,0.15625,0.52500004,3.275,5.45,8.25,10.012501,3.2333333,1.15625,0.2916667,0.09375,0.008333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03125,0.09166667,0.083333336,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.26875,1.8666667,3.6562502,4.3500004,10.243751,20.091665,16.43125,5.575,1.375,0.18125,0.27500004,0.31250003,0.008333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.33125,0.025,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016666668,0.26875,0.025,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.09166667,0.9375,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08888889,0.99166656,2.3777778,6.466666,14.455556,18.475,12.355556,6.783333,3.1444445,2.688889,5.4,6.7222223,7.5000005,6.544445,9.483334,15.311111,17.688889,6.725,3.877778,3.5583334,6.0333333,4.6916666,8.444445,10.808333,7.8999996,5.1888885,2.3666668,3.4000003,4.858333,4.3444443,6.0499997,5.577778,4.5555553,5.241667,9.633333,10.316667,8.333334,5.891667,4.322222,4.533334,5.2083335,5.7555556,6.1666665,6.3333335,12.191668,17.733334,9.650001,2.4666667,1.6777778,1.1166668,0.6222222,0.3083333,0.34444445,0.49166667,0.71111107,1.4000002,1.9333334,2.6666667,2.8249998,3.5666668,4.2166667,4.122222,2.8333333,1.9111112,1.0,0.6333333,0.31111112,0.125,0.12222223,0.10000001,0.099999994,0.22222222,0.40833336,0.6111111,0.475,0.25555554,0.0,0.0,0.0,0.20833336,0.5222222,1.3166667,2.2666667,3.3833334,3.9444444,4.7333336,5.3777776,5.944445,8.516667,13.333334,18.175,17.233334,8.250001,3.3777778,2.2444446,1.4416666,0.48888892,0.40000004,2.1666667,4.85,5.2333336,3.8500001,2.7555554,2.3555558,2.0083332,1.5666666,2.0,3.0666666,4.7500005,4.911111,4.6000004,4.6333337,4.188889,4.0,3.3555555,4.3333335,2.1333334,0.7777778,0.058333337,0.0,0.0,0.0,0.0,0.0,0.0,0.022222223,0.4666667,4.3,7.2222223,4.3083334,1.8000001,0.24166666,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14444444,1.6333334,3.6222222,3.7500002,2.5666666,0.99166673,0.4,0.26666668,0.7111111,0.6888889,0.30833334,0.011111111,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.55,0.51111114,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.0333333,3.6333334,4.7222223,8.308332,10.1,9.308333,4.8444448,3.058333,2.1444445,1.5333334,8.891666,20.022223,22.150002,21.166666,16.133333,33.31111,27.88889,2.7166667,2.9333334,8.366667,13.533333,14.008333,17.044445,17.191666,13.922222,9.0222225,5.8333335,4.8444443,3.0666668,2.0666666,3.358333,4.5666666,11.288889,27.208334,33.088894,25.416668,10.277778,4.1416664,2.6333332,3.5777779,4.1333337,4.6333337,5.1,7.9000006,9.15,8.1888895,5.5416665,2.8999999,2.0333333,1.0500001,0.24444446,0.116666675,0.32222223,0.38333338,0.6,0.47777778,0.9416667,1.9333334,4.383334,4.544444,4.866667,3.677778,2.8416667,2.1111114,1.4555557,0.6000001,0.16666669,0.8333334,0.5222222,0.13333334,0.18888889,0.24444446,1.3,1.7222223,0.875,0.14444444,0.13333334,0.0,0.0,0.0,0.022222223,0.125,0.43333334,0.9833333,1.2222221,2.3583333,4.522222,6.2666664,7.2666664,10.311111,18.866667,25.500002,22.308334,13.277778,5.388889,2.2666667,2.9222221,6.2083335,8.155556,6.1749997,8.011111,7.3083334,5.333333,4.3333335,3.5499997,3.1222222,2.2916667,1.488889,1.8750001,3.3111112,5.9555554,10.208334,7.4666667,6.0249996,4.6666665,3.2166667,2.7222223,1.2777779,0.30833334,0.0,0.0,0.0,0.116666675,0.6000001,0.075,0.1,0.0,0.05,0.53333336,0.77500004,0.7222222,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.1333334,10.555556,4.7666664,2.9777775,2.9333332,0.5555555,0.125,0.022222223,0.011111111,0.025000002,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016666668,0.22222224,0.14166668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025000002,0.28888887,0.21111113,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.2916667,0.45000002,0.90833336,7.6187506,10.716667,8.568749,5.925,5.7374997,7.25,1.9416665,8.09375,15.349999,14.5125,19.025,10.500001,17.266666,8.891666,4.76875,8.416667,13.250001,23.983335,35.7125,33.75833,22.2875,14.033334,11.925,7.95625,3.9,3.00625,7.9916673,20.1625,28.858334,36.08334,41.175,29.350002,15.1625,8.225,7.2875,6.575,7.3000007,9.900001,12.775001,15.606251,17.883333,16.118752,13.366667,12.04375,11.05,5.541667,2.7625,0.15,0.081250004,0.058333337,0.11250001,0.35833335,0.53333336,1.8687501,4.3083334,6.33125,6.666667,5.2312503,3.841667,2.6374998,2.15,1.75,1.0875001,1.675,4.3375,0.9333334,0.13750002,0.325,0.67499995,1.6624999,2.6583333,2.0375,0.39166668,0.15625,0.20833333,0.43333334,1.0374999,1.5583334,1.78125,1.9666667,3.18125,3.4916668,2.8875003,1.775,1.3666667,2.925,4.1916666,8.462501,13.808333,14.856251,9.825,6.8,6.6187506,10.799999,10.650001,9.05,7.51875,8.841667,9.2375,8.450001,7.766667,7.4625,5.8999996,5.26875,3.516667,1.9187499,1.3083334,2.85,5.2062507,5.3250003,4.54375,3.6250002,2.525,3.45,3.3083332,1.5562501,0.5583334,0.0,0.06666667,0.05,0.0,0.24375,0.275,0.0,0.425,0.85,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.4916667,0.78125,0.19166668,0.39375,0.60833335,0.18750001,0.033333335,0.041666668,0.05,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03125,0.025,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.033333335,0.06666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.17777778,5.3166666,10.822222,8.816668,6.166667,6.1,15.233334,4.233333,11.016667,20.288889,18.758335,12.811111,2.9833333,0.13333334,0.022222223,0.0,1.6888889,5.166667,16.622223,41.391666,54.944447,33.6,12.922223,8.266666,5.0916667,4.8,5.8999996,11.566668,13.758334,12.0666685,14.400002,14.666667,9.988889,8.733334,10.388889,13.783333,14.733334,17.244444,22.45,14.022223,13.983334,11.433334,7.2083335,5.355556,3.9499996,1.7444446,1.0111111,1.1166667,0.14444445,0.3,0.47777778,1.5333334,2.4444444,3.0777779,3.1166668,2.7444444,2.9833333,2.6444445,2.0416667,1.8444446,1.8833334,2.1777775,3.0444446,4.6333337,3.2666667,0.7916666,0.033333335,0.025000002,0.13333334,0.44444445,1.5833331,2.377778,3.025,1.5555555,0.9666667,1.011111,0.9,1.0916667,1.1222222,1.7,2.5444446,6.5916667,9.711111,8.216667,3.9111114,1.6555556,1.3416667,2.088889,4.4333334,6.1444445,6.933334,5.777778,4.577778,5.9416666,6.7666664,6.6,6.0000005,7.05,12.288888,14.783333,14.211109,12.333334,12.300001,11.033334,9.016666,7.5,6.2000003,6.577778,6.633333,5.375,4.488889,3.8000004,1.7333333,2.9166667,7.3555555,7.4111114,1.2416668,0.0,0.0,0.0,0.0,0.033333335,1.2750001,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.6666667,1.2916667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011111111,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05,0.2,3.7062497,9.341667,6.2437506,4.3916674,2.25,10.499999,6.4333334,7.9749994,9.15,3.25625,2.1499999,0.57500005,0.016666668,0.0,0.0,0.28333333,3.825,13.225001,28.16875,25.291666,17.918749,12.258334,8.366667,8.831251,14.950001,16.075,11.458333,5.025,2.275,1.6250001,2.8374999,6.4666667,8.975,13.625,18.29375,14.708333,12.958335,11.831251,9.416666,6.606251,3.15,0.98749995,0.38333336,0.32500002,0.15833333,0.3416667,0.6125,0.75,0.98125005,0.125,0.33125,0.6,0.6166667,0.43124998,0.85,4.24375,3.0249999,2.6187503,3.7000003,5.1875,11.625001,22.85,20.06875,4.858333,1.3249999,0.083333336,0.6187501,1.7583334,2.075,2.5375,3.25,4.3875,5.7166667,7.7125006,7.6749997,9.858335,8.94375,8.308333,5.1124997,4.025,4.975,4.608333,4.1187506,3.55,3.658333,2.7625,1.85,2.9812498,6.6916666,9.868751,7.4249997,5.3,6.2312503,6.200001,6.7375,7.0999994,5.1375003,8.849999,11.1875,11.5,10.275,8.53125,7.8166666,7.8500004,8.433334,10.81875,14.666667,16.083334,17.15625,16.875,13.825,10.258333,7.3062506,3.6666665,1.3083334,0.77500004,0.5,1.09375,0.5416667,0.0,0.05,0.22500001,0.93333334,0.7,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.20833334,0.31875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.7250001,9.422222,4.6083336,1.7444445,1.1833333,2.311111,2.8000002,1.5333333,1.1666667,2.8750002,1.1111112,0.73333335,0.0,0.0,0.0,0.022222223,0.725,4.488889,6.9083343,9.422222,11.216668,9.722221,9.222223,18.691666,22.166664,14.483333,7.1,4.516667,1.0777777,0.7555555,3.0749998,5.6222224,5.908334,5.8222227,6.4750004,8.3,13.044445,13.908334,6.1555557,1.9416668,1.3,1.9666667,4.0222225,4.141667,2.9888887,3.277778,3.1333334,1.5333333,0.35833332,0.044444446,0.0,0.0,0.0,0.23333333,0.9111111,3.7666667,4.1555557,5.341666,7.1,8.2,14.111111,25.677776,16.358334,3.2,0.47500002,0.5,1.8333333,2.411111,3.8777776,3.2916667,4.422222,7.391667,9.811111,14.65,14.944445,9.466666,7.5666666,8.277778,8.85,9.1,9.283334,7.633334,6.583333,5.455556,3.7444444,2.2333333,1.9,2.9916668,6.311111,8.866668,5.377778,3.6,2.9666665,1.1333333,3.3666663,2.411111,1.0,1.2111112,2.9083335,4.5111113,4.366667,4.791667,6.955556,9.075,11.833334,14.525002,14.844444,15.8,18.058332,17.322224,20.550001,25.377777,24.383335,20.222221,14.466666,8.625,14.533333,4.0750003,0.0888889,0.30000004,0.0,0.16666667,0.022222223,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.425,3.1125002,6.6083336,3.2187498,1.0333335,0.69375,0.1,1.2416667,1.11875,0.50000006,2.3812501,2.5833335,1.1187501,0.116666675,0.0,0.09375,1.0833333,5.31875,2.3,2.44375,3.2583337,5.1875005,6.508333,7.075,5.8750005,6.533333,4.5937505,3.8916667,4.5874996,3.0833333,2.5166667,2.5875,2.575,2.5062501,4.3750005,6.5,6.1499996,5.7333336,3.0062501,2.875,2.99375,3.4833333,8.9375,11.033334,6.4624996,8.266666,6.45,4.1437507,1.7666669,0.125,0.0,0.056250002,0.19999999,0.71666664,3.2312505,3.3916667,5.0000005,2.0916667,0.75,1.6166667,2.6499999,3.9333336,5.266667,3.50625,1.05,0.275,0.6166667,1.3625,2.2166667,2.275,1.6812502,2.5249999,4.46875,6.691667,9.15,11.625,10.025,8.712501,9.225,12.474999,15.2,17.625002,18.275002,18.631252,19.975,21.358334,15.15,12.966667,8.443749,7.616667,8.231251,10.233334,15.691666,15.49375,13.008335,11.518751,5.766667,6.125,5.325,4.70625,4.2166667,3.9833333,4.99375,7.233333,7.21875,8.3,9.35625,9.424999,9.991666,11.525,10.516667,8.88125,11.091666,17.225002,28.950005,31.533333,21.962498,9.733334,2.6999998,0.025,0.0,0.0,0.125,0.2,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016666668,0.11111111,1.25,2.0666666,0.8833334,1.0333334,0.7583333,0.15555556,1.2,1.3083334,0.8333333,0.5,1.4666668,0.22500001,0.0,0.72222227,2.3083334,0.43333337,1.3499999,0.42222223,0.525,2.7777777,3.4916668,1.7111111,0.3,1.5666666,4.9222226,7.7000003,10.622222,15.891665,13.355557,9.233334,8.650001,8.588889,6.4333334,3.3,0.8166668,0.40000004,1.9222223,5.0,9.611111,19.233334,29.155558,27.283335,30.655554,21.7,16.555555,9.400001,2.7416668,0.2111111,0.125,0.07777778,0.7416667,1.9222224,2.2444446,3.2333333,5.9666667,7.5249996,0.8,0.025,0.14444445,0.925,1.0666666,0.4888889,0.16666667,0.14444445,0.525,0.88888884,1.0916667,1.3222222,1.8333334,3.7416666,7.5111117,12.616667,14.744444,11.741668,7.122222,7.988889,8.3,6.622223,8.191668,10.955556,18.708334,24.97778,33.125,43.166668,59.8,69.10834,75.53334,60.00834,34.77778,17.858334,13.244444,21.666668,33.591667,30.766666,26.25,15.4,8.858334,4.6222224,3.6916666,1.8777778,1.1888889,2.375,4.2222223,4.125,3.3444448,2.6,2.8777778,4.0222225,5.0750003,5.7000003,5.216667,4.711111,3.4666667,2.5444443,5.1888885,9.108332,3.7444446,0.23333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016666668,0.0,0.0,0.13125001,0.09166667,0.10625,0.275,1.4916667,1.03125,0.69166666,0.625,1.3583333,0.4125,0.16666667,0.9916666,2.30625,0.0,0.1,0.26666665,0.19375,0.8000001,0.43125004,0.7333333,1.3750001,4.325,9.441667,14.81875,19.725,25.393747,28.816666,35.758335,33.31875,20.81667,10.725,3.9166667,0.85624987,0.3416667,1.8416667,12.34375,24.675,36.53125,47.783333,50.225002,45.575,34.06875,20.949999,13.058333,4.1375,0.5583334,0.73125,1.0250001,1.18125,1.6416669,1.0500002,0.38124996,0.41666666,0.225,0.0,0.0,0.20833333,1.0562501,0.6833334,0.24166663,0.71875,1.4666667,1.5,0.725,0.49375004,0.44166666,0.7666667,2.54375,6.5583334,10.49375,11.65,9.825001,9.041667,11.991667,18.25,24.008335,26.68125,27.066666,24.09375,32.175003,41.518753,50.100002,55.45,59.887497,62.05,56.262505,45.725002,32.068752,22.208334,22.333336,26.893753,26.4,20.287498,16.625,13.09375,8.025,5.3750005,5.575,5.408334,6.2999997,6.291667,5.3937497,5.791667,5.35,4.7416673,3.9166665,2.9437501,5.0083337,4.18125,2.4,2.1125,1.2833333,0.575,0.31875,0.5916667,0.16875002,0.26666668,0.13125001,0.058333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.21666667,0.45555556,2.4555557,0.425,0.044444446,1.3666667,0.7333333,0.0,1.6000001,1.25,0.64444447,0.6555556,1.8249999,1.5333333,0.3166667,0.0,0.35000002,0.6777778,1.9444447,1.525,0.31111112,0.116666675,0.22222224,0.14166668,0.044444446,0.0,0.044444446,0.2777778,2.825,6.311111,10.266667,14.177778,21.241667,27.066668,30.18889,31.924997,16.355555,6.3000007,2.0222223,2.475,3.4222221,6.8444443,19.733334,39.98889,43.408333,48.622223,41.308334,28.366669,17.066666,6.733333,3.377778,1.3083334,0.8333334,0.99166656,0.9666667,2.0333333,4.3555555,5.5444446,2.0166667,0.46666673,0.041666668,0.0,0.0,0.0,0.0,0.0,0.1777778,1.0749999,2.588889,2.1166668,0.2777778,0.275,0.36666667,0.3888889,0.45833334,0.59999996,0.78333336,1.4111112,2.3583333,3.6333332,5.6666665,12.466667,19.944445,23.541668,23.722223,16.591667,15.755555,21.041666,27.033333,22.022223,17.191668,17.41111,16.150002,16.444445,21.125,25.077778,24.977777,29.8,29.022223,25.816668,19.433334,10.358334,5.0222225,3.9583333,5.0111113,5.8444448,8.674999,10.533333,9.65,6.7444444,6.383333,6.8333335,5.7222223,2.5166664,0.2777778,0.06666667,0.0,0.116666675,0.20000002,0.07777777,0.016666668,0.2888889,0.0,0.0,0.0,0.011111111,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.8916667,7.1000004,17.077778,32.39167,11.211111,9.141666,10.1,3.2333338,2.1666667,15.541668,30.666668,12.388889,0.7250001,0.5888889,1.1750001,0.3222222,1.125,0.3555556,2.3777776,3.4833333,2.3777778,0.21666668,0.044444446,0.075,0.0,0.0,0.0,0.19999999,1.4083334,3.977778,6.8166666,11.444445,17.583334,27.277779,29.511112,15.200001,2.9888887,0.825,0.8777777,2.2083333,4.877778,13.744444,24.716667,33.98889,32.300003,27.255556,17.158333,8.088889,3.5583334,0.81111115,1.0111113,0.64166665,2.222222,4.1666665,6.3555555,6.791667,5.466667,3.088889,1.475,0.25555554,0.24166667,0.2777778,0.73333335,0.70000005,0.5083334,0.18888889,0.32222223,1.65,2.088889,1.3166666,0.5,0.55,0.4333333,0.35555556,0.975,1.3555555,1.2,1.4000001,1.4583333,1.2555555,0.96666664,0.7916666,0.7777778,1.4666666,2.222222,0.90833336,0.7,1.3,3.0222223,4.4555554,6.9333334,3.5555556,3.1416667,2.9222224,5.391667,7.122223,11.066667,16.85,20.377779,19.2,16.044445,13.333332,11.4,8.900001,7.7777786,6.9333334,9.0,10.3555565,10.791667,12.266667,13.316668,11.511112,7.4222226,2.3916667,0.18888889,0.15833335,0.0,0.0,0.0,0.011111111,0.34166667,0.13333334,0.0,0.0,0.0,0.044444446,0.22500001,0.10000001,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.28750002,0.0,0.0,0.0,0.0,0.0,0.0,0.26875,4.3500004,13.983333,22.787502,12.725,9.0,8.858334,9.0,11.858334,33.1625,61.033333,52.65,12.93125,2.125,1.46875,0.6833334,0.7125,0.775,1.4333333,2.525,2.1416667,0.6187501,0.35833335,0.57500005,0.31666666,0.13750002,0.0,0.05,0.61249995,2.3333335,5.2812505,12.308333,19.20625,18.683334,12.366668,4.5750003,0.69166666,0.23125,0.15,1.5250001,13.658333,27.250002,37.49375,42.025,31.175001,19.1,8.143749,1.6416667,0.118750006,0.05,0.8250001,1.0625,2.8583333,3.04375,2.9666667,2.0625,0.575,0.075,0.00625,0.35833335,1.7750001,3.5833335,3.74375,1.7999998,0.825,0.28333336,0.47500002,0.3125,0.058333337,0.1875,0.7333333,0.7750001,0.78333336,4.108333,1.1875001,0.083333336,0.93125,1.9250001,4.24375,0.7083334,0.108333334,0.84375006,2.7,1.5,0.025000002,0.0,0.13333334,0.65,3.0083334,4.691667,6.1812496,13.924999,10.075001,1.9333333,1.8125,2.2666667,2.4416668,4.5,5.141667,6.1875,13.238637,20.71875,15.491667,7.9687495,3.8833337,3.1416664,4.55625,7.758333,7.93125,7.0166664,7.337501,5.433333,3.2333333,1.43125,0.725,0.34375,0.0,0.0125,0.033333335,0.05,0.0125,0.0,0.0,0.0,0.0,0.49166664,1.025,0.7583333,1.625,0.34375,4.3083334,0.28750002,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.20833333,0.89374995,0.083333336,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.266667,0.0,0.22222222,0.0,0.0,0.0,0.0,0.0,1.4222223,8.255556,7.333333,2.0,2.1750002,1.5888889,3.5,11.522222,33.716667,51.21111,57.96667,54.525,8.811111,1.4333334,1.2222222,0.09166667,0.044444446,0.0,2.1583333,2.0555553,0.3,1.3888888,1.0333333,0.13333334,0.06666667,0.0,0.0,0.325,2.6444445,13.333333,71.52222,30.525,7.6666675,2.6111112,0.7916667,0.16666669,0.35000002,1.5666666,5.675,13.933334,24.944445,37.016666,39.799995,31.175,17.277779,7.125001,1.9111111,0.94166666,2.3111112,5.555556,4.125,6.788889,3.4833333,0.55555564,0.4583334,0.9888889,0.75555557,0.062121212,0.0,0.23333336,2.977778,0.8916666,0.011111111,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016666668,0.36666667,1.9,0.041666668,0.0,0.15833333,0.36666667,2.2166667,0.85555553,0.0,0.23333335,2.8222222,2.675,0.42222223,0.050000004,0.21111113,0.33333334,0.43333334,2.688889,7.7083335,9.9,7.908333,6.7111115,7.991667,9.955557,12.455556,12.733333,4.288889,2.975,11.255555,17.074999,12.244445,5.458333,2.1666667,2.0222223,3.5,2.8999999,2.4416666,1.5666667,1.175,1.7,1.8111112,2.425,1.3333333,0.9166667,0.36666667,0.16666669,0.5555555,0.6666667,0.75,0.7444445,0.60833335,2.911111,3.216667,1.0333333,1.3583333,1.1444445,1.6444445,2.05,2.7222223,0.25,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.95000005,0.2777778,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.35,2.5833333,3.4083333,0.0,0.0,0.056250002,0.24166666,0.35,0.40833333,1.4166667,3.8687499,1.1083333,0.44375002,0.116666675,2.3437498,5.4583335,27.487501,52.058334,63.00833,50.95,25.25,3.49375,2.391667,2.1687498,0.4083334,0.23333333,1.05625,1.525,0.9687501,1.4000001,1.7375,0.21666668,0.09375,0.008333334,0.08333334,0.84375,3.525,32.225,51.733337,20.44375,4.25,0.6000001,0.575,2.3083334,4.48125,7.55,14.2875,26.466665,40.5,52.4875,43.858337,31.65625,11.241667,2.1437502,0.93333334,1.375,1.55,1.1666665,1.09375,1.95,2.55,0.47499993,2.5266666,5.0249996,1.2166667,0.06666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.075,0.33333337,0.375,2.4750001,0.33875,0.2916667,1.3687499,1.4749999,1.7249999,0.9083333,0.31666666,0.1875,0.15,0.68125,1.8083333,3.0000002,4.9000006,5.366667,2.7187502,1.3083333,2.40625,3.1757574,1.0733334,0.80833334,1.7875,1.6833334,1.0583334,0.9875,1.625,0.47499996,0.15833335,0.34375,0.37500003,0.6166667,1.675,1.7583334,2.0,2.391667,0.8,0.55833334,0.5416667,0.91875,1.6166668,2.59375,4.175,10.325001,8.083333,2.5375,1.7333333,2.2999997,4.6562505,1.5666668,0.00625,0.0,0.099999994,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.087500006,0.5416667,0.1625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,6.6000004,6.6444445,0.0,0.0,3.7666667,3.4888892,3.416667,2.8777778,0.06666667,0.25,0.6888889,1.25,0.2,0.0,1.7555556,8.633333,35.255558,67.46667,55.983334,43.5,18.683334,3.411111,2.4,1.4888889,0.9777778,0.85833335,0.14444445,1.3166667,4.211111,2.9166665,0.0,0.0,0.0,0.14444445,2.533333,3.855556,21.566666,46.38889,40.608334,1.8888887,2.6222224,5.441667,11.011111,10.291667,8.866667,16.158333,29.866667,30.622223,28.791666,24.044443,16.475,3.1999998,1.1666666,1.1555555,1.5250001,2.666667,1.7333333,2.5333333,0.3111111,0.9000001,0.011111111,0.008333334,0.43333334,0.0,0.0,0.044444446,0.016666668,0.0,0.0,0.0,0.0,1.2888889,0.055555556,0.16666667,0.24444444,0.20833333,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.31250003,0.41666666,0.0,0.0,0.0,0.075,0.08888889,0.0,0.0,0.0,0.083333336,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.23333333,0.47777775,0.6666666,1.7666667,5.4250007,7.744445,5.1222224,1.8500001,0.13333334,0.29999998,0.4333333,1.1166667,0.6888889,0.18888889,0.16666669,0.8444444,1.3166667,2.1666667,2.1166668,0.48888886,1.2111111,0.95,0.7555555,1.575,4.266667,4.9416666,7.9111114,8.325,10.788889,13.388889,6.508333,0.53333336,0.016666668,0.0,0.28333333,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.48333332,0.12222222,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,3.4333334,15.650001,15.312502,0.0,4.6,4.241667,3.3562498,3.183333,0.5833333,0.2875,0.0,0.23750001,0.125,0.0,0.0,0.325,5.7666664,25.941666,29.26875,31.974997,30.78125,12.150001,5.6000004,3.1666667,1.5083333,0.3375,0.15833335,0.65625,2.0416665,1.125,0.0,2.34375,2.4833336,2.5333333,1.275,0.54999995,3.8375006,49.450005,33.699997,7.1833334,16.091667,31.74375,28.141668,23.45,13.825001,18.4125,27.283337,30.783333,14.262501,10.383334,5.4875,4.7333336,2.65625,2.5833333,1.8375001,1.6712121,1.3083332,0.10000001,0.09166667,0.056250002,0.0,1.0237501,0.85833335,1.05,4.7125,4.7833333,0.55,0.0,0.0,0.058333337,0.2375,0.6,1.0749999,0.34375,0.0,0.0,0.0,0.0,0.0,0.35833335,6.075,1.8083334,0.6625,0.13333334,0.0,0.0,0.04,0.09375,0.026515152,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05,0.15,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.087500006,0.21666667,1.85625,5.6083336,7.5037875,6.48125,3.875,2.9750004,4.1916666,5.1562495,3.9250002,3.0583334,1.4062501,0.5083333,0.425,0.80833334,1.1625,0.65,4.1499996,4.8125,1.3583333,1.275,2.625,1.8937501,1.425,7.9375005,17.875002,16.141668,7.9937506,0.8166667,0.0,0.0,0.025,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03125,0.06666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,22.644445,37.191666,6.9333334,1.025,2.0,0.52500004,0.36666667,2.3333335,1.9916668,0.3,0.17500001,0.10000001,0.14166668,0.2777778,0.075,0.32222223,2.2111113,7.1333337,10.644445,18.783335,13.866667,7.4083323,0.71111107,0.61111116,1.8750001,0.51111114,0.40833336,1.2777778,2.4916668,0.31111112,1.4583333,1.8000002,2.2111113,0.78333336,0.33333337,1.4083335,6.8000007,10.041668,18.7,63.11111,64.691666,63.266666,47.516666,28.955555,28.333334,36.63333,32.755554,10.733334,2.6777778,0.25000003,0.0,0.0,0.022222223,0.038333334,0.0,0.0,0.025000002,0.0,0.016666668,0.58888894,4.45,1.0777777,1.3111112,2.3166666,3.2111113,2.7166667,0.5555556,0.041666668,0.39999998,1.3166666,2.6222224,2.8444443,0.55,0.033333335,0.0,0.0,0.0,0.044444446,0.06666667,2.2,14.888889,9.933333,2.4333334,0.675,0.34444448,0.54305553,0.729293,1.3313493,0.8333334,0.8555556,0.025000002,0.0,0.0,0.0,0.0,0.0,0.0,0.7166667,1.0,1.1583333,0.6666666,0.3333333,0.06666667,0.0,0.0,0.0,0.0,1.3555555,2.5833337,2.3,3.0079367,4.0333333,3.295238,3.8083339,6.6555557,11.291666,8.977779,8.033334,4.841667,1.7777779,0.48333338,0.24444443,0.3166667,0.34444445,1.8666668,8.766666,5.988889,2.6333334,4.4444447,4.366667,0.93333346,4.425,7.1,6.111111,3.2583332,0.5777778,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05,0.0,0.8000001,2.8333335,3.8222222,0.0,0.0,0.0,0.0,1.6222222,2.725,3.5333335,5.1333337,1.1666666,0.8083334,0.6555556,0.0,0.15555556,0.25555557,1.0166667,4.5111113,11.266667,14.655555,4.775,1.1555556,1.1777779,1.1499999,0.24444446,0.6833334,1.9000001,2.3583333,3.3444443,5.7749996,7.5444446,3.4666667,1.5749999,1.3111112,5.3583336,8.1,18.058332,29.122223,63.5,47.45,49.12222,34.858334,23.11111,23.933334,19.97778,12.433333,5.2166667,0.67777777,0.041666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.033333335,0.16666667,0.125,0.022222223,0.1888889,1.8833334,4.133333,6.041666,1.8,0.025000002,0.42222226,1.6416667,3.3888888,5.7111115,8.424999,0.044444446,0.016666668,0.2,0.99999994,1.3000002,0.25555557,0.058333337,0.9111112,1.75,1.0333334,0.35833335,0.16666667,0.15555556,0.26666668,2.4333334,1.8666668,0.10000001,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06666667,0.32222223,0.7166667,0.7111112,0.36666667,0.108333334,0.0,0.0,0.022222223,0.075,1.6444446,4.783334,4.7666664,4.5319448,6.241667,7.2444444,7.716666,10.344444,10.333333,6.7888894,7.6666665,6.916667,4.0111113,2.35,0.8444445,0.32500002,0.2888889,0.4888889,2.026515,3.2111113,1.2916666,1.0222223,5.4666667,2.4222224,5.0333333,11.311111,12.488888,4.05,0.4666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0375,0.0,0.0,0.00625,0.008333334,0.025,0.0,1.35,1.8000001,2.375,1.2937499,4.35,12.13125,8.966666,3.53125,0.8000001,0.0,0.0,0.0,0.16250001,1.5333334,5.4687505,8.066668,5.8,1.25,0.9083334,0.0,0.058333334,0.21875,1.3916665,0.1875,2.7,6.05,5.591667,3.958333,2.95625,5.958334,18.6875,18.075,20.087502,26.925,36.2,31.825,30.175,23.275002,19.158333,14.393749,8.141666,3.9833336,1.3562499,0.70000005,0.0,0.0,0.0,0.033333335,0.075,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.16666667,0.58124995,0.65833336,0.6875,0.9083333,0.13125,0.12500001,0.59374994,1.4166665,2.5583334,3.2250001,0.8166667,0.075,0.0,0.112500004,0.11666667,0.058333334,0.475,3.1833332,4.65,5.0833335,3.2625,1.2083334,0.57500005,0.09375,0.09166667,0.13125,1.6750001,1.0312501,0.55833334,0.1375,0.275,0.0,0.0,0.0,0.09375,0.38333333,0.575,0.075,0.0,0.0,0.0,0.0,0.025,0.29190478,1.6083333,3.81875,5.991667,5.766667,4.4375,5.95,9.912499,13.741668,13.906251,10.983334,7.575,9.512501,9.249999,4.3375,1.6750001,0.47666666,0.8166666,0.6083334,0.08125,1.4083334,1.31875,1.6,2.3875,10.816667,17.9,37.916668,31.158333,17.86875,4.3916664,0.075,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.008333334,0.13333334,0.17500001,0.0,0.0,2.4,2.2666667,0.17500001,0.13333334,4.9249997,20.877779,15.208335,0.0,0.0,0.0,0.0,0.116666675,0.56666666,0.17500001,0.5555556,1.4749999,0.36666667,0.24444446,0.016666668,0.11111111,1.3833332,3.4888892,0.275,0.35555556,4.0916667,2.788889,0.2777778,11.966668,22.633335,14.533334,10.299999,18.25,21.477777,28.6,18.275,14.888889,11.216667,7.644444,4.703788,2.5888891,1.3888888,0.43333334,0.13333334,0.025,0.0,0.0,0.24444444,0.225,0.0,0.0,0.083333336,0.06666667,0.22500001,0.18888889,0.31666666,0.7222222,0.0,0.0,0.0,0.0,0.5333333,2.6833334,2.3777776,1.0416667,0.3333333,0.0,0.0,0.0,1.45,5.3111115,7.0583334,4.433334,1.7333333,0.20833334,0.06666667,0.5916667,1.3666667,0.9750001,0.7666667,1.0777779,2.0833333,2.2347224,2.5178032,2.386111,0.6166667,1.1333334,0.52500004,0.6888889,0.033333335,0.0,0.0,0.008333334,2.3222222,0.7416667,0.20000002,0.06666667,0.0,0.2888889,0.5274242,2.081389,11.483334,19.21111,11.758333,6.0555563,6.788889,3.9333334,3.222222,4.275,6.3777785,9.683334,9.255555,6.8777776,6.3666663,13.2,11.666667,4.677778,2.8333333,3.0555556,2.7444448,3.025,4.9888887,6.225001,6.188889,4.35,39.044445,46.225,71.76666,94.08888,62.875,13.7,0.7,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.14375,0.0,0.0,0.0,0.05,0.0125,0.025,0.075,1.0,0.88333344,0.0,0.0,0.0,14.966667,17.1375,0.0,0.0,0.0,0.0,0.0,0.008333334,0.0,0.0,0.0375,0.083333336,0.116666675,0.0,0.35,0.98125005,1.2,0.96250004,1.3666667,0.82500005,0.033333335,1.2583334,22.15,17.966667,3.4812503,2.7833333,8.437501,7.133333,5.216666,4.55,6.466666,2.6546211,1.7264069,0.4925,0.39166668,0.25,0.06875,0.0,0.0,0.0,0.0,0.083333336,0.0,0.0,0.0,1.2125,1.2416666,3.7187502,0.53333336,2.1437502,1.4583335,0.0,0.0,0.0,0.54375,6.341667,16.15,17.708334,9.675,3.6833334,1.0166668,0.112500004,0.0,0.75625,3.4916666,6.0625,4.196819,2.025,1.5875001,1.0416667,2.2375,3.0416667,2.0500002,0.9749999,0.43333334,1.4,1.9000001,1.4653409,2.265,2.2625,0.18333334,0.0375,0.15,0.0,0.075,0.28333333,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.50625,7.7916675,12.7325,17.199999,18.78125,12.708334,10.841667,11.200001,10.625001,8.61875,6.3166666,2.7375002,2.3166666,2.5166667,2.9812503,6.375,13.45,13.400001,12.093751,8.208333,4.1666675,2.3875,3.025,5.98125,8.1,12.75625,49.60833,91.76875,126.59167,154.39168,127.006256,40.033333,5.3375,0.050000004,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.67499995,0.0,0.0,0.0,0.033333335,0.22499998,0.13333334,0.0,0.0,0.022222223,0.0,0.0,0.0,0.22222221,4.391667,3.8222225,0.20000002,0.0,0.0,0.0,0.0,0.0,0.22222224,0.27500004,0.0,0.0,0.0,0.13333334,0.9916667,0.044444446,1.2916667,0.5888889,0.7416667,0.044444446,0.2888889,3.525,2.0777779,0.7750001,1.5333334,10.883334,4.388889,3.7861109,0.889394,0.32083333,0.0,0.0,0.05,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0888889,3.8166668,2.2444446,2.3583336,0.0,0.15,0.0,0.0,0.23333335,0.0,2.1333332,13.611111,37.383335,61.600006,39.300003,10.744445,5.2666664,2.8166666,5.944445,3.625,1.8666667,6.1,4.288889,3.838889,6.3410606,4.6444445,1.0583334,0.4180556,0.09166667,0.0,0.0,0.016666668,0.011111111,0.0,0.0,0.0,0.0,0.0,0.8555556,0.82222223,0.67499995,1.8666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.5666666,5.5111117,9.008333,9.466667,10.800001,7.5916677,10.722222,7.0166664,4.288889,4.5666666,0.24444446,0.0,1.7833334,3.2666667,10.408334,12.900002,7.6916666,3.866667,2.3333335,1.075,1.2444445,2.4166667,3.2333336,15.841667,27.511112,61.84167,85.66667,112.44444,111.216675,65.78889,15.983334,0.45555553,0.375,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,3.4624999,0.17500001,0.0,0.0,0.0,1.9875001,0.0,0.0,0.0,0.033333335,0.15625,0.10833334,0.28125,0.45,0.025,0.875,0.71875006,0.0,0.0,0.0,0.0,0.0,0.23333333,0.67499995,0.125,0.099999994,5.70625,7.425,1.2875001,1.4916668,1.31875,1.125,0.89375,1.4083333,1.125,0.51250005,0.041666668,0.025,1.355303,6.728757,0.8208334,0.21666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.74166673,0.0,2.6000001,1.6666667,0.087500006,0.0,0.0,0.0,0.0,0.65625006,0.41666672,5.7375,31.108335,37.987503,27.658335,34.85,23.69167,19.266666,11.4,6.925,7.73125,13.333334,13.762501,10.483334,8.575001,4.896369,4.7855554,5.587143,5.8583336,1.13125,0.2,0.725,3.7375002,2.0166667,0.0625,0.0,0.0,0.0,0.0,0.65,0.60833335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.045,1.3306565,10.108333,21.616665,25.2375,25.375002,24.016668,5.5437503,3.3083334,6.0625005,3.9,3.825,1.225,1.3,4.3125,5.9666667,5.85,5.941667,2.29375,0.625,0.14166668,0.85,0.38333333,0.40625,0.75000006,2.30625,4.158334,30.79375,45.825,53.066666,64.49375,35.949997,13.26875,3.4166667,0.275,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,10.783333,0.4888889,0.15555556,0.1,6.8666673,26.816666,6.4444447,0.0,0.0,0.0,0.06666667,0.011111111,0.9333333,3.8666668,0.41666666,0.7666667,0.9916668,0.0,0.0,0.0,0.0,0.0,0.0,0.5,0.5777778,1.5,10.1,16.98889,1.4916666,1.2222223,2.2583334,3.3222225,4.8083334,4.0,2.3222222,1.5166667,0.36666667,0.7583334,0.011111111,0.11468254,0.2952381,0.0,0.0,0.0,0.008333334,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011111111,0.008333334,0.11111111,0.0,0.8166667,3.666667,0.4666667,0.0,0.0,0.0,0.0,0.17500001,0.98888886,10.725,20.077778,9.766667,9.9777775,21.525,28.0,20.122221,14.583332,4.644445,1.3916667,11.433333,9.549999,1.0888889,3.277778,20.274998,29.886108,7.7916665,1.7777778,0.3,1.9777778,1.0666666,4.633333,0.18888889,0.0,0.0,0.0,0.0,1.4583333,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.4916666,11.166667,16.191666,6.3861113,4.6916676,11.533334,18.141665,30.688889,25.633335,19.608332,8.511112,7.0750003,2.788889,4.2083335,6.6000004,5.088889,14.450002,13.0222225,8.833333,7.711111,4.683333,3.5666668,0.9,0.0,0.0,0.016666668,0.0,0.26666665,0.5666667,10.108334,25.755554,23.3,22.958334,11.877777,1.4250001,0.1,0.025,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.008333334,0.022222223,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,3.5416667,0.0,0.51111114,3.7750003,16.311111,23.125002,4.0777783,0.10833333,0.0,0.0,0.0,0.0,0.0,3.3222222,1.3250002,0.3,0.77500004,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.033333335,0.35555556,1.5333334,7.211111,3.5083334,1.888889,4.0666666,5.833333,6.9,4.577778,3.0111113,1.675,0.0,0.0,0.0,0.0,0.0,0.0,0.24166667,0.14444445,0.016666668,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.0,0.022222223,1.7166667,3.0222225,0.083333336,11.711111,3.2500002,1.2333333,0.23333335,0.0,0.37777779,3.758333,12.388889,1.1416667,4.522222,10.366667,17.08889,5.855555,0.42500004,1.2777778,0.5416666,3.5333333,10.675,4.3,1.9111112,14.858333,23.955557,14.966668,0.0,0.0,0.24444446,0.8333333,1.1500001,0.2,0.0,0.14444445,0.7916667,0.8555556,0.45833334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.3333333,1.9222223,10.108335,26.033333,29.933334,12.169445,19.183332,13.844445,21.849998,30.144444,19.866667,24.066668,7.955556,5.3666663,3.7111113,3.9583335,5.677778,4.8,14.191667,19.755554,21.349998,17.088888,3.8166666,4.5555553,4.5555553,0.15833335,0.0,0.0,0.0,0.0,0.40000004,13.516667,23.733334,23.433334,27.208334,17.377777,4.3916664,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.075,0.17777778,0.12222223,0.05,0.011111111,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13333334,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.35,0.0,0.0,3.1375003,8.016666,7.6375,3.1333334,0.10625,0.0,0.0,0.0,0.0,0.0,0.68333334,0.89375,0.92499995,1.8312501,0.075,0.0,0.0,0.0,0.01875,0.025,0.0,0.0,0.20000002,0.91249996,1.9666668,5.7937503,3.4166665,2.8937502,3.9833333,6.3499994,4.133333,0.91666675,0.26250002,0.0,0.0,0.0,0.0,0.0,0.0,0.375,0.14166668,0.0,0.0,0.0,0.0,0.0,0.00625,0.0,0.0,0.0,0.0,0.0,0.57500005,2.2416668,0.008333334,1.25,1.6916667,0.7375001,0.8916667,0.38125002,0.32500002,0.075,0.0,0.7166667,0.23125,4.616667,2.61875,2.716667,3.95,5.8916664,8.05,5.20625,7.058334,3.2187502,1.6333333,7.825,7.7000003,6.816667,3.53125,4.3999996,0.59999996,2.3750002,0.8625,3.6916666,11.033333,11.49375,8.133332,3.26875,1.7568182,0.5046591,0.8541666,0.0,0.0,0.0,0.9204167,2.3166666,0.17500001,1.1166667,2.6875,1.3180952,1.8742427,4.8770237,8.168679,7.619167,3.0151517,3.2749999,4.675,1.9750001,2.525,3.1166666,4.24375,0.85833335,3.00625,2.9750004,5.7062497,11.650001,10.408333,8.2,9.683333,7.625,8.95,3.9912503,4.324091,2.0083332,1.3499999,0.36666667,0.1375,0.0,0.03125,0.38333333,0.58750004,6.450001,21.108335,38.2125,38.175003,21.8375,1.3666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.5625,1.25,0.85833335,0.23750003,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016666668,0.06250001,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0375,0.05,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,6.5833335,6.455556,6.783334,0.61111116,0.06666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,5.111111,3.3666668,1.2888889,0.14444445,0.075,0.0,0.30000004,0.21111113,0.09166667,0.0,0.0,0.0,1.5,3.6916668,4.4111114,3.2583332,1.5666667,1.5583334,0.41111112,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.1555556,0.0,0.0,1.6333334,1.1500001,0.0,0.0,0.0,0.0,0.0,0.31111112,2.1333334,0.13333334,1.0,3.3222222,9.633334,3.0333333,1.1444445,0.0,0.0,1.9750001,1.2,5.2916665,23.188889,19.699999,7.158334,5.7222223,5.5,8.511112,5.7500005,5.9333334,5.0,5.9833336,13.555555,10.683333,5.15,1.3625542,1.0640874,0.0,0.0,2.2777777,4.941667,8.698414,3.6128788,0.4488889,2.3348486,5.672222,4.943056,1.6939393,1.6819443,2.5499995,1.0291667,0.1,0.0,0.0,0.0,0.20000002,0.8416667,1.0888889,0.44166666,0.93333334,0.0,4.0888886,8.311111,6.758333,8.411112,4.808334,6.0666666,11.516666,9.777779,1.4777778,0.75,1.1666667,0.0,0.0,0.0,0.0,0.0,1.1444445,7.411111,25.224998,36.755554,23.341667,5.5,0.7083333,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.5555556,3.541667,10.566667,5.844444,0.97499996,0.044444446,0.28333333,0.16666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06666667,0.06666667,0.0,0.0,0.0,0.13333334,0.15555556,0.016666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.875,1.5000001,0.7333333,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.3,2.625,0.96875,0.22500001,0.0,0.0,0.0,0.0,0.13333334,0.27500004,0.16666667,0.13749999,5.4833336,6.14375,3.475,0.9666667,2.2250001,4.2166667,7.7750006,1.8000001,0.25,0.18333334,1.8833332,0.4125,0.0,0.72499996,1.2333333,1.1437501,0.083333336,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.8916667,1.0812501,0.0,0.28750002,0.28333333,3.36875,0.0,0.0,4.99375,35.36667,51.26875,4.0,3.29375,8.033334,5.691667,4.1,3.3333335,18.5875,12.425001,6.55,6.8333335,1.8000001,0.39999998,1.4833333,9.4125,3.3416667,2.69375,1.215909,0.09464286,1.3090909,0.0,0.8125,3.125,4.2125,1.2583334,0.50625,2.3212123,2.0510607,0.40666667,0.1,1.15625,0.6,0.3,1.2000002,0.60625005,0.016666668,0.0,0.30625,1.5250001,4.65,4.908334,1.20625,0.49166667,0.7,1.3750001,5.8583336,7.30625,8.408333,4.9812503,5.3507576,4.383333,5.9375,6.7333336,1.6625,0.0,0.0,0.0,0.0,0.26666665,1.8833332,3.1375,8.075001,16.4375,9.133335,2.9562497,0.24166667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.37500003,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.106249996,3.3750002,11.324999,28.0,15.058334,2.7875,0.38333333,1.7625002,1.0749999,0.099999994,0.4,0.14166667,0.09375,0.025,0.59375,0.57500005,0.0,0.0,0.0,0.0,0.0,0.16250002,0.20000003,0.0125,0.008333334,0.043750003,0.025,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.108333334,3.9125001,9.425,10.066667,0.5875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.09166667,0.6333334,7.05,2.6555557,1.5222223,8.458333,10.766665,19.991667,8.255556,2.141667,2.8777778,3.8222222,4.3500004,0.7444444,0.058333337,0.044444446,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,7.6416664,13.48889,2.65,0.0,0.16666667,11.200001,43.655556,72.81667,2.6000001,1.2,0.0,0.0,1.6833335,0.0,9.583334,4.788889,6.55,7.5999994,4.1,2.1916668,0.53333336,0.025000002,0.033333335,0.2916667,0.17222223,3.625758,6.4125,0.0,0.0,0.0,0.0,0.22222222,0.16666667,2.6222224,3.388889,2.051515,1.1444445,0.65,0.0,0.40000004,0.8000001,0.28333336,0.0,0.0,0.0,3.1555557,9.708334,7.6555557,3.575,2.0777779,2.5222225,1.6166667,0.57777774,3.9500003,3.9,7.7583337,7.484722,12.215277,16.80606,23.400002,7.466667,2.9333334,0.5,0.0,0.0,0.07777777,1.6333333,3.7833335,8.755555,10.683334,8.044444,4.575,2.0222223,1.3333333,0.6666667,0.0,0.0,0.0,0.0,0.0,1.2916666,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.18888889,1.3166666,9.688889,23.708336,41.866665,23.666668,7.166667,3.0777779,2.8666668,1.8000001,1.6166667,1.5555556,1.4111111,0.9583333,0.67777777,1.8583332,2.0222223,1.175,0.6,0.22222224,0.116666675,0.011111111,0.0,0.0,0.0,0.0,0.05,0.022222223,0.0,0.0,0.0,0.0,0.0,0.23333333,0.12222222,0.36666667,0.275,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.5222222,5.6000004,13.7,17.099998,5.1666665,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.40625,0.9166667,0.89166665,5.00625,11.016666,13.49375,11.708334,6.8375006,5.9249997,12.783333,23.452084,18.991669,3.4499998,0.008333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.075,0.70000005,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.88124996,2.1333334,0.0,0.0,0.0,0.58125,0.28333333,0.0,0.0,0.0,0.0,0.0,0.0,1.7583333,2.28125,0.0,5.7437506,1.875,2.5,3.0062501,0.0,0.0,0.36666664,0.65,0.925,0.28333336,0.8643939,0.18888889,0.22756413,0.0,0.3125,1.0833334,0.5327381,2.8959093,4.5,4.125,6.0492425,1.425,0.0,3.675,2.0,0.0,0.0,0.0,1.7437501,6.1666665,5.6625,9.966667,9.58125,12.791667,5.183333,1.1125001,0.3,4.60625,10.558334,7.998333,10.708333,23.557577,35.51875,42.175003,12.950892,3.6833334,2.0625,0.4,0.15,0.0,0.275,3.3000002,6.8250003,9.706249,10.616668,7.6625004,7.4583335,1.7750001,1.30625,0.0,0.0,0.0,0.025,0.0,0.22500001,0.20000002,0.30833334,0.15,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.31666666,3.06875,17.183332,39.59375,44.474995,27.85,17.1625,13.699999,5.75625,4.7083335,12.175001,10.466667,9.475,6.9437504,4.4750004,3.8125002,3.925,4.2562504,3.8666668,1.4583335,0.53125006,0.14166667,0.10625,0.22500002,0.31875002,0.058333337,0.043750003,0.041666668,0.0,0.0,0.0,0.0375,0.025,0.325,0.46666667,0.39166668,0.59374994,0.6666666,0.29999995,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,4.7749996,11.516666,10.291667,5.3625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06666667,0.08888889,0.0,0.49166667,3.8111115,7.008333,11.722222,4.6500006,3.3777776,6.211111,17.475,9.344445,0.55,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,4.758333,0.0,0.0,0.0,2.8749998,3.9555557,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.044444446,0.1019192,1.1888889,2.275,8.744444,6.4888887,2.8504043,6.276389,9.630357,2.648016,3.9583335,5.381944,5.7583337,5.0249996,8.0222225,4.0333333,1.2666667,1.8000002,2.2666667,1.3833333,0.16666667,0.34444445,10.241667,12.511112,9.016667,10.6,13.258333,7.988889,2.188889,5.241667,1.288889,2.3166666,7.355556,6.4000006,3.5555558,5.055556,9.800002,10.922223,8.558334,4.4333334,2.7083335,5.8555555,0.7416667,0.0,0.0,0.34166667,6.1222224,14.283334,17.444443,15.883334,13.01111,7.7555556,5.3250003,0.14444445,1.4916667,0.22222224,0.6333333,0.0,0.050000004,0.48888892,0.9,0.40000004,0.0,0.0,0.0,0.0,0.033333335,0.1,0.041666668,0.055555556,0.0,0.26666668,3.8166668,21.244446,50.891674,43.13333,32.9,30.366669,30.277779,11.858334,9.4,25.358334,26.133335,27.077778,27.858335,21.61111,14.799999,10.288889,12.5,12.988889,4.7000003,2.975,2.777778,2.075,0.95555556,0.9083333,0.13333333,0.025000002,0.033333335,0.0,0.0,0.0,0.0,0.0,0.70833325,0.5888889,0.16666667,0.008333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.041666668,0.06666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.008333334,0.033333335,0.17500001,0.68888885,1.0111111,0.4916667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.5,0.6,0.0,1.2,0.40000004,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01875,0.33333334,4.8,23.041666,9.5,2.466667,1.7083335,2.0875,7.641667,3.8062503,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0375,3.5583334,0.8249999,0.0,0.0,0.0,0.0,0.0,0.0,0.16875,1.2249999,4.0583334,4.03125,0.23333335,0.0,0.0,0.08125,0.325,0.20833334,0.0,0.0,0.0,0.0,0.01875,0.0,0.0,0.0,0.0,0.0,0.0,0.0375,0.5683983,1.9542208,2.5439396,3.132222,4.435,3.5583334,4.9178934,1.2358333,6.32375,7.8949995,3.2333333,1.5875,13.508333,6.575,5.7305555,1.4864287,0.61666673,1.425,5.3250003,10.816668,54.256256,57.883335,13.2875,7.583334,6.40625,8.066667,4.3083334,2.59375,2.9083333,2.05,4.0000005,1.68125,4.4500003,3.6166663,4.04375,9.833333,8.193749,10.108333,6.5687504,2.775,0.76875,0.0,0.0,0.0,0.40833336,5.5625005,13.541666,16.1,16.900002,14.925,6.49375,10.516666,15.031249,5.9583335,1.1624999,0.35000002,0.84375006,0.55,0.06666667,0.0125,0.0,0.21875,0.47500002,0.6125,1.4083334,2.6333332,1.34375,1.4583333,0.5,0.48333335,4.1062503,21.058334,49.137497,36.3,25.100002,29.175,38.666668,23.8625,21.983334,32.75625,30.333332,38.35,55.074997,54.833332,41.831253,37.074997,31.86875,21.416666,12.316668,12.018751,13.891666,8.45625,2.8000002,1.08125,0.36666664,0.10625001,0.0,0.0,0.275,1.0,0.9375,1.0916667,1.59375,1.1,0.65,0.46250004,0.5916667,0.47500002,0.38333333,0.34375,0.26666668,0.275,0.075,0.008333334,0.04375,0.125,0.16875002,0.14166668,0.0375,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.008333334,0.15,0.23333335,0.075,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01875,0.108333334,0.14999999,0.075,0.0375,0.008333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.75,0.0,1.3111112,1.9666667,0.0,0.0,0.0,0.0,0.0,0.0,1.2,0.40000004,0.0,0.0,0.0,0.0,0.5,4.422222,1.8666668,0.016666668,0.0,4.4666667,32.833336,23.091667,5.077778,0.95555556,0.4916667,0.0,0.0,0.0,0.0,0.0,1.9083333,1.5888889,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.3333333,0.82222223,0.083333336,0.0,0.0,0.0,0.0,0.0,1.2916667,1.8111113,4.4666667,4.508333,1.3000001,0.0,0.0,0.0,0.10000001,1.1,2.8833334,1.5333334,0.20000002,0.13333334,1.2083335,3.3666668,0.26587301,0.108333334,0.35555556,0.5555556,0.32420635,0.5924243,2.1055555,1.6916666,1.8222222,1.2111111,2.15,0.0,0.19,0.22222224,2.625,4.1888885,2.4301589,1.95,4.8333335,6.3500004,6.8777776,5.0666666,7.1,7.5833335,33.4,25.211111,34.141666,52.43333,29.300001,9.355556,8.408334,11.244445,10.6,5.366667,5.7333336,6.3833337,4.0666666,4.55,8.222222,8.377778,7.5916667,7.533334,13.425001,15.4,7.3999996,5.577778,3.6000001,0.0,0.0,0.0,0.0,0.5416667,4.0555553,9.191667,13.822223,17.188889,11.125,18.1,23.808334,16.266666,0.9083333,0.0,0.625,0.47777778,0.0,0.0,0.06666667,0.425,0.33333334,0.47500002,0.6555555,1.4444444,0.7583334,2.8666668,2.7416666,1.3000001,6.0,20.922222,44.749996,24.38889,21.855556,27.45,47.444443,41.208332,30.333332,33.883335,25.977777,20.366667,52.674995,54.655556,53.966663,48.31111,44.149998,32.82222,28.866669,28.475,22.9,16.183332,8.266667,2.916667,2.6222222,3.1666667,3.5000002,2.877778,2.8166668,3.0555556,3.2916667,4.9333334,5.925,4.5111113,3.5,2.5750003,2.2444444,2.2833333,2.288889,2.2833335,2.1111112,1.45,0.7888888,0.6444444,0.5166667,0.3111111,0.35000002,0.37777776,0.6333333,0.26666668,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.058333334,0.8111112,1.4583334,1.4444444,1.7166667,1.3555555,0.9,0.36666667,0.12222222,0.025,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.1666665,0.44444448,0.13333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,5.55,17.822222,23.6,1.9999999,0.0,0.0,0.75555557,3.666667,2.5333333,0.8222223,2.05,0.0,0.0,0.0,0.0,0.0,0.041666668,0.011111111,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.275,0.12222222,0.0,0.0,0.0,0.0,0.075,0.32222223,0.5222222,0.34166667,0.06666667,0.0,0.06666667,1.2916666,0.22222224,0.0,2.8333335,4.966666,1.5416667,0.8888889,0.49166664,2.3111112,1.2111111,0.90000004,1.7291667,1.8499999,0.4,0.42500004,0.011111111,0.35833335,0.2777778,0.022222223,0.0,0.0,0.0,0.0,0.036363635,0.84444445,2.6333334,0.1,1.1111112,0.83333325,2.777778,2.7333333,5.688889,3.6750002,9.633334,1.388889,5.6666665,18.066668,11.15,6.977778,10.375,10.666667,18.844444,10.958333,12.766665,12.374998,6.288889,1.1166667,3.4888892,5.3333335,11.133334,13.677777,13.691668,9.966667,3.6916666,4.455556,2.3916667,0.0,0.0,0.0,0.0,0.0,0.2,5.4666667,9.677778,14.233332,15.166667,13.544445,23.675,19.988892,3.2083335,2.0444443,2.266667,2.1111112,1.1777778,2.7666667,2.1666667,0.81666666,1.1666667,0.225,0.43333334,0.26666668,0.53333336,3.4333334,7.0,7.322222,11.991667,23.022223,38.850006,44.11111,23.655558,29.725,47.18889,41.633335,33.011112,32.625,23.1,12.377779,29.475002,30.200003,33.74167,35.22222,34.675,30.399996,31.011112,25.450003,25.68889,29.483332,31.83333,31.591667,22.300001,12.300001,6.077778,5.5444446,3.5833333,4.2999997,4.5166664,5.6444445,6.3166666,5.622222,4.8555555,4.308334,2.944445,2.325,1.9666667,2.5083334,2.1555557,1.6083333,1.1,0.8888889,1.4916668,1.0,1.9166666,2.911111,4.8250003,3.2222223,1.2222223,0.6166667,0.48888892,0.5083333,0.7777778,0.60833335,0.35555556,0.18888889,0.18333334,0.6333333,0.725,0.57777774,0.9916667,0.8333333,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06666667,0.044444446,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.09166667,0.51111114,0.74999994,0.65555555,2.9000003,4.111111,2.7833333,1.3111112,0.3777778,0.09166667,0.044444446,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,10.50625,2.05,0.9333334,1.15,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,4.3437495,18.783333,24.733334,8.71875,0.0,0.0375,0.025000002,0.61875,0.0,0.008333334,0.3375,0.0,0.0,0.0,0.0,0.0,0.0,0.016666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.050000004,2.01875,0.40000004,0.0,1.36875,1.7916667,0.24208334,0.0,0.058750004,0.28030303,4.9416666,7.725,5.200001,4.4812503,5.241667,7.70625,6.483333,3.7875001,3.3500001,1.25,0.0,0.0,0.0,0.0,0.17500001,0.5939394,3.8704548,6.10625,3.5749998,1.3589286,0.71666664,0.725,3.1833336,3.7,4.383333,6.0083337,3.2062502,3.591667,7.1875,6.2333336,5.2437506,6.4416666,13.566668,22.612501,14.625001,6.6812496,3.4,0.24375002,4.2083335,10.825001,13.94375,7.45,4.5125,11.3,4.8062496,1.4250001,0.73125,0.16666669,0.26666668,0.17500001,0.0,0.0,0.0,0.9062501,3.4250004,6.6499996,10.5375,12.474999,14.706249,14.5,11.012501,7.025,9.243751,9.008333,6.966666,3.5499997,2.5416667,2.54375,3.0583334,1.46875,0.7416667,1.2833333,2.13125,6.858333,10.93125,16.475,13.206251,20.1,25.3375,53.11667,23.725,33.78125,35.416668,32.31875,30.824999,28.606247,23.150002,11.116667,12.525,12.424999,11.93125,12.65,14.887501,16.316668,16.066666,23.375,37.241665,49.70625,48.608334,42.45,32.4,22.31875,20.591665,22.1,23.2125,18.475,10.9,8.716666,12.099999,15.391666,16.725,18.050001,16.8,13.925,12.675001,11.143751,12.658333,9.95625,8.9,10.608334,11.556251,12.883334,14.1,17.25,17.4875,16.824999,12.891667,8.8625,7.3250003,4.34375,5.3583336,6.1500006,4.05,6.7250004,6.4937506,4.2250004,2.4875,2.5416665,3.8125002,4.825,3.66875,1.8750001,1.5916666,0.44375002,0.016666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0125,0.0,0.0,0.0,1.6750002,3.6833334,3.3374999,1.675,0.21666667,0.01875,0.058333337,0.0,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,7.75,13.477779,13.933333,2.666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,7.0666676,7.6916666,0.0,2.0583334,10.411112,13.177777,4.3333335,0.0,0.45000005,0.67777777,1.1833334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,3.0777779,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.041666668,0.12222223,0.016666668,0.06666667,2.1777778,4.391667,3.7555556,1.8533335,0.02777778,4.608333,6.2222223,2.455556,6.325,7.8777776,6.283334,13.433334,16.416666,15.722223,23.675003,17.044445,5.1444445,0.0,0.6777778,0.0,1.7402779,1.8338889,1.2222223,8.177778,13.542424,6.1914682,5.215152,2.3,6.4583335,11.311111,13.258334,16.08889,22.022223,9.433333,0.93333334,0.0,1.2444444,3.9000003,1.9444444,1.0222223,4.9500003,8.0,3.9666667,0.0,0.18333334,0.40000004,0.47777778,1.0666666,0.3888889,0.0,6.3333335,1.9333332,0.31111112,0.9666666,1.2888889,0.6666667,0.0,0.0,0.0,0.0,0.0,0.57777774,2.277778,7.8833327,7.266667,8.191667,13.088888,13.5,9.111112,10.466667,11.033334,10.233334,5.6,4.7444444,5.0583334,3.4444447,0.80833334,1.2222222,2.911111,3.6083333,8.766666,10.166666,15.299999,6.858333,8.522223,30.141666,44.033337,23.177778,39.175003,34.61111,30.483334,29.588886,25.575,21.111115,15.022224,9.666667,6.833333,5.383333,7.2222233,8.816668,13.277779,22.844444,34.691666,45.066666,53.55,57.022224,58.691666,49.966667,39.350002,39.85556,42.422222,40.7,30.966667,17.816666,11.988888,12.291667,17.022223,18.9,20.683334,20.255554,18.558336,18.911112,17.425,17.522223,16.141668,16.688889,18.466667,24.358334,28.466667,30.783335,26.6,25.933334,27.011112,27.822224,27.483334,25.611113,22.866669,19.6,18.2,17.4,18.077778,20.058332,19.133335,15.650002,13.744445,15.3,15.411111,14.866667,11.688889,8.144444,3.6583333,0.0,0.13333334,0.22222222,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.6111111,0.53333336,0.05555556,0.22500001,0.2,0.06666667,0.1,0.9111111,1.2333332,0.7222222,0.39166668,0.18888889,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,28.675,31.075,17.016666,1.36875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.2916667,4.24375,3.333333,9.456249,6.525,2.4666667,0.0,0.0,0.7125001,0.94166666,0.25625002,0.41666666,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.89166665,0.0,0.0,0.0,0.0,0.0,2.475,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.081250004,0.44166666,0.17500001,0.0,1.6666667,3.3187504,0.59999996,0.9875,1.9500002,1.8562499,2.9833336,0.9333334,1.7875,2.175,2.11875,14.308334,4.4375005,9.866667,12.64375,3.7333336,3.4750001,0.49999997,0.0,0.0,0.38333333,1.0250001,0.0,3.625,5.4875,1.2916667,0.7937499,1.4674243,6.3312507,14.708334,17.800001,14.316667,10.508334,10.0,7.883333,1.85,0.0,0.4,0.40000004,0.5333333,2.3249998,1.1666666,0.86249995,0.26666668,0.2,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.31875002,0.33333337,0.0,0.0,0.0,0.0625,0.083333336,0.53125,1.1916667,1.7916666,2.275,5.1916666,7.58125,8.766666,9.4625,7.483333,9.15,8.25,6.316667,6.6875005,9.508334,8.9875,4.641667,1.8375,2.233333,1.4416667,2.08125,10.408335,9.64375,13.541667,4.525,11.283334,21.943754,22.125,26.958332,44.875,36.183334,37.99375,38.100002,29.612501,20.758337,18.95,12.20625,9.058333,11.275001,16.708334,15.968751,15.975,25.733334,36.124996,44.55834,47.199997,50.69167,49.73125,44.633335,39.10625,38.358334,39.11667,40.13125,27.2,19.3375,15.875,14.968751,15.791667,16.199999,15.5375,15.066667,14.931251,17.316668,20.44375,23.933334,28.98125,32.708332,33.9,36.33125,42.108334,47.96875,51.750004,44.875,39.216667,44.91667,50.4875,53.058334,52.35,47.50833,39.90625,34.60833,36.666664,39.68125,42.858337,37.23125,36.425,37.88125,33.06667,26.600002,19.958332,15.45,11.8625,8.349999,4.53125,1.5500001,0.00625,0.108333334,0.14166667,0.03125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.3125,1.1833334,0.0,0.0,0.075,0.15,0.016666668,0.14375,1.6833332,3.20625,2.5666666,1.4374999,1.0083333,0.2,0.025,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05,17.183334,11.011111,2.1666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.022222223,1.6000001,6.9999995,9.550001,4.633333,0.5,0.016666668,0.9333334,1.3666667,1.3666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.51111114,0.65833336,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.22500001,0.7,4.3416667,8.211111,3.0416665,0.044444446,0.5777778,4.9166665,4.6,1.3916667,14.233334,43.975,29.1,12.258332,4.422222,4.2000003,2.4500003,0.0,0.0,0.0,2.6666667,4.444444,0.88888884,0.0,0.0,3.0600002,0.3,0.7448485,5.744445,14.208334,8.4777775,2.5666666,4.3083334,4.688889,10.333333,0.0,0.0,0.0,0.0,2.2749999,5.422222,2.6999998,0.48888892,1.15,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.041666668,0.22222222,0.20833333,0.5666667,0.6666667,1.6333334,3.1555557,3.6333334,4.1444445,5.2,3.0555558,3.2500002,4.111111,3.5333333,7.016667,11.044445,10.941667,6.544445,6.6499996,6.7000003,8.400001,11.525002,12.155555,10.058333,14.711112,7.5749993,10.422223,13.549999,25.833334,39.13333,41.85,29.455557,30.116669,36.155556,27.100002,18.955557,16.677778,11.075001,11.144445,8.741666,8.900001,6.666667,6.755555,9.733334,10.558333,12.555554,18.55,22.566668,17.558334,17.500002,24.641666,30.68889,36.044445,37.733334,30.366667,29.533335,23.244446,25.683334,26.544447,27.544443,27.575,29.166668,33.3,43.98889,55.941666,68.78889,79.208336,88.0,95.255554,95.09167,91.433334,88.0,82.08889,72.78334,62.377777,67.56667,75.10834,77.67778,74.64167,70.82223,58.283333,50.000004,46.18889,46.875,55.13333,60.791664,59.32222,48.966667,43.944443,37.083332,32.066666,27.81111,21.358334,14.844445,8.225,3.588889,1.0250001,1.0,0.67777777,0.15833336,0.08888889,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.75555557,2.25,0.21111111,0.0,0.0,0.0,0.0,0.0,0.12500001,0.23333332,1.3666667,2.1666667,1.3583333,0.6888889,0.5444445,0.041666668,0.0,0.0,0.0,0.033333335,0.0,0.0,0.0,0.0,0.0,0.13333334,0.27500004,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.35,1.05,1.0875,1.0000001,2.84375,4.733333,5.066667,1.8678571,1.1416667,1.3312501,0.20000002,0.0,0.0,0.0,0.0,0.10000001,0.0,0.0,0.0,0.20000002,0.15,0.43333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.90625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.075,0.6,1.5,0.0,0.0,0.0,0.0,0.0,0.0,0.88125,0.625,0.0,0.0,0.0,0.0,0.48787883,1.3687501,1.4250001,1.38125,7.275,10.549999,7.6,0.058333337,2.7562501,13.799999,32.35,17.975,4.125,0.07878788,0.0,0.84375,2.25,0.5625,0.5500001,0.3375,0.31666666,0.8,0.20208335,0.0,0.0,0.0,0.125,2.025,2.5875,0.125,1.9583333,4.9500003,4.4166665,3.0125,0.7166667,0.6,0.3,0.7,1.5187501,1.8083335,0.175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.043750003,0.058333334,0.13125001,0.45,0.65,0.675,0.57500005,0.8249999,1.1083333,4.3187504,7.566667,8.96875,9.291667,12.656249,16.65,22.766665,21.406252,19.5,20.737501,20.816666,17.487501,15.95,18.2375,22.466667,25.466665,21.53125,19.508333,23.0125,18.09167,13.743751,11.883334,13.124999,10.44375,9.541667,7.8749995,6.65,5.8625,5.441667,4.25,3.84375,2.875,3.8687503,8.316667,14.187501,19.825003,19.425,24.741667,31.058334,36.15,40.083336,42.7625,32.741665,31.40625,23.975,22.6,21.743752,32.316666,42.631252,50.258335,65.65,83.816666,96.075,104.375,108.325,110.04375,103.350006,97.75,90.175,82.875,76.68333,77.75,83.15625,85.274994,81.087494,73.625,63.175007,54.16667,52.46667,56.84375,65.86667,74.4,67.02501,52.05625,44.008335,41.381252,37.375,36.041664,29.418749,18.824999,13.49375,10.316667,3.48125,1.7500001,1.2416667,0.76875,0.50000006,0.39375,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.48750004,1.4666668,0.15625,0.0,0.0,0.0,0.0,0.06666667,1.9083335,0.63125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.108333334,0.14999999,0.0,0.0,0.0,0.0,0.075,0.32500002,0.28125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.5083334,3.2444444,6.625,4.6000004,0.13333334,0.67777777,3.022222,5.25,1.9222223,0.275,0.0,0.0,0.0,0.0,0.0,0.13333334,0.0,0.0,0.116666675,0.0,0.0,0.5555556,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.25833333,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.7416668,0.0,0.2,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,5.1,10.6888895,14.600001,10.533334,2.5333333,2.0500002,5.9555554,7.891667,14.1444435,7.15,2.711111,0.0,0.0,0.0,0.75,0.0,0.24166667,3.1000001,4.1,0.30833334,0.0,0.0,0.0,0.0,0.033333335,0.29999998,0.4,0.0,0.0,1.3333333,0.0,0.53333336,0.70000005,0.4666667,0.5555556,4.8416667,3.2444444,0.175,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.20833334,0.16666667,0.0,0.06666667,0.42222223,2.0833335,2.4444444,3.833334,6.7333336,9.883333,13.066668,15.444444,17.941666,18.322224,18.958336,18.98889,19.333334,19.166666,16.891666,13.388889,12.422222,11.983335,14.0,14.3916645,10.433332,8.85,9.5,9.788889,8.825001,7.288889,5.7916665,4.7555556,5.5499997,5.788889,8.8555565,7.8083334,9.1,10.091666,13.944445,17.541668,14.755557,21.375,22.47778,22.011112,21.850002,28.366667,18.883335,25.644445,18.15,14.41111,14.166666,16.041666,25.177778,38.24167,57.155552,70.89167,78.94444,88.98334,93.78889,92.33333,93.725,93.53334,93.35834,90.299995,85.208336,82.27778,79.87778,76.78333,72.744446,66.558334,62.31111,59.233337,56.65556,62.355553,73.99167,68.8,55.433334,47.566666,37.875,28.466667,23.183334,22.055557,23.200003,24.09167,17.577778,14.766666,13.222223,6.408334,7.5000005,6.9555554,3.5916662,3.0555556,2.0916667,0.08888889,0.016666668,0.022222223,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.022222223,0.45833337,0.055555556,0.0,0.0,0.0,0.0,0.46666667,1.6777778,1.1444445,0.0,0.0,0.0,0.0,0.0,0.07777777,0.0,0.0,0.0,0.0,0.17777778,0.025,0.14444445,0.22222222,0.0,0.0,0.23333335,0.30000004,0.375,0.0,0.0,0.0,0.0,0.0,0.3416667,0.0,0.0,0.0,0.0,3.3250003,7.077778,3.1,13.011111,8.1,3.5777779,0.0,4.0,3.5333333,1.675,0.0,0.0,0.0,0.2,0.0,0.0,0.0,0.0,0.0,0.0,0.23333335,0.17777778,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.6888889,0.51666665,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.62222224,0.9666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.5999999,1.9444444,2.4,0.9888889,1.1166667,3.4111114,2.5833335,5.611111,6.5249996,5.5777774,0.6333334,0.85833335,0.011111111,0.0,0.0,0.016666668,1.0888889,1.6666669,0.0,0.0,0.0,0.25555557,5.0249996,7.9,17.408335,2.5888891,0.0,0.0,0.79999995,0.5,1.9555557,0.2,0.48888892,1.4555557,3.3333333,5.0444446,0.81666666,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.033333335,0.49999997,0.075,0.3111111,0.725,2.1222224,4.375,6.411112,6.4888887,7.750001,9.833334,12.341667,12.511112,11.916667,13.366668,11.124999,11.511111,10.033334,9.6,9.3555565,11.066667,9.477778,10.825,8.566667,7.333333,6.0833335,4.922222,4.7000003,5.9666667,5.4500003,5.3,7.3111115,7.666666,8.744445,12.691667,14.322223,15.308333,18.755558,23.791666,22.044445,24.066666,16.133333,22.98889,17.558332,15.388891,12.716667,15.322223,15.755557,20.516668,27.21111,39.433334,47.36667,52.925003,57.466667,63.083336,68.05556,67.488884,65.5,62.73333,62.833336,63.04445,60.816666,56.3,53.855556,54.475,56.28889,56.783337,59.81111,64.01666,69.22222,70.46667,78.433334,79.67779,59.15,44.777775,37.433334,24.266668,19.533335,15.48889,15.388889,18.233334,14.511112,13.900001,13.511111,9.266667,11.655556,11.222223,8.383334,7.4555554,6.083333,2.4333332,1.6500001,0.11111112,0.008333334,0.0,0.011111111,0.0,0.0,0.0,0.0,0.016666668,0.0,0.0,0.025,0.0,0.0,0.0,0.0,0.0,0.24166667,0.033333335,0.0,0.0,0.0,0.0,0.0,0.20833333,0.0,0.0,0.0,0.0,0.016666668,0.0,0.016666668,0.5222222,0.12222222,0.0,0.06666667,0.27500004,0.17777778,0.1,2.54375,0.2916667,1.4977274,0.05,3.0750003,3.6874998,5.1416664,1.15,4.2,6.7666664,6.7624993,20.256664,9.375,12.191666,3.1237502,1.2499999,0.20625001,2.3484848,1.1212121,2.375,1.1,0.25625002,0.0,0.075,0.0,0.0,0.0,0.15,1.28125,0.5333333,0.0,1.125,1.73125,2.0416667,1.5416667,0.775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.6333333,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.7083334,4.94375,0.0,0.23750001,0.050000004,0.15625,0.23333335,0.17500001,0.98749995,1.7416667,1.975,0.85,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.9312499,7.508333,11.85625,9.016666,6.0500007,7.1583333,6.6499996,7.0833335,11.858334,14.306251,11.658334,5.83125,1.7939395,0.78124994,0.35833335,0.13333334,0.0,0.0,0.025,0.8386364,2.8750002,3.8000002,2.6875,1.5833333,4.65,3.8125,6.833334,7.1250005,3.575,2.7562501,0.65,0.06666667,0.6,2.7333333,2.225,1.3583333,0.1375,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.16250001,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.041666668,0.03125,0.15,0.21875,0.47500005,1.275,2.3999999,4.4250007,4.7062497,4.4166665,4.7500005,4.7583337,3.9187503,4.841666,6.9500003,5.34375,4.7166667,6.593749,6.341667,6.6875,5.0416665,3.1333334,2.06875,2.7416668,5.21875,5.6916666,2.8249998,2.4083333,3.4833333,3.15,3.0,5.2187495,7.7000012,7.58125,9.491667,12.8625,13.941666,13.691667,14.4375,16.291668,16.962502,19.216665,25.631248,28.783335,31.800001,41.0,44.39167,45.631252,44.94167,45.462505,48.158333,48.90625,48.375,44.941666,42.98125,39.86667,39.7875,40.866665,41.59375,43.208336,45.725002,44.59375,42.891666,46.06875,52.508335,55.3125,58.21667,61.075,67.381256,70.083336,66.04375,60.466663,57.062504,46.458336,41.88125,37.075,32.275,28.862503,24.899998,21.05,17.058334,14.725001,14.366666,14.258333,14.30625,12.725,11.9625,10.183333,5.8812494,1.8916668,0.85625005,1.0,0.4166667,0.23750004,0.34166667,0.34375,0.32500005,0.22500002,0.050000004,0.05,0.1875,0.3,0.16874999,0.074999996,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05,0.075,0.0625,0.0,0.0,0.0,0.008333334,0.15,0.6166667,0.82500005,0.25833336,0.06666667,0.15625001,0.25833336,0.09375001,0.016666668,0.0,1.3,2.9666667,4.3366666,0.9333333,5.633333,3.8,0.0,0.075,2.2583332,9.938889,7.8021536,12.853453,3.525,4.4874997,3.2616668,4.133333,1.8000002,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.033333335,1.2204545,0.0,0.9583333,0.6666667,0.2916667,0.0,0.34444445,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.0916667,0.055555556,0.0,0.16666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.175,2.788889,2.125,0.06666667,0.375,1.5444444,1.4666667,0.0,0.5,0.9750001,0.76666665,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.3,1.7333333,4.588889,7.966667,7.288889,4.025,3.4444444,3.2,4.208333,6.611111,4.2416663,2.511111,2.75,2.4555554,1.4777778,0.43333334,0.0,0.0,0.0,0.0,0.0,0.0,2.288889,7.366667,7.3166666,4.1666665,2.5583334,1.9333334,0.37500003,0.0,0.44444448,2.45,4.822222,3.625,2.6555557,0.975,0.044444446,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.75000006,1.511111,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14444445,0.56666666,0.7916667,0.16666667,0.15833333,0.16666667,0.24166667,0.88888896,2.9416668,2.6444445,3.4111114,2.3249998,1.4,1.6083333,0.6888889,0.9000001,0.62222224,0.8888889,1.7583334,2.4666665,2.05,1.2,0.725,1.1,1.7555555,0.9000001,0.2888889,0.5583334,1.6111112,2.325,4.211111,6.116667,7.066667,8.333333,11.366667,17.955557,21.233335,20.288889,21.525,27.655558,36.63333,46.00834,44.755554,39.550003,36.311115,35.283333,36.322224,36.21667,34.5,31.655556,28.533333,26.433334,23.15,21.288889,19.858332,19.88889,20.900002,23.783335,27.811111,31.616667,37.166664,39.61667,40.58889,44.155556,49.108334,55.17778,59.316666,56.444447,58.125,57.41111,58.60833,59.988888,55.911106,49.466667,43.055557,35.916668,27.222223,20.625,18.833332,16.711113,16.9,18.733334,18.099998,18.777777,15.15,10.888888,6.4833345,3.188889,1.688889,1.8333334,1.9777778,1.5333333,1.6444445,1.8583333,1.8777779,2.4666667,3.2250004,2.8444445,1.3833334,0.43333334,0.025,0.0,0.0,0.0,0.0,0.0,0.07777778,0.09166667,0.011111111,0.0,0.0,0.0,0.0,0.22222222,0.95000005,1.6,0.98333335,0.36666664,0.3888889,0.43333337,0.022222223,0.0,0.0,0.18333334,0.225,0.98333335,0.3416667,0.57125,0.31060606,0.555,1.7083335,0.1625,1.7972223,1.15,0.0,1.3486363,0.85309064,0.5,1.3125,6.608333,3.8937502,1.3833333,0.0,0.0,1.8,0.61875004,0.225,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.17500001,0.4375,0.0,1.3916667,0.0,0.0,0.0,0.0,0.0,0.0,0.15833333,1.36875,0.68333334,0.09375,0.7083333,0.09375,0.375,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.175,0.39374998,0.0,0.0,0.0,0.0,0.1375,0.5166667,0.21875,0.7166667,0.125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016666668,0.375,1.1486363,1.875,4.2250004,6.5750003,4.4000006,1.3668182,0.87916666,0.41666666,0.99375004,1.8962122,3.8812501,4.1916666,2.5416667,0.63124996,0.025000002,0.0,0.0,0.0,0.0,0.0,0.95000005,1.425,0.09375,0.083333336,0.4625,0.058333334,0.0,0.18333334,0.51666665,0.40000004,0.24166669,0.7625,0.8333334,0.3125,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.19166668,0.275,0.0,0.0,0.15625,0.36666667,0.46249998,0.625,0.65625,0.35000002,0.3,0.20625001,0.008333334,0.1125,0.29166666,0.45624998,0.59999996,0.8916667,1.1625,0.84166664,1.26875,1.05,0.53749996,0.6916667,0.6666667,0.46875,0.64166665,0.51250005,0.7083333,1.16875,2.025,2.4812498,2.8083334,3.7583334,4.625,6.8666673,9.0625,10.25,10.90625,12.550001,16.675,23.1375,23.841671,20.349998,16.916668,18.112501,21.491667,23.06875,22.866665,21.500004,18.706253,16.133333,14.73125,11.466667,9.88125,10.349999,12.341666,14.524999,16.366667,17.925001,21.641665,24.318748,26.558332,30.508333,37.562504,47.933334,57.518753,66.083336,65.043755,62.666668,63.29375,68.825005,69.274994,63.268753,56.69167,47.6375,38.241673,29.38125,23.308334,19.75,19.4875,21.716667,23.65625,24.775002,26.61875,25.891666,21.05625,14.6,8.291666,5.4874997,4.775,5.3187494,5.7916675,5.7937503,3.6666667,2.3416667,4.3937507,9.083333,10.743751,7.3750005,3.275,0.61666673,0.0,0.0,0.0,0.01875,0.033333335,0.0,0.0,0.0,0.0,0.016666668,0.1,0.4,0.66250014,0.625,0.83124995,0.52500004,0.2,0.09375,0.0,0.0,0.3,0.17500001,0.8666666,0.0,0.0,0.0,1.1111112,0.0,0.0,0.0,0.0,0.0,2.0044446,3.9611113,4.4958334,9.445833,7.437778,4.688889,1.4416667,0.3222222,0.0,0.0,0.6097222,0.25,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13333333,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.325,0.0,0.0,0.0,0.0,0.0,0.0,0.025000002,0.24444443,1.7416668,1.6888889,0.6583333,0.06666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.008333334,0.05555556,0.4378788,1.1222222,1.7458333,3.1476188,3.3113098,4.866667,4.1375003,4.25,4.6222224,2.0416665,0.14444445,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.1555555,1.5833335,2.4333334,0.3916667,0.15555556,0.0,0.0,0.022222223,0.18333334,0.033333335,0.041666668,0.15555556,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025,0.4,0.475,0.61111104,0.41111112,0.4666667,0.36666667,1.0166667,0.9333333,0.65000004,0.90000004,0.6555556,0.2,0.15555556,0.15833333,0.10000001,0.275,1.0444444,1.9666667,2.1777778,2.511111,3.0166667,4.111111,4.791667,4.022222,3.275,2.811111,3.1666667,4.4000006,5.5777774,6.1499996,6.488889,7.3,8.51111,9.441667,10.677778,10.166668,9.4,8.411112,8.283333,8.233334,9.575001,11.822222,14.4,16.349998,17.57778,17.916668,19.377779,21.724998,23.955553,26.111115,27.741667,34.800003,49.81667,59.02222,57.6,56.288887,56.625,57.933334,59.86667,59.108337,57.57778,54.49167,49.300003,39.55,30.2,23.666668,21.058334,20.622223,22.241667,21.133333,21.316666,23.544445,26.341665,27.588888,26.422222,21.516666,16.788889,15.183332,15.444447,15.391667,13.68889,11.0222225,12.550001,16.922222,18.316668,13.3,5.7083335,1.6666669,0.675,0.44444445,0.40000004,0.18333335,0.033333335,0.11666667,0.22222222,0.19166666,0.13333334,0.20000002,0.06666667,0.07777778,0.75833327,0.6999999,0.36666667,0.07777778,0.10000001,0.025,0.0,0.22500001,0.07777778,0.10000002,0.25625002,1.4083334,0.38333333,1.725,1.175,1.1375,0.8416667,0.45000002,0.0,0.0,0.0,0.0,0.3543269,2.4568183,2.25,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.09375,0.25,0.0,0.0,0.0,0.0,0.325,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.8749999,1.2083333,1.53125,3.1083333,0.41666666,0.0,0.0,0.0,0.0,0.0125,0.025000002,0.025,0.0,0.016666668,0.12142858,0.5866667,1.5658333,2.85,3.0875,1.0,0.28333336,0.325,0.13333336,0.025,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.8250001,0.17500001,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.081250004,0.016666668,0.0,0.008333334,0.0,0.0,0.016666668,0.0875,0.275,0.47500002,0.71666676,0.73333335,0.29375002,0.108333334,0.5812501,0.9166667,1.1375,1.2750001,1.3562499,1.1916668,1.1583334,1.2250001,1.125,0.89375,0.57500005,0.41875005,0.48333332,0.45000005,0.45000005,0.5416666,0.78125006,0.8416667,0.84375,1.675,2.7624998,3.0833335,3.1583333,4.51875,5.7833343,6.8374996,7.541666,8.19375,9.658334,11.416666,13.012501,16.775002,17.843752,19.933334,23.693752,26.708332,29.258335,35.21875,37.125,34.46875,37.56666,42.0875,46.25,48.425003,47.933334,47.83334,47.6375,48.225002,50.3875,50.10833,44.71875,38.15,33.275,31.39375,31.358335,31.21875,30.258335,27.006252,23.983334,23.35625,24.866667,26.091667,25.756252,24.233334,24.568748,25.608334,20.81875,14.35,12.658333,17.3875,22.216667,22.181252,17.800001,10.36875,4.916667,2.1687498,1.0500001,0.76666665,1.11875,1.725,1.93125,1.8500001,1.6624999,1.1666667,0.91666675,0.625,0.15,0.24375002,0.275,0.16875,0.025000002,0.0,0.06875,0.14999999,0.38125002,0.36666667,0.025,0.3416667,0.0,0.0,0.6833334,0.45555556,0.0,2.488889,0.0,1.1555556,0.0,0.0,2.3733332,0.0,0.0,0.9133333,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.70000005,0.47777778,0.09166667,1.2,1.6583333,0.0,0.0,0.0,0.2,0.08333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.4333333,2.125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016666668,1.5666666,1.6833334,5.1666665,8.466667,0.725,0.0,0.041666668,0.28888887,0.9166667,0.31111112,0.06666667,0.20833334,0.24444444,0.23333335,0.3,0.4166667,1.4555556,2.175,0.9666667,0.11111112,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06666667,0.32222223,0.225,0.044444446,0.0,0.11111111,0.28888887,0.25000003,0.24444446,1.0083333,1.2333333,1.0083334,0.7666667,0.8666668,0.9888889,0.6444445,0.52500004,0.43333337,0.47500002,0.47777778,0.5416667,0.4666667,0.3888889,0.43333334,0.53333336,0.5833334,0.44444448,1.4166665,3.011111,1.925,1.1777778,0.97777784,2.4916668,3.6000001,4.45,4.8555555,4.466667,5.1666665,7.766667,9.608334,13.78889,18.399998,20.766668,27.291666,32.399998,39.622223,46.591663,51.3,50.19167,44.34444,43.274998,41.08889,39.591667,38.61111,39.033333,42.11667,46.877777,51.466667,51.855553,44.933334,40.677776,39.600002,41.36667,49.744446,56.975,56.300003,52.550003,46.800003,39.516666,34.266666,30.099998,27.650002,23.122221,19.7,21.533335,18.725002,15.833334,13.822224,12.983334,16.444445,18.908333,18.233334,13.283334,7.4000006,3.4583335,1.7666668,2.0,2.8416667,3.266667,2.5500002,1.9555557,1.575,1.1555556,0.8666667,0.51666665,0.35555556,0.8416667,0.41111112,0.17500001,0.07777778,0.06666667,0.41666666,0.7,0.31666666,0.0,0.0,0.0,0.0,0.79999995,0.0,0.0,0.0,0.0,0.3125,0.8666667,3.4166667,3.5464287,2.4016666,1.5604167,0.0,0.78882796,0.69595957,0.0,0.0,0.0,0.0,0.4416667,5.8932695,0.09166667,0.0,0.825,4.083333,5.0375004,1.3583333,1.3625,0.6666667,0.925,1.275,1.775,3.1916666,3.6833334,0.84375,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.3000001,1.5875001,5.541667,4.3416667,2.6187499,0.54999995,0.03125,0.016666668,0.9812499,2.433333,2.725,1.7249999,0.9666667,0.48125002,0.38333336,1.10625,1.6999998,1.53125,0.46666667,0.0,0.10625,0.2,0.125,0.89166665,0.4875,0.2,1.5583334,0.05,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.25,0.71250004,0.84166676,4.1937504,1.1333333,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.11250001,0.5,0.5375,0.16666669,0.1375,0.16666667,0.0,0.01875,0.033333335,0.18750001,0.3166667,0.23750001,0.13333334,0.14375001,0.20000002,0.19166668,0.2625,0.80000013,1.5374999,1.5250001,1.08125,0.75000006,0.65000004,0.68125,0.8666667,1.06875,1.0666667,1.5937501,1.8499999,1.9750001,1.3750001,1.0916667,2.0687501,2.641667,2.5562499,2.7166667,2.625,2.4833333,3.7833333,5.5750003,12.166668,18.4375,23.54167,30.812502,37.44167,49.533337,65.625,65.96667,54.94375,43.816673,33.26875,26.425,24.162498,23.966667,23.633333,24.71875,27.966667,32.043747,34.79167,34.537502,30.775002,31.716667,37.831253,50.55833,65.06875,72.458336,71.3375,66.566666,59.55,51.183334,47.583336,44.693752,41.25,37.362503,34.958332,28.7,21.800003,16.25,14.0375,15.783334,18.95625,21.816668,18.13125,10.75,5.5375,2.6666665,2.7083335,4.1875,4.375,3.4499998,2.841667,2.1125002,1.2916667,0.89166665,0.50625,0.53333336,0.9875,0.49166667,0.38125002,0.9416667,0.8833333,0.6625,0.083333336,0.09375001,0.06666667,0.075,0.0,0.0,0.0,0.0,0.0,0.0,0.9444445,1.9416667,0.0,0.0,3.375,0.0,3.112619,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.6888889,0.0,0.0,4.0444446,8.599999,4.7,4.3500004,1.6222222,0.59999996,1.7888889,1.6666666,1.9111112,0.48888892,0.20000002,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025000002,1.0,4.116667,5.633333,0.8666667,0.0,0.0,0.0,0.044444446,1.2916667,1.888889,4.1,2.6000001,0.9111111,0.275,0.13333334,2.3,3.4333332,3.1333334,2.483333,1.0777779,0.48333338,0.26666668,1.0916669,3.3111112,1.8083333,0.044444446,0.0,0.058333337,0.12222223,0.9250001,8.455556,1.9499999,0.08888889,1.7333333,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.022222223,0.083333336,0.3111111,1.6,0.6,0.025,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07777778,0.38333336,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.008333334,0.15555556,0.25833336,0.08888889,0.23333333,0.07777777,0.044444446,0.16666667,0.022222223,0.125,0.34444445,0.7083333,0.9666667,0.58333325,0.3888889,0.08888889,0.12500001,0.26666668,0.18333334,0.10000001,0.14166668,0.2777778,0.4444445,0.70833325,0.9666666,1.3666668,1.8444444,1.8499999,1.5888889,1.7833333,2.1,1.5,0.65000004,0.44444442,0.7916667,1.1444445,1.3000001,1.9000001,2.6222224,3.9666667,8.722221,13.483332,18.044447,25.808332,30.733332,35.188892,43.900005,48.133335,41.499996,32.822224,26.483335,22.41111,20.533335,20.688889,21.455557,22.908335,25.788889,25.850002,21.866667,21.458334,19.833336,19.055557,21.300003,34.73333,55.291664,69.62222,69.71667,65.31111,65.0,61.477776,56.077778,53.683334,48.755558,43.13333,38.72222,32.683334,24.233334,19.433332,18.375,20.655556,23.350002,23.444443,21.058334,16.566668,11.825001,7.0888896,6.633333,10.750001,13.677778,12.858333,10.333334,8.175,5.8222218,4.2222223,2.5666666,1.6111112,1.0583334,0.34444445,0.2,0.4,0.033333335,0.083333336,0.06666667,0.1,0.2,0.20000002,0.0,0.0,0.0,0.0,0.0,0.26666668,0.73333335,0.0,0.6555556,0.0,2.1,0.0,1.7722223,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.6222223,12.025,12.711111,2.3416665,0.12222223,0.29999998,0.39999998,0.275,0.12222223,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.12222223,0.9583334,4.055556,5.722223,0.29166666,0.0,0.0,0.0,0.0,1.5555557,5.1222224,4.5249996,1.3222222,0.05,0.22222222,1.6666666,6.1444445,5.7666664,3.0416665,0.88888884,0.041666668,0.033333335,0.34166667,0.9888889,0.80833334,0.0,0.0,0.0,0.0,0.19166666,0.7222222,0.075,0.0,0.0,0.05,0.5,1.4833335,6.700001,1.5083333,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.033333335,0.25,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.45000002,0.2,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011111111,0.05,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.055555556,0.12222223,0.16666667,0.5777778,0.23333335,0.0,0.0,0.0,0.0,0.0,0.0,0.016666668,0.24444446,0.5083333,0.15555555,0.033333335,0.044444446,0.06666667,0.23333333,0.32222223,0.33333334,0.26666668,0.10833335,0.0,0.044444446,0.083333336,0.11111111,0.15833333,0.2777778,0.4416667,0.51111114,0.6,0.5888889,0.68888885,0.75,0.6888889,1.8499999,2.9333334,2.5666668,2.5666666,3.177778,3.8,6.3555555,8.65,12.155557,17.616667,22.511108,26.433334,28.916666,27.833334,24.858335,23.46667,23.216665,20.944445,20.541664,21.244444,23.355556,25.8,28.777779,27.600004,23.566668,23.708334,24.722223,25.255556,27.358334,36.57778,51.08334,58.733337,58.433334,58.411114,60.283337,58.677776,54.466667,48.791668,47.300003,47.358334,44.18889,36.725,26.288889,20.91111,21.283333,22.58889,24.991665,25.411112,22.641668,18.855556,15.208334,12.48889,11.755556,12.275001,14.588891,15.800001,13.711113,10.641665,7.977778,7.044444,4.3250003,2.333333,0.7416667,0.38888887,0.19166668,0.13333334,0.17777778,0.116666675,0.17777778,0.22500002,0.24444446,0.28333336,0.0,0.0,0.0,0.0,0.29999998,0.425,0.0,2.4625,5.1166663,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.4106061,3.2247376,0.0,0.0,0.0,0.0,0.20000002,2.3333335,3.8375,9.416666,3.3374999,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.46250004,0.35,0.52500004,0.041666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025000002,0.69375,2.2250001,2.60625,0.8833333,0.0,0.20833334,0.45833337,3.2062502,3.4416666,4.4304166,1.6666667,3.775,8.266666,7.158334,4.7000003,1.5749999,0.04375,0.0,0.0,0.116666675,0.7625,0.10000001,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.09166667,0.05,0.45,0.56875,0.64166665,0.68333334,0.46875,0.13333334,0.050000004,0.033333335,0.0,0.0,0.0,0.0,0.0,0.056250002,0.7666667,0.13125,0.0,0.15,0.21875,0.8333334,1.56875,0.39166668,0.7875001,0.30000004,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.34166667,0.18333334,0.0,0.0,0.0,0.0,0.125,0.35000002,0.53333336,0.7375,0.6916666,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016666668,0.00625,0.008333334,0.0,0.0,0.0,0.0,0.0,0.025,0.016666668,0.0,0.0,0.050000004,0.108333334,0.17500001,0.25833333,0.33333334,0.45,0.70000005,1.76875,2.8083334,2.8625,2.6333332,2.8333335,3.4625,5.0249996,6.2062497,7.8166666,10.912498,12.558333,15.541665,17.16875,18.783335,18.09375,17.641668,19.575003,19.658333,19.750002,22.308336,25.683334,29.018751,30.150002,30.025003,27.874998,26.331251,25.741667,27.533335,33.781246,42.658337,51.325005,52.925,50.95,50.108334,50.856247,53.641663,51.908333,50.84375,49.975,49.475002,48.708336,44.618748,40.141663,32.86667,27.7875,26.81667,29.8,30.24167,26.874998,23.341667,21.118752,19.158333,14.433334,10.712501,10.225,10.125,8.375,6.693751,5.6000004,3.75,2.5125,1.6916667,1.91875,1.4166667,1.0625,0.95000005,0.82500005,0.65625,0.5583334,0.55,0.45000002,0.34375,0.0,0.0,0.0,0.0,0.39999998,0.6833334,0.39999998,1.05,2.7999997,0.18888889,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.125,0.0,0.0,0.0,0.05,0.75555557,1.4555556,1.1416667,0.24444444,0.5333333,0.0,0.0,0.0,0.0,0.11111113,0.6222222,0.91666675,0.45555553,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.09166667,1.2111111,1.6166666,0.98888886,0.0,0.0,0.0,0.016666668,0.011111111,0.0,0.0,0.008333334,0.06666667,0.033333335,0.0,0.0,0.0,0.6111111,2.7583332,2.9666667,0.90000004,0.0,0.0,0.0,0.2888889,2.891667,9.844444,10.316668,7.7888894,6.8777785,4.183334,1.9111111,0.19166669,0.0,0.0,0.0,0.39999998,0.13333334,0.0,0.0,0.0,0.0,0.3,0.108333334,0.033333335,0.022222223,0.016666668,0.0,0.016666668,0.055555556,0.7000001,1.8222222,1.675,0.7888889,0.47777775,0.19166668,0.17777778,0.05,0.0,0.0,0.0,0.06666667,0.008333334,0.0,0.008333334,0.22222222,0.19166668,0.41111115,0.94444454,1.0666667,0.9888889,0.41666672,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.40833333,0.4666667,0.0,0.0,0.0,0.85555553,0.5555556,0.38333336,0.0,0.0,0.1,0.175,0.5555556,1.8555557,0.43333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.075,0.15555555,0.12222222,0.0,0.0,0.0,0.0,0.016666668,0.044444446,0.041666668,0.07777777,0.1888889,0.4666667,0.9333334,1.7416667,1.7333335,1.7083333,2.0444446,2.3888886,2.8583333,3.6,4.375,4.9222217,5.1916666,6.822222,10.533333,13.308335,14.711112,16.041668,16.411114,17.308334,17.677776,18.208334,20.677776,22.266666,23.191668,23.744444,24.34167,22.877779,21.925001,23.211111,25.52222,31.933336,40.06667,45.333336,45.822227,45.61667,44.47778,43.933334,44.11111,44.41111,46.199997,48.577778,52.125,52.67778,54.01667,55.67778,54.122223,49.041664,44.32222,40.750004,38.37778,36.666668,32.911114,28.391666,26.11111,24.633335,20.575,15.555556,12.558334,11.111111,9.458334,7.6444454,5.8888893,5.041667,5.477778,5.3916664,4.366667,2.9333334,1.8666667,1.6111112,1.2833335,1.2555556,1.1083333,0.9555556,0.68333334,0.0,0.0,0.275,0.45,0.033333335,0.0,0.0,0.64375,4.5666666,3.45,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05,0.25,1.2250001,1.6249999,0.45000002,0.0,0.0,0.0,0.0,0.0,0.0,0.008333334,0.24166667,0.81875,1.3833333,0.2375,0.22500001,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.25,1.0375001,2.1000001,3.2187502,4.0333333,1.20625,0.025000002,0.0,0.0125,0.125,0.01875,0.0,0.0,0.13333334,0.46875,0.17500001,0.14166667,0.025,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.49166667,0.30625004,0.7666667,1.1624999,1.2583331,1.1833333,0.8187499,0.35833335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025,0.50624996,1.25,0.36249998,0.09166667,0.06666667,0.01875,0.0,0.23750003,0.9583334,1.5624999,0.86666673,0.15625,0.0,0.0,0.0,0.0,0.0,0.05,0.1375,0.25833336,0.9833333,1.5874999,1.4166667,1.625,1.1250001,0.4875,0.5916667,2.5000002,0.48750004,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.16875,1.375,0.3,0.97499996,0.19375001,0.51666665,0.60833335,1.125,0.7916666,0.125,0.058333337,0.03125,0.6916666,3.25,3.6937501,0.59999996,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.058333337,0.30625004,0.76666677,1.3374999,1.6666665,1.9,2.5166667,2.9916666,3.6812499,4.0583334,4.0125,4.2250004,4.7812505,5.2166667,8.016666,11.043751,12.45,14.7375,15.358335,16.04375,18.216665,21.575,25.066666,24.683332,24.2625,23.466667,22.137499,20.141668,20.956251,23.2,25.916668,31.837502,40.225,44.46875,46.249996,46.8875,47.416664,47.200005,46.116673,46.458336,45.85625,45.933334,49.5625,51.89167,52.981255,53.683327,56.000004,56.15625,54.233334,51.3375,48.283337,47.4375,45.174995,40.55625,35.133335,33.0,34.756252,36.541668,34.062504,27.824999,23.118752,19.033333,15.883333,12.662499,11.608335,12.6125,8.733333,6.14375,4.216667,3.4916668,3.3062503,3.1083336,2.7875001,2.1833334,1.5875,0.0,1.9999999,0.0,0.29999998,0.0,0.0,0.45555556,1.8166666,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05555556,0.275,0.33333334,0.17777778,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.1999999,2.3444445,2.3000002,2.488889,3.233333,0.8666667,0.022222223,0.0,0.011111111,0.1,0.0,0.0,0.4222222,1.2666667,0.9444445,0.36666664,0.1,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.7111112,0.6750001,0.0,0.083333336,0.022222223,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.022222223,0.116666675,0.08888889,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.4,3.9250002,1.2333333,0.72222227,1.625,1.6555556,1.7916666,1.8333335,3.3916667,4.2000003,4.866667,4.4333334,3.6,1.3416667,0.31111112,0.075,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.45555556,0.40000004,0.6444444,0.0,0.6,0.055555556,0.21666668,0.95555556,0.11666666,0.0,0.0,0.5888889,6.1000004,12.45,2.2555554,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05,0.011111111,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.033333335,0.25,0.66666675,1.5583333,2.5111113,3.3083332,4.0888886,4.533334,5.2583337,5.4111114,4.8750005,4.711111,5.0333333,4.1777782,4.444444,6.191667,9.0222225,12.833334,16.7,20.433332,23.099998,25.6,26.777779,26.57778,28.291666,27.355555,24.583334,22.28889,22.216665,25.655556,32.2,38.833336,43.58889,47.683334,50.377777,51.44166,51.95556,51.716667,49.93333,50.0,49.400005,46.455555,48.583336,50.8,52.875004,53.52222,54.422222,53.175003,51.86667,52.891666,53.02222,52.44166,51.41111,48.91667,45.800003,43.98889,43.908333,46.72222,51.708336,52.288895,47.375,41.344444,35.72222,29.45,24.755556,22.958334,17.833334,15.991668,11.766667,9.455556,7.9833336,7.0,6.7166667,6.2,5.5249996,0.0,0.7916667,0.19166668,0.01875,0.008333334,0.54375005,0.38333333,0.25,1.0833334,2.1,0.0,0.0,0.0,0.0,0.0,0.0,1.2375,0.0,0.0,0.0,0.0,0.11761905,0.20833334,0.0375,0.21666667,0.28333333,0.0375,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.30833334,1.8875002,2.5583334,1.9000001,2.025,1.4333334,0.0,0.0,0.0125,0.09166666,0.05,0.108333334,0.41875,0.9499999,1.4166666,1.4625,0.59166676,0.04375,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06875001,0.041666668,0.0,0.0,0.041666668,0.2125,0.2916667,0.05,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016666668,0.03125,0.29166666,0.25833336,0.50625,0.0,0.0,0.0,0.01875,1.95,2.99375,1.3136363,1.125,2.48125,3.4750001,3.01875,3.6166666,4.03125,4.616667,3.2583334,2.0812502,1.1583333,0.32500002,0.04166667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.17500001,0.17500001,0.0125,0.0,0.0,0.016666668,0.0,0.0,0.1,0.03125,0.0,0.00625,0.24166667,3.7250001,8.618751,1.4666667,0.0,0.0,0.0,0.0,0.06666667,0.25,0.23333332,0.081250004,0.008333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.075,0.3416667,0.525,1.0000001,1.7416667,2.8812501,4.0583334,5.2,5.916667,5.95,6.34375,7.041667,6.6187496,6.3416667,6.23125,5.616667,5.3500004,6.0499997,7.3,10.318749,14.5,18.281248,21.583334,24.39375,27.900002,30.25,31.956253,29.883335,26.412502,24.208334,25.443752,31.491669,38.641666,43.71875,45.94167,46.4,45.375004,45.350002,45.450005,46.418755,45.666664,44.808334,42.443752,40.816666,42.81875,45.43334,47.637497,49.175,51.775,54.356243,54.949997,53.818752,54.666668,59.362495,63.183334,64.725006,63.483334,61.00834,58.95625,57.29167,58.75,59.425,57.631252,55.633335,51.816666,47.20625,43.63334,35.7125,30.008333,24.3375,19.616667,15.85,11.775,9.183333,8.306251,7.8500004,7.0062504,0.0,0.0,0.0,0.3416667,0.0,1.0250001,1.2777778,2.5749998,3.0444446,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14166668,0.26666665,0.083333336,0.6666667,1.0444444,0.7166667,0.022222223,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06666667,0.26666668,0.7666667,0.8916666,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.3,1.8555557,2.6166663,1.6888889,2.266667,0.6166667,0.3222222,0.14166668,0.06666667,0.083333336,0.06666667,0.008333334,0.0888889,0.4888889,1.2249999,1.7888889,1.0666666,0.11111111,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.41111115,1.0,0.85555553,0.25833336,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016666668,0.22222224,0.64444447,0.9583334,0.42222226,0.058333337,0.0,0.0,0.0,0.008333334,0.06666667,0.48888892,2.0333333,3.5111115,2.6666667,2.211111,1.9666668,1.4777778,1.0666667,0.53333336,0.1,0.016666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.4166667,0.0,0.0,0.0,0.0,0.0,0.0,0.058333337,0.41111112,0.0,0.0,0.0,0.13333334,1.8888891,2.3416665,0.28888887,0.0,0.0,0.06666667,0.48888892,0.67777777,0.23333333,0.0,0.0,0.0,0.0,0.044444446,0.016666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06666667,0.33333334,0.5777778,1.0166667,1.8444445,2.8083334,3.4333334,3.8166666,4.366667,4.311111,4.4916663,5.322222,5.825,6.2111115,5.9916663,4.988889,5.3444443,7.116667,8.400001,10.733335,13.377777,15.933333,17.811111,20.95,23.366665,25.011112,26.65,27.000002,25.7,25.666668,30.8,35.555557,38.322224,41.375004,44.18889,43.125004,41.4,40.275,40.36666,40.958332,40.488888,38.966667,36.541664,35.377777,35.783337,38.166664,41.649998,45.444443,49.711113,55.13334,60.511112,63.61667,63.877777,63.908333,69.42222,72.683334,68.88889,67.77778,68.333336,62.17778,61.14167,64.688896,64.60834,62.822224,61.28889,56.333336,48.61111,39.949997,30.744446,24.791668,19.9,17.333332,13.65,11.299999,9.383333,8.311111,8.168182,0.82500005,0.25555557,1.1444445,0.0,0.39999998,1.3666667,0.9666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.126515,0.0,0.0,0.0,0.425,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.041666668,0.33333334,1.4916668,4.055556,4.4833336,3.1111112,0.64444447,0.058333337,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.4,0.6,0.18333334,0.0,0.0,0.15555555,0.25833336,1.3000001,1.2444445,1.0,0.46666667,0.79999995,0.44444445,0.34166667,0.08888888,0.008333334,0.0,0.0,0.17500001,0.47777778,1.0416667,0.8888889,0.1,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.43333334,1.4916668,0.67777777,0.25833333,0.7,1.2416668,0.7555555,0.17777778,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016666668,0.26666665,0.0,0.0,0.0,0.06666667,0.65833336,1.7222223,1.5222223,1.6666667,3.8555555,2.5333333,0.37777779,0.40833333,0.3,0.19999999,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.108333334,0.1,0.008333334,0.0,0.0,0.011111111,0.13333334,0.15,0.033333335,0.0,0.0,0.3083333,0.24444446,0.06666667,0.0,0.0,0.0,0.07777777,0.44166666,0.34444442,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1,0.08888889,0.13333334,0.19166666,0.54444444,1.0666667,1.9555557,2.5666666,2.8000002,3.0666666,4.041667,5.5111113,6.2916675,6.855556,6.7749996,5.7444444,4.9333334,6.0166664,7.677778,9.8,12.9,16.133333,18.322224,19.441668,20.222221,21.38889,23.0,22.788889,23.56667,29.066666,33.925003,35.899998,37.711113,42.86667,44.38889,44.191666,44.333336,43.625,44.444443,43.316666,41.711113,40.6,39.95001,40.255558,38.516666,39.7,42.000004,43.677776,45.233334,49.54167,54.88889,56.900005,56.577778,56.083332,59.011112,62.91667,66.0889,62.86666,58.55,52.81111,50.391666,54.544445,54.999996,52.822224,50.533333,43.141666,36.355556,32.841667,29.522223,28.21667,25.588888,21.266668,17.133335,13.677778,10.475,8.388888,7.7833333,0.91875005,0.0,0.0,0.0,0.0,0.0,0.0,0.28750002,0.9583333,1.05,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.6375,0.90833336,0.2916667,0.087500006,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.008333334,0.16875002,0.9666667,2.3874998,3.1833334,2.75625,2.1416667,2.4083333,0.96875,0.1,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025000002,0.54999995,0.78749996,0.0,0.0,0.0,0.0,1.1500001,2.8083332,2.4,1.375,0.79375,1.0833334,0.6375,0.4666667,0.225,0.058333337,0.0,0.0,0.016666668,0.13125,0.116666675,0.0375,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0375,0.29166666,0.78750014,0.39166668,0.7062501,1.6250001,1.6687502,0.7666667,0.23333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.28125,1.525,0.15,0.18333334,1.00625,2.1333332,2.825,1.73125,2.0583334,1.6875002,0.20833334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00625,0.07500001,0.17500001,0.49374998,1.0333333,1.4125,1.2,0.2875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.17500001,0.8375,0.72499996,0.5833334,0.35625002,0.36666667,0.49375,0.7416666,1.25,1.7750001,2.458333,3.25625,3.7166667,4.8249993,6.025,6.75625,5.658334,4.3083334,4.9812503,6.283333,8.66875,11.550002,15.05625,18.2,19.381252,19.133333,19.533333,22.393751,27.550003,33.625,38.74167,42.1375,40.483334,38.916668,39.262505,41.783333,45.48125,47.7,50.1125,51.016666,47.5625,45.741665,46.35,48.2625,49.875004,46.862503,46.649998,46.61875,45.141666,45.683334,46.9625,50.241673,50.95625,52.975002,52.125,48.81667,46.143745,47.166668,47.375,45.350002,40.383335,37.231255,38.625,39.287502,37.708336,33.50833,29.00625,26.508333,28.58125,28.508335,28.20625,26.258335,23.933332,20.631248,15.991667,13.512501,10.674999,12.942499,0.0,0.39999998,0.39999998,0.79999995,0.39999998,0.6833334,0.0,0.0,0.0,0.5555555,0.0,1.1555555,0.0,0.0,2.0916665,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14444445,0.93333334,1.6444445,0.83333343,0.13333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.16666666,0.85,1.0555556,0.36666667,0.46666664,0.11111111,0.016666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.033333335,0.37500003,0.0,0.0,0.0,0.0,0.0,0.8666667,2.3083334,2.1111112,1.2583333,0.57777774,1.1666667,0.7222222,0.7666667,0.44444445,0.08888889,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05555556,0.21666667,0.25555557,0.26666668,1.0444444,0.7083334,0.3,0.022222223,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.075,0.6,1.075,1.6444445,4.183334,2.4444444,1.8888891,1.0500001,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08888889,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.022222223,0.1,0.42499998,0.92222226,1.1583333,0.35555556,0.033333335,0.1,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011111111,0.016666668,0.055555556,0.30833337,0.8555556,1.4666667,2.1666667,2.6666665,3.9416666,4.1888895,4.2833333,5.2777777,5.1000004,5.1083326,5.888889,6.674999,8.455556,11.55,14.411111,15.425,17.244446,20.477777,27.416668,37.233334,42.291664,43.1,42.233334,39.322224,39.95556,41.925,45.92222,52.116673,57.06667,59.54167,57.833336,53.141674,50.36666,52.133335,52.416668,50.722225,51.10833,50.377773,48.766666,48.022217,47.833336,47.583332,47.46667,46.9,46.32222,45.6,41.844448,40.0,40.72222,39.86667,37.625,33.733334,34.541664,34.88889,35.56667,33.2,30.344444,27.408337,25.044443,26.258335,27.033333,28.083332,26.988892,24.966667,22.716665,19.644445,17.075,15.688889,15.875,0.0,0.3416667,0.0,0.0,0.0,0.48125,0.3416667,0.0,0.0,0.0,0.76875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08125,0.18333332,0.04375,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.075,0.69166666,1.9875001,1.3083334,0.57500005,0.49166664,0.0625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.056250002,0.6333333,0.50000006,0.16875,0.0,0.0,0.0,0.0,0.0,0.0,0.4,2.6666665,2.2500002,0.9666667,0.7875001,1.1000001,1.0812501,0.81666666,0.47500002,0.44375002,1.1416667,0.38124996,0.083333336,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.22500001,0.38333333,0.18749999,0.108333334,0.1375,0.075,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.008333334,0.38125,0.9916667,0.38125002,0.075,0.82500005,0.475,0.23333333,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.8166667,0.48125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.008333334,0.033333335,0.275,0.51666665,0.13125,0.0,0.4125,2.1833334,2.6374998,0.24166667,0.05,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14166667,0.0,0.0,0.0,0.0,0.0,0.0,0.041666668,0.05,0.36875,1.0666668,2.0500002,3.3666668,4.462499,5.9500003,7.533334,8.89375,9.991668,11.1625,12.716666,13.937499,15.158334,15.4375,15.191668,15.066668,16.29375,19.35,27.2,32.933334,38.40625,41.483334,44.350002,46.612503,51.225002,57.0625,64.25,65.775,62.925,57.83125,53.808334,50.899998,50.431248,48.824997,46.4875,43.941666,42.64375,42.625004,42.199997,42.999996,41.691666,40.068752,39.600002,37.83125,36.375,36.100002,37.108334,37.008335,32.55625,35.616665,37.36875,37.691666,36.73125,34.966667,35.375,34.61875,32.791668,32.662502,31.550003,30.96875,30.741669,26.816668,22.293753,17.408333,14.275,11.766666,10.50625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.29999998,0.0,0.45555556,0.76666665,0.71111107,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.20833333,0.4,0.13333334,0.0,0.0,0.0,0.2777778,0.44166666,0.3,0.25833336,0.11111111,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.2,5.0000005,10.48889,7.2083335,3.8555555,2.7416668,0.53333336,0.055555556,0.0,0.0,0.0,0.0,0.0,0.0,0.25833336,1.6111112,1.6333333,0.57500005,0.26666668,0.058333334,0.46666664,0.09166667,0.0,0.42222223,3.5,2.0,0.78333336,2.5555553,1.1333333,0.13333334,0.22500001,0.22222221,0.33333334,0.40833336,1.1222222,3.1333337,1.4444445,0.20833334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025000002,0.25555554,0.30833334,0.15555556,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.275,1.0888889,0.8777778,1.1166667,1.2888889,0.90000004,0.6666666,0.46666667,1.0111111,1.2166666,0.3888889,0.2888889,0.008333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016666668,0.011111111,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06666667,0.7111112,4.0,7.611111,1.975,0.2777778,0.3,0.06666667,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.21666668,0.18888889,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.09166667,0.17777778,0.45,1.3111111,2.4666667,4.2444444,6.377778,9.158333,12.322223,15.816667,18.177778,19.216667,19.633335,18.425,18.244444,17.555557,16.616665,15.011111,15.141667,19.066668,24.758333,32.688892,40.36667,44.558334,48.055557,53.983337,57.844448,59.225,56.622227,52.733334,52.955555,53.72222,51.80833,47.344448,43.591667,40.31111,38.300003,37.511112,36.81111,36.5,36.233334,34.683334,33.233334,30.875,26.322224,24.816668,24.366667,24.533333,24.625,25.666668,30.108334,35.86667,37.433334,38.933334,38.333336,40.258335,39.855553,36.758335,31.722221,31.125002,28.722221,28.444445,25.350002,19.333334,15.575001,12.655556,11.283333,2.2625,0.10833333,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.041666668,0.20000002,0.45,0.7250001,0.95625,2.3166666,2.75,1.1166668,0.65000004,0.21666667,0.05625,0.008333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.38125,3.0666666,8.7875,12.325001,9.45625,5.116667,2.141667,0.34375,0.0,0.0,0.0,0.0,0.0,0.0,0.016666668,0.20000002,0.58750004,0.51666665,0.20000002,0.4416667,0.25625002,0.06666667,0.15833333,1.0750002,1.2666667,0.26250002,0.525,0.69375,0.725,0.3,0.0,0.06666667,0.16875,0.18333334,0.54375005,0.55,0.61875004,0.15833333,0.016666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00625,0.09166667,0.056250002,0.041666668,0.081250004,0.058333337,0.03125,0.016666668,0.025000002,0.075,0.15,0.23750001,1.0666666,2.575,3.7083335,4.7166667,5.2250004,6.05,4.65625,3.5833335,3.25,3.1999998,2.2562504,0.9416667,0.34166667,0.0125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0375,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025,0.24375,0.7916667,1.6750001,2.7333336,3.0375,1.6166667,0.48125002,0.41666672,0.4,0.1875,0.025,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.008333334,0.0625,0.1,0.15,0.15,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.043750003,0.34999993,0.81875,1.5083334,2.475,4.1499996,6.1500006,8.7625,10.924999,13.156252,16.075,19.362503,22.316668,23.925001,23.10625,19.391668,15.968752,15.450001,18.243752,20.991665,26.683334,32.275,34.908333,33.250004,35.24167,39.4375,41.508335,43.287502,46.258335,48.266666,47.918755,45.583336,40.9875,36.633335,33.79375,31.008333,29.075003,27.656252,26.983334,26.887503,26.341667,25.83125,24.55,23.693748,23.283335,23.433334,25.731253,26.883335,28.500002,32.441666,32.24375,33.675,35.516666,38.518753,40.51667,41.28125,37.61667,36.193752,35.458336,34.541668,34.024998,30.308334,27.706251,24.708334,20.2,4.633333,2.211111,0.22222222,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016666668,0.033333335,0.033333335,0.06666667,0.2,0.55,2.788889,3.9750001,0.90000004,0.30833334,0.08888889,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.21666665,2.5444443,6.408334,10.011111,7.3333335,3.8083336,0.74444443,0.16666667,0.0,0.0,0.044444446,0.10000001,0.033333335,0.044444446,0.26666668,0.64444447,0.2916667,0.2666667,0.23333335,0.2777778,0.988889,0.6,0.7666667,0.39166662,0.0,0.85833335,1.6333336,0.7083334,0.08888889,0.6,1.1166667,0.5222223,0.5,0.1,0.7166667,0.9666667,0.48888892,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025000002,0.2888889,0.19999997,0.10000001,0.0,0.0,0.0,0.0,0.0,0.0,0.022222223,0.033333335,0.033333335,0.075,0.33333334,0.5,0.2916667,0.6,0.5916667,0.75555557,0.7,0.64444447,0.2,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.23333332,0.7555555,1.2166666,1.4333335,1.1166667,0.8222222,0.2833333,0.24444446,0.18333335,0.10000001,0.07777777,0.1,1.2000002,2.216667,3.8888888,1.9333332,0.3888889,0.08888889,0.20833334,0.044444446,0.0,0.0,0.0,0.0,0.05,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025,0.13333334,0.22500002,0.6777777,1.1555555,1.5833333,1.9333333,2.2,3.322222,5.05,6.9666667,9.475,12.033334,14.411111,17.233332,20.044445,20.566668,19.222225,18.241667,17.144445,16.622223,16.491667,17.211113,20.583334,22.733335,26.816668,28.933332,32.808334,34.855556,37.344444,39.475,39.6,38.73333,37.199997,35.525,33.37778,30.455559,28.166666,25.122225,22.500002,20.199999,18.5,18.244446,19.475,20.0,20.877777,24.025,29.266666,34.441666,36.055557,33.175,33.6,33.1,34.891666,37.6,42.76667,45.988888,47.233337,48.0,47.755554,44.641663,37.41111,32.216667,29.366667,23.066666,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.4166667,0.8444444,0.975,0.6222222,0.5,0.0,0.78888893,0.18333334,2.477778,2.3333337,1.5888889,0.19999999,0.0,0.033333335,0.058333337,0.11111111,0.275,1.2111111,3.7500002,3.1111112,1.1833334,0.34444445,0.22222224,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.1666667,3.5222225,7.733334,9.908334,6.255555,2.0583334,0.8,0.1,0.10000001,0.65000004,0.9333334,0.44444445,0.31666666,1.1666667,1.3666668,0.06666667,0.041666668,0.14444445,0.4,0.375,0.07777778,0.20000002,0.06666667,0.9166666,4.2444444,3.5083334,2.1555557,2.0555556,1.3666667,1.0555556,0.7166667,0.13333334,0.0,0.0,0.14444445,0.116666675,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.058333334,0.15555555,0.19166666,0.055555556,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016666668,0.1888889,0.4,0.44166666,0.26666668,0.12500001,0.0888889,0.075,0.08888889,0.43333337,1.1666666,1.8111111,2.3333333,7.7,12.783334,9.6,3.625,0.8777778,0.5111111,1.1166667,1.9,0.91666675,0.42222223,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.022222223,0.016666668,0.033333335,0.0,0.20833334,0.3888889,0.4166667,1.1222223,2.9916668,5.2000003,5.5,5.888889,6.1666665,8.066667,10.044445,13.25,16.999998,18.266668,18.7,20.577778,23.016666,23.222223,20.333334,17.51111,16.725,20.055555,24.175001,29.211111,33.788887,36.841667,36.58889,35.308334,33.31111,30.933334,29.633335,29.177778,27.633333,24.666666,21.991665,19.266668,16.591667,14.422223,14.1,14.877777,15.733333,19.550001,23.711111,26.750002,26.8,24.133331,23.07778,23.877779,27.16667,33.48889,35.74167,37.76667,39.699997,43.733334,43.988888,44.041668,40.63333,36.458336,31.177778,23.775,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.125,0.13333333,0.4875,1.2333333,1.475,0.9916667,0.76875013,0.225,0.008333334,0.0375,0.0,0.0,0.20833334,0.08125,0.22500001,0.1,0.10625,0.14166667,0.28750002,0.7916667,1.1304166,3.5219696,3.2437496,1.9166665,2.1916666,0.75,0.075,0.01875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.2916667,1.7750002,4.40625,6.716667,5.9000006,1.7333332,0.45625,0.0,0.25625,1.0333334,1.0833335,0.20000002,0.13333334,0.43125,0.5416667,0.28125,0.0,0.0,0.0,0.0,0.01875,0.0,0.275,1.175,0.55625,0.67499995,0.5416667,0.51874995,0.28333333,0.19375001,0.0,0.0,0.0,0.041666668,0.11250001,0.09166667,0.01875,0.0,0.0,0.0,0.0,0.025,0.1,0.175,0.041666668,0.00625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.008333334,0.20000002,0.8083333,0.9916667,0.49375004,0.0,0.0125,0.05,0.0375,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.008333334,0.025,0.025000002,0.33125004,0.90833336,1.2625,1.1333333,1.2416667,1.6312501,2.0333333,3.3249998,1.9000001,1.3125,0.88333344,1.2416667,3.6,1.2500001,0.73125005,0.3,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.083333336,0.3375,0.975,1.5937501,2.0916667,2.3666668,2.96875,3.9000003,4.7875,6.0833335,7.70625,9.183333,10.758333,14.612501,19.583334,22.343752,23.350002,22.462502,19.583334,17.09375,18.491667,22.033333,27.843748,31.225,32.43125,32.125,29.86875,28.641668,25.933334,23.806252,22.066668,20.21875,19.191668,16.79375,15.541668,15.231249,16.108332,16.116667,18.037502,20.850002,22.54375,20.116667,20.856249,23.574999,26.375,29.275,31.891668,34.487503,37.883335,40.318752,40.225002,38.333336,35.737503,35.291668,33.318752,32.475,29.4875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011111111,0.67499995,3.4222221,0.16666667,0.0,0.0,0.0,0.0,0.0,0.0,0.083333336,0.011111111,0.0,0.0,0.0,0.0,0.0,0.0,0.22222222,1.5672619,3.6458335,3.8555558,2.3666668,0.88888896,0.17500001,0.022222223,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.40000004,0.90000004,1.8666667,2.0555556,0.6916667,0.06666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1,0.2,0.0,0.0,0.0,0.0,0.0,0.0,0.62222224,1.875,0.8444445,0.0,0.0,0.011111111,0.1,0.3,0.5416667,0.22222222,0.0,0.0,0.0,0.06666667,0.20000002,0.2916667,0.28888887,0.083333336,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.099999994,0.4,0.6111111,0.43333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06666667,0.24999997,0.28888893,0.31666666,0.4333333,0.35555556,0.25833333,0.40000004,0.5083333,0.47777778,0.15833335,0.07777778,0.044444446,0.06666667,0.06666667,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13333334,0.22500001,0.44444448,0.77500004,1.2111112,1.7833333,2.2444446,3.0222223,4.45,7.622222,13.083334,20.755558,23.008333,21.5,19.225,17.111113,17.744444,21.675001,22.566668,24.383333,25.955557,26.483334,26.822222,26.444443,25.716667,23.177776,20.908333,19.1,17.85,16.766668,16.266666,17.822224,19.555557,21.399998,22.344446,24.741667,26.766666,26.908335,25.333334,28.555557,30.4,32.666668,34.241665,35.08889,36.100002,35.4,35.633335,30.025002,26.622223,23.641666,23.366667,22.516666,0.025,1.7166667,0.30833337,0.4375,0.0,0.056250002,0.0,0.0,0.0,0.0,0.0,0.0,1.10625,3.0416667,1.6437502,0.6333333,0.0375,0.1,0.0,0.0,0.0,0.0,0.0,0.28125,0.25,0.15,0.075,0.025,0.00625,0.0,0.0,0.0,0.10708334,0.1448052,1.3710316,2.1812496,1.9750001,0.64375,0.15833335,0.0125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.31875,1.5916668,1.40625,0.55,0.6625,0.20000002,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025,0.26250002,0.9250001,0.5124999,0.1,0.0,0.0,0.0,0.0,0.10000001,0.20625,0.0,0.0,0.0,0.20000002,0.6,1.1666666,1.35625,1.5666668,1.45625,0.7666667,0.24166666,0.0375,0.09166667,0.15625,0.36666664,0.65625006,0.65000004,1.03125,1.2916667,0.8416667,0.6625001,0.5833334,0.39375,0.28333336,0.25,0.075,0.083333336,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0625,0.058333337,0.025,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025,0.06875,0.016666668,0.0,0.0,0.025,0.0,0.016666668,0.00625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025,0.075,0.2,0.3416667,0.69166666,1.39375,2.15,3.3374996,5.533334,8.787499,13.375,15.849999,17.000002,19.966667,24.056252,25.441668,25.225002,25.474998,25.5,25.358334,27.724997,28.55625,28.125,27.35,25.433334,23.243752,21.358334,19.906252,18.89167,18.408333,21.024998,24.375,25.45,25.466665,27.325,31.383333,33.183334,34.831253,37.524998,37.475,37.1,37.36875,36.425,32.4,27.46875,23.599998,21.775,23.5,23.89375,0.0,0.0,0.033333335,0.0,0.07777778,2.1416667,1.7222222,0.1,1.5666668,1.4444445,1.2333333,3.8666668,3.525,6.7333336,3.7583334,0.43333337,0.116666675,0.0,0.0,0.18333334,0.8333334,0.48333335,0.18888888,0.19166666,0.36666667,1.0333333,0.14166667,0.08888889,0.008333334,0.0,0.0,0.0,0.0,0.0,0.0,0.5464286,1.7984127,0.7583334,0.34444445,0.083333336,0.0,0.0,0.05,0.033333335,0.0,0.0,0.0,0.0,0.0,0.1,0.8222222,2.1166668,0.75555557,0.0,0.0,0.0,0.0,0.0,0.0,0.011111111,0.13333334,0.044444446,0.0,0.0,0.0,0.0,0.0,0.53333336,1.0888889,0.5250001,0.7,0.22500002,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.19166668,0.76666665,1.7250001,2.888889,3.4916668,2.1111112,1.1555556,0.59999996,0.31111112,0.49166664,0.65555555,0.6333334,0.40000004,0.22500002,0.22222224,0.54444444,0.73333335,0.5333333,0.6333333,0.54444444,0.6333333,0.5555556,0.2,0.05,0.31111112,0.4083333,0.2777778,0.15,0.16666667,0.24999999,0.4,1.0222223,1.4583335,1.3555555,0.7750001,0.21111111,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13333334,1.625,2.5444443,2.2333333,1.7166667,1.0888889,0.39166668,0.11111112,0.041666668,0.044444446,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.033333335,0.20000003,0.53333336,0.99166673,1.2777778,3.241667,4.6666665,6.183333,7.5888886,10.611112,14.516667,19.733334,25.208332,29.48889,30.650002,32.166664,32.18889,33.475002,32.600002,32.283333,29.922222,28.400002,27.788889,27.783333,26.833332,25.322224,24.975002,25.488888,26.658333,28.177778,30.191666,31.688889,34.28889,35.091663,36.88889,37.850002,37.98889,39.591667,39.211113,36.622223,29.616667,26.8,23.55,26.211111,25.825,0.0,0.0,0.0,0.04375,0.32500002,0.96875,0.7583333,0.118750006,0.49621212,5.4916673,10.612501,9.775001,7.5750003,6.4416666,2.5687501,1.2055554,0.46249998,0.2666667,0.23333335,1.7812501,6.4833336,5.4125,1.1,0.043750003,0.025,0.041666668,0.043750003,0.008333334,0.03125,0.0,0.0,0.0,0.0,0.0,0.02,0.04107143,0.029166669,0.42067307,0.25,0.0625,0.0,0.0,0.01875,0.2,0.4,0.2,0.0,0.0,0.0,0.0,0.23333333,1.3000001,1.0,0.12499999,0.0,0.0,0.0,0.0,0.0,0.008333334,0.28125,0.15833333,0.0,0.0,0.0,0.0,0.77500004,10.868752,7.5333333,2.24375,0.425,0.44375002,0.13333334,0.016666668,0.0,0.13333334,0.46250007,0.42500004,0.0125,0.0,0.0,0.0,0.041666668,0.24374999,0.98333347,1.4499999,1.225,1.5083334,1.8937501,1.825,1.5875001,1.3583333,0.9812499,0.64166665,0.325,0.25833336,0.16666667,0.5875,2.1916668,1.9,1.3333334,1.3875,1.7583333,1.6333332,2.2499998,2.5,2.30625,1.8583335,1.8437501,1.7083334,1.325,1.1500001,1.0166668,0.9375001,0.5,0.1375,0.008333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.175,0.06666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.1166667,4.425,7.1333337,7.1625,6.158334,5.1333337,3.8312502,2.5666666,1.34375,0.80833334,0.4875,0.32500002,0.2,0.17500001,0.06666667,0.15625,0.15,0.05,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025000002,0.15625,0.22500002,0.39374998,0.65000004,1.0625,1.7250001,3.0625,4.458333,5.616667,7.9812493,10.033333,13.650001,19.15,23.687504,26.758335,29.991669,31.581247,32.14167,30.7625,29.44167,28.650002,30.141666,31.775002,33.241665,33.033333,34.0375,36.191666,36.012505,36.058334,37.80625,41.308334,43.63333,46.712498,48.100002,46.268753,46.591667,45.34375,43.800003,36.666668,29.481249,25.808334,28.806248,33.216667,31.306253,0.18333334,0.45555556,0.38888893,0.083333336,0.6222222,0.625,0.23333332,0.041666668,0.2611111,0.88611114,3.6541667,2.3944445,2.0907648,1.7375001,2.3083334,1.7222223,1.5550001,0.8888889,0.41111112,1.5,2.6666665,1.4416666,0.7666667,0.48484856,0.14444445,0.06666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.15555556,0.05,0.0,0.0,0.0,0.0,0.0,0.0,0.39166668,0.25555557,0.60833335,0.0,0.0,0.0,0.0,0.25,0.44444445,0.19999999,0.0,0.0,0.0,0.0,0.18333334,0.12222223,0.008333334,0.0,0.0,0.0,0.0,0.0,0.0,4.366667,1.9,1.6666667,0.18888888,0.48333335,0.76666665,0.14444444,0.0,0.85555565,1.5833335,1.0333333,0.18333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14444445,0.47500002,0.6666667,0.40833333,0.4,0.5,0.788889,1.2583334,0.97777766,0.7777778,0.79999995,0.57777774,0.24166667,0.23333335,0.075,0.16666667,0.27777776,0.33333334,0.32222223,0.18333334,0.07777778,0.041666668,0.011111111,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.8666667,5.625,10.333334,12.583334,11.555556,10.750001,10.622221,10.377778,9.675,8.01111,6.116667,4.7444444,2.9833336,1.5444444,0.72222227,0.25,0.0,0.0,0.13333334,0.26666668,0.5,0.25,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.033333335,0.13333334,0.33333334,0.5222223,0.75000006,0.88888884,0.90000004,1.2,2.3333333,3.4333334,4.855556,6.866667,9.144444,11.666666,14.844444,15.733334,18.591667,22.377777,25.025,26.533333,27.741665,29.68889,32.433334,35.32222,36.56667,38.133335,40.622223,41.11667,41.82222,41.758335,42.3,45.422222,46.225006,47.18889,47.158333,47.81111,46.708332,41.58889,34.666668,28.708336,27.577778,29.366665,31.433336,31.141668,0.0,0.26666668,0.40833333,0.58750004,0.0,0.1875,0.0,0.0,0.058333334,0.59015155,0.175,0.29000005,0.25285715,0.63750005,1.1569444,1.9981601,3.2632575,3.2566664,3.195,1.2345835,1.980303,0.65000004,0.5833334,0.68125004,0.30833334,0.21666667,0.10000001,0.008333334,0.0,0.0,0.0125,0.8,0.16875,0.2,0.3416667,0.38125,0.275,0.0875,0.0,0.0,0.008333334,0.008333334,0.23125002,0.42499998,0.23750001,0.22500001,0.99999994,0.9166667,0.92499995,2.5375004,2.8500001,0.625,0.033333335,0.01875,0.48333335,0.125,0.45833334,0.0,0.01875,0.93333334,1.13125,0.39166665,0.01875,0.0,0.0,0.0,0.0,0.0,0.0,0.76250005,1.2583333,0.9062501,0.88333344,0.44166666,0.26874998,0.3,0.94375,0.575,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.008333334,0.05,0.016666668,0.0,0.083333336,0.7125001,0.9666667,0.8666667,0.8562499,0.5,0.35625002,0.6916666,0.6750001,1.6499999,2.3249998,2.25625,1.6583333,0.99375,0.6083333,0.29375002,0.07500001,0.00625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.375,14.166667,15.0375,15.325001,15.062502,18.083334,20.075,22.183332,23.175001,23.2,21.408335,17.762499,13.283333,9.225,5.6916666,3.425,1.8625,1.0666666,0.8125,0.7083333,0.77500004,0.80833334,0.67499995,0.13333334,0.29999998,0.11875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00625,0.041666668,0.30625,0.8166667,1.125,1.225,1.7333335,2.26875,3.2416668,4.9,6.0833335,6.9499993,9.225,12.3,14.46875,18.641666,22.587502,26.908333,31.787502,35.283333,36.391666,37.69375,38.350002,40.33125,41.225002,40.95,41.275,44.11667,46.781254,47.033333,48.05,47.333336,47.53125,44.666664,35.766663,28.168753,28.625,29.237501,26.966667,26.6875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.15,0.65555555,0.8666667,0.73333335,0.9666667,1.6659092,0.93333334,2.0666668,3.4000006,3.5227273,2.7222223,1.2111111,0.6833334,0.5222222,0.8666667,2.1444445,1.7750001,0.70000005,0.25555557,0.14166667,0.022222223,0.0,0.0,0.016666668,3.4555557,2.766667,2.2333333,2.2,1.2833335,1.5111113,2.2083335,1.7111111,0.37500003,0.022222223,0.24444446,1.2666667,2.0555556,1.1833334,0.8,0.5833334,1.7444444,1.8555555,4.916667,1.8666668,0.6166667,0.15555556,0.016666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.23333335,0.4916667,0.688889,1.5555556,2.116667,0.67777777,0.57500005,0.44444445,0.116666675,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08888889,0.4333333,0.875,0.44444448,0.6666667,0.9777778,0.09166667,0.0,0.3333333,0.12499999,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08888889,0.8833333,0.53333336,5.541667,24.966665,32.56667,24.583334,30.244446,36.925,41.5,40.791668,37.800003,34.566666,29.491669,25.011112,19.833336,14.555555,10.375,7.666667,6.2555556,5.775,4.7000003,3.825,4.2111115,3.5749998,3.6000001,2.775,2.488889,3.7444446,1.9583334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.022222223,0.12500001,0.51111114,0.6,0.7083334,0.88888896,1.3166666,1.3777778,1.2333333,1.6111112,2.1777778,2.9583337,3.8222225,5.7833333,9.844445,13.149999,14.822222,16.800001,20.72222,25.811113,30.3,33.600002,36.3,38.655552,38.550003,38.87778,38.455555,39.69167,42.65556,46.058334,47.688892,45.758335,40.522224,37.32222,31.533333,30.133333,34.141663,33.177776,32.06667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13333334,0.125,0.033333335,0.30833334,0.35555553,0.56666666,1.6666667,4.416667,3.7111108,1.9777777,0.68333334,1.2666667,0.6166667,0.51111114,1.9,2.0888891,1.6000001,0.36515152,0.033333335,0.175,0.0,0.025,0.0,0.43333334,2.3222222,3.1333332,3.6666667,3.0222223,1.5500002,2.788889,3.4916668,1.3777777,0.22222222,1.0166667,2.3222225,6.5083327,4.7111115,11.391668,7.6000004,2.211111,3.4833336,3.4444444,1.85,0.81111115,0.108333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.30833334,0.25555557,0.1,0.0,0.0,0.0,0.025,0.13333334,1.4444444,2.8499997,1.7555556,1.1083333,0.67777777,0.525,0.57777774,0.022222223,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.033333335,0.5,0.35833335,0.34444445,0.375,1.0111111,0.24166667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.044444446,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.1666667,5.833334,12.411112,17.275002,30.766666,40.755554,61.541668,64.57778,61.308342,61.155556,53.025,43.288887,35.522224,29.425001,24.555555,19.183332,14.500001,10.641668,7.666667,6.855556,5.908334,4.4333334,3.791667,5.2666664,6.0666666,5.1555557,5.716667,7.5555553,8.677778,4.0499997,0.5222222,0.26666665,0.7888889,0.32500002,0.11111111,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.022222223,0.07777778,0.5,1.1444445,0.9916667,0.6333334,0.2,0.4777778,0.68888885,1.4583333,2.6666667,3.0333335,3.455556,5.8416667,9.877777,11.049999,12.466667,15.300001,18.7,22.466667,26.666668,29.644444,32.566666,35.96667,37.600002,37.941666,37.67778,36.566666,37.766663,38.966667,36.622223,33.077778,24.891666,21.866667,29.775002,40.533333,39.316666,0.0,0.0,0.0,0.0,0.0,0.0,0.15,0.00625,0.083333336,0.2,0.3375,0.64166665,1.3500001,2.3249998,2.4125,2.2083333,3.5437498,3.3500001,2.8000002,1.3375,3.1583333,1.50625,0.9416667,0.45625,0.56666666,1.0166667,1.3499999,0.6111111,0.14375,0.3,0.38125002,1.1219698,1.96875,1.8833334,2.2083333,3.4375,4.425,5.3437505,3.05,1.6249998,2.125,1.5083333,0.28750002,0.8,2.9625,7.1,8.912499,7.2499995,6.508333,3.6374998,5.258333,4.7749996,2.1750002,1.6312499,1.1416668,0.17500001,0.0,0.0,0.0,0.083333336,0.17500001,0.016666668,0.0,0.0,0.0,0.6125,3.5166667,4.9000006,0.29166672,0.06875,0.0,0.0,0.0,0.075,1.19375,2.1,2.2875001,3.1083333,1.14375,0.5083333,0.24166666,0.025,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.43125004,0.075,0.025,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.33125,0.21666668,0.16874999,0.0,0.0,0.0,0.0,0.0125,0.125,0.23125,0.39166665,0.51666665,0.64374995,0.7333334,0.95,1.475,6.2499995,20.625,28.500002,39.725,53.575,68.5,70.81667,62.249996,56.19167,51.993755,43.941666,33.566666,24.262499,17.933334,13.80625,10.324999,7.2999997,5.208334,4.2583337,3.36875,2.1999998,1.83125,2.1416667,2.8874996,5.0333333,6.8812504,9.591667,8.049999,3.6687496,3.5333335,4.675,4.0333333,1.9937501,0.43333334,0.05,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.008333334,0.016666668,0.20625001,0.9250001,1.6875,2.6416667,3.13125,4.116667,7.012501,9.325,10.225,11.475,14.166667,20.556252,23.9,26.03125,28.1,29.658333,31.63125,32.11667,31.54375,29.375,29.468752,29.125,28.900002,27.100002,24.324999,19.43125,22.091667,33.518745,0.041666668,0.055555556,0.0,0.0,0.0,0.0,0.0,0.0,0.07777778,0.07777778,0.058333337,0.033333335,0.16666666,0.22222222,1.7416667,1.6666666,1.0083333,1.0555556,1.4555557,0.92499995,2.9222221,1.9666667,1.9666667,1.2333333,1.0111111,0.74444443,0.47500002,0.4222222,0.25,0.31111115,1.2083333,2.3222222,3.6750002,5.0333333,6.888889,6.2499995,4.366667,4.6916666,7.522222,6.4333334,1.9555557,0.85555565,0.5416666,0.38888893,1.2083335,1.0444444,2.5166667,3.3444445,4.711111,6.741667,7.244445,6.625,5.7555556,3.6833334,1.7555557,0.3166667,0.0,0.0,0.0,0.033333335,0.22500002,0.98888886,0.41666666,0.22222222,0.0,0.0,1.0555556,1.875,0.87777776,0.14166668,0.022222223,0.0,0.0,0.022222223,0.5083334,1.6666667,1.9666667,1.6777778,1.275,1.2222223,0.6,0.425,0.022222223,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.008333334,0.044444446,0.058333337,0.11111111,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05,0.22222221,0.34166667,0.011111111,0.2,0.06666667,0.0,0.0,0.0,0.0,0.033333335,0.11666667,0.17777778,0.25555557,0.3,0.35555556,0.7,1.488889,8.733333,19.811113,36.749996,50.45556,62.31111,64.99168,59.2,52.44167,43.555557,39.125004,31.288889,20.933332,14.216666,9.866667,7.3666673,5.5222225,4.3583336,3.677778,3.2555556,2.5583334,1.511111,1.3583333,1.3000002,1.575,1.8333334,2.8666668,3.8444443,2.5222223,2.9083335,6.1000004,7.266667,6.444444,3.8583333,1.2444444,0.51111114,0.14166667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.058333337,0.34444442,0.8333334,1.3777778,2.0,2.711111,3.6666665,5.8222227,8.3,9.700001,10.466666,11.474999,16.366667,21.449999,24.566668,24.711111,23.208334,22.544445,22.683334,22.333334,21.641666,22.955555,23.133333,24.85,23.833334,25.341667,21.011112,23.533333,0.00625,0.008333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.008333334,0.55625,1.5166667,3.1624997,1.975,0.725,0.3,2.1333334,0.75625,1.0333333,1.40625,1.2333333,0.7,0.53125,0.24166669,0.43750006,0.35,0.31875002,1.125,3.1562502,6.333333,8.45,9.95,9.725,7.18125,5.675,3.8437505,5.116667,2.6916666,0.40000004,0.3166667,0.7375,1.4916664,0.93125004,0.39166668,0.6416667,3.4437501,5.916667,5.1375,4.958333,5.775,4.9583335,1.5625,0.69166666,0.025,0.0,0.0,0.35625,0.14166667,0.21374999,0.058333337,0.0,0.0,0.0,0.9625001,0.7083334,0.025,0.0,0.0,0.0,0.0,0.23125002,0.7083334,1.0500001,2.4750001,1.09375,0.9166666,0.9583334,1.34375,2.2166667,0.48125,0.0,0.0,0.0,0.0,0.0,0.0,0.8125,1.3916667,0.67499995,0.9333334,1.13125,1.1166667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025,0.5083334,1.29375,2.1416667,2.8000002,3.60625,4.491667,4.69375,3.1166668,7.45,16.416668,25.0125,29.8,38.316666,40.800003,33.124996,30.00625,24.783335,20.45625,14.349999,10.066666,4.9125,2.8,4.0,5.425,6.79375,7.125,7.1833334,4.8187504,3.6750002,2.1187499,1.3083334,1.2687498,1.5166668,1.4625,1.125,1.1499999,1.71875,4.691666,4.6625,4.0833335,4.4875,4.358333,2.3000002,0.5125,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.50625,0.083333336,0.33749998,0.7583333,1.38125,1.9583334,2.64375,3.866667,5.25,7.2999997,9.208334,9.78125,10.5,11.7,15.299999,18.325,19.1625,19.433334,18.11875,17.091667,16.3125,15.241665,15.758333,18.39375,21.916668,22.525,21.016666,17.762499,0.041666668,0.06666667,0.022222223,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.3888889,1.4166666,1.5000001,2.588889,2.0,1.9000001,0.55833334,1.0555557,2.291667,2.5333333,1.6666667,1.3916667,0.7555556,0.41666672,0.44444445,0.53333336,0.43333334,1.3500001,3.6888885,4.9222226,8.099999,10.6888895,10.641666,9.888889,6.416667,2.788889,2.1666667,1.5166667,0.6666667,1.1,0.6666667,0.54166675,0.23333335,0.06666667,0.46666664,1.8333334,2.3166666,3.1555557,2.4833333,3.7555556,3.2749999,0.7,0.7777778,0.0,0.0,0.0,0.43333334,0.06666667,0.1,0.07777778,0.0,0.0,0.35,1.7333335,0.016666668,0.0,0.0,0.0,0.0,0.16666667,0.0,0.3166667,1.2555556,2.6000001,1.5888891,1.2555557,0.9083333,1.0888889,1.0083334,0.0,0.033333335,0.055555556,0.022222223,0.033333335,0.0,0.0,0.011111111,0.18333334,0.08888889,0.22500001,0.48888892,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.044444446,0.25833333,1.0,2.1916668,3.5888891,4.5444446,5.65,6.877778,6.0666666,8.066667,14.558333,18.722221,16.358334,14.822223,17.544443,18.941666,18.277775,13.266667,8.544445,8.041667,6.6333337,6.7111115,8.425,15.233334,17.9,13.722221,6.225001,3.688889,1.4222223,1.05,1.1666666,1.95,1.8333333,0.9666667,0.22222224,0.0,0.0,0.44444448,1.1166667,1.8555555,2.891667,5.9444447,5.6999993,2.2444446,0.8444445,0.13333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.20833333,0.5222222,0.4916667,0.42222226,1.3833333,2.3777778,3.3,5.258333,6.7777777,8.333332,8.966666,9.483334,10.033333,10.277778,11.400002,12.066667,13.108334,12.588888,12.625,13.411112,12.98889,11.375,11.444445,14.166666,16.055555,14.658336,1.1625001,0.8583334,0.3166667,0.19375002,0.24166669,0.38125002,0.3916667,0.1,0.041666668,0.09166667,0.050000004,0.06666667,0.06875,0.4416667,1.0375001,1.3833334,1.4312501,0.56666666,1.4999998,2.0375,1.5916667,0.55,0.8416667,0.86875,1.2499999,1.6416665,2.35625,3.1750002,3.4687502,3.3333333,1.6437502,1.1666667,1.53125,1.5749999,2.3666666,3.5374997,3.2416666,5.68125,6.166666,6.787501,4.3333335,1.7583334,0.9937499,1.5083334,2.0375,2.2916665,0.68125004,0.016666668,0.008333334,0.03125,0.29999998,1.2391666,0.8781818,0.78166664,0.40833333,0.33125,1.55,0.28333333,0.15,0.0,0.0,0.0,0.175,0.05,0.041666668,0.00625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.087500006,0.5166667,3.0124998,7.058334,3.4666667,1.29375,0.05,0.00625,0.083333336,0.03125,0.08333334,0.21666665,0.40000004,0.14166667,0.0375,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.056250002,0.17500001,0.7875,1.2916666,1.46875,2.1000001,2.6666665,3.3687499,5.341667,3.6249998,3.1916666,6.8125,6.950001,10.012501,20.95,29.933336,32.743755,27.599998,16.575,7.391667,5.96875,7.216667,8.85,8.793751,5.1833334,5.5187497,6.333333,1.93125,0.20000003,0.116666675,0.0,0.0,0.03125,0.12500001,0.17500001,0.14166668,0.0125,0.016666668,0.26666668,0.75625,1.275,2.1750002,2.7666671,1.75,0.75833327,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.041666668,0.09375001,0.041666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0625,0.13333334,0.28125003,0.65833336,0.82500005,1.1166667,2.0416667,3.75,5.9833336,8.087501,9.283333,9.01875,9.041666,9.333333,9.85,10.116667,10.36875,9.858334,7.8250003,6.7333336,7.6583333,8.375,8.833333,9.418751,10.150002,10.93125,3.55,4.3666663,4.9888887,3.4916668,1.8777777,1.4749999,0.92222226,0.65,0.36666667,0.44444442,0.16666669,0.07777778,0.108333334,0.28888887,0.9083333,0.7777778,1.0999999,1.3,3.0555558,1.4166667,0.79999995,1.1166667,1.1777778,0.875,0.5222222,0.6666667,1.7333333,3.6222224,7.275,10.922223,11.191667,7.088889,3.4,2.9333334,1.7777779,2.25,2.411111,1.4234848,1.2333333,2.4,1.5222223,1.2,2.225,4.0333333,2.4083333,2.266667,1.4083334,0.24444444,0.011111111,0.0,0.022222223,0.19166669,0.3888889,0.35000002,0.26666668,0.25,0.08888889,0.1,1.0333333,0.6,0.0,0.0,0.016666668,0.14444445,0.0,0.008333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.7166667,1.5888889,4.475,4.766667,2.2222223,1.7916667,2.9555554,0.425,0.033333335,0.17500003,0.18888889,0.70000005,2.2500002,1.1,0.050000004,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025,0.22222222,0.51666665,0.8333333,1.1083333,1.3666667,1.6111112,2.25,2.0555556,4.5,9.755555,8.683332,8.388889,10.811111,16.408333,14.48889,9.141666,4.411111,4.516667,10.222221,17.216667,26.655556,35.077778,38.11667,35.13333,29.516668,22.88889,26.983334,24.344442,21.300001,14.633333,4.922222,1.4916668,1.8777778,1.1583333,0.18888889,0.32222223,0.24166669,0.2,0.1,0.044444446,0.016666668,0.0,0.0,0.022222223,0.3555556,1.2333333,1.7555556,1.4916667,0.67777777,0.675,0.45555556,0.28888887,0.35,0.32222223,0.2,0.18888889,0.09166667,0.011111111,0.0,0.0,0.0,0.016666668,0.044444446,0.008333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.12222223,0.19166668,0.6555555,0.8166666,0.97777784,1.3777779,2.3833334,4.0555553,5.908334,8.055555,9.733334,10.677777,10.300001,9.75,9.377777,8.95,7.5444446,5.908334,4.788889,3.988889,4.2583337,5.233333,5.6916666,5.377778,6.0416665,2.4333334,2.3666668,1.5777777,3.9166667,3.4444444,2.1583333,0.8777778,0.9833334,0.73333335,0.9888889,0.5333333,0.41111112,0.34166667,0.5111111,0.6583333,0.7666667,0.92499995,2.388889,6.4777775,5.508333,2.977778,2.825,1.8666668,2.25,2.4888887,2.7333333,4.366667,7.8444448,10.183333,14.911111,18.841667,19.500002,14.075,8.066667,4.588889,2.6666665,1.6999999,1.0472223,0.48055553,0.4027778,0.14444445,0.18888889,0.2439394,1.6222222,8.833334,7.188889,0.8833333,0.58888894,0.36666664,0.10000001,0.0,0.23333335,0.0,0.04166667,0.13333334,0.05,0.044444446,0.0888889,0.116666675,0.46666667,0.0,0.0,0.0,0.0,0.022222223,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.008333334,0.3,1.4666668,2.5111113,3.4166667,3.2111115,2.711111,2.0333333,1.3111112,1.3416667,0.1777778,0.04166667,0.35555556,1.1111112,0.99166673,1.2222222,0.55,0.13333334,0.033333335,0.0,0.0,0.0,0.0,0.0,0.044444446,0.083333336,0.11111111,0.15833333,0.06666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05,0.3111111,0.84166676,1.6888887,2.4666667,3.366667,4.522223,5.5750003,5.0888886,6.6250005,12.966668,13.375001,11.855556,13.055556,17.650003,12.555556,7.083333,4.288889,3.8416667,7.2666664,12.875002,23.655556,38.144444,54.450005,61.733337,61.366665,52.966667,42.15,32.233334,23.811111,14.141667,6.111111,4.141667,3.2333333,1.9250001,3.688889,5.077778,4.566667,3.733333,3.1000004,2.277778,1.3249999,0.7,0.40833336,0.45555562,0.87777776,1.2166667,0.87777776,0.8,1.8444446,3.9916663,4.133333,3.3888888,2.4833336,1.4555556,1.05,0.8444445,0.625,0.37777779,0.24166669,0.08888889,0.022222223,0.0,0.0,0.0,0.0,0.0,0.11111112,0.2777778,0.23333333,0.13333334,0.14166667,0.54444444,0.7583334,1.0111111,1.1666665,1.3222224,1.3000001,1.525,2.1333334,3.0333335,4.5333333,5.9916663,8.055555,9.48889,9.558334,8.322222,7.0166674,6.5777783,5.416667,4.4333334,3.5555558,3.4750001,3.6777778,4.158334,4.177778,4.15,4.025,4.9083333,5.116667,5.50625,4.9833336,4.5750003,2.1666665,2.31875,2.8750005,3.8666668,4.55,5.4333334,5.5062504,4.583333,2.71875,1.4583334,1.0375,2.3583336,4.841667,3.1374998,1.7333333,1.60625,1.075,1.63125,3.2083335,4.4500003,6.45625,9.349999,11.45,12.575,16.7875,25.125002,32.68125,29.658335,20.658335,11.550001,5.143182,2.0770833,0.83500004,0.27272728,0.043181818,0.016666668,0.043750003,0.59166664,1.5812498,1.4583333,1.2187499,2.15,2.725,2.3375,1.4583335,8.81875,9.325001,0.20000002,0.1,0.0,0.016666668,0.075,0.01875,0.23333333,0.80625004,1.1666667,1.6875,0.76666665,0.4166667,0.056250002,0.05,0.14375,0.033333335,0.0,0.0,0.0,0.0,0.0,0.09375,0.6583334,1.34375,2.3,3.10625,2.675,2.9083333,2.81875,2.6583333,1.35,0.4333334,0.14375001,0.25,1.95,3.0625002,3.9333334,3.53125,2.4833333,2.1937501,2.2,1.7,0.96666676,0.56666666,0.21250002,0.116666675,0.17500001,0.25833333,0.36875,0.21666667,0.19166668,0.28125,0.1,0.025,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025,0.10000001,0.325,0.53124994,0.6833332,1.0083334,1.3374999,1.7749999,1.8812499,1.4333334,2.5625,3.9333332,4.5583334,3.50625,1.6166667,2.9,3.15,4.0125,5.283333,7.6625,12.358333,24.525002,36.43125,40.458332,44.85625,44.799995,33.875004,21.958334,14.349998,8.73125,6.1,7.8375,12.291666,12.443749,21.933334,28.5,24.65625,17.166668,13.137501,9.558334,5.85625,3.2833335,1.9437503,0.9833333,0.675,0.35000002,0.55833334,0.56875,0.73333335,0.99375004,1.5333333,1.9416668,2.3249998,3.4666667,2.8125,1.4416666,1.4562501,1.4833333,1.35625,1.2083334,1.0083333,0.90625006,0.8666667,0.86875,0.96666664,0.43750003,0.275,0.22500001,0.84375,1.1166667,0.95625,0.7833334,0.5375,0.59999996,0.79375,0.85,0.9166666,1.2375001,1.1916668,1.3875,1.7916667,2.5437503,3.9750001,5.1916666,6.65,6.9249997,6.0375004,5.1833334,4.762501,4.116667,3.6583333,3.3625002,3.4416666,3.7625,3.7916665,3.21875,2.325,3.5,2.788889,3.5916667,4.7777777,5.708333,3.288889,3.6583335,5.4333334,7.9333334,10.325,13.400001,21.591665,26.611113,17.183332,8.244445,6.3666673,4.9888883,3.1444447,0.5,0.07777778,0.050000004,0.08888889,0.55833334,1.7444444,3.3222222,6.9250007,12.766666,13.391666,11.622223,9.166666,11.9,26.900003,40.144444,37.155556,26.708336,16.9,8.558332,4.077778,0.9765152,0.331746,0.2793651,0.17045456,0.33333334,0.7250001,1.0,1.975,4.088889,4.266667,5.0666666,3.4333334,2.7416668,0.8777778,0.25000003,0.28888887,0.025000002,0.0,0.0,0.016666668,0.022222223,0.6166667,1.6777778,2.6750002,3.2999997,2.1333332,0.7833333,0.5777778,0.79999995,0.25555557,0.016666668,0.0,0.0,0.022222223,0.0,0.0,0.0,0.19166669,1.4666667,3.8500001,4.822222,3.5333333,1.2416667,2.8444445,3.2000003,2.0555556,0.57500005,0.0,0.5555556,0.5750001,2.7333336,8.041666,7.3,6.4333334,3.8555555,1.9083335,0.77777785,0.2777778,0.07500001,0.011111111,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.116666675,0.022222223,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016666668,0.06666667,0.1,0.0,0.0,0.0,0.10000001,0.46666664,0.78888893,0.73333335,2.5888891,5.65,10.4777775,16.016666,24.177776,23.622221,17.058332,14.744445,20.708332,21.07778,12.258333,9.1,9.1888895,9.608334,12.977778,15.541666,18.744444,30.291668,51.799995,73.86667,74.90835,55.08889,51.300003,48.02222,31.825,15.98889,7.2999997,3.3444443,1.6888889,1.6333333,2.3666668,2.225,2.288889,1.7416668,2.4222221,3.8555555,4.508333,6.8888893,7.266667,4.7777777,4.0166664,5.577778,6.4083333,5.0111113,4.1333337,3.15,1.6555555,0.4416667,0.36666667,0.49166667,0.0,0.0,0.116666675,0.38888887,1.1916667,1.188889,0.65833336,0.82222223,1.0916666,0.9222223,1.0777779,1.2333333,1.1666667,1.3000002,1.3444445,1.2750001,1.6333334,2.8000002,4.475,5.8888893,6.108333,5.433334,4.45,3.6222224,3.0444446,2.791667,2.9444447,2.7583332,2.311111,2.4666667,1.6750001,0.9,2.6000001,2.4812498,3.3583333,5.35625,6.65,11.099999,11.733334,11.608334,11.337501,10.183333,9.075001,9.4,7.3937497,5.3,7.95,10.241667,8.975,9.2875,6.308334,3.0500002,1.0333334,0.71875006,1.1833333,2.1750002,5.25625,11.175,10.2875,9.875,7.637501,7.5250006,14.150001,28.766666,35.883335,32.125,19.141668,11.587501,8.55,6.3875,4.525,3.5583332,1.6920832,0.95833325,0.34375,0.13333334,1.9062501,3.8083334,5.1250005,4.7000003,3.1,0.47500002,0.0,0.48125002,0.40000004,0.1875,0.0,0.016666668,0.0,0.0,0.10625,1.3166666,3.2625,5.683333,5.5083337,1.50625,0.5083333,0.88125,1.3083334,0.50625,0.025,0.0,0.116666675,0.28333336,0.46875,0.11666667,0.03125,0.22500001,1.54375,3.8916667,6.1083336,3.4562502,1.275,2.28125,4.483333,2.7625,1.1166667,0.18333334,0.2375,0.43333337,1.2062501,1.5333334,1.5812501,1.3916665,0.5124999,0.27499998,0.09166667,0.00625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05,1.525,1.91875,0.2916667,0.18333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.20833334,0.5875,0.38333333,0.0625,0.0,0.0125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.125,1.2187501,2.8083334,5.2125,6.5666666,12.09375,19.091667,25.475,19.19375,13.124999,6.73125,7.0000005,13.3125,20.350002,27.091665,37.15,33.866665,26.6625,34.399998,62.906254,108.86668,111.03334,106.08125,92.450005,78.52501,62.783337,51.274998,40.24167,25.2625,11.750001,6.1333337,3.8875003,4.083333,3.8562498,3.8166666,3.4624999,3.016667,2.625,2.1000001,2.0416667,2.575,3.525,3.275,2.6499999,2.46875,1.9416666,1.6499999,1.5874999,0.91666675,0.26875,0.0,0.14375003,0.225,0.30833337,0.1875,0.116666675,0.76875,1.25,0.95625,1.2666665,1.5874999,1.4250001,1.5166667,1.75,1.6916667,1.30625,1.3916668,1.4000001,1.6,2.1000001,3.0750003,4.908334,6.125,5.55,4.1,3.2000003,3.1750002,3.7875001,4.0416665,4.1375003,4.7999997,4.24375,2.7250001,1.7333333,0.98888886,2.9999998,5.733334,6.675,6.3444448,7.733333,6.9222217,5.355555,6.8166666,6.166667,7.1749997,9.722221,6.6083336,8.266667,8.833334,13.711112,10.066667,10.191666,19.5,10.766667,5.211111,1.775,0.98888886,1.4666667,2.55,4.4,9.658334,6.333334,6.1749997,8.066668,5.708334,11.933332,25.277779,28.983334,20.822224,9.6,8.233334,7.575001,7.8666663,8.033334,5.5666676,1.1666666,0.48333335,0.37777779,0.325,2.1333334,3.9222221,3.4500003,3.588889,0.6916667,0.0,0.26666665,0.33333334,0.47500002,0.033333335,0.15555556,0.16666666,0.033333335,0.0,0.8333334,2.9083333,6.433333,7.6,3.2000003,0.7111111,0.825,2.2222223,1.3166667,0.3,0.13333334,0.07777778,0.3888889,0.975,1.2,0.8416667,0.32222223,0.41666672,1.5666668,3.3111115,5.2333336,4.088889,1.5583335,1.1444445,1.9333334,2.377778,1.9666668,0.7083333,0.11111111,0.10000001,0.07777778,0.016666668,0.011111111,0.0,0.0,0.11111111,0.058333337,0.044444446,0.008333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.6888889,2.4833336,6.9999995,1.8416667,0.7222222,0.17777778,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.041666668,0.0,0.0,0.0,0.0,0.0,0.54444444,0.5083333,0.36666667,0.0,0.022222223,0.15000002,0.8333333,0.15555555,0.0,0.0,0.0,0.0,0.0,0.055555556,0.025,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.4888889,2.6,5.6777773,10.366666,13.122221,22.616669,39.58889,54.644447,58.05,56.411114,53.425,45.922222,42.86666,36.95556,29.944447,22.225002,18.711111,25.508331,40.577778,70.65,94.877785,99.00001,96.10833,87.68889,81.01666,71.85556,64.54167,59.533333,43.841667,25.933334,14.633334,10.991667,9.244446,5.675,7.4555554,12.900002,9.988889,5.8,2.1250002,3.5,13.075001,12.011111,9.016668,5.0666666,1.1500001,0.24444443,0.0,0.0,0.0,0.0,0.0,0.0,0.033333335,0.33333337,0.8416667,1.1666666,1.3583333,1.4444444,1.2,1.7666667,3.125,3.5666668,3.455556,3.1000001,3.0333335,2.2666667,1.588889,1.4166667,1.6222223,1.8777778,2.5416663,3.8888888,5.3083334,5.9444447,5.133333,3.9,3.4333332,3.875,4.0555553,4.241667,5.3444443,4.7166667,9.34375,7.0,5.158333,3.53125,3.641667,6.1499996,6.95,7.3875,6.791667,4.075,5.19375,5.8250003,7.325,5.3083334,3.4,3.4916666,6.500001,6.958334,4.283334,4.35,7.241667,7.31875,6.391667,3.8250003,0.7416667,0.35833332,0.78125006,1.4833333,4.1,4.3416667,3.2125,4.7833333,3.5187502,3.05,10.108334,19.3125,14.95,8.84375,4.391667,4.6062503,6.658333,8.099999,8.35625,5.2916665,2.09375,3.5,2.475,2.5249999,3.0416665,2.375,2.7833333,0.88124996,0.008333334,0.08125001,0.21666668,0.7375,0.041666668,0.4166667,0.57500005,0.20833334,0.0125,0.075,2.0375001,5.3916664,10.05,5.79375,2.05,0.9625,1.6333334,2.2625,1.3666666,0.64375,0.33333334,0.033333335,0.3375,0.9833333,1.5875001,1.9333334,2.0062501,1.2166668,0.9499999,1.8875,1.8666668,2.5874999,1.2333333,2.025,3.1666667,1.2666668,0.35,0.1,0.0,0.0,0.0,0.0,0.0,0.025000002,0.3,0.15625001,0.09166667,0.0125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13333334,0.0875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06666667,0.081250004,0.0,0.0,0.0,0.0125,0.25,0.38333333,0.35625,0.116666675,0.0,0.22500002,1.0875001,2.175,0.21666667,0.0125,0.05,0.3125,0.125,0.28125,0.05,0.0,0.28333333,0.91666675,0.2875,0.0,0.075,0.66666675,0.49374998,0.2,0.033333335,0.03125,0.0,0.125,0.62499994,1.53125,4.7166667,10.0625,32.325,45.500004,44.6,26.19167,37.156246,41.600002,29.0125,21.550003,27.683334,37.125,43.099995,53.55,44.966667,42.918747,59.125004,73.96667,79.387505,81.725006,75.91875,66.625,64.0375,57.50833,47.4375,34.574997,29.366667,29.987501,32.125,29.743748,20.350002,12.193751,6.1083336,3.4666667,2.3187501,1.375,2.4875,4.2,3.0937502,3.3666666,2.90625,2.7,1.4000001,0.25625,0.175,0.175,0.125,0.10625,0.083333336,0.06666667,0.118750006,0.5416666,1.4562501,2.1666667,2.4875,2.3583333,2.6125002,3.3333335,3.5916667,3.1875,2.4333334,1.7250001,1.4166666,1.49375,1.7333335,1.7166667,1.9250001,2.5333335,3.86875,4.258333,4.4875,3.85,3.0249999,3.2937498,4.3,5.2562504,5.625,5.6687503,16.025,13.566667,10.900001,8.95,7.9666667,7.25,8.266666,9.366667,9.088888,5.1333337,5.1916666,5.4,5.450001,4.877778,3.5916672,3.1000001,1.8666667,1.3888888,3.022222,2.1333332,2.288889,0.97499996,0.32222223,0.15,0.0,0.0,0.0,0.0,0.0,0.9222223,1.7583334,2.677778,2.9916668,1.7,2.2555556,8.625,10.58889,8.008334,3.7666667,2.5916667,4.7000003,6.4333334,10.075001,8.8111105,5.5500007,15.033333,13.25,7.177778,2.5444446,1.8333333,1.6444446,1.0250001,0.044444446,0.016666668,0.044444446,0.7083334,0.11111111,0.2111111,0.76666665,0.8555556,0.108333334,0.011111111,0.94166666,3.2888887,5.0111113,4.0750003,1.1555556,0.35833335,1.3,3.0749998,2.3,1.8833334,0.40000004,0.0,0.008333334,0.055555556,0.81666666,2.2555556,2.625,2.7555554,1.2888889,0.625,1.3222222,1.0416666,0.18888889,1.1916667,1.7111112,2.311111,1.6833334,0.24444444,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08888889,0.008333334,0.0,0.0,0.0,0.05,0.12222223,0.12222224,0.13333334,0.0,0.033333335,0.48888892,3.5916667,1.7111111,0.6,0.5083334,0.9555556,0.45000002,0.81111115,0.22500001,0.0,0.075,0.1,0.022222223,0.016666668,0.0,0.50833327,2.7444446,2.0916667,0.4222222,0.6,1.8166667,1.0333334,1.225,2.6555555,4.966666,8.577778,16.033335,30.955555,40.544445,47.324997,34.988888,35.408333,43.955555,53.024998,55.422226,58.35556,49.850006,32.13333,35.000004,44.77778,91.41666,109.577774,101.77778,80.666664,64.477776,55.591667,57.62222,59.274994,53.555557,40.508335,31.300001,26.02222,23.041666,23.211113,29.45833,20.488888,11.133333,7.5,7.588889,6.8833337,3.4666665,1.2833334,0.7777778,1.7,3.5666666,5.9833336,6.5,4.5222225,4.8083334,5.7222223,5.008333,3.7,3.341667,2.7555556,2.5555556,1.7750001,0.77777785,1.4999999,2.577778,3.8166668,4.055556,3.641667,3.3666666,2.9555557,2.2416666,1.1777778,0.67499995,0.5888889,1.0333333,1.6777779,1.5555557,1.0666666,0.9,1.0083334,1.8444445,2.2416668,2.9666667,3.2444444,3.9583333,6.0222225,8.383332,10.566667,10.591667,12.25,16.266668,15.222222,12.466667,8.744444,7.95,4.977778,8.875,7.922222,5.933334,6.5916667,8.9777775,9.200001,8.911112,6.191666,1.1,0.47500002,0.90000004,1.3444444,1.4166666,1.0,0.058333337,0.17777778,0.23333335,0.25555554,0.26666668,0.18333334,0.13333334,0.0,0.98888886,3.4583335,5.088889,3.4333334,2.6222222,3.8222222,3.7250001,8.266666,8.408333,5.977778,4.2000003,5.5333333,7.3,12.65,13.677777,7.9500003,8.2,12.058332,2.7222223,1.6777778,2.0416667,1.0333334,0.69166666,0.044444446,0.033333335,0.06666667,0.041666668,0.0,0.011111111,0.9333334,1.1111112,0.39166668,0.044444446,0.16666667,0.5888889,0.92222226,1.7833332,0.7444445,0.083333336,1.1,2.8000002,1.3111111,0.43333337,0.22222221,0.044444446,0.0,0.0,0.09166667,0.8222223,3.375,3.6444445,2.266667,1.9916668,0.9333334,0.34166673,0.0,0.14166668,0.6777778,1.5111111,1.3916667,2.2666664,1.275,0.6,0.008333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.022222223,0.041666668,0.033333335,0.06666667,0.13333334,0.15555556,0.13333334,3.2888892,2.5750003,0.76666665,1.1333333,1.5333332,1.1888889,0.51666677,0.7777778,0.0,0.0,0.125,0.0,0.6333333,0.55,0.7888889,0.116666675,1.611111,2.7499998,0.06666667,1.5000001,3.9916668,2.5888886,2.3416665,4.3000007,7.3583336,12.688889,27.033333,52.0,75.399994,94.575005,86.700005,51.29167,40.922226,42.36666,41.34444,42.977783,41.458332,33.9,29.775002,32.755554,51.55,51.6,42.788887,33.925,35.355556,33.608334,36.744446,38.716667,36.4,27.28333,24.111113,20.644445,18.141666,18.466667,20.983332,22.355556,21.341667,15.377778,10.6888895,7.216666,3.1444445,0.9833333,0.41111112,0.6666666,1.1222223,1.7750001,3.1000001,5.0111117,7.450001,8.8,7.7916665,6.177778,5.0666666,4.111111,3.0555556,2.4,1.588889,1.7916667,3.3222222,5.275,6.166667,6.4083333,6.0222225,5.1111116,3.7833333,2.3000002,1.5666667,1.3111112,1.2083335,0.788889,0.98888886,1.1583334,1.3666667,1.4083334,1.5777777,2.1833336,3.4444447,4.2777777,3.9916666,5.211111,6.6416674,8.933332,10.341667,8.44375,6.0583334,8.183333,4.8,2.9666667,1.7562501,0.68333334,0.45000002,1.4166667,2.6666665,4.3499994,9.191667,9.481251,7.2666664,3.7500005,0.65833336,0.0625,0.033333335,0.0,0.03125,2.6583333,2.0500002,4.9166665,7.6875,6.2583327,3.3583336,1.9625001,1.6833334,3.0187502,2.7583334,3.9937499,6.6,6.0874996,5.5250006,3.325,4.674999,5.591667,8.1625,7.4833336,5.61875,5.491667,8.841667,14.343751,18.041666,14.581249,7.091666,3.05,0.041666668,0.38333336,1.3,2.25,0.58125,0.09166667,0.0375,0.14166668,0.0375,0.0,0.0,0.9000001,1.2916667,0.75624996,0.13333334,0.0,0.0,0.058333337,0.78124994,0.3416667,0.0375,0.40833333,0.7687501,0.7833333,0.21875,0.0,0.0,0.3375,0.35833335,0.2125,0.69166666,3.2875001,3.1333334,1.9250001,1.6874998,4.05,1.225,0.34166667,0.0,0.38333336,0.19166666,0.30624998,0.33333337,0.82500017,0.38333333,0.0125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.008333334,0.0,0.0,0.008333334,0.10000001,0.20833336,1.7500001,2.4333334,0.45,0.5416667,0.88333327,0.96875,0.45000002,0.51250005,0.125,0.18125,1.025,1.0875001,0.55,2.0666666,1.9875002,0.47500002,0.4125,1.95,0.9125,1.3,3.9999998,5.7,3.6583338,6.33125,12.216667,20.03125,30.516668,41.025,51.7,58.46667,63.212505,54.38333,36.349995,22.508331,17.59375,15.974999,22.133335,23.18125,21.808334,17.95625,17.9,32.2625,40.049995,34.775,29.937502,24.725002,20.85625,18.483334,16.26875,16.591667,14.087502,11.341667,11.916666,14.09375,16.25,18.46875,21.808336,24.406248,23.241667,16.066666,7.0625005,2.1166666,0.93750006,1.2416666,2.4437501,3.0,3.54375,4.391667,3.7750003,3.99375,3.5499997,2.5125,2.425,2.59375,2.65,2.8083332,2.3749998,3.9333334,4.45625,5.1166677,5.6125,6.3416677,6.793751,6.5750003,6.3,5.8875003,4.8250003,4.00625,3.2916667,3.08125,2.7416666,1.8166667,1.3875002,1.1250001,0.7875001,0.9000001,1.48125,2.8083334,4.833333,5.2124996,6.0666666,6.9125,7.7333336,9.362499,9.941667,6.244445,8.466666,5.4166665,2.577778,2.3,2.411111,2.0083332,0.7444445,0.31111112,1.1916667,2.2444446,4.6833334,4.0,2.5666666,2.3333335,0.7916667,0.44444445,0.36666667,0.375,0.1,0.16666667,1.7111112,2.5833335,2.311111,1.0666667,0.44166672,0.07777778,0.14166668,0.0,0.26666668,1.0444446,3.9166665,11.933333,13.58889,6.4416666,5.677778,6.891667,7.588889,5.4833336,4.988889,9.955556,15.45,19.27778,13.841666,7.4333334,4.0000005,0.34444442,0.0,0.65000004,3.7555554,2.1916668,0.36666667,0.025000002,0.14444445,0.09166667,0.0,0.0,0.5083333,1.3666666,2.708333,0.2,0.033333335,0.0,0.0,0.025,0.0,0.0,0.13333334,0.5833334,0.0,0.0,0.0,0.0,0.0,0.11111111,0.575,0.65555555,1.5916667,0.73333335,1.1222223,0.15833333,1.4777778,2.5166667,1.777778,0.0,0.9777778,0.0,0.0,0.0,0.07500001,0.15555556,0.025000002,0.18888889,0.025000002,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.2777778,0.2,0.14444445,0.0,0.0,0.033333335,0.12500001,0.18888889,0.46666664,0.10000001,0.083333336,0.11111112,0.24444446,0.058333334,0.0888889,0.058333334,0.3111111,0.7666667,1.077778,0.5916667,0.05555556,0.7777778,0.75000006,0.41111112,1.3500001,2.8222222,5.0250006,10.155556,11.455557,7.883333,2.0333333,2.3666668,3.8444448,6.675,8.1,15.925,22.211111,25.455557,25.091667,20.244446,12.166667,5.9555554,4.458334,6.055556,9.855556,10.016666,19.377777,24.558334,28.177776,21.983332,20.355555,20.455555,22.508331,22.377777,23.75,21.933334,21.991667,18.366667,12.483334,7.5888896,5.388889,7.1416674,8.122223,8.341667,9.044445,11.524999,13.433334,11.844445,5.6166663,3.1666667,4.9666667,6.7444444,7.133333,15.711112,22.666668,19.98889,13.98889,9.55,7.988889,7.125,5.5222225,2.4833336,1.2,1.1111112,1.45,1.7333333,3.2833328,4.755555,4.3333335,5.3777776,5.2083335,4.7333336,4.4555554,4.633333,4.7666664,4.925,4.6555557,4.166667,4.411111,4.0222225,2.95,3.0666668,3.0333333,2.1888888,1.3583333,2.7666667,4.677778,5.5250006,6.466667,6.241667,6.7000003,6.2583337,5.8624997,3.791667,2.4,3.3500004,5.383334,4.59375,2.1666665,0.88750005,2.625,10.958332,10.243751,9.575,6.9125004,4.108333,1.6249998,0.7583334,1.54375,3.1416671,4.8583336,4.43125,2.9833333,0.925,0.73333335,0.83124995,0.65000004,0.34166664,0.12500001,0.10833334,0.112500004,0.108333334,0.23124997,0.6500001,2.2625,6.0416665,9.891667,11.356251,7.9333334,10.19375,8.450001,5.3,7.041667,12.408334,15.975,18.166668,10.831251,7.116667,3.1,0.65000004,0.125,0.1,3.1916668,4.7999997,2.025,0.25,0.16666667,0.25625002,0.025,0.0,0.21875,0.74999994,1.38125,0.36666667,0.28750002,0.0,0.0,0.0,0.0,0.0,2.1833334,1.86875,0.20000002,0.0,0.0,0.0,0.0,0.0,0.03125,0.71666676,0.9125001,0.825,0.8083334,0.043750003,0.0,0.04375,0.30833337,0.2,0.0,0.0,0.00625,0.058333337,0.43750006,0.625,0.1375,0.22500001,0.01875,0.4416667,0.108333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.9312503,0.5083333,0.15625001,0.14166668,0.041666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025,0.37499997,0.9416667,0.78125006,0.43333334,0.05,0.0,0.05,0.09375001,0.025,0.00625,0.016666668,0.0,0.0,0.0,0.2375,0.54999995,1.01875,1.2166667,0.51875,0.13333334,0.03125,0.116666675,0.875,0.74375004,0.425,0.95625,1.9083333,2.89375,9.941666,10.774999,5.9125,4.7250004,6.2249994,12.025,18.5,24.666668,24.59375,19.025002,15.241666,12.231249,7.333334,2.7124999,4.8500004,11.993751,27.416668,27.333332,15.174999,16.391665,22.850002,24.058336,18.95,15.291667,18.46667,13.793751,14.558332,15.699999,13.900001,11.03125,9.025,7.1749997,4.233333,3.3583336,3.6312504,2.3999999,1.20625,0.625,1.04375,1.4583334,1.5166667,1.3625001,1.725,3.6875,6.8,7.64375,13.6,28.800001,30.841665,22.783333,17.450003,22.641666,21.225,13.066666,6.8,3.5416665,2.5333333,2.3625,1.9833333,1.425,2.5583334,4.9000006,5.35,5.0750003,4.95,4.5,3.6875,3.5499997,3.9249997,4.8,5.01875,4.658333,3.891667,3.0062501,2.1999998,1.6625001,1.1166668,0.65625,0.6333334,1.75,3.6125,5.641667,5.8312497,6.583334,7.4500003,0.9416667,1.8666668,2.7666667,2.15,1.5444444,1.15,0.88888896,3.008334,7.7444444,14.3111105,14.741667,12.922221,10.150001,4.2444444,0.89166665,0.24444446,0.17500001,0.84444445,2.666667,6.491667,12.844444,14.65,7.2222233,1.6999999,0.32222223,0.06666667,0.016666668,0.0,0.058333337,0.15555556,0.4666667,0.5888889,2.125,6.3555555,8.266666,12.541666,14.3555565,21.783335,19.388887,11.866667,9.433333,10.777778,16.666668,14.777777,9.758333,6.544444,2.7999997,0.47777778,0.13333334,0.016666668,0.97777784,3.8500001,2.9000003,0.97499996,0.9666667,1.0833335,0.5222222,0.06666667,0.0,0.0,0.016666668,0.0,0.0,0.0,0.0,0.0,0.0,0.041666668,4.6,7.1416674,0.8888889,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.0666667,2.5444443,1.3444445,0.058333334,0.011111111,0.0,0.31111112,2.0416665,0.8,0.0,0.0,0.0,0.5416666,1.3000001,0.8083334,0.2888889,0.083333336,0.2777778,1.2444445,0.4583333,0.3,0.083333336,0.011111111,0.0,0.0,0.0,0.0,0.0,0.0,0.044444446,0.7416667,0.25555557,0.18333334,0.13333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.044444446,0.12222223,0.9250001,1.0444444,0.8666667,0.14444445,0.0,0.0,0.0,0.091666676,0.11111113,0.17500001,0.08888889,0.083333336,0.22222224,1.2555556,3.2,1.8666667,1.5166667,0.77777785,0.025,0.0,0.0,0.033333335,0.11111112,0.15833333,0.14444445,0.8083333,1.7555556,3.0416667,5.777778,4.377778,3.9166667,8.444445,18.441668,22.311113,23.09167,24.488888,27.450003,27.477777,23.011112,15.233335,10.033335,5.5166664,2.8,4.675,8.411111,10.933334,9.875,14.322223,17.716667,20.58889,21.7,23.177776,23.822224,13.616668,10.366667,5.2583337,2.3,1.6583333,0.011111111,0.45833334,0.18888889,0.011111111,0.125,0.11111111,0.0,0.0,0.0,0.0,0.0,0.225,1.1666667,2.5499997,3.1555557,6.65,17.58889,28.316666,34.066666,28.699999,18.916668,24.277779,31.533335,19.677776,7.675,2.877778,2.188889,1.6666665,1.1555555,0.9583333,0.8111111,1.9833332,4.5333343,4.375,4.933334,4.8333335,3.916667,3.6777778,3.6416667,3.5333333,3.8500004,3.9,3.4444447,2.9666667,2.3,1.4333334,0.5222222,0.22500002,0.38888887,0.3888889,1.1916666,2.3666666,4.2250004,5.888889,8.058334,0.95000005,3.5666666,3.7416666,1.5312501,0.825,2.49375,7.408334,9.53125,14.0,17.433334,13.731251,6.491667,5.3187504,5.891667,4.94375,0.4583333,0.0,1.5833333,4.375,5.64375,11.108334,18.11875,10.608334,4.26875,1.7999998,0.41666663,0.28125,0.083333336,0.25,0.008333334,0.06875,0.6833334,2.3625002,3.8,10.575,15.618752,19.824999,25.81875,27.066664,20.775002,13.291667,7.8166666,12.73125,11.483334,8.987499,5.841667,2.24375,0.38333333,0.025,0.0,0.20000002,2.11875,3.3,1.8812499,3.1999998,5.606251,2.3083334,0.40833336,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0125,0.40000004,0.48125,0.31666666,0.0,0.0,0.0,0.0,0.0,0.0,0.025,0.1,0.09166667,0.016666668,0.05,0.016666668,0.0,0.075,1.5374999,3.375,1.45,0.25625,0.025,0.112500004,0.17500001,0.118750006,0.025,0.0375,0.23333332,0.36666664,0.18125,0.108333334,0.03125,0.008333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0125,0.2,0.48333335,0.6750001,0.42499998,0.31249997,0.0,0.0,0.0,0.17500001,0.3,0.05,0.56874996,0.32500002,0.21249999,1.5166667,1.5999999,2.04375,2.7166665,1.70625,0.3333333,0.2125,0.06666667,0.0,0.28333333,3.1083333,1.3625001,0.108333334,0.3125,0.5166667,3.94375,3.3,0.8083334,2.85,9.608334,16.55625,18.275,27.856253,15.691668,14.55,22.141666,26.458334,12.237499,6.1583333,6.3812504,7.3666663,4.2000003,5.791667,12.491667,14.112501,11.575,7.34375,6.1583333,6.175,7.291667,5.808333,3.0875,2.2083335,0.0625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0375,0.52500004,1.2125001,5.2166667,10.95,19.733334,29.81875,33.100002,31.866667,20.14375,12.2,15.556251,14.666667,9.2125,4.233333,1.9333333,0.4625,0.033333335,0.03125,0.5833333,0.7625,0.81666666,2.0062501,2.9250002,3.933333,4.4187493,4.5999994,4.55625,4.025,3.0375,2.9583335,2.7583332,2.4937499,2.2916667,2.84375,2.8583333,2.03125,1.6083333,0.7916666,0.68125004,2.1999998,4.7562504,5.6583333,7.0875,0.18333334,0.65555555,1.388889,3.8916667,4.8444443,7.1083336,12.166666,9.175,5.5,4.977778,5.7833333,5.1666665,5.9333334,7.966666,3.4666672,1.1444445,0.55,0.48888892,5.4444447,11.983334,11.622223,10.075,5.577778,6.775,1.5777779,0.055555556,0.0,0.44444445,0.8416667,0.4222222,1.0,3.2333336,5.475,10.766666,17.222223,20.066666,23.844444,24.625,22.588888,16.408335,11.733334,6.122223,9.258332,8.055555,6.033333,3.266667,1.1833334,0.12222222,0.0,0.0,0.08888889,1.25,2.7222223,6.275,8.933334,14.333334,14.066667,2.4444444,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.15833335,1.1555555,1.0416666,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.18333334,0.0,0.0,0.0,0.0,0.0,0.033333335,0.058333334,1.7444445,4.0555553,15.425,3.8666668,0.14166667,1.2333333,2.075,1.2666667,0.050000004,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05,0.0,0.033333335,0.016666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016666668,0.044444446,0.0,0.0,0.075,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016666668,0.0,0.041666668,0.16666669,0.41111112,0.20000002,0.07777778,0.083333336,0.0,0.0,0.0,0.42222223,0.7916667,0.9111111,0.75000006,0.37777779,0.20833334,1.9555556,2.7,2.45,3.522222,3.0916667,2.4222224,1.4416668,1.0555556,0.058333334,0.011111111,3.7555556,4.241667,0.0,2.1333332,7.7222223,7.725001,5.377778,4.388889,6.3666663,5.0222225,3.8750002,7.5111113,9.583335,7.1111116,6.383333,16.5,25.011112,26.108335,21.811111,14.808333,12.133333,6.2250004,4.5222225,7.0888886,8.983334,6.1888885,5.15,3.8000002,4.091667,3.8111112,3.2333333,1.9166667,0.73333335,0.083333336,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.26666668,1.7777778,4.9083333,5.0222225,3.0888886,1.3333334,0.82222223,1.45,3.5333338,4.375,2.777778,1.488889,0.46666664,0.07777778,0.0,0.11111111,0.85,1.5444446,1.7666667,3.3222222,4.0444446,5.3333335,5.188889,5.091667,5.1666665,4.0666666,2.8222222,2.2555559,2.45,3.9888892,4.6666675,4.4777784,3.6166666,3.0111113,2.1333334,1.7833333,1.9000001,2.666667,4.2333336,5.6333337,0.118750006,1.0666666,4.125,6.118749,4.708333,4.36875,3.641667,2.75,3.2916663,5.475,7.35625,5.8000007,3.3999999,3.525,2.3812504,3.7000003,1.5187502,3.1916668,8.416668,17.324999,13.208333,6.5000005,3.6249998,5.2124996,2.1333332,0.016666668,0.0,0.0,1.00625,2.5583334,3.30625,5.8250003,9.25,14.733335,19.025,21.525,22.158335,21.212502,16.008335,9.837501,8.416667,4.466666,6.25,5.783333,3.7687497,2.1999998,1.0375,0.016666668,0.0,0.01875,0.28333333,1.04375,2.7500002,5.9187503,14.641666,13.637501,3.6750002,0.33333334,0.0,0.016666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.25625,3.8249998,3.9250004,0.25,0.3125,0.0,0.0,0.0,0.21666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00625,0.20000002,1.175,6.1312504,8.725,0.88750005,3.3916664,13.700001,8.075,0.37500003,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.16250001,0.083333336,0.23333333,0.0625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0375,0.13333336,0.0,0.0,0.24374999,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.20625001,0.15000002,0.03125,0.1,0.17500003,0.075,0.0,0.0625,0.0,0.0,0.0,0.5166667,0.8937501,0.6916667,0.9375,0.43333337,0.6500001,1.475,1.9750001,0.9250001,1.9000002,2.7937498,2.7916665,1.2437501,3.625,0.28125,0.0,0.0,0.4125,0.0,1.375,4.8083334,2.6812499,4.616667,2.4750001,3.85,5.133333,6.13125,9.483334,9.606249,8.074999,10.012501,20.525002,25.091667,18.893751,17.675001,19.83125,20.833336,18.462502,12.400001,7.525,2.2312498,1.5166667,2.88125,1.275,0.56875,0.23333335,0.2,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025,0.14375,0.041666668,0.0,0.0,0.0,0.01875,0.050000004,0.14375,0.10000001,0.050000004,0.025,0.0,0.0,0.0,0.0,0.52500004,3.5437503,7.175,7.2666674,6.45,5.133333,4.5375,4.9333334,4.69375,3.2166667,1.8749998,2.95,4.375,4.4374995,4.2,3.4437497,3.2583334,3.241667,3.0375001,2.0833333,1.25625,1.5833335,2.1625,1.8416666,4.588889,4.266667,0.36666667,0.24444444,0.33333334,0.6333333,2.6416664,5.4222226,16.255556,20.466665,7.566666,1.7833334,1.0888889,1.9333334,1.7666667,0.8666667,3.8222222,9.677777,16.341667,9.788889,5.025,1.3444444,0.6916666,1.2555556,0.93333334,0.10833334,0.0,1.0083333,2.6111112,4.65,7.588889,12.45,15.888889,16.755556,17.533333,16.355556,12.991666,7.088889,5.6916666,5.6222224,2.3333335,3.2583337,3.3666668,1.8000002,2.1222224,1.4333334,0.0,0.011111111,0.59166664,1.0111111,1.2166667,1.8333333,4.3583336,10.177778,10.908334,4.411111,0.42222223,0.033333335,0.08888889,0.0,0.0,0.06666667,0.17777778,0.0,0.033333335,0.5888889,1.1416668,5.3888884,3.6583335,0.033333335,0.525,0.033333335,0.1,1.45,2.6222224,0.0,0.0,0.0,0.08888889,0.41111112,0.0,0.0,0.1,3.4444447,1.4083333,0.5333333,0.16666667,0.4083333,2.0777779,1.9583333,1.4555554,0.425,0.61111116,0.22500001,0.022222223,0.0,0.0,0.0,0.48333335,0.988889,0.016666668,0.033333335,1.8333335,1.5250001,0.64444447,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.033333335,0.0,0.0,0.0,0.0,0.0,0.15833335,0.18888889,0.0,0.0,0.27499998,0.12222222,0.23333335,0.4777778,0.39999998,0.041666668,0.16666667,0.0,0.0,0.0,0.0,0.0,0.0,0.011111111,0.016666668,0.06666667,0.2916667,0.1777778,0.06666667,0.22222224,0.36666667,0.15833333,0.14444444,0.16666666,0.0,0.0,0.0,0.5,0.18333334,0.13333334,0.5,0.2,0.5083333,0.44444448,0.26666668,0.175,2.4444447,1.6333334,1.0,1.0083333,1.2777778,1.1750001,0.6888889,0.0,0.0,0.23333333,3.4583335,7.922222,1.5416665,1.0333334,1.8111112,1.0833333,2.0444446,8.891666,15.211109,16.183334,14.555555,13.799999,11.455556,25.4,24.099998,23.555557,25.083332,19.188889,22.391666,20.455557,14.233334,1.2333333,0.08888889,0.98333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.25833333,0.65555555,0.40000004,2.4,9.355556,11.558333,7.3333335,4.275,6.0333333,8.4,5.755556,4.0,5.0916677,4.9444447,3.9916668,3.8,3.725,4.211111,4.7333336,4.4,3.0222225,1.7166666,0.8,0.7333334,0.49166667,2.1777778,4.233333,1.5166667,0.022222223,0.42499998,1.5333334,1.2,2.7777777,13.533334,14.916666,7.066667,5.0583334,2.1666665,0.90000004,2.3,3.5750003,1.9777777,5.3888893,9.858334,6.088889,3.325,0.0,0.0,1.3888888,2.8222222,1.0666667,0.06666667,0.65000004,2.811111,6.5583334,8.777779,11.666668,13.1,15.922222,12.558332,11.08889,6.1833334,4.3444443,4.5499997,3.4666667,1.1222222,1.6249999,1.9444444,1.1166667,1.6666667,1.1999999,0.05555556,0.15555556,1.2166667,1.488889,1.9083334,2.0333335,5.425,13.455556,12.916666,6.333333,0.47777778,0.1,0.11111111,0.0,0.0,4.383333,4.133333,0.0,0.26666668,1.0444446,1.175,3.2555552,1.2166667,0.0,0.041666668,0.0,1.2555556,1.7583334,0.3,0.0,0.0,0.0,2.1,1.5000001,0.0,0.0,0.0,1.1555556,3.516667,3.3666668,0.57777786,0.15833333,0.022222223,0.37499997,0.4222222,0.058333337,0.16666667,0.5083333,0.33333334,0.044444446,0.0,0.0,0.0,0.08888889,0.16666667,0.0,0.0,0.0,0.0,0.0,0.12222222,0.725,0.68888897,0.11666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.3222222,0.016666668,0.06666667,0.016666668,0.0,0.0,0.48333338,0.1,0.0,0.0,0.24166666,0.033333335,0.116666675,0.54444444,0.37777773,0.15833335,0.47777775,0.008333334,0.0,0.0,0.0,0.0,0.0,0.10000001,0.16666667,0.46666664,0.4416667,0.37777779,0.058333337,0.14444445,0.6333333,0.3,0.47777778,0.175,0.0,0.0,0.0,0.0,0.016666668,0.044444446,0.34166667,0.54444444,1.1583334,0.41111112,0.0,0.4166667,1.1111112,1.6916666,1.7444444,1.7250001,1.4888891,2.2083335,4.3444448,0.6333333,1.2666668,0.3,4.8333335,11.011111,5.058334,0.0,2.111111,1.2666667,4.1444445,15.433334,25.055557,21.625,11.388889,5.416667,1.9000001,7.1333337,7.8499994,11.833334,14.741667,6.044445,7.325,15.322224,12.922223,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.15555555,0.48333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.57777774,1.125,1.2666667,1.7,4.633333,8.477778,6.191667,11.077778,15.308332,11.933332,8.822223,6.75,5.4111114,4.6416664,4.677778,5.1416664,6.3888893,7.5999994,7.25,6.1555557,4.7750006,2.977778,2.2083333,0.50625,1.7083333,3.1833336,1.40625,0.275,0.4875,0.5416667,0.63124996,2.4583335,6.975,7.7437506,6.6916666,12.0875,7.866667,6.2437506,6.0916667,2.075,0.5916667,1.7416668,7.5999994,6.708334,0.76874995,0.125,0.75625,0.19166668,4.633333,2.2625,0.6,0.85,2.4333334,5.90625,7.0,8.78125,10.416666,10.583334,7.09375,4.0250006,2.1000001,3.266667,5.23125,2.6583333,1.8000001,1.7312502,2.1833334,1.28125,1.6916666,1.0687499,0.43333334,0.675,2.59375,3.9416668,3.025,3.016667,6.31875,16.508333,13.668751,9.791667,1.9583335,0.15000002,0.016666668,0.0,0.0,4.025,2.9416666,0.1,2.5125,3.8416665,1.1187501,0.35000002,0.275,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.116666675,0.9125,1.9333334,0.24166667,0.0,0.0,0.0,0.0,1.26875,5.3583336,2.6375,0.26666668,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.5083333,5.075,4.741667,1.1312499,0.0,0.0,0.0,0.0,0.0,0.0,0.0375,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1875,0.6333333,0.1,0.45833334,0.125,0.033333335,0.13333334,0.6999999,0.016666668,0.0,0.0,0.0625,0.11666666,0.0375,0.21666668,0.35833332,0.51250005,1.05,0.04375,0.0,0.0,0.0,0.0,0.05625,0.11666667,0.18750001,0.52500004,0.74375,0.35,0.087500006,0.21666668,0.6,0.19375,0.06666667,0.0,0.0,0.0,0.0,0.0,0.0,0.16666669,0.81875,0.82500005,0.9875,1.1416667,0.7166667,0.45000002,0.93333334,2.7937503,3.8166668,3.0375001,1.1166666,2.825,10.625001,3.6333337,0.4625,2.35,2.05,5.191667,2.60625,0.016666668,0.116666675,0.24375002,5.0000005,14.387502,27.283333,26.06875,10.025001,4.44375,0.7583333,0.38333336,0.3375,0.29999998,2.1875,0.36666667,0.48125,0.9583334,0.5833333,0.03125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.35,0.9625,0.09166667,0.0,0.0,0.0,0.0,0.0,0.0,0.13333334,0.55,0.8916667,1.13125,1.8,2.55,3.3124998,3.6916664,4.84375,10.466667,18.73125,15.391666,10.091666,6.4750004,5.75,6.2749996,6.5083337,7.4062495,8.6,7.841667,6.15,5.533334,5.5750003,4.5416665,4.2937503,1.0333334,1.3777778,2.5333335,0.48333335,0.0,0.25,1.2333335,3.0000002,3.0000002,8.9777775,9.858334,9.122222,8.408334,4.766667,4.091667,3.4555557,0.0,2.0444443,0.7222222,1.5583334,2.1666665,0.6833334,0.13333334,1.8583333,2.0444446,0.055555556,1.3499999,1.0222223,1.0000001,2.5,4.1666665,5.111111,5.733333,6.5777783,5.866667,3.0166667,1.9888887,2.4166667,2.5333333,4.3999996,6.244445,3.1666667,2.925,2.8444445,1.8666668,2.1222222,1.4833332,1.0222222,1.5666667,4.158334,6.1777782,4.9,3.8111112,5.9416666,16.966667,16.25,10.444445,1.7,0.35833335,0.0,0.0,0.0,0.041666668,0.11111111,0.7444445,1.8333334,0.6111111,0.29166666,0.54444444,1.1999999,0.8222222,0.09166667,0.0,0.0,0.0,0.0,0.05,0.0,0.375,0.26666668,0.0,0.0,0.0,0.0,0.0,0.033333335,0.08888889,2.166667,0.74166673,0.0,0.0,3.222222,12.525001,21.855556,12.566666,1.5,0.1,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.3583333,1.9666667,0.30833334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.44166666,0.0,0.16666667,0.18888889,0.16666667,0.0,0.0,0.45000002,0.0,0.025,0.0,0.0,0.0,0.0,0.0,0.41111112,0.38333338,1.6444445,0.325,0.0,0.0,0.0,0.0,0.033333335,0.25555557,0.19166669,0.23333336,0.7,0.48888892,0.058333337,0.16666667,0.07777778,0.041666668,0.33333334,0.25,0.055555556,0.0,0.0,0.022222223,0.025,0.41111112,1.65,1.0777777,0.9666667,2.9,3.6555557,1.0500001,3.2777781,6.5916667,6.755555,3.6583335,1.8777776,0.4583333,2.8333335,1.2555555,2.8333335,6.0222225,3.325,0.14444444,0.0,0.0,0.055555556,0.2,6.0666666,5.0916667,7.1777773,9.141666,6.8111115,3.025,0.85555553,0.21111111,0.0,0.033333335,0.40000004,1.0333334,1.425,0.64444447,0.5222222,0.24166667,0.3888889,0.50000006,0.62222224,0.6000001,0.35555556,0.18888889,0.016666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011111111,0.60833335,0.45555556,0.22500002,0.055555556,0.0,0.0,0.0,0.008333334,0.34444442,1.0666668,1.0555556,1.625,1.7444444,1.9666667,2.8333335,2.9555554,2.5499997,2.3888886,7.841666,15.444444,12.633334,9.458333,8.755556,9.3,9.533334,10.033334,9.111111,7.8111115,6.758333,6.8999996,6.6916666,5.0333333,5.675,5.4249997,3.7333336,1.875,0.03125,0.083333336,0.075,0.23333335,2.55625,6.025,7.308334,9.531249,7.158334,5.89375,1.3499999,0.73125005,0.95833343,0.12499999,0.825,6.0750003,10.2125,2.8666666,3.0625,0.31666666,3.4125004,8.183333,2.675,4.175,0.68333334,2.825,6.1833334,3.94375,4.475,3.84375,3.108333,3.3416667,3.0687501,2.9666667,4.9812503,3.9500003,3.775,5.0,6.5,5.4937496,4.0083337,2.3937495,2.125,1.7875,2.0,2.4416666,6.6374993,5.2833333,5.05,4.75,6.875,14.733334,15.98125,9.791667,1.5916667,0.38749996,0.14166668,0.1375,0.22500001,0.4875,0.36666667,1.5583334,3.15,0.425,0.06875,2.391667,3.5749998,1.5083334,0.63125,0.0,0.025,0.0,0.15,0.9375001,1.1416667,4.3062496,3.083333,0.125,2.8125,6.9333334,0.0625,0.0,0.0,0.0,0.0,0.0,0.0,0.0875,2.7083335,6.36875,3.0666668,1.3687501,0.25,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1,4.40625,2.3583333,0.13125001,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.18125002,0.0,0.1375,0.16666666,0.125,0.0,0.0,0.025,0.0,0.34375,0.25,0.0,0.0,0.0,0.025,0.96666676,0.9125,0.79999995,0.59375006,0.0,0.0,0.0,0.0,0.0125,0.108333334,0.16250001,0.36666667,0.64374995,0.3,0.0,0.008333334,0.008333334,0.47500002,0.89166665,0.71874994,0.041666668,0.0,0.0,0.13333334,0.16250001,0.70000005,1.5375,1.2583334,2.64375,4.2000003,1.5,0.44375002,3.6166666,4.1250005,5.283333,1.075,1.0583334,1.35,1.5583334,0.9833334,1.38125,4.5666666,8.512501,7.1666665,8.225,5.9666667,2.7416668,1.8187499,1.1583334,10.125,9.9,15.087501,24.75,17.487501,7.533334,3.3666668,2.68125,2.0,4.70625,5.3166666,3.04375,1.3583333,1.825,2.00625,3.0166667,3.4000003,2.6166663,1.8625,0.7333334,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.175,0.8625001,1.375,1.05625,0.6583333,0.35833335,0.18125,0.05,0.13750002,0.20000002,0.29999998,0.5416666,0.75625,1.1333334,1.825,2.5625,3.266667,3.40625,2.6750002,4.10625,7.3916664,10.008333,13.18125,13.441667,10.975,9.558333,8.575001,7.408334,7.175,6.95,7.1,6.3375,6.541667,6.6812506,11.558334,8.5,3.8777776,1.25,1.1777779,0.13333334,0.044444446,0.98333335,4.0666666,7.7222223,8.7,8.422222,5.9416666,1.3777778,0.05,0.3,1.1500001,6.033334,14.233334,13.041666,5.9444447,5.116667,1.4777777,4.4583335,13.200001,12.111111,6.825,1.3444445,5.333333,7.1444445,7.541667,5.2999997,4.8166666,3.9333336,4.588889,5.05,7.688889,9.433333,6.422222,6.583334,7.866667,9.444445,8.891666,6.1111107,3.3500001,2.4444447,2.0916667,3.2111113,3.7222226,8.325001,7.877777,5.4583335,4.577778,6.116667,10.655557,11.508334,7.1222215,1.7333333,0.5916667,1.2666668,0.29166666,1.388889,3.1000001,1.4125,1.977778,1.0916667,0.23333335,0.39166668,2.7555554,2.8833334,0.44444448,0.016666668,0.0,2.1666667,1.3416667,3.6,2.9583335,0.46666667,1.5500001,0.6,0.0,0.15833335,3.9555557,0.041666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.008333334,0.08888889,0.5083333,0.16666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.35,1.0666667,0.050000004,0.0,0.0,0.0,0.0,1.0,0.54444444,0.0,0.0,0.0,0.14444444,1.7666667,1.5000002,0.5666667,0.17500001,0.12222223,0.09166667,0.0,0.0,0.0,0.0,0.008333334,0.1,0.016666668,0.0,0.0,0.0,0.033333335,0.59166676,0.8,0.36666667,0.0,0.0,0.0,0.0,0.3,0.95555556,0.55833334,1.0555556,1.7833334,1.7555555,2.1555555,0.9083334,1.1666667,1.8000001,1.5111113,1.1333333,4.1666665,4.25,5.9888887,8.466667,5.983333,2.511111,15.558332,7.955556,7.491667,5.5000005,11.222222,10.891667,10.311111,17.758335,21.122223,19.291666,18.655556,15.066668,10.211111,6.555556,6.325001,15.555556,30.116669,27.7,13.233334,3.8444448,1.0777777,0.22500002,0.3,0.20833336,0.17777778,0.05,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.26666668,0.0,0.0,0.016666668,0.13333334,0.77500004,2.1777778,2.6,2.4111114,1.2444445,0.26666668,0.1,0.24999999,0.2777778,0.108333334,0.25555557,0.70000005,1.7222223,2.5666668,3.3583336,3.588889,3.6083336,3.8000002,3.9916668,4.311111,5.2555556,11.275,13.633333,10.725,8.48889,7.6916666,6.866667,6.7999997,6.4083333,5.4999995,5.766667,6.811111,6.933334,12.106249,8.624999,1.8750001,0.9312501,0.5,0.01875,0.47500002,1.5000002,1.9166666,5.1916666,11.593751,11.091667,6.2749996,3.2166665,0.5375,0.38333336,0.85,3.8916667,7.091667,6.10625,6.866667,5.7062497,4.4000006,5.95625,19.916668,11.466666,8.000001,3.716667,5.9,6.450001,8.03125,9.85,10.90625,10.424999,13.766666,15.725,13.424999,23.224998,13.533334,10.137501,11.383333,14.216667,12.43125,8.775001,5.6749997,3.6833334,2.2375002,3.858333,4.508334,7.3312497,8.650001,11.3875,4.766667,2.8187501,4.666667,5.8375006,1.766667,0.6833333,1.1625001,1.4833332,0.81875,2.6416664,3.7312498,2.0533333,1.2,0.9875001,0.68333334,1.03125,3.2583332,3.0708332,0.033333335,0.67875004,3.0166664,3.8416667,2.3875,5.575,4.9312496,2.225,0.48416665,0.36666667,0.0,0.0,0.0,0.14375001,0.85833335,0.025,0.0,0.0,0.0,0.225,1.23125,1.5333333,0.17500001,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00625,0.10000001,0.30624998,0.1,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1,0.025,0.0,0.0,0.0,0.0,0.16250001,0.35000002,0.00625,0.0,0.0,0.0,0.09166667,1.4625001,0.5583333,0.075,0.083333336,0.01875,0.10833333,1.9916668,2.25,2.1750002,0.14375,0.175,0.13125,0.0,0.1,0.056250002,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06666667,0.34374994,0.425,0.043750003,0.0,0.0,0.0,0.041666668,0.25625002,0.6499999,0.8374999,1.3333333,1.1374999,0.575,2.275,2.25625,2.25,2.25,1.8083334,2.00625,3.116667,2.91875,2.9166665,1.1916668,1.0125,1.5083333,6.4875,5.1749997,2.10625,1.4833333,1.4916667,5.5249996,8.583333,8.74375,7.591666,7.0249996,5.833333,4.025,2.4083333,2.0583334,4.43125,10.816668,17.768751,16.691668,8.65,2.8666668,0.6916666,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0125,0.06666667,0.0,0.0,0.0,0.00625,0.15833335,0.53749996,1.5250001,2.8125,2.6916668,1.65,0.6875,0.31666666,0.11250001,0.041666668,0.26875,0.9833334,1.5937502,2.65,3.6166668,4.2749996,4.55,5.14375,4.7916665,5.4000006,5.491667,5.35,7.4875,9.233334,12.225,11.066667,8.2375,6.541667,6.325,6.1124997,6.2249994,7.26875,7.5,7.475,7.1499996,3.4222221,1.6444443,0.53333336,1.1222222,1.5333333,1.7666667,2.2583337,3.7555554,3.9555554,7.108334,10.2,14.450001,10.922222,1.1833333,1.0333333,0.5833333,0.6666667,1.1,1.9250001,2.8222222,2.8,7.866667,16.158333,21.199999,10.488889,6.525,10.300001,10.916666,13.877778,18.216667,15.544445,20.166666,17.377777,20.211111,20.475,15.588889,25.516668,19.744446,14.299999,18.622223,20.98889,14.483332,7.8444448,5.408334,3.8555555,2.141667,1.9000001,4.0555553,4.375,6.1666665,11.758334,3.0777776,1.1999999,0.8444445,0.7749999,0.6444444,0.6111111,0.70000005,2.1888888,3.7583332,5.166667,4.041667,3.2666667,1.4555557,0.95,1.4444445,4.4416666,4.6222224,1.1166667,0.2,2.2250001,6.3416667,1.3767858,1.9083333,4.2000003,2.6916666,2.266667,1.2189394,0.48888892,0.0,0.0,0.0,4.05,7.7777777,0.4416667,0.0,0.0,0.0,5.1555557,5.1250005,5.9444447,3.2749999,0.57777774,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06666667,0.57500005,0.7888889,0.25,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.6333333,0.225,0.0,0.0,0.0,0.0,0.025,0.0,0.0,0.06666667,0.2,0.16666667,0.0,0.875,0.9111111,0.050000004,0.11111112,0.2,0.06666667,1.4111111,1.7083334,1.3333334,0.116666675,0.0,0.0,0.0,0.32222223,0.45,0.0,0.0,0.0,0.025,0.011111111,0.0,0.0,0.033333335,0.14166668,0.15555558,0.0,0.0,0.0,0.0,0.07777778,0.09166667,0.43333334,0.775,0.54444444,0.4,0.06666667,0.72222227,2.358333,1.5777777,2.2083333,1.5,2.1166668,2.5,2.1500003,2.2555556,0.6,0.275,0.0,0.125,1.2777779,5.0250006,9.6,6.111111,0.74166673,2.9444447,3.1083333,1.2444446,1.3083333,4.4333334,5.4083333,7.288889,7.7000003,7.0,5.4,2.8249998,1.511111,3.3833332,2.8333335,0.06666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.18888889,1.075,1.1000001,0.125,0.011111111,0.2777778,0.041666668,0.0,0.175,1.0222223,2.95,3.4,1.8555557,2.1333332,0.8666667,0.3,0.5888889,1.2249999,2.611111,3.3833332,4.333333,5.111111,5.2833333,5.3111115,5.458333,6.255556,5.983334,5.1555557,4.977778,6.541667,9.144444,9.758333,9.344445,8.016667,9.833333,10.122222,8.816668,7.8,6.641667,6.188889,4.95,7.95,6.6333337,4.288889,1.2166667,2.411111,2.3000002,2.4222224,2.35,2.3333333,3.6777778,8.691667,11.266668,9.425,8.822222,8.591666,11.5222225,10.266667,6.255556,2.788889,0.7166667,0.3777778,2.2583332,3.3666666,4.383333,3.177778,5.2666664,9.291667,16.588888,24.65,32.31111,32.025,15.122223,16.383331,15.68889,16.177778,23.025002,15.088889,17.85,18.322224,18.391666,19.91111,18.122223,11.641667,6.133333,4.7416663,1.8222222,0.25833336,0.18888888,1.811111,2.6416667,6.3,10.016666,1.9444444,1.0749999,0.68888885,0.45,0.54444444,2.0555556,4.3083334,7.5666666,7.7,6.8555555,4.1083336,2.9555554,1.8000001,2.6333332,4.8555555,5.0666666,3.1888888,1.4416667,0.2777778,2.8530302,11.915874,6.0666666,5.6583333,5.0,2.6340907,1.0027779,1.9916667,0.76666665,0.0,0.0,0.0,0.33333334,0.5222222,0.0,0.0,0.0,0.31666666,7.388889,4.3083334,17.78889,14.916666,2.0111113,0.10000001,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016666668,0.11111111,0.083333336,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.64166665,0.25555557,0.0,0.0,0.0,0.0,0.0,0.0,0.21111111,0.0,0.0,0.0,0.6666667,0.26666668,0.0,0.0,0.0,0.42222223,0.075,0.044444446,0.0,0.24444446,0.53333336,0.9499999,0.21111111,0.06666667,0.57777786,0.33333334,0.18888889,0.69166666,0.08888889,0.4888889,0.90000004,0.40000004,0.20833333,0.033333335,0.0,0.42222223,0.16666666,0.4666667,0.08888889,0.0,0.0,0.016666668,0.2777778,0.0,0.022222223,0.0,0.008333334,0.022222223,0.0,0.0,0.0,0.0,0.0,0.0,0.08888889,0.25000003,0.0,0.041666668,0.055555556,0.08888889,3.8333335,4.7222223,2.5166667,1.1666667,2.6833334,3.3333335,4.0583334,6.333334,4.7,1.825,0.53333336,0.3,1.0666667,5.741667,10.200001,5.9222226,1.95,1.0000001,1.1,0.0,0.016666668,1.8555555,3.5916667,2.5777779,1.9555557,1.3666667,0.0,0.0,0.0,0.08333334,0.11111112,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011111111,0.058333337,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011111111,0.24166667,0.6222223,1.6833334,1.8888888,1.2416666,0.2777778,1.0555556,0.4916667,0.13333334,0.325,1.8333334,1.0833334,1.3777777,1.5444444,2.1166668,0.6666667,0.4416667,1.7444444,2.6833334,3.9333334,4.7499995,5.388889,6.3555555,6.5249996,6.6222224,5.4833336,5.3555555,6.1,5.200001,5.4,7.175,7.611111,8.166667,6.577778,7.7333336,10.788889,9.466667,6.208334,5.455556,4.6083336,2.4222224,1.3166667,2.4125001,0.6,0.50000006,0.79375005,1.0166668,0.53749996,0.30833334,0.5,0.44166666,1.8083335,3.725,6.741667,10.431251,10.241668,11.9375,13.108335,10.1125,4.5333333,2.0500002,1.43125,1.2666667,1.1875001,2.0833335,3.85625,5.4500003,8.041667,6.575001,7.258333,18.5625,31.21667,28.868752,14.141666,14.475001,12.358334,14.091666,23.5,16.925001,19.550001,24.091667,23.462502,14.591667,10.841667,7.36875,5.6333337,5.1312504,1.1416667,0.33124998,0.19999997,0.59166664,0.45,3.1166668,4.08125,0.66666675,0.6,0.34166667,2.0625,4.358333,5.4249997,7.4937496,8.25,7.2375,6.533333,4.9937506,5.083333,5.7999997,6.4375,6.6916666,5.2375,2.4916666,0.53125006,1.0833333,3.2937503,7.066667,6.958334,5.1983337,2.625,1.4937501,0.90833336,0.43124998,0.083333336,0.15833335,0.0,0.0,0.29999998,0.0,0.0,0.0,0.0,0.0,0.57500005,1.6187501,4.791667,2.00625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0125,0.13333334,0.13125,0.041666668,0.0,0.0,0.0,0.0,0.0,0.29999998,0.90833336,0.03125,0.0,0.0,0.0,0.0,4.3562503,9.941667,0.7125,0.0,0.0,0.0,0.0,0.0,0.14166667,0.0,0.0,0.0,0.108333334,0.06875,0.0,0.0,0.0,0.09166667,0.10000001,0.0,0.0,0.15833335,0.40000004,0.4625,0.40833336,0.18124999,0.2833333,0.13125,0.13333333,0.53125006,0.4166667,0.3166667,0.41875005,0.26666668,0.44375002,0.41666666,0.45625,0.16666667,0.25,0.0,0.0,0.025,0.35833335,0.087500006,0.64166665,0.325,0.15,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.125,0.23333333,0.7062501,2.1333334,1.0500001,1.9666666,1.73125,3.8000002,2.4625,2.825,2.3166668,2.9250002,3.4750001,3.13125,3.3166666,4.53125,6.3916664,3.6916666,3.26875,3.2,0.68125004,1.6500001,1.325,0.0,0.39375,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.008333334,0.125,0.3,0.28125003,0.09166667,0.00625,0.0,0.0,0.325,0.26666668,0.28750002,0.49166662,1.6062499,2.4416666,3.3625002,2.6166668,2.1833332,2.4437501,1.1333333,1.0125,1.5,0.74375004,0.55833334,0.975,1.7625,1.325,1.2,2.1833334,3.7124999,4.5083337,4.775,5.475,5.858333,6.1937504,6.05,5.6687503,6.9000006,5.825,4.7583337,4.925,5.6750007,5.4,5.1625,4.775,4.0125,3.691667,3.833333,3.50625,2.525,1.5687499,0.45000005,0.32500005,5.766667,3.8333335,3.3,1.8916667,0.47777778,0.45000002,0.34444445,0.18333332,0.11111111,1.9777778,2.525,4.7000003,8.766666,3.7777777,1.5333333,0.5222222,1.3833332,2.9666667,5.777778,4.65,2.5666666,1.3583332,1.5444443,1.3833334,2.5444446,3.711111,3.375,5.977778,12.008333,18.300001,20.591667,15.955556,14.733334,15.5,20.355556,22.574999,19.788889,21.208332,16.055557,11.700001,7.8555555,6.5,4.291667,3.5444443,2.175,0.21111111,0.025,0.0,0.0,0.36666667,1.0222223,0.7,0.18888889,0.6583333,1.8333333,3.125,3.977778,5.4888887,5.625,5.6888885,6.4,6.7222223,7.55,7.5111113,7.233333,6.991667,4.6111107,1.9166665,0.42222223,0.13333334,0.35555556,2.5416667,5.333333,5.788889,2.8583336,2.177778,0.87500006,0.06666667,0.050000004,0.24444446,0.6666667,0.26666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.050000004,0.61111104,0.041666668,0.0,0.0,0.0,0.0,0.7583333,5.977778,1.8,0.0,0.0,0.0,0.0,0.0,0.0,0.21666667,1.8333334,1.9916666,0.21111113,0.36666667,0.31111112,0.0,0.0,0.0,0.016666668,0.0,0.0,0.0,0.14444445,0.1,0.12222222,0.0,0.0,0.51666665,0.5333333,0.9083333,0.43333334,0.7555555,0.55833334,0.50000006,0.13333334,0.15555556,0.83333325,0.7555555,0.055555556,0.016666668,0.0,0.108333334,0.71111107,0.30833334,0.3888889,0.8666667,0.1,0.13333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05,1.2888889,1.1583333,0.6,1.1833334,0.25555557,0.6666666,1.9111111,1.9888889,1.475,2.7666667,4.075,2.9555554,2.4083333,2.3222222,2.388889,2.225,2.3555555,0.68333334,0.37777779,1.0,0.2777778,0.8666667,0.055555556,0.38888887,0.13333333,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.044444446,0.10833335,0.15555556,0.125,0.31111112,0.25833336,0.77777785,0.76666665,0.675,0.82222223,0.875,0.8666667,0.25000003,0.06666667,0.13333334,0.15833336,0.27777782,0.28333336,0.22222224,0.8833333,2.8333335,4.4583335,4.6444445,3.5111113,4.5583334,4.322222,4.2333336,2.1555557,2.2666664,2.088889,2.3222222,3.191667,3.6000001,3.0749998,3.1555552,4.7083335,5.3333335,4.825,5.422222,5.766667,5.633333,6.3666663,5.3166666,6.411111,5.875,4.477778,3.7555554,4.2,3.9555554,4.741667,4.644445,3.1000001,2.1777778,1.5,1.5416666,1.0555556,0.26666668,0.022222223,0.13333334,2.0187502,1.5583334,2.2333336,3.1374998,2.1499999,1.8625002,1.491667,0.625,0.36666667,0.775,2.48125,4.4249997,4.225,1.875,2.8125002,3.65,4.20625,3.7499998,3.016667,2.8687499,2.8333335,2.60625,4.008333,8.837501,11.874999,9.2,5.2187495,4.9833336,9.268749,13.358334,22.75,20.125002,12.518751,11.683334,13.075001,17.393751,11.733334,10.01875,7.916667,5.3125,3.5416665,2.9166665,1.41875,0.8000001,0.3,0.016666668,0.0,0.0,0.125,0.21875,0.26666665,0.125,0.325,0.64375,2.25,3.925,4.683334,5.0166674,5.09375,6.375,6.4125,7.433333,7.3250003,5.45,4.75,3.6375,1.6916667,1.1634614,0.41904762,1.1962501,1.2333333,3.3625,3.8400002,1.8416668,0.5396978,1.0145454,0.40625003,0.0,0.0,1.05,1.6500001,1.35,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.13125,4.241667,2.5500002,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.625,0.86875004,0.5083333,0.49375004,0.65,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00625,0.0,1.175,0.0,0.03125,0.31666666,0.19375001,0.59999996,0.5833333,0.8875,0.28333336,0.25,0.0,0.40000004,0.5666667,0.2,0.01875,0.033333335,0.0,0.3,0.14375001,0.06666667,1.10625,0.19166666,0.041666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0125,0.30833334,0.73125005,1.3166667,0.55625,0.091666676,0.31249997,2.1416667,2.4833333,0.7687501,0.275,2.31875,3.2499998,4.16875,2.1333332,1.9083333,3.43125,4.85,4.05,4.5333333,4.525,2.0666666,2.075,0.875,1.575,0.2625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.058333337,0.5875,2.3416667,3.0312502,4.458333,5.3125,5.8250003,6.9750004,6.5874996,5.1750007,4.6375003,3.3083334,2.05,1.2083333,0.50000006,0.5125,0.31666666,0.28124997,0.72499996,1.7874999,2.6083336,5.2625,5.708334,5.1333337,5.45,6.6916666,7.2375,6.9000006,6.2875,5.5666676,4.7250004,4.818751,5.408334,5.075001,5.1749997,4.9375,5.1,4.6375003,5.208334,5.2583337,6.0499997,6.266667,6.8124995,8.208333,7.0875006,4.6749997,3.45,3.30625,3.3500001,3.5374997,3.9333334,3.6937501,3.483333,3.0083337,2.50625,0.78333336,0.00625,0.0,0.025,3.2,1.9222223,2.1666667,0.5083334,0.23333333,0.45833334,0.47777775,0.3916667,0.6333333,0.72222227,2.1,2.4555554,1.5333333,2.0444446,4.383333,5.177778,8.525,11.588889,11.633334,9.458335,4.2333336,4.6833334,8.9777775,8.55,6.9,5.2555556,2.5916667,1.6555555,1.1916666,1.8888888,10.308334,8.966667,6.208333,3.0333333,3.2444446,2.525,1.9555554,1.9333335,2.3444443,2.2,0.75555557,0.16666667,0.18333332,0.84444445,0.25833333,0.0,0.0,0.0,0.16666667,0.20833334,0.21111111,0.18333334,0.8888889,1.6999999,2.3888888,4.3,5.833334,7.0444446,6.991666,6.633333,6.0916667,5.422222,4.0166664,3.5333333,3.8222227,2.7,1.7666667,2.4083335,5.211111,5.1666665,2.2666667,1.3666667,0.8688493,0.50277776,0.04,0.51111114,0.69166666,0.59999996,0.10000001,0.50000006,1.4000003,0.5999999,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.29166666,3.511111,5.0750003,0.5888889,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016666668,0.14444444,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.675,0.2,0.0,0.24444444,0.041666668,0.7777778,1.1777778,1.2833334,0.11111111,0.4,0.4666667,0.14166667,0.45555556,0.44444445,0.20833333,0.32222223,0.13333334,0.3333333,0.34166667,0.15555556,0.5833334,0.42222223,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.008333334,0.2777778,0.74166673,0.64444447,0.35000002,0.47777775,0.016666668,0.7444445,1.6666665,1.0916667,0.34444445,0.8333334,1.4111111,1.5083333,2.3444445,2.6777778,2.2500002,4.2222223,5.35,6.044445,4.575,9.444445,4.575,1.4777777,1.6666666,0.4083333,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07777778,1.475,3.0333335,2.3,3.8555555,5.3999996,7.7666664,9.211112,9.275001,8.666667,7.758333,6.433334,6.808333,7.4,5.655556,3.091667,2.4222221,3.7416666,4.3444448,4.6833334,4.411111,5.991667,5.8888884,5.7333336,6.8500004,8.577778,9.466666,9.455557,9.8,7.6,6.577778,5.8833337,5.5111113,5.7833333,5.833334,4.925,4.0666666,4.6666665,6.6444445,6.0555553,4.975,5.2333336,6.333334,7.611111,8.025,6.7000003,4.211111,2.5333333,2.766667,2.8500001,2.6666667,1.9083333,2.8333335,3.6444445,2.3083334,1.0666667,0.008333334,0.0,0.0,1.3062501,1.6,1.9833333,2.3625002,2.4833333,2.6875,2.1666667,1.775,1.5583333,0.8666666,2.21875,3.6666667,7.3687496,12.783334,17.893751,21.050001,21.1625,19.774998,18.375,14.837501,7.966666,6.58125,6.9666667,6.8625,3.5916667,1.7833334,0.5875,0.04166667,0.18125,1.4583334,11.35,17.100002,9.775002,4.4416666,0.99166673,2.59375,3.2833333,1.9125,2.8583333,1.8062501,0.40833336,0.43333337,0.20624998,0.5333333,0.075,0.0,0.0,0.0,0.116666675,0.49375004,0.43333337,0.90625006,0.9083332,1.21875,3.0583334,7.70625,12.016667,12.141668,11.76875,10.591666,6.950001,3.891667,2.0000002,2.0583334,1.7166667,2.13125,3.3333333,7.0812507,7.6833334,4.6687493,3.0666668,1.8950001,0.829394,0.09469697,0.575,1.2833333,1.3715476,3.9583333,2.84375,0.8333334,0.93333334,0.31875002,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.55,2.6625,0.29999998,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.4,1.30625,3.3416667,0.68125,0.45833334,0.0,0.10833334,0.32500002,0.0,0.0,0.0,0.14166667,0.0,0.06666667,0.15,0.13333334,0.23333333,0.0625,0.0,0.075,0.59166664,0.35625002,0.40833333,0.18333334,0.30625,0.18333334,0.112500004,0.1,0.38124996,1.1583333,0.64375,0.35,0.24166666,0.025,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00625,0.23333333,0.33125,0.35833332,0.10000001,0.425,0.175,0.0,0.19166666,0.20625001,0.34166667,0.81250006,1.0916667,1.1625001,0.71666664,0.7916666,1.75,1.125,0.90625,1.6583334,0.775,1.2333333,1.7562501,0.84999996,0.8416667,0.25,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.050000004,0.6416667,4.25625,7.175,2.9562502,1.7166667,3.9875002,6.8333335,8.266666,9.50625,9.566668,10.1,10.083332,9.212502,9.349999,8.516667,7.9437494,7.3083334,6.9375,8.191668,6.762501,6.5416665,7.03125,5.4666667,6.2,7.6499996,9.241667,10.575,10.508334,10.75,9.933333,8.150001,6.99375,5.8166666,5.9124994,6.1583333,4.2562504,3.941667,6.15625,6.308334,5.383333,5.3624997,5.891667,5.80625,4.9666667,4.8124995,3.4499998,2.4333334,2.1874998,0.675,0.51250005,0.7916667,1.25,1.275,1.9083335,1.4125001,0.0,0.0,0.0,0.0,3.358333,2.4666667,1.5444444,0.82500005,0.74444443,1.2166667,1.0888889,0.5083333,0.66666675,1.4555557,3.8583336,7.9888887,11.191668,12.488889,14.108334,15.755556,16.333334,16.033333,20.211111,15.599999,9.377778,9.45,9.655555,6.4333334,7.977778,8.1888895,4.6083336,3.8999999,1.725,2.1777778,4.4750004,11.98889,19.458336,13.544445,8.455556,14.108334,10.98889,8.450001,8.155556,4.2750006,0.4555556,0.38888893,0.11666667,0.0,0.0,0.0,0.0,0.0,0.31111112,0.7083334,0.5888889,1.5333334,1.1777779,3.925,8.622223,14.325002,17.311111,15.233334,12.683332,10.611112,5.408333,2.088889,1.9500002,1.888889,2.0555556,3.516667,6.077778,7.175,6.3111115,4.7750006,2.1333332,1.2666668,0.06666667,0.0,0.69166666,2.0666666,2.7250001,5.6,3.916667,1.4444445,2.5111113,0.98333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.22222222,1.0333334,2.1777778,2.2583334,0.9444445,3.4444447,0.33333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.055555556,0.61666673,0.9111111,0.5222222,0.26666668,0.35555556,0.44166666,0.055555556,0.125,1.4777777,1.3333334,0.23333335,0.05555556,0.06666667,0.13333334,0.15,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.23333332,0.19999999,0.11666667,0.044444446,0.033333335,0.0,0.0,0.0,0.055555556,0.0,0.0,0.25833333,0.6666667,0.11111112,0.05,0.022222223,0.0,0.0,0.0,0.26666668,2.15,0.22222224,0.0,0.68333334,0.0,0.0,0.0,0.0,0.0,0.06666667,0.22500001,0.0,0.0,0.0,0.0,0.0,0.0,0.008333334,0.0888889,0.25,0.42222223,1.1999999,4.666667,7.025,9.566668,10.2,9.466668,7.3444443,6.8500004,7.2333326,7.5333333,8.311111,8.711111,8.6,7.3222227,6.75,5.877778,5.4,6.6000004,5.9999995,5.5666666,7.5333333,10.891667,11.222223,10.900001,10.6,10.250001,11.0,10.555555,8.825001,7.288889,7.4583335,6.0555553,5.158334,6.2111106,8.849999,10.6888895,8.255555,5.975,4.5888886,3.9583337,2.766667,2.8500001,2.911111,1.3,0.53333336,0.36666664,1.0833334,2.4666667,2.1583333,1.3666667,1.5333333,0.50000006,0.0,0.1,0.20000002,0.058333334,5.8125,6.275,6.2666664,4.7312493,4.916667,5.5437503,6.1083336,6.88125,7.4833336,9.291667,12.0625,15.408334,16.4,9.075,6.1937504,8.4,8.599999,9.491667,11.133335,13.2125,4.0,2.03125,2.3,7.825,6.4583335,5.8416667,2.26875,0.66666675,1.0625001,1.6833334,2.9625,10.683333,17.5625,19.258335,17.050001,18.2,8.283334,4.75,5.9666667,0.98749995,0.725,0.48333335,0.03125,0.033333335,0.01875,1.1166667,0.21875,0.0,0.06666667,0.29375002,1.1666667,1.7875003,3.5166671,7.09375,10.158333,11.44375,9.466667,9.858334,9.2,7.0333333,3.36875,2.4666667,1.74375,2.4916668,2.9583335,6.21875,9.241667,9.725,7.7666674,4.3812504,0.66666675,0.17500001,0.3,3.0583332,7.775,13.741667,19.90625,16.816666,10.31875,3.2833335,1.3,0.3,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.15,0.033333335,0.0,0.0,0.16250001,1.0666666,4.033333,8.0375,1.8583333,0.65000004,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.125,0.5062501,0.0,0.1375,0.18333334,0.13333334,0.18124999,0.525,0.91875005,0.2,0.25625,0.53333336,1.2875,0.47500002,0.25833336,0.38125002,0.108333334,0.22500001,0.3166667,0.0,0.083333336,0.13333334,0.025,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.11666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.17500001,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.28333336,0.3375,0.19166666,0.40625003,0.0,0.0,0.0,0.09166667,0.0,0.0,0.0,0.075,1.24375,4.2500005,6.950001,7.6833334,8.283333,6.8312497,6.091667,6.21875,7.5,10.925,13.741667,13.916667,12.675001,12.191668,9.762501,5.6000004,6.6249995,10.358333,10.0,9.666667,10.341667,13.9625,13.683334,12.062499,11.591666,11.856251,12.325001,11.000001,9.86875,9.616668,9.6875,8.6,7.0687504,7.3166676,8.125,10.65,10.991667,8.756249,5.1083336,2.2687502,1.6999999,2.7500002,1.5666666,1.7416667,1.21875,0.46666664,0.23125,0.8166667,0.41875,0.23333335,0.7250001,0.33125,0.0,0.1375,0.46666664,0.2,4.6333337,1.7222222,1.2666668,4.1,7.5000005,10.95,11.644444,12.624998,11.933333,11.244444,7.750001,4.511111,2.2333336,1.9222223,2.2250001,4.5333333,8.908334,12.322223,11.866667,5.741667,2.288889,1.6333334,4.0888886,3.5249999,3.0888886,1.3444445,1.1916667,2.6777778,3.5333333,2.7777777,3.7,5.488889,6.9333334,13.088889,19.233334,14.483334,2.766667,1.3916667,0.61111116,0.725,2.7555556,2.5888891,0.6666667,0.35555556,0.14166667,1.2444444,0.47500002,0.0,0.0,0.18333334,1.2,3.5916667,5.0555553,7.783334,7.4666667,8.891666,12.011112,12.966667,9.099999,4.633333,3.4,2.7666667,4.683334,4.8444448,6.2333336,9.291667,12.2,9.675001,6.0111113,3.6583335,0.9666667,1.6666667,3.8777778,14.6888895,26.775002,37.944447,42.23333,41.11111,24.466667,13.466667,4.422222,2.9,2.6999998,0.5666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14444444,1.2833334,0.24444446,0.0,0.0,0.0,0.0,0.34444445,4.783333,7.6555557,4.8083334,1.0222223,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.033333335,0.0,0.0,0.06666667,0.36666664,0.38333336,0.9777778,0.85833335,0.53333336,0.275,0.15555556,0.36666667,0.3,0.23333335,0.76666665,0.51111114,0.2916667,0.18888889,0.0,0.022222223,0.3,0.21666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.18888889,0.13333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06666667,0.97777784,2.2583334,2.7000003,5.0000005,4.641667,3.7555556,5.1416664,7.0000005,12.316668,16.466667,15.544445,15.041666,13.988889,12.841667,9.811111,8.583334,11.177778,13.5,12.422223,12.733334,14.325,12.955556,13.383334,13.177778,13.991667,13.433334,11.677777,11.299999,11.8555565,11.033334,9.211111,7.3500004,7.2777777,7.991667,4.811111,5.9111114,5.733334,1.8333333,0.5,0.06666667,0.099999994,0.31111112,0.33333334,0.87499994,0.6111111,0.35833335,0.95555556,1.8166666,0.57777774,0.033333335,0.0,0.0,0.0,0.0,0.0,3.1833334,3.0333333,1.8333333,2.0,2.4222221,4.383333,5.7444444,5.6583333,5.5666666,4.933334,3.7916665,2.2444446,1.5083333,1.5111111,3.4583335,6.9888887,11.966668,15.555556,15.822223,12.741666,8.988889,6.841667,5.7222223,5.158334,2.5666666,2.666667,4.0833335,5.6000004,4.8500004,3.0777779,1.7166668,2.2333333,6.3749995,14.3,16.177778,12.583334,7.5,3.391667,6.0000005,7.2250004,7.422222,4.6555557,1.25,0.17777778,0.25833336,0.15555556,0.041666668,0.08888889,0.36666667,1.65,2.1222222,4.591667,9.3111105,12.241667,14.666666,15.208334,14.3,10.966667,7.008333,3.6222222,3.0083332,3.9111114,3.8249998,5.777777,8.077778,10.983334,10.077778,7.2916665,3.1000001,1.8083335,2.3111112,6.716667,10.0222225,13.077778,31.375002,33.800003,39.108334,42.96667,31.183334,18.055555,8.777779,5.725,3.9999998,3.05,1.4555556,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.044444446,1.4833332,1.2333333,0.075,0.0,0.0,0.0,0.0,0.058333334,2.6333334,5.566667,4.177778,0.25,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.022222223,0.26666668,0.22500001,0.7444445,0.7583333,0.5222222,0.3,0.22222222,0.5083333,0.62222224,0.44444448,0.70000005,1.0888889,0.49166667,0.044444446,0.0,0.0,0.06666667,0.13333334,0.055555556,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05,0.044444446,1.3749999,2.2222223,2.2333333,3.4000003,3.4111116,4.3916674,5.988889,6.1583333,6.6000004,11.466666,16.133333,17.033333,14.558334,12.266666,9.808333,11.744444,14.808333,12.644445,11.833333,13.558332,14.3,14.466667,13.544444,13.208333,13.3,12.811111,12.483334,12.522222,11.216666,8.444445,7.5166664,6.8888893,5.241667,5.5000005,3.5666666,1.9166667,0.8111111,1.1083333,2.5222223,2.983333,3.311111,0.82222223,0.9416667,0.6666667,0.225,0.3,0.27499998,0.044444446,0.022222223,0.0,0.0,0.0,0.0,0.0,0.0,0.016666668,0.016666668,0.03125,0.06666667,0.19375001,0.5166667,0.9625,1.1833334,1.2333332,0.83125,0.51666665,0.44375005,1.475,3.7937496,5.9416666,8.525,12.275001,18.866667,20.325,17.225002,10.90625,4.9166675,2.4562502,2.5166667,2.6416664,3.3249998,3.15,2.0750003,1.4416667,2.95625,5.466666,9.125001,11.55,10.208334,8.24375,11.583333,16.956251,21.041666,11.093751,5.608333,1.8583332,0.78125,1.0500001,1.5812501,2.2166667,0.6750001,0.075,0.375,2.7,6.4999995,10.3,17.966667,20.349998,18.558334,13.793751,7.8333335,4.175,4.0562496,5.166667,4.00625,3.2416668,4.1687503,6.8250003,8.766667,9.668751,7.700001,3.1875002,1.15,2.3625,4.391667,7.7875004,12.833333,12.658334,19.0,18.866669,19.48125,24.425001,20.606249,8.558333,4.0583334,1.7437502,0.375,0.16250001,0.25,0.118750006,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.2625,1.7666665,1.1125,0.058333334,0.0,0.0,0.0,0.0,0.0,0.5,2.35,1.13125,0.058333334,0.0,0.0,0.55,0.0,0.0,0.0,0.0,0.0,0.0,0.1,0.0625,0.083333336,0.1,0.375,0.39375,0.075,0.025,0.13333334,0.6333333,0.5875,0.84166664,0.8249999,0.15,0.025,0.0,0.0,0.0125,0.008333334,0.0125,0.0,0.0,0.0,0.0,0.01875,0.05,0.0125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.033333335,0.1375,0.4166667,0.7624999,1.4166667,1.1500001,0.91249996,1.65,3.1125004,3.6083336,2.83125,3.6,4.816667,8.256249,12.025,13.500001,12.475,10.362499,8.841667,10.14375,12.2,13.058333,15.381249,15.199999,12.637501,10.616667,9.112499,7.1333337,6.6499996,9.099998,8.750001,5.45,4.4750004,4.64375,4.5,3.9375,2.6000001,2.7083328,2.91875,2.2583334,3.5125,4.7583337,4.475,1.375,2.766667,2.0125003,1.2333335,0.7750001,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011111111,0.16666669,0.2166667,0.19999999,0.3,0.35555556,0.43333337,0.6666667,0.26666668,1.0833334,1.0000001,2.141667,2.2222223,3.175,4.9777775,6.35,8.288889,11.066667,15.458333,11.900001,3.4083335,0.9666667,1.0583334,0.8111111,0.73333335,0.325,0.31111112,0.89166665,2.588889,4.1833334,5.0333333,4.708333,5.7555547,5.555556,15.566668,16.4,16.050001,10.322222,7.316666,5.044444,2.1666667,1.4916668,1.0,0.075,0.0,0.06666667,0.7444445,2.5000002,6.2416673,9.744445,12.85,15.633334,15.224999,11.48889,6.15,4.2222223,3.5888891,2.5,1.6999999,2.75,4.911111,4.6916666,5.688889,6.6111107,5.9666667,3.8333333,1.875,2.5,1.2916667,1.6555556,7.8083334,17.999998,33.822224,40.150005,30.211113,26.258333,18.055553,10.875,2.9222224,0.41111115,0.108333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.11111112,0.5083333,0.44444445,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.13333333,0.8000001,0.06666667,0.0,3.2444444,2.2333333,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06666667,0.041666668,0.0,0.0,0.0,0.11111111,0.3333333,0.2888889,0.14166667,0.31111112,0.425,0.08888889,0.011111111,0.083333336,0.12222223,0.075,0.0,0.0,0.0,0.0,0.025000002,0.15555555,0.25833336,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.033333335,0.14166668,0.2,0.45555553,2.1083333,2.977778,2.8500001,3.0777776,1.7083334,1.0777777,2.1222222,4.941667,8.566667,11.208333,14.955556,15.791666,12.388889,11.658334,12.266666,10.888888,10.775001,9.855556,11.358334,12.500001,9.208332,7.744445,6.666667,6.216666,5.488889,4.691667,4.5,2.9416666,4.4444447,2.8,0.9111111,1.7444445,6.733333,5.3555555,3.4833333,0.95555556,3.1750002,3.8444448,3.266667,2.6833334,0.9777779,0.4,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.025,0.13125,0.075,0.225,0.26666668,0.59999996,0.51875,0.6333334,1.9,4.3833327,2.7,1.4083333,0.96875,0.5083333,1.8416668,2.78125,2.825,2.35625,2.3916667,2.7,2.0,1.65,2.2,3.5416667,5.15625,7.458334,6.4499993,4.4916663,3.475,7.0333333,7.575,13.94375,15.058332,13.3625,10.35,7.75,3.1499999,0.675,0.03125,0.0,0.0125,0.033333335,0.475,2.0416667,4.2583337,6.8500004,7.858333,12.6375,18.308336,15.80625,8.416667,5.2625003,2.8,1.85,1.7562501,3.1250002,4.6625,4.4999995,4.3062496,5.4749994,5.8,4.1875,4.9500003,3.175,2.9166667,4.3437505,8.075,22.55,47.575,51.958336,65.725,66.47499,46.94375,28.583334,22.831251,2.6750004,0.16666667,0.15625,0.016666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1,0.0,0.0,0.0,0.0,0.0,0.0625,0.025000002,0.0,0.0,0.0,0.0,0.11666667,0.275,0.17500001,0.0125,0.0,0.225,0.0,0.0,1.7375001,0.15833333,0.15625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.10625,0.0,0.0,0.0,0.0,0.00625,0.05,0.087500006,0.06666667,0.0125,0.26666668,0.0,0.00625,0.083333336,0.21250004,0.27499998,0.112500004,0.0,0.06666667,0.0625,0.14166668,0.64375,0.60833335,0.0625,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.033333335,0.43333334,0.7312499,0.6416666,1.625,3.9833336,2.5687501,1.5333333,1.3166668,2.3125002,4.3166666,6.8562493,8.841666,8.849999,9.575001,10.7125,9.825001,9.450001,13.868749,14.883334,12.94375,10.233334,9.374999,9.05,8.849999,9.062502,9.366667,7.125001,6.7666664,6.1312504,7.3500004,6.6937494,2.9499998,2.875,5.7000003,5.05,4.5875,3.7416666,2.5875,3.125,1.7416668,0.31875002,0.1,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.7687501,4.091667,2.21875,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.5833333,0.19999999,2.125,3.5222225,2.2333333,2.7416666,1.3222222,0.68333334,1.3555555,2.0583334,2.2333333,7.7777777,18.875,22.033335,18.316668,11.9,5.3083334,2.8333333,4.6583333,7.788889,12.844445,19.416668,14.5,9.783335,2.5111113,0.5500001,0.06666667,0.0,0.0,0.0,0.05,0.33333334,1.475,2.733333,3.5444446,6.4333334,11.588889,13.825001,17.38889,11.200001,4.5666666,1.6833334,0.5666667,0.9666667,3.2166667,4.7,4.4833336,4.7333336,4.4333334,4.5222225,4.8333335,6.341666,5.377778,4.125,5.2444444,13.016667,11.122223,41.833332,62.055553,62.944443,104.675,104.055565,64.875,50.466663,45.083332,5.4444447,4.788889,6.258333,5.5222225,2.8833334,0.59999996,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.083333336,0.0,0.0,0.0,0.0,0.041666668,0.19999999,0.0,0.0,0.0,0.0,0.0,0.041666668,0.32222223,0.19166669,0.011111111,0.0,0.0,0.0,0.0,0.0,0.28333333,0.38888887,0.0,0.0,0.0,0.0,0.0,0.033333335,0.13333334,0.116666675,0.0,0.0,0.0,0.0,0.016666668,0.044444446,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13333334,0.41111112,0.5583334,0.2888889,0.2777778,0.34166667,0.2,0.116666675,0.055555556,0.0,0.0,0.0,0.0,0.0,0.14999999,0.022222223,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.033333335,0.35000002,0.62222224,0.20833336,0.0,0.0,0.033333335,0.24444444,0.0,0.022222223,0.20833334,3.4333336,4.4,2.0666668,1.388889,0.8666666,2.522222,4.9333334,4.566667,5.0,7.7000003,9.366667,10.911111,10.811111,11.333333,12.233334,10.1,7.733333,8.075,8.433333,7.9666667,10.316667,7.988889,6.416667,5.1777782,4.3166666,3.6,2.7416668,1.4111111,2.3333333,3.4499998,4.0777774,3.4083333,0.7,0.0,0.0,0.0,0.1,0.06666667,0.0,0.0,2.6000001,0.44444445,0.0,0.0,0.0,0.0,1.0222223,0.17500001,0.0,0.116666675,0.15,0.050000004,0.075,0.043750003,0.058333337,0.00625,0.0,0.0,0.0,0.0,0.03125,0.058333337,0.55625,2.2083335,5.4812503,5.8749995,6.558334,5.81875,2.1916666,3.10625,4.083333,7.8812504,14.633333,21.250002,21.231247,14.083332,6.16875,2.4166665,2.5375001,3.4500003,6.7375,10.599999,9.858335,7.5937505,3.1500003,0.74375004,0.19166668,0.05,0.3166667,0.21666667,0.125,0.0,0.15,0.44166666,1.2125001,2.2083335,4.841666,12.724999,16.316668,15.76875,9.341667,3.6249998,1.1166668,1.0,2.4,3.241667,3.95,4.0083337,4.45,4.8416667,5.2625,4.241667,4.116667,4.8937507,2.225,4.8625,11.475,17.937498,20.600002,64.75625,76.49167,88.441666,132.50626,125.89167,59.908035,63.19167,48.924995,8.249999,6.925,5.6062503,4.5583334,2.8500001,0.975,0.081250004,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.29166666,0.43124998,0.0,0.0,0.0,0.0,0.0,0.033333335,0.075,0.0,0.0,0.0,0.0,0.0,0.0,0.043750003,0.033333335,0.0,0.0,0.0,0.0,0.0,0.65,3.1083333,0.8125,0.0,0.0,0.0,0.0,0.05,0.175,0.43125004,0.26666665,0.0,0.0,0.0,0.0,0.0,0.10625,0.0,0.0,0.0,0.0,0.0,0.0,0.00625,0.075,0.54375005,0.56666666,0.20833334,1.01875,1.5166667,0.43749997,0.05,0.0125,0.28333333,0.45000005,0.16666667,0.0,0.38750002,0.5166667,0.056250002,0.025,0.0,0.033333335,0.13333334,0.025,0.05,0.118750006,0.25833333,0.175,0.05,0.025,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1,1.5000001,2.525,2.125,1.2062501,0.675,2.025,1.9416666,3.3937502,5.483333,6.0374994,6.9833336,9.841666,13.15,17.46667,13.3875,8.958333,6.06875,5.0000005,5.0916667,3.7312498,2.2000003,1.7062502,2.0416665,1.4937501,0.95,0.05,0.16666667,1.8166668,1.8125,1.1083333,0.41250002,0.0,0.0,1.9000001,4.0583334,1.0125,0.0,0.0,1.1,0.225,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.19166666,0.43333334,0.34444445,0.24166667,0.21111111,0.1,0.08888889,0.033333335,0.0,0.0,0.0,0.0,0.06666667,0.44444445,2.0333333,7.988889,13.625001,9.333335,6.1555552,2.7583332,2.2888892,8.416667,16.811111,19.84167,16.91111,9.288889,4.4333334,1.8444445,1.2666668,2.4777777,3.575,4.811111,6.2666674,4.3555555,2.6222222,1.0083333,0.5555556,0.54999995,0.35555553,0.17500001,0.13333334,0.0,0.0,0.0,0.13333334,0.38888893,2.1583333,7.088889,11.555556,14.266666,14.433332,9.758333,5.0555553,2.525,1.3666668,1.7916666,2.7444446,2.9,3.8333335,4.4666667,5.4416666,5.9111114,5.5750003,4.3111115,4.2888885,2.5416665,3.8777778,8.883334,15.311111,24.191666,27.677778,62.266666,66.888885,87.888885,104.49167,105.22221,49.274998,55.233334,32.841667,4.377778,2.8888888,0.8833333,0.24444446,0.15833335,0.11111112,1.1916666,0.56666666,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.033333335,0.025,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.33333334,0.94166666,0.044444446,0.0,0.0,0.06666667,0.14999999,0.3333333,0.23333333,0.6888888,0.05,0.0,0.0,0.0,0.0,0.0,0.08888889,0.23333335,0.15555556,0.0,0.0,0.044444446,0.07500001,0.5777778,0.5416666,1.0666666,1.8444445,1.8916668,2.8333333,2.225,0.28888887,0.016666668,0.19999999,0.116666675,0.7333334,0.65555555,0.60833335,1.388889,0.34166667,0.1777778,0.2916667,0.044444446,0.23333333,0.275,0.44444442,0.15,0.6666666,1.3083334,0.9888889,1.1833334,0.36666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.033333335,0.125,0.10000001,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.22500001,0.6666667,0.25833336,0.0,0.05,0.73333335,1.3444445,1.3249999,0.33333334,0.26666668,1.2333333,3.825,8.866667,10.833333,9.555555,7.7555566,6.308333,7.244444,9.033334,9.377778,7.8500004,3.6999998,3.011111,0.52500004,1.6777779,1.1166667,0.35555553,0.525,0.8333334,1.0250001,4.477778,3.0777779,0.0,0.0,0.025,0.16666667,0.22499998,3.3333337,6.1,1.0416667,0.0,0.0,1.5111111,1.1333333,0.0,0.7444445,1.1166668,0.0,0.0,0.0,0.0,1.9666667,3.655556,3.9555557,2.7166667,1.8888891,1.4166667,0.7111112,0.42500007,0.022222223,0.0,0.0,0.0,0.0,0.033333335,0.3166667,2.4222224,2.4833333,0.37777779,0.16666667,1.6833334,7.544445,15.233334,19.6,13.625,6.1555552,2.7666667,0.975,0.99999994,1.6083333,1.9444444,3.45,3.2222223,2.2083335,2.2555559,1.5111113,0.6,0.8333334,0.21666667,0.1,0.0,0.0,0.0,0.0,0.13333334,1.1000001,3.1777778,5.366667,8.5,11.977778,13.075,8.444445,7.7833343,5.0666666,2.6666665,2.6333332,2.7833333,3.2555556,3.9444442,4.6916666,4.688889,4.3083334,3.7222223,2.6666667,5.3777785,4.0222225,3.0,8.388889,17.525,27.777777,38.550003,38.08889,56.833332,58.533337,61.055553,59.766666,54.333336,30.05,26.933334,11.458335,1.9666665,0.92222226,0.075,0.0,0.0,0.111111104,1.6416668,0.18888889,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.083333336,0.8333333,0.0,0.0,0.033333335,0.38333336,0.44444445,0.41666666,0.07777777,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.10000001,0.044444446,0.0,0.0,0.05555556,0.25,0.6666666,0.5416666,0.41111112,0.6666667,1.8166666,3.0222225,3.5500002,2.3000002,1.1833335,0.64444447,0.33333334,0.6,0.6333334,1.5166668,1.2888889,0.8833334,0.8333334,1.175,1.2,0.2111111,0.22500001,0.32222223,0.2916667,0.4888889,1.8083334,4.133333,3.0666664,3.2888892,1.0444444,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.51111114,1.3666668,0.85833335,0.11111112,0.0,0.0,0.0,0.0,0.0,0.011111111,0.0,0.60833335,2.6888888,1.1500001,0.033333335,0.1,0.3777778,0.5555555,0.5666667,0.11111111,0.016666668,0.26666668,1.2333333,3.3333335,5.6166663,4.6222224,2.7000003,1.0500001,0.25555554,0.42499998,1.0666667,5.4666667,10.055555,5.966667,3.6666665,2.7777777,4.35,1.9555557,0.90000004,1.0777777,0.74166673,3.3333335,2.7222223,0.0,0.0,0.05,0.13333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.7444445,1.1166668,0.0,0.0,0.0,0.0,0.50625,2.25,2.5333335,1.4250001,1.625,0.7562501,0.7250001,0.21874999,0.025,0.0,0.0,0.0,0.0125,0.025000002,0.22500002,0.85833335,1.1750001,2.1166668,3.625,5.7625,8.475,11.41875,11.891668,6.5437503,2.7416666,1.0333333,0.9562501,1.7416668,2.4250002,2.2083335,1.73125,1.0583334,0.60625,0.25,0.033333335,0.0,0.0,0.0,0.0,0.0,0.016666668,0.06666667,0.38125002,1.4833332,3.30625,6.0333333,8.818749,13.691668,12.291667,8.175001,6.625,6.618749,3.7166667,2.36875,1.8833332,4.9937496,5.866667,5.291667,3.8875,2.4916668,1.08125,0.68333334,1.4374999,3.5333335,4.075,10.537499,24.333334,40.74375,59.125,70.59375,62.949997,52.112503,54.35,32.55833,32.3375,21.250002,10.8125,6.55,1.275,0.15,0.025000002,0.0,0.0,0.075,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.42500004,0.68125004,3.1333337,1.0583334,0.0,0.0,0.1,0.13333334,0.0,0.025,0.0,0.0,0.0,0.0,0.25833333,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.2625,0.5500001,0.6312501,0.6666666,0.84166664,1.375,1.8083333,5.7125,9.325,5.03125,2.175,2.19375,2.2833333,1.7083334,1.4000001,1.5833334,0.65000004,0.52500004,2.50625,3.7916667,3.358333,1.2500001,0.8333334,1.6000001,0.94166666,1.7812501,3.3583333,5.04375,3.6499996,2.3833332,0.70625,0.84166676,0.06875,0.0,0.0,0.0,0.5,0.5625,0.0,0.0,0.0,0.0,0.20833336,0.28333333,0.01875,0.0,0.0,0.0,0.1,0.0,0.0,0.06666667,0.28333333,0.32500002,0.7083334,0.74999994,0.19999999,0.01875,0.5916667,0.59999996,0.33124995,0.25833333,0.075,0.0,0.0375,0.016666668,0.0,0.0,0.116666675,0.2875,0.44166666,0.6875,0.18333335,0.00625,1.0333333,1.1166667,1.6250001,1.6000001,0.32500002,0.3,0.76875,0.26666668,0.125,0.6666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.84166664,1.7437501,0.46666667,0.23750001,0.1,0.05,0.0,0.0,0.0,0.0,0.0,0.0,0.033333335,0.1,0.26666668,0.36666667,0.20000002,0.13333334,0.008333334,0.022222223,0.1,0.27500004,0.4,0.35833338,0.51111114,1.075,0.9777778,2.9666667,4.977778,7.3444448,8.25,5.3333335,3.0,1.1444445,0.9083334,0.54444444,0.41111112,0.15833335,0.41111115,0.23333333,1.9111111,4.1833334,2.0222223,0.8000001,0.42222223,0.7666667,0.125,0.07777778,0.041666668,0.0,0.0,0.0,0.7111112,3.6000004,7.055556,9.508333,12.155556,12.358334,9.844444,7.355555,4.233334,2.3333333,3.3999999,1.7222223,1.1250001,3.211111,4.958334,4.588889,4.166667,2.8166666,0.8666667,0.5500001,0.8777778,5.9083333,7.711111,12.5222225,26.008333,47.38889,63.408333,74.26666,72.808334,50.022224,36.86667,35.466663,13.0,16.908333,8.422222,2.1083333,0.47777778,0.083333336,0.0,0.0,0.0,0.0,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.36666667,3.5750003,4.966666,6.377778,0.65833336,0.0,0.0,0.0,0.0,0.06666667,0.3333333,0.11111111,0.0,0.0,0.22222222,0.0,0.0,0.0,0.06666667,0.15555556,0.083333336,0.011111111,0.06666667,0.5888889,0.8666667,0.9555557,0.9444444,1.15,2.0333333,3.2416666,5.933334,7.1416664,3.388889,1.1416667,1.8555557,1.1777778,1.4166666,1.6777779,1.2,1.0333333,1.1333333,2.877778,3.8888893,4.3,2.4222221,3.0083332,3.6111112,2.35,3.666667,3.3666666,3.1444445,3.022222,2.1166668,1.8111111,0.95000005,0.6666667,0.70000005,0.11111112,0.022222223,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.083333336,0.74444443,1.3000001,0.24444446,0.0,0.0,0.022222223,0.06666667,0.011111111,0.0,0.0,0.0,0.0,0.07777778,1.0500001,1.9333334,2.1916666,2.6111112,0.76666665,0.26666668,0.23333335,0.0,0.0,0.16666669,0.08888888,1.0833333,2.7555556,0.44166666,0.17777778,0.35555556,0.2,0.8000001,0.5666668,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.6222222,3.9583333,2.488889,1.4000001,0.4888889,0.13333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.116666675,0.4375,0.7083334,0.57500005,0.225,0.0375,0.016666668,0.4083333,0.89374995,1.5833333,1.7187499,1.8666666,1.925,2.05,2.2875,2.4416666,4.116667,5.21875,4.741667,3.86875,2.3416665,1.30625,0.6416666,0.35833335,0.04375,0.0,0.18125,0.083333336,0.33125,0.0,0.0375,0.09166667,0.18333334,0.0,0.0,0.0125,0.36666667,0.94375,1.9833333,3.666667,6.7437496,9.125,9.775,8.141666,6.64375,4.7999997,3.1166666,2.4374998,2.6666667,1.78125,1.8583331,2.1,2.6833334,2.2124999,1.275,0.90000004,0.89375,0.43333334,0.32500002,2.6416667,6.8687506,15.258333,25.941668,40.2,49.258335,49.7625,45.608337,39.574997,28.325,17.28125,14.425,14.283334,6.9375,1.65,0.4375,1.1666666,0.075,0.0,0.0,0.0,0.0,0.0,0.0,0.0625,0.7,0.16666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.4666667,4.0875,7.0,11.108334,1.2,0.0,0.0,0.0,0.0,0.11666667,1.1187499,1.2416666,0.21666667,0.056250002,0.0,0.0,0.18333334,0.7875,0.15,0.18333334,0.36249998,0.24166667,0.15000002,1.0666666,1.3499999,1.1333333,1.0916667,1.0625,1.425,1.3875,1.4833335,3.1937501,3.9750001,1.225,0.825,1.1583333,1.89375,3.4166665,2.9312496,2.2250001,1.71875,2.4750004,3.7250001,3.5937502,3.8333335,3.5187497,3.6999998,4.1875,6.5416665,4.6500006,3.091667,3.0583334,1.9312501,1.6,1.9749999,1.4583333,1.875,2.1250002,1.6916666,0.31875,0.525,0.89374995,0.52500004,0.13125001,0.43333334,1.1833334,0.41250002,0.025000002,0.0,0.0,0.48125,0.033333335,0.01875,0.29166666,0.6583333,0.14375,0.3,0.61875,0.09166667,0.0,0.0,0.0,0.66875,1.2499999,1.8749999,2.2583334,7.6812496,9.325,6.0,0.8916667,0.0,0.0,0.0,0.056250002,0.0,0.0,0.0,0.0,0.0,0.075,0.1125,0.05,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.3000001,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.011111111,0.17500001,0.5777778,0.97499996,0.92222226,0.45,0.07777778,0.022222223,0.041666668,0.08888889,0.21666667,0.5,1.1333333,1.8555557,2.2416666,2.7444446,3.8777778,2.5666668,1.4111112,0.66666675,0.56666666,0.3666667,0.011111111,0.17777778,0.3166667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08888889,0.4666667,1.0,1.3833334,1.9555557,2.788889,4.0666666,4.322222,2.85,1.8666667,3.1750002,4.5,3.266667,3.0416667,2.8555558,3.0416667,2.0,0.9,0.41111112,0.51666665,0.3555556,0.14444445,1.1750001,1.5222222,2.541667,7.7000003,15.05,23.577778,27.177778,28.308334,26.11111,22.108335,19.800001,17.691668,14.144445,8.608334,4.0111113,6.266667,3.3916667,1.2666668,0.38333336,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08888889,0.044444446,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13333334,0.2916667,0.33333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.058333334,0.0,1.225,9.155556,5.911111,1.4166666,0.0,0.0,0.0,0.0,0.0,0.23333333,0.8444445,2.177778,0.8416666,0.06666667,0.06666667,0.4,0.06666667,0.0,0.07777777,0.9083333,0.5,0.13333334,1.4444444,1.7416667,1.2999998,1.3222222,1.0250001,1.0555557,0.975,0.7666667,1.1999999,2.3222222,1.1500001,0.17777778,0.8111111,0.9333334,1.6111112,3.7166667,3.188889,2.841667,3.2777777,3.6444445,2.466667,1.9333334,1.7916666,1.2555556,4.166667,7.366667,3.9833333,3.1444445,2.9444444,1.475,1.1333334,0.8666666,1.5555557,3.7166667,4.2555556,3.7111113,2.4,2.877778,4.075,3.0666668,1.8416667,2.6555557,4.111111,4.375,2.2666667,1.7333333,0.044444446,0.0,0.13333334,0.22500001,1.0111111,3.911111,3.9916668,2.522222,1.85,2.7444444,1.6166668,0.9222222,0.29999998,1.5416667,1.4000001,3.8583336,3.3555555,0.33333334,1.3555555,1.9833332,2.2333333,6.2444444,9.125,2.888889,1.1166667,0.45555556,0.008333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1625,0.4166667,0.23333335,0.075,0.083333336,0.0625,0.008333334,0.0,0.0,0.0,0.05,0.0,0.0,0.0,0.0,0.0,0.0,0.125,0.4333333,0.7875,1.0500002,1.3249999,1.5166667,0.81250006,0.85,0.8583333,0.75624985,0.9166667,1.3125,2.7749999,3.53125,4.1166673,3.0749996,2.0062501,0.79166675,0.46875,0.8333333,1.55,1.7166667,2.4125,2.9583335,3.0666668,4.9249997,5.491667,10.55,16.816666,17.69375,20.616667,21.1,27.112501,29.783333,22.10625,14.416667,12.493751,7.016667,3.60625,0.4583333,0.3,1.1249999,1.2249999,0.53125006,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.7416667,1.8000001,2.4333332,0.92499995,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.043750003,0.52500004,0.16250001,2.1166668,5.825,2.85625,0.0,0.0,0.0,0.0,0.0,0.03125,1.3666667,5.383333,5.887501,0.85,0.0625,0.0,0.0,0.075,0.11666667,0.05,0.3333333,0.625,1.7249998,2.0937498,1.975,1.9333333,1.6437501,1.7250003,1.4625002,0.9333334,0.99375,0.8500001,1.2875,0.42500004,0.275,0.54375,0.99166673,0.85625005,0.81666666,1.7375,2.2583334,2.8249998,1.3625,0.28333336,0.21875,0.6166667,3.6,10.208334,5.7875,1.9833333,2.7916667,2.025,0.5083334,0.0,2.2416668,2.9625,2.9083333,1.9416666,1.65625,1.3750001,4.7999997,5.5666666,4.1625,4.9333334,6.4250007,7.4750004,4.1666665,2.25625,1.5416667,1.55625,2.3083334,0.4875,0.9333333,2.975,3.11875,2.1916668,3.7937496,3.25,2.9875,1.15,0.96666676,1.7562501,2.8916664,5.15625,4.25,2.74375,2.4333332,5.0375004,2.3916667,1.916667,4.1687503,5.166667,5.6562505,4.9833336,1.09375,0.59166664,0.025000002,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.43333334,0.36666667,0.13333334,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13333334,0.19999999,0.3222222,0.32222217,0.4333333,0.67777777,1.0333333,0.8777778,0.70000005,0.43333334,0.9888889,1.9583333,3.1222224,3.241667,3.1333334,1.1500001,0.32222223,0.26666668,0.29166666,1.3111111,2.325,6.877777,9.941668,10.788888,12.666667,18.38889,17.644444,26.283333,33.266666,42.05833,45.444443,45.716663,48.34444,45.78889,37.44167,31.966665,20.266666,11.422223,7.016667,2.266667,1.6333333,0.0,0.44444448,0.7166667,0.95555556,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.4333334,7.3666673,1.1888889,0.27500004,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.22500001,0.28888887,0.0,0.0,1.2555556,1.8916667,0.0,0.033333335,0.0,0.0,0.26666668,0.5333333,0.62222224,2.477778,6.3583336,3.7944443,0.2348485,0.033333335,0.0,0.0,0.0,0.016666668,0.24444444,1.3500001,1.988889,2.5000002,2.4,2.711111,2.7083335,2.7444444,2.2583334,1.3444445,1.5416667,1.3888888,0.775,1.0111111,0.5555556,0.575,0.8666667,0.94166666,0.48888886,0.94999987,1.8,2.2555556,1.8333335,0.59999996,0.56666666,0.62222224,1.7333332,6.5444446,3.8166664,2.2555556,2.4222221,2.125,0.54444444,0.125,0.67777777,1.25,1.3666667,1.3333334,1.9333333,1.8555555,3.0333333,6.166667,4.925,5.2333336,2.9444447,2.775,3.3555555,5.4333334,6.533334,6.375,4.5777774,1.4,0.46666664,0.51111114,2.3166666,4.177778,3.95,3.188889,6.2833333,4.4333334,2.8,2.0,0.62222224,3.025,7.255556,8.583333,4.9222226,2.0166667,1.9555556,2.5111113,8.05,8.2,3.9333334,0.7222222,2.0083332,1.2888888,0.033333335,0.28333333,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1,0.041666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.9250001,1.4333334,1.0777779,0.52500004,0.11111111,0.016666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.033333335,0.10833335,0.16666667,0.3,0.38333336,0.48888886,0.5583334,0.64444447,0.7916667,1.7111112,3.111111,3.975,3.0444446,1.7666667,0.81111115,0.4666667,0.6,1.3444446,2.9083335,3.8555555,8.983334,16.866667,23.875,31.98889,44.54167,55.333336,55.822224,55.44167,55.800007,53.341663,52.055553,50.233337,43.944447,33.7,22.616665,14.711111,6.7000003,2.5777779,2.3500001,1.0,0.32500002,0.0,0.08888889,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.21111113,6.191667,6.5,0.48333335,0.4666667,1.2583333,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.3166667,0.0,0.125,0.08888889,0.0,0.13333334,0.1,0.0,0.65555555,2.5416665,3.1444445,0.71666664,0.25555557,0.2,0.022222223,0.0,0.108333334,0.26666668,0.40000004,1.3777776,2.2916667,2.7,3.2444444,3.1416664,2.9444444,2.8416665,1.9777777,1.7333333,1.5333335,0.95000005,0.88888896,0.34444442,1.275,2.3555555,1.9083333,0.3111111,0.6416667,0.46666667,1.3,1.775,0.5888889,0.625,0.42222223,0.39999998,1.8888888,4.1416664,5.677778,4.588889,1.9916666,1.2888889,1.4333333,1.6222223,2.3583333,2.1777778,1.5333333,2.9416666,3.211111,4.4583335,3.8999996,2.4,3.2333333,2.8444445,3.0333333,4.444444,4.6833334,4.2000003,3.6416664,2.477778,5.45,4.0222225,0.43333334,0.40833336,1.3444445,3.9583337,2.1111112,1.8416668,3.1555555,6.1111107,5.0583334,0.92222226,1.5583334,4.0222225,4.516667,2.511111,2.5250003,5.9555554,6.755556,4.55,2.911111,0.68333334,1.5111111,1.5916669,2.0555556,1.6333334,1.0666667,0.25555557,1.8416667,2.7666667,3.9583335,3.5222223,1.3166666,1.7777779,2.8555555,3.4083335,1.7222222,0.775,0.35555556,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0125,0.29999998,0.75000006,0.93125004,0.6583333,0.33750004,0.06666667,0.0125,0.0,0.0,0.0,0.06666667,0.10625,0.63333327,0.08125,0.0,0.0,0.0,0.0,0.087500006,0.15833333,0.025,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016666668,0.15000002,0.2166667,0.18333334,0.22500001,0.6,1.65,2.4,2.425,2.7583334,2.6166666,1.5187502,0.8250001,0.40625,1.6916668,2.6625,7.2166667,11.383333,19.98125,29.208334,48.343754,57.575005,65.875,67.59167,56.787502,51.641666,42.9,38.6625,35.7,33.65625,30.099998,20.143751,13.691668,8.866667,2.7812502,1.1750001,0.36874998,0.2,0.73749995,0.6583333,0.081250004,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.083333336,1.2,2.0666668,1.54375,0.47500002,0.075,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14999999,0.29166666,0.0,0.033333335,0.0625,0.0,0.18333334,0.53125,0.725,0.34375,0.25833333,0.18125,0.125,0.1,0.10625,0.20833334,0.30625004,0.25833336,1.0187498,1.55,2.1333332,3.0500002,2.9083338,3.2375002,2.7083335,2.1125,0.82500005,0.7125,0.35,0.0,1.4000001,3.5500002,4.5437503,1.8916667,1.98125,1.6499999,0.85833335,0.71874994,0.84999996,2.1625,2.0166667,0.73125,1.0083334,4.60625,4.2583337,3.2,1.3062499,2.25,3.1687503,4.375,3.175,3.2083335,2.516667,3.575,3.9749997,6.0687494,7.5250006,5.275,3.2583337,2.3083332,3.90625,4.866667,2.74375,2.0666666,3.1374998,2.2333336,3.8125,1.5500002,0.6416667,0.19375001,0.38333336,0.5375,0.050000004,0.35625,2.8666666,5.258333,5.30625,6.1916666,5.6812496,2.5,3.23125,1.8666667,2.125,7.7416663,7.283334,3.1625,2.5666666,3.05,4.983333,8.3,8.066667,8.35,7.35,4.666667,6.7374997,8.275001,8.9,8.675,5.2124996,3.2583334,2.1833336,1.5124999,2.2749999,3.13125,3.0250003,1.46875,0.25833333,0.6166666,0.575,0.425,0.48125,0.21666667,0.118750006,0.016666668,0.0,0.0,0.0,0.0,0.0,0.0,0.23333333,0.42222223,0.43333334,0.9583334,1.8777778,2.3083334,1.2333333,0.25833336,0.0,0.0,0.3,0.15555556,0.6833333,0.54444444,0.54999995,0.5,0.36666667,0.13333334,0.13333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.05,0.0,0.016666668,0.11111111,0.13333334,0.15833335,1.0000001,1.9250002,1.9000001,1.8583335,1.7444444,2.4444444,2.9,6.1,7.625,16.611113,20.25,33.988888,43.555553,52.64167,54.533337,51.25833,49.93333,36.100002,27.400002,19.416668,16.333334,14.355556,11.775,9.777778,7.241667,4.877778,1.6333334,0.7,0.5888889,0.275,0.51111114,0.80833334,2.3000002,2.2,0.5111111,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.21666667,0.16666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06666667,0.06666667,0.016666668,0.1,0.27499998,0.40000004,0.0,0.525,0.23333332,0.34166667,1.3222224,0.52500004,0.9,0.32222223,0.3416667,0.67777777,0.2916667,0.3666667,0.75000006,1.0888889,2.2444444,2.2416668,2.3777778,2.3833334,3.4,2.2933333,1.0611111,0.475,0.1888889,0.0,0.94166666,2.9888892,5.8583336,2.3222222,1.9833335,3.1666667,2.1,0.68333334,0.22222222,1.8583333,2.2666667,0.65833336,0.11111111,2.466667,4.311111,2.533333,0.725,1.2888889,3.5000002,4.2444444,3.0333335,3.977778,5.866667,5.0750003,4.577778,6.2500005,10.655556,10.275,5.533334,2.8333335,3.1166668,3.0888886,3.3916667,4.1222224,2.8666666,3.2444446,3.016667,0.5555556,1.5333333,2.0166667,1.0444446,0.075,0.0,0.16666667,1.2777777,1.9444444,4.041667,4.088889,2.3166668,1.3,2.8833332,2.4222224,2.3583333,6.3,4.955556,2.8416667,3.4666667,1.5083334,2.8111112,9.008333,9.866667,12.233334,17.558334,16.077778,7.258333,3.4,4.275,4.7666664,4.4833336,1.0444444,0.9888889,0.9,2.2888892,3.5749998,3.6444445,0.7416667,0.20000002,0.32222226,0.24166667,0.16666667,0.12500001,0.10000001,0.008333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.1437501,1.9083334,2.025,2.2375,2.9583333,3.5125003,3.2083333,1.9125001,0.825,0.6666666,1.8125,2.3083334,2.8374999,1.9750001,1.5875,1.575,0.9562501,0.38333333,0.29166672,0.025,0.0,0.0,0.0,0.0,0.38333336,0.16666667,0.35000002,0.5,0.46249998,0.48333335,0.40625003,0.35833335,0.31875002,0.35,0.275,0.61875004,1.2916667,2.9812498,4.4,6.2875004,8.191668,10.008333,11.1875,20.091667,25.868752,37.925003,45.081253,50.316666,50.149994,39.5125,35.391666,20.706251,14.508335,7.45625,4.0833335,1.28125,1.4000001,1.7916667,1.8437502,1.2750001,0.7125,0.6333333,0.7625,0.95,1.125,1.70625,3.8583336,3.86875,2.391667,0.93750006,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.00625,0.0,0.0,0.0,0.175,0.5083333,1.175,2.54375,1.425,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.125,0.2,0.0,0.0,0.0,0.0,0.0,0.087500006,0.15,0.075,0.35833335,0.23125,0.32499996,0.27499998,0.0,0.05,0.41875,3.1000001,8.075,7.2250004,2.9916668,3.4437501,2.098485,0.35000002,0.7583333,1.325,2.591667,4.991667,6.9500003,7.0166664,8.71875,6.560606,4.261607,2.338889,0.31420454,1.0583333,0.375,1.71875,2.1,4.15,2.775,6.93125,8.791667,7.2666674,3.61875,0.77500004,1.4124999,1.5666668,0.46249998,0.0,1.13125,4.991667,4.4083333,1.2750001,1.1916666,1.7375,3.9916668,3.35,2.7416668,4.7250004,5.79375,6.441667,3.4062498,5.15,11.96875,7.8166666,2.3833334,2.93125,3.5749998,1.7624997,3.016667,4.85625,6.0,4.6312504,2.7333333,3.4416666,3.19375,3.25,1.9562498,1.9416667,2.5,3.575,6.5,6.9249997,2.4916668,3.13125,3.3833334,2.74375,3.1416667,3.1062498,3.8416667,2.825,2.00625,2.9500003,1.7625,2.8,3.29375,4.2250004,2.1833334,2.7312498,2.5666666,1.29375,1.4083333,2.1937501,2.6583333,1.5687499,1.0833334,1.2416666,1.05,1.1750001,0.30625004,0.30833334,0.15,0.38333336,0.55,0.6437501,0.8,0.39375,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.5666666,2.488889,3.5333335,3.1416667,1.8444446,1.2750001,1.0444443,0.9,1.4333334,2.3777778,2.4833336,1.4333334,0.79999995,0.36666667,0.7083333,0.26666668,0.18333334,0.0,0.0,0.0,0.0,0.0,0.0,0.15,0.97777784,2.1777778,2.516667,1.688889,1.0000001,0.93333334,0.6,0.59999996,0.45000002,1.1,1.4222221,3.5749998,7.166667,11.791666,14.8111105,21.233334,20.655556,24.911112,32.816666,46.388893,51.108334,50.266666,39.575005,33.61111,24.288889,12.8,8.744446,4.5083337,1.1555557,0.74166656,0.7,0.025,0.17777777,0.033333335,0.40000004,0.76666665,1.125,1.7111113,2.4083335,3.3666663,6.5111113,4.6416664,4.0333333,1.2333333,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.23333335,0.2166667,0.011111111,0.0,0.0,0.09166667,0.36666667,1.9444445,3.716667,3.4777777,0.52500004,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06666667,0.24166666,0.18888889,0.033333335,0.0,0.0,0.0,0.0,0.0,0.43333334,0.20833334,0.055555556,0.0,0.0,0.0,0.0,0.0,1.3833333,8.655556,14.216666,11.955556,7.166667,2.5583334,2.2111113,3.15,2.4,1.7333333,2.7666667,4.8111115,9.491667,13.044444,15.433333,10.577777,11.75,10.366668,2.1166668,1.3111112,1.1,2.8666668,2.1555557,6.8,6.2333336,11.349999,14.044445,12.022223,9.016666,3.988889,3.2833335,1.9777777,0.37500003,0.0,0.5,2.9000003,2.4444447,1.8000002,2.7444444,1.7083334,1.5666666,1.55,0.35555553,1.1222223,2.7666667,5.2666664,5.508333,5.4444447,8.733334,10.244445,7.377778,2.8583333,2.1000004,1.2500001,1.7,2.9,4.5222225,3.4500003,2.7333336,3.6,5.016667,4.811111,1.8166666,0.9555556,0.20833334,1.1000001,2.6666665,3.625,2.8888888,2.6916666,2.6222222,4.875,4.2222223,6.1000004,7.422222,7.666667,5.9500003,8.155556,9.458334,6.5666666,2.25,0.53333336,0.8888889,1.6666667,0.6888889,0.14166668,0.33333334,0.44166666,1.3777778,3.0833333,4.5333333,4.255556,5.5333333,6.1444445,4.766667,4.711111,2.7333333,0.54444444,0.22222222,0.52500004,0.26666668,0.15,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,3.9250002,3.8333335,3.6833334,2.8062499,2.1666667,1.58125,1.2,0.6875001,0.425,0.46666667,0.13125001,0.125,0.24374999,0.36666667,0.225,0.008333334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.22500001,0.5,0.61666673,1.075,2.3833334,1.8062502,1.2166667,1.0875,2.7416666,3.55625,5.9416666,8.400001,15.06875,19.908333,24.51875,25.550001,23.743752,25.824999,29.558334,35.037502,40.333336,38.256252,30.758333,23.737501,18.108332,13.891666,8.375,4.8916664,2.2749999,1.1416667,0.9125,0.8249999,0.63125,0.39166668,0.675,0.89375,1.0666667,2.0187497,3.4916668,4.1125,5.200001,4.866667,1.5625,0.075,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.03125,0.49166667,0.0375,0.0,0.0,0.0,0.033333335,0.40000004,0.94166666,0.29999998,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0125,0.0,0.0,0.0,0.0,0.0,0.083333336,0.4375,0.29166666,0.0125,0.0,0.0,0.06666667,0.033333335,0.21875,1.7166667,11.868751,18.341667,12.83125,4.875,2.2833335,2.04375,3.2083335,4.2937503,4.416667,2.9375,1.8416668,2.691667,4.8,8.849999,11.55625,12.091667,10.44375,12.275758,5.2312503,1.4833333,2.1666667,4.0562496,8.458334,8.50625,5.25,6.4624996,13.15,14.733334,7.1187506,8.25,5.6374993,4.1,1.8062501,0.5,0.36875,2.1833334,1.2166668,0.81875,2.125,3.45625,4.941667,3.69375,1.8333335,1.15,1.46875,3.8,4.075,2.8249998,2.56875,5.1083336,7.2666664,5.6187496,5.2499995,4.5125003,4.5583334,3.8062499,2.125,1.3500001,0.9416667,1.1666667,3.1125002,2.2916667,1.05625,0.116666675,0.10625,0.975,1.8166668,2.125,1.6416667,0.96875,2.05,4.05625,5.625,8.431251,8.625,8.116667,7.5625,8.55,10.112499,8.791666,7.23125,6.2250004,5.3166666,2.7437499,1.85,2.2625,2.8583333,3.3687499,4.516667,2.0749998,1.4000001,1.8166667,5.2375,9.775,8.349999,3.8166666,3.06875,0.5833333,0.40833336,0.79375005,1.2416668,1.525,0.35,0.112500004,0.3166667,0.45000002,0.0625,0.0,0.0,0.0,0.0,6.625,5.7000003,5.2000003,4.533333,3.3111115,1.5916667,0.8,0.8416667,0.64444447,0.6666666,0.48333332,0.1888889,0.15,0.08888889,0.116666675,0.23333335,0.32500005,0.31111112,0.73333335,0.125,0.11111112,0.13333334,0.42222223,1.0999999,0.5777778,0.8888889,0.88333327,1.1666667,1.4333334,2.211111,4.208334,5.344445,9.550001,13.622223,16.88889,23.499998,26.655558,26.499998,25.322224,25.833332,26.855556,32.38889,35.300003,39.666668,39.49167,35.81111,27.041666,19.577778,16.455553,10.016667,6.4000006,3.5,2.4555554,1.1916667,0.57777774,0.125,0.0,0.0,0.0,0.099999994,1.1166668,0.8111112,0.5416667,0.26666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.20833334,0.24444446,0.075,0.0,0.0,0.0,0.0,0.28333333,1.3555555,0.9083333,0.07777778,0.0,0.0,0.0,0.075,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13333334,0.2777778,0.06666667,0.0,0.0,0.0,0.033333335,0.25555554,0.9777778,5.0916667,11.822224,18.266666,20.400002,11.383333,4.088889,0.98888886,1.3083334,2.0888886,5.625,7.2555556,5.9999995,2.8000002,2.2333333,2.3750002,5.922222,9.483334,11.000001,8.049999,8.0,6.933334,6.1666665,6.711111,7.8916664,8.622222,5.450001,3.7555559,3.7583332,10.433334,15.677777,5.216666,7.4888887,6.825,4.555556,3.8416667,1.3222222,1.1583334,1.3666667,0.61111116,0.4166667,1.0000001,1.7666667,6.766666,8.366667,3.6666667,2.5555558,2.85,6.6777782,5.2249994,3.0666666,3.5083332,3.2,2.766667,3.6499999,1.9555556,1.3333335,1.9333335,2.5916667,3.311111,2.125,1.9222221,2.8333335,1.85,1.2888889,1.6666667,2.8333335,3.4750001,5.333333,6.955556,7.4333334,4.688889,3.65,4.322222,4.3666663,6.7666664,7.833333,5.7666674,5.833334,6.408334,6.422222,7.5750003,8.988889,9.375,5.644444,3.7444444,3.6749997,4.3444448,4.2583337,3.7555554,3.4499998,2.677778,1.6916667,0.7,0.15555558,1.4416667,2.1111112,2.2083333,1.2222222,0.20833334,0.0,0.0,0.016666668,0.4666667,1.05,0.9333334,4.841667,5.6555557,3.2666664,0.65,0.0,0.0,0.0,0.0,9.024999,8.25,7.716666,6.7374997,5.55,4.51875,4.533334,4.45625,3.7833333,3.3666668,2.53125,2.0833333,1.6624999,1.3416667,1.11875,1.1916666,1.60625,1.5166667,1.4583334,1.4125,1.7166667,1.35,1.0583334,0.8875,0.575,0.28333333,0.26250002,0.3,1.04375,3.15,6.41875,12.233335,20.506252,31.791668,42.583332,45.306248,45.583336,42.068752,41.108334,46.30625,57.616665,65.34167,64.293755,60.81667,48.725006,37.00833,27.6375,20.525,14.308333,8.475,2.35,1.45,0.24166667,0.09375,0.18333334,0.03125,0.0,0.0,0.0,0.0,0.1375,0.1,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03125,0.125,0.23125,0.0,0.0,0.0,0.0,0.112500004,0.85833335,0.46250004,0.5333333,0.24374999,0.025,0.0,0.06875,0.083333336,0.0,0.0,0.0,0.0,0.0,0.0,0.33333334,0.58750004,0.5416667,0.20625001,0.0,0.0,0.0,0.06666667,0.00625,0.0,0.0,0.0,0.0,0.125,0.84374994,3.966667,13.141666,21.7,24.441666,21.706253,13.283334,4.3999996,2.4583333,2.275,1.7125001,2.0666666,3.0000002,5.308334,3.6875002,2.7749999,1.8666668,1.3625,5.125,7.8062506,8.225,5.08125,4.85,9.56875,9.325001,8.925001,6.4937506,3.666667,2.0625002,1.7416664,1.8062501,7.5083327,11.1,4.1000004,6.058334,14.25,7.725001,1.9250002,2.5166667,5.6000004,3.5583334,1.0833334,1.3499999,2.341667,0.65,2.1499999,3.825,3.8666668,3.1750002,2.4125,3.3500004,5.1875005,5.383333,2.9062498,2.9666667,1.0500001,1.30625,1.3333334,2.35,2.4416666,3.29375,3.8166668,1.8687499,1.4749999,1.1916666,1.125,1.45,2.8750002,4.3083334,3.9624999,2.841667,2.975,3.35,3.9250004,4.3875003,5.1000004,3.8625002,4.225,4.625,5.2833333,6.025,7.5,8.808333,9.812501,9.066667,8.1875,6.333333,4.4666667,2.1625,1.4083334,2.85,4.6749997,5.11875,3.8833332,6.725,8.591668,7.0666666,4.4687505,3.9333336,3.45625,2.1333332,1.86875,1.7250001,1.2583333,1.60625,4.533334,10.418751,9.966666,6.2999997,2.9083335,1.0416667,0.51875,0.18333334,0.0,0.0,0.0,6.3750005,6.3888884,6.3222218,6.6250005,6.5555563,6.7666674,7.2333336,7.0083337,6.333333,5.966667,5.5416665,5.033334,4.4916663,3.9111114,3.6666667,3.3333335,2.5416667,1.6666667,1.6,1.375,1.2666667,1.5416665,0.7111111,0.7083333,0.5444445,0.31111112,0.24166669,0.51111114,2.7083337,7.0666666,12.100001,19.644445,35.483334,42.355556,47.144444,40.425,36.511112,36.8,42.41111,49.125004,64.1,72.18889,63.708332,60.477783,52.666668,34.86667,25.966667,18.07778,9.111111,3.3500001,1.2222223,0.025000002,0.0,0.075,0.1,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016666668,0.033333335,0.008333334,0.0,0.0,0.0,0.0,0.0,0.13333334,0.4,0.28888887,0.79166675,0.5,0.0,0.0,0.033333335,0.1,0.1,0.0,0.0,0.0,0.055555556,0.2888889,1.125,1.1,0.30833334,0.5222223,0.33333334,0.23333332,0.18888889,0.625,0.29999998,0.175,0.23333332,0.425,2.1444445,6.4083333,13.111112,17.277779,22.041666,22.099998,10.933334,2.7777777,2.0833333,2.5000002,3.5,2.4333332,0.93333334,0.8666666,2.0111113,1.3666667,1.1444445,1.2555556,1.45,4.577778,5.9,4.5111113,2.975,5.366667,7.908334,8.611112,10.311111,7.666667,2.7000003,2.491667,1.5777777,2.1583333,4.566667,4.811111,2.8666668,3.3222225,11.933334,10.544445,2.4833333,7.977779,14.149999,9.277778,3.2333333,2.425,2.0666666,0.45,1.6111112,3.9333332,3.3444445,2.4111114,2.6916668,1.6222222,2.7416666,6.588889,5.6416664,6.3444443,3.0888891,2.4166665,2.288889,3.3583336,4.911111,5.758334,3.0,1.8666667,1.9555554,2.4888887,2.4583333,1.1111112,0.9083334,1.0888889,0.4916667,0.13333334,0.0,0.16666667,1.0777777,2.9583333,3.2888892,2.1416664,3.4888892,4.3166666,5.588888,7.6444445,8.45,11.2,13.125001,12.766666,7.641667,4.3333335,7.0333333,5.575,4.377778,4.708333,1.8444445,0.95000005,1.2,3.4916668,5.122222,3.2555556,5.3666663,9.555555,9.016666,6.966666,6.0666666,7.6999993,9.433333,8.733333,5.0111113,5.1833334,1.7222223,1.3833334,3.3555555,1.6333333,0.3,0.0,0.0,0.0,0.0,3.3916664,3.3,2.8,2.2749999,2.5666666,3.475,3.0888891,2.7833333,3.311111,4.233333,4.366667,4.277778,3.775,3.6777778,2.1416667,1.5555556,1.5416666,1.388889,1.2777778,0.76666665,0.74444443,1.25,1.0777779,1.0083333,1.2888888,0.9555556,0.91666675,2.6111114,7.9416666,13.21111,18.791668,25.18889,29.491669,32.86667,33.711113,31.916668,33.100002,36.191666,40.47778,43.133335,46.38889,49.255554,40.483334,33.41111,27.233334,17.955557,9.1,4.2222223,2.1333334,0.9916667,0.38888887,0.025,0.27777776,0.74166673,0.62222224,0.075,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.008333334,0.0,0.0,0.0,0.0,0.0,0.022222223,0.16666667,0.33333334,0.44166666,0.22222224,0.3416667,0.36666667,0.033333335,0.05,0.57777774,0.51666665,0.16666667,0.025,0.15555556,0.116666675,0.26666665,1.5111111,1.625,2.1333332,2.575,4.1888885,3.9416668,3.2222223,3.411111,3.6250002,2.6222222,3.4833336,5.122223,8.158333,12.622223,15.833334,15.711112,14.877778,12.533333,8.277778,2.775,1.5111111,2.6583333,3.0666668,3.8111112,1.5583334,0.5888889,0.7083334,0.21111111,0.8083333,0.90000004,1.2,1.925,3.5222225,2.9,3.0666668,4.775,7.1444445,10.116666,9.388889,7.888889,6.8916674,3.4666667,2.225,1.6999999,2.275,4.166667,3.8111115,1.8083334,1.588889,3.9583333,4.922222,4.333333,11.288889,14.116667,10.644445,5.3555555,4.116667,3.4444444,1.125,1.1222223,1.95,1.6555557,1.1333334,2.7416668,2.0222225,1.3333334,4.3333335,10.325001,11.555555,6.333333,4.716667,5.266667,5.9083333,9.1444435,8.3,4.1444445,3.6916668,3.7555554,3.0333333,1.5666668,0.6888889,0.31666672,0.39999998,0.5166667,0.4666667,0.15555556,0.36666664,0.7444444,1.6416668,3.722222,4.425,5.722222,7.375,7.0777774,7.6,6.6583333,5.5,5.841667,5.5888886,4.958333,3.5222228,2.5333333,3.391667,3.1111112,3.7166667,2.4444447,1.0500001,1.8222222,3.9500003,2.522222,0.8777778,2.0416667,3.6777778,2.358333,0.7666667,0.6916667,1.9555554,3.5888891,2.5833333,1.011111,0.875,0.5666667,2.308333,3.3333333,2.8000002,1.2416666,0.0,0.0,0.0,0.0,0.71875006,0.40000004,0.4,0.32500005,0.49166673,0.45000005,0.57500005,0.75625,0.95000005,0.93333334,1.2812501,1.0333333,0.8687501,0.53333336,0.45625,0.56666666,0.58750004,0.625,0.8,1.0875,1.2083334,1.9375,2.2916667,1.80625,1.825,1.8833333,3.08125,7.3833337,13.55625,14.666665,18.45,22.041666,26.25625,31.983335,37.958336,37.24375,38.29167,37.725002,40.941666,41.9375,41.666668,36.683334,27.7625,17.516666,11.8125,9.25,6.15625,2.1416667,2.125,0.90625006,0.033333335,0.4875,1.1333333,1.4062499,0.525,0.03125,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14999999,0.44374996,0.116666675,0.01875,0.0,0.0,0.0,0.0,0.0,0.016666668,0.0125,0.0,0.0,0.0,0.03125,0.14166667,0.53333336,0.52500004,0.30833334,0.3,0.32500002,0.35625,0.44166666,0.53125,0.9,2.2333333,3.55625,5.05,8.375,8.433334,8.400002,9.641668,7.641668,4.98125,8.208334,13.68125,17.291666,19.8875,18.166668,15.293751,11.233333,8.816667,3.3750005,1.6083333,1.5312501,2.0083334,2.7812502,2.3,1.3416667,0.7562501,0.75,1.1187499,0.675,0.28125,0.35,0.71666664,2.0874999,2.3666668,1.9812499,4.375,7.89375,8.625,7.4375005,4.333334,3.35,5.5625005,3.0083332,2.2750003,1.6666666,1.7125001,3.3166668,2.0416665,1.6312499,1.7916666,2.1374998,2.9916668,5.1937504,9.883332,9.181251,12.741668,8.875,5.3187504,6.283333,5.1062503,2.2416666,1.0687499,0.6666667,0.9666667,0.6874999,0.92500013,1.4187499,1.6916667,3.56875,7.124999,5.841667,8.793751,15.6,17.418753,12.283334,7.781251,6.275,4.84375,4.516667,1.5166667,0.11875,0.016666668,0.50624996,2.5916665,1.15,0.34166667,0.25000003,0.55,0.61666673,0.9312499,2.6583333,3.3812501,2.4166667,1.9687501,1.5916667,1.2750001,0.84374994,0.40833336,0.25,0.18333334,0.2125,0.0,0.1,0.15,1.0833334,2.6,1.7916666,0.6625,0.075,1.35625,3.2500002,5.85,6.3812494,2.9,1.9875001,0.55833334,0.54375005,0.43333334,0.7166667,1.1625,0.69166666,0.0,0.06666667,0.58124995,0.5416667,0.3,0.0,0.0,0.13749999,0.06666667,0.0,0.008333334,0.022222223,0.033333335,0.008333334,0.0,0.0,0.45555556,0.125,0.26666668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.1,0.44444445,0.6666667,0.5777778,0.84999996,1.388889,1.8333333,2.777778,4.188889,8.775,12.1,15.475,17.833334,23.608334,33.166664,36.26667,33.722225,34.2,36.233334,35.45556,34.333332,29.011112,30.591667,34.68889,33.722225,38.61667,39.66667,19.316666,5.5666666,3.2416668,0.3888889,0.13333334,0.108333334,0.38888887,0.6333334,0.7,0.19166666,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.32500002,0.0,0.0,0.033333335,0.0,0.0,0.0,0.0,0.13333334,0.05,0.0,0.08888889,0.06666667,0.0,0.083333336,0.099999994,0.0,0.0,0.66666675,1.7833332,2.1333334,1.0250001,0.22222224,0.32500005,0.33333337,1.0583333,1.5,2.4222224,4.5750003,6.2555556,7.1333337,9.422222,10.041668,6.9222226,6.4111114,9.658333,17.07778,23.091667,17.9,10.0,7.3555555,6.333333,4.0444446,1.2777777,0.89166665,1.3444445,1.8833332,1.7666665,1.0166667,0.25555557,0.988889,1.3666668,1.0,1.1833334,1.2333333,0.57500005,0.45555556,0.7111112,2.625,3.7222223,2.75,4.788889,8.075,6.622222,2.3249998,0.7111112,1.7666667,3.6916666,1.2111112,1.1416668,2.1333332,1.3666667,2.5,2.0555556,1.1750001,0.91111106,0.96666676,1.7111111,2.4583335,3.2555556,5.633333,12.1888895,10.366666,8.641667,10.3,10.616668,6.0222225,2.4666665,1.7777778,0.93333334,0.30000004,0.47777778,0.31666666,1.1333333,1.6416669,1.7111112,2.4,4.1416664,8.28889,9.641666,5.288889,3.1916668,1.9222223,4.2083335,3.7333336,2.7555556,3.7916667,3.0777779,1.9000001,2.6333334,5.125,5.1,3.011111,0.96666676,0.45555556,0.47500002,0.25555557,0.24166666,0.24444446,0.20833333,0.12222222,0.044444446,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.9083333,2.8444445,1.525,0.13333334,0.22500001,1.5444444,2.9777777,4.116667,1.7,3.1166668,3.6555557,2.641667,2.8333337,1.2666668,0.7833333,1.0666667,1.1333334,0.033333335,0.0,0.2,0.33333334,0.0,0.0,0.0,0.0,0.041666668,0.31250003,0.23333335,0.19166668,0.15000002,0.43333334,0.22500001,0.31666666,0.01875,0.0,0.0,0.0,0.0,0.0625,0.38333336,0.7875,0.90833336,1.05,1.2,0.625,0.70624995,0.7416667,0.35625,0.8166667,3.0,6.408334,7.5166664,12.418751,15.5,17.800001,20.258331,23.3,28.916664,27.33125,21.508331,20.425,21.181252,18.8,18.80625,20.224998,21.487501,22.283335,26.883335,24.018753,22.966667,17.9,5.633333,1.13125,0.75,0.93333334,0.9562501,0.6666667,0.34375003,0.06666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.075,0.075,0.0,0.1375,0.074999996,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.22500001,0.80833334,1.6666669,2.1312501,1.3416667,0.88125,0.69166666,0.475,0.14166667,0.09166667,0.43125,1.4000001,0.94375,0.26666668,0.28125,1.7666668,1.6000001,2.9750001,3.4583335,1.5500001,1.4916668,3.0687494,3.908333,4.625,5.2749996,7.7249994,11.6875,13.066668,8.575,6.191667,6.6625004,8.508334,3.2062502,0.24166669,0.21666667,0.61875,1.05,0.9812499,0.5333333,0.0625,0.06666667,0.375,0.50625,0.35,0.7874999,1.7750001,1.5374999,0.50000006,0.6500001,1.3562502,1.8500004,1.85625,3.2583332,4.51875,3.75,1.5187501,0.7750001,0.95833325,1.10625,0.46666667,0.60625005,1.3583333,2.875,3.6833334,1.875,0.7875,0.45000005,0.39375004,1.0583334,1.7499999,2.5583334,5.90625,10.1,10.191667,10.806251,10.866666,11.556251,8.500001,3.75625,1.0416666,0.24166667,0.15625001,0.050000004,0.0,0.12500001,0.63125,0.9583334,2.5083332,4.9187503,5.0333333,5.3999996,4.1,1.1500001,0.69166666,1.0625,1.7083334,4.0083337,4.8250003,6.9083333,6.38125,8.866667,8.04375,6.1749997,4.183334,1.1375,1.9916666,3.3062503,2.9583335,1.0125,0.28333333,0.30624998,0.25833333,0.033333335,0.0,0.0,0.0,0.0,0.0,0.0,0.025,0.25625002,0.94166666,3.2499998,4.2083335,12.10625,18.933334,19.362501,17.291668,15.041666,9.35625,4.6583333,2.3375,3.5166667,4.61875,2.8749998,1.4416666,1.8125,0.9083333,0.23125,0.0,0.0,0.0,0.0,0.375,0.1,1.025,2.9416666,4.2875004,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0;
 } 
