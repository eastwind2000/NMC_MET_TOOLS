netcdf QPE_CPC_CMORPH.2018072700{
dimensions: 
 lat = 180; 
 lon = 281; 
variables:  
float lat(lat) ; 
   lat:long_name = "latitude" ;
   lat:units = "degrees_north" ;
   lat:standard_name = "latitude" ;
float lon(lon) ;
   lon:long_name = "longitude" ;
   lon:units = "degrees_east" ;
   lon:standard_name = "longitude" ;
float APCP_24(lat, lon) ;
   APCP_24:name = "APCP_24" ;
   APCP_24:long_name = "Total Precipitation" ;
   APCP_24:level = "A24" ;
   APCP_24:units = "kg/m^2" ;
   APCP_24:_FillValue = -9999.f ;
   APCP_24:init_time = "20180726_000000" ;
   APCP_24:init_time_ut = "1532563200.0" ;
   APCP_24:valid_time = "20180727_000000" ;
   APCP_24:valid_time_ut = "1532649600.0" ;
   APCP_24:accum_time = "240000" ;
   APCP_24:_FillValue = -9.99e8 ;
   APCP_24:accum_time_sec = 86400 ;
 // global attributes: 
 :_NCProperties = "version=1|netcdflibversion=4.4.1.1|hdf5libversion=1.8.12" ;
	:FileOrigins = "CPC_CMORPH_DAILY_PRCP" ; 
	:MET_version = "V7.0" ;
	:Projection = "LatLon" ;
	:lat_ll = "15.125 degrees_north" ; 
	:lon_ll = "70.125 degrees_east" ; 
	:delta_lat = "0.250000 degrees" ;
	:delta_lon = "0.250000 degrees" ;
	:Nlat = "180 grid_points" ; 
	:Nlon = "281 grid_points" ; 
data:
lat = 15.125,15.375,15.625,15.875,16.125,16.375,16.625,16.875,17.125,17.375,17.625,17.875,18.125,18.375,18.625,18.875,19.125,19.375,19.625,19.875,20.125,20.375,20.625,20.875,21.125,21.375,21.625,21.875,22.125,22.375,22.625,22.875,23.125,23.375,23.625,23.875,24.125,24.375,24.625,24.875,25.125,25.375,25.625,25.875,26.125,26.375,26.625,26.875,27.125,27.375,27.625,27.875,28.125,28.375,28.625,28.875,29.125,29.375,29.625,29.875,30.125,30.375,30.625,30.875,31.125,31.375,31.625,31.875,32.125,32.375,32.625,32.875,33.125,33.375,33.625,33.875,34.125,34.375,34.625,34.875,35.125,35.375,35.625,35.875,36.125,36.375,36.625,36.875,37.125,37.375,37.625,37.875,38.125,38.375,38.625,38.875,39.125,39.375,39.625,39.875,40.125,40.375,40.625,40.875,41.125,41.375,41.625,41.875,42.125,42.375,42.625,42.875,43.125,43.375,43.625,43.875,44.125,44.375,44.625,44.875,45.125,45.375,45.625,45.875,46.125,46.375,46.625,46.875,47.125,47.375,47.625,47.875,48.125,48.375,48.625,48.875,49.125,49.375,49.625,49.875,50.125,50.375,50.625,50.875,51.125,51.375,51.625,51.875,52.125,52.375,52.625,52.875,53.125,53.375,53.625,53.875,54.125,54.375,54.625,54.875,55.125,55.375,55.625,55.875,56.125,56.375,56.625,56.875,57.125,57.375,57.625,57.875,58.125,58.375,58.625,58.875,59.125,59.375,59.625,59.875;
lon = 70.125,70.375,70.625,70.875,71.125,71.375,71.625,71.875,72.125,72.375,72.625,72.875,73.125,73.375,73.625,73.875,74.125,74.375,74.625,74.875,75.125,75.375,75.625,75.875,76.125,76.375,76.625,76.875,77.125,77.375,77.625,77.875,78.125,78.375,78.625,78.875,79.125,79.375,79.625,79.875,80.125,80.375,80.625,80.875,81.125,81.375,81.625,81.875,82.125,82.375,82.625,82.875,83.125,83.375,83.625,83.875,84.125,84.375,84.625,84.875,85.125,85.375,85.625,85.875,86.125,86.375,86.625,86.875,87.125,87.375,87.625,87.875,88.125,88.375,88.625,88.875,89.125,89.375,89.625,89.875,90.125,90.375,90.625,90.875,91.125,91.375,91.625,91.875,92.125,92.375,92.625,92.875,93.125,93.375,93.625,93.875,94.125,94.375,94.625,94.875,95.125,95.375,95.625,95.875,96.125,96.375,96.625,96.875,97.125,97.375,97.625,97.875,98.125,98.375,98.625,98.875,99.125,99.375,99.625,99.875,100.125,100.375,100.625,100.875,101.125,101.375,101.625,101.875,102.125,102.375,102.625,102.875,103.125,103.375,103.625,103.875,104.125,104.375,104.625,104.875,105.125,105.375,105.625,105.875,106.125,106.375,106.625,106.875,107.125,107.375,107.625,107.875,108.125,108.375,108.625,108.875,109.125,109.375,109.625,109.875,110.125,110.375,110.625,110.875,111.125,111.375,111.625,111.875,112.125,112.375,112.625,112.875,113.125,113.375,113.625,113.875,114.125,114.375,114.625,114.875,115.125,115.375,115.625,115.875,116.125,116.375,116.625,116.875,117.125,117.375,117.625,117.875,118.125,118.375,118.625,118.875,119.125,119.375,119.625,119.875,120.125,120.375,120.625,120.875,121.125,121.375,121.625,121.875,122.125,122.375,122.625,122.875,123.125,123.375,123.625,123.875,124.125,124.375,124.625,124.875,125.125,125.375,125.625,125.875,126.125,126.375,126.625,126.875,127.125,127.375,127.625,127.875,128.125,128.375,128.625,128.875,129.125,129.375,129.625,129.875,130.125,130.375,130.625,130.875,131.125,131.375,131.625,131.875,132.125,132.375,132.625,132.875,133.125,133.375,133.625,133.875,134.125,134.375,134.625,134.875,135.125,135.375,135.625,135.875,136.125,136.375,136.625,136.875,137.125,137.375,137.625,137.875,138.125,138.375,138.625,138.875,139.125,139.375,139.625,139.875,140.125;
APCP_24 = 0.32999998,0.28,0.53999996,1.15,1.11,1.42,0.84,0.16,0.01,0.0,0.0,0.01,0.099999994,0.26,1.27,0.14999999,0.08,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02,0.25,0.69,1.1899999,1.4399999,1.36,1.23,1.05,0.87,0.48,0.26999998,0.19999999,0.08,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.099999994,0.39999998,0.11,0.03,0.0,0.0,0.07,0.06,1.26,3.1599998,5.85,14.66,26.47,34.82,44.2,36.46,25.71,23.97,15.299999,10.889999,7.69,3.05,1.1899999,1.86,2.02,0.77,0.24,0.97999996,0.95,0.16,0.7,2.25,3.04,0.85999995,0.32999998,0.62,0.93,0.84999996,1.74,8.46,8.53,10.01,3.99,8.17,33.25,3.11,4.06,5.73,12.2,15.849999,12.09,14.34,10.76,12.69,10.08,10.929999,17.4,11.79,1.35,0.01,0.0,0.0,0.76,0.52,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.5,6.3999996,9.0,9.26,13.63,11.71,13.679999,14.179999,10.84,19.359999,20.93,14.49,4.64,4.71,7.5499997,11.4,19.73,31.769999,33.2,8.389999,0.0,0.0,0.0,0.0,0.93,1.4499999,6.08,1.54,0.39,0.53999996,0.0,0.0,0.0,0.0,0.0,0.26,1.5999999,4.15,7.8999996,2.59,1.49,0.0,0.71999997,1.9599999,2.04,1.3299999,0.44,0.0,0.0,0.0,0.0,0.0,0.14999999,0.39,0.59999996,0.64,0.65,0.63,0.52,0.90999997,2.95,4.23,4.5499997,1.78,0.13,0.0,0.0,1.4,4.45,2.33,0.08,1.11,1.7199999,5.3199997,3.46,0.71999997,0.94,0.0,0.0,0.0,0.0,0.81,5.43,4.0,2.31,2.02,1.0799999,0.65999997,0.22,0.089999996,0.03,0.19999999,0.0,0.0,0.0,0.0,0.0,0.19,0.35999998,0.65,3.27,0.44,0.37,0.32999998,0.39999998,1.01,1.73,2.12,0.94,0.19,0.01,0.0,0.0,0.0,0.69,2.11,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06,0.48,1.04,1.5,1.75,1.8299999,1.18,0.65,0.25,0.22999999,0.29,0.14999999,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.0,0.02,0.14,0.19999999,0.03,0.03,0.13,0.08,0.13,0.96999997,3.06,13.2699995,30.599998,45.809998,59.719997,43.809998,22.81,22.93,14.15,6.0299997,4.16,2.62,1.1899999,1.4599999,1.91,1.3399999,0.63,0.65,1.24,1.11,1.66,2.09,1.5899999,3.05,2.2,1.6899999,0.41,1.28,1.5899999,5.99,10.01,7.48,5.16,7.02,20.18,5.68,4.08,4.7799997,13.059999,12.73,13.139999,13.96,14.5,12.09,6.6499996,9.91,11.2699995,5.41,0.0,0.0,0.0,0.0,0.08,8.15,2.05,1.99,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.39999998,3.6,1.81,1.37,3.32,5.15,9.429999,14.48,11.4,8.03,11.34,6.02,3.56,2.11,2.58,1.79,3.09,10.62,20.64,36.57,46.6,31.929998,10.87,0.75,0.0,0.0,0.0,0.0,0.37,1.9599999,0.32,0.089999996,0.14999999,0.0,0.0,0.0,0.0,0.72999996,1.9499999,3.57,21.82,17.8,0.55,1.11,0.089999996,0.53,0.93,0.96999997,0.32999998,0.0,0.0,0.0,0.0,0.0,0.0,0.16,0.57,0.61,0.24,0.11,0.099999994,0.17,1.4399999,3.04,5.97,3.46,0.66999996,0.0,0.0,0.0,1.7099999,3.26,1.61,1.23,2.0,1.89,7.95,4.37,1.41,1.5799999,2.9199998,3.1799998,1.49,0.0,0.22999999,2.12,0.93,0.45,0.5,0.16,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.16,2.6,0.19,0.63,3.9199998,5.21,0.68,0.38,0.19,0.04,0.22,0.89,1.63,1.8299999,1.99,0.97999996,0.17,0.07,0.089999996,1.11,1.49,0.0,0.0,0.0,0.0,0.04,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.11,0.04,0.0,0.0,0.0,0.0,0.0,0.13,0.51,1.04,1.43,1.29,0.9,0.57,0.26,0.17999999,0.11,0.04,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.049999997,0.11,0.47,1.54,1.24,2.4099998,5.0899997,0.77,0.22999999,0.90999997,1.2099999,0.59999996,0.84,2.49,10.91,28.189999,45.43,61.53,38.44,17.85,17.92,11.83,2.99,1.79,2.23,1.79,1.41,1.3299999,1.6899999,1.23,1.05,0.87,2.23,3.29,3.8,5.1,3.9599998,2.56,2.6599998,1.0699999,3.29,3.52,7.58,14.059999,8.05,7.81,9.4,15.559999,9.5,6.96,7.0,10.8,12.55,15.849999,12.509999,13.28,11.87,5.25,4.38,5.43,0.17999999,0.0,0.0,0.0,0.0,0.08,18.05,10.2699995,10.32,1.8299999,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.53999996,1.3199999,0.59999996,0.26999998,1.01,3.79,9.7699995,17.55,16.68,7.2,7.5899997,7.1,1.51,1.26,1.43,1.0799999,2.4299998,7.08,25.65,41.7,51.87,13.389999,4.58,1.3299999,1.78,0.0,0.0,5.41,3.83,0.93,3.62,4.56,0.0,0.0,0.0,0.0,0.03,0.35,1.8,6.1099997,13.719999,6.43,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.93,2.45,2.3999999,2.53,2.95,0.52,0.02,0.14999999,0.90999997,1.5,0.9,8.7,8.11,1.8499999,3.6699998,7.0,5.24,2.87,4.97,14.07,13.46,4.7,0.66999996,0.17999999,0.42999998,0.099999994,0.02,0.0,0.0,0.0,0.11,0.02,0.0,0.0,0.0,0.0,0.0,1.39,2.6399999,2.3799999,3.3,6.83,9.33,0.31,0.48,0.39,0.14,0.11,0.53,1.0699999,1.74,2.72,2.69,2.22,1.26,0.65,0.42999998,0.51,0.0,0.0,0.0,0.0,0.049999997,0.13,0.17,0.17999999,0.099999994,0.089999996,0.01,0.01,0.0,0.0,0.0,0.06,0.13,0.22999999,0.31,0.22999999,0.26999998,0.39,0.099999994,0.0,0.0,0.0,0.0,0.0,0.0,0.02,0.21,0.16,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.099999994,0.08,0.13,0.13,0.099999994,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.19,0.08,0.39999998,2.56,5.0,2.3,7.47,4.0299997,1.9,1.18,2.33,2.98,3.3999999,7.1299996,15.089999,25.23,45.76,49.16,29.06,17.64,15.91,12.69,3.85,1.53,1.0699999,1.39,2.08,1.73,3.4199998,2.1399999,1.88,1.39,1.9699999,6.35,5.38,9.21,6.98,4.0,4.11,4.0,6.3999996,8.21,12.559999,18.08,12.08,11.41,14.719999,17.51,16.26,10.0199995,10.82,14.32,12.92,16.01,10.54,13.07,10.12,5.7,2.18,0.69,0.26999998,0.19999999,0.0,0.0,0.06,0.44,5.42,6.98,7.37,2.33,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.45,5.02,8.889999,6.15,2.03,1.16,3.3,1.41,3.3999999,1.39,0.39999998,0.29,1.8399999,15.969999,32.48,22.98,6.73,8.3,20.47,31.41,14.5,27.96,2.23,0.11,1.74,5.69,6.0,0.0,0.0,0.0,0.0,0.0,0.0,0.26,1.8499999,2.03,0.39999998,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.45999998,0.35,0.0,0.0,0.0,0.0,0.0,0.34,0.72999996,0.32999998,2.75,4.0899997,0.53,0.07,0.29999998,0.9,0.71,0.82,1.9,2.08,3.62,5.79,4.96,6.21,2.49,2.9199998,10.86,9.57,1.1,0.0,0.14999999,0.71,0.06,0.0,0.0,0.0,0.0,0.0,0.02,0.29999998,0.58,1.48,0.53,0.049999997,0.64,0.58,0.65999997,2.47,4.58,6.97,0.25,0.099999994,0.71999997,1.02,0.45999998,0.45,0.52,1.01,1.9799999,2.53,3.37,2.79,2.95,1.17,0.42,0.11,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.01,0.0,0.0,0.0,0.02,0.04,0.049999997,0.07,0.19999999,0.38,0.29999998,0.45999998,0.48999998,0.19,0.12,0.089999996,0.049999997,0.049999997,0.0,0.06,0.08,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06,0.08,0.11,0.28,0.29,0.78999996,2.4099998,3.09,1.7199999,1.63,0.35999998,0.24,2.61,5.67,7.6499996,11.19,18.4,26.13,43.149998,43.67,31.88,22.789999,17.039999,16.07,4.7,1.6899999,0.84999996,0.71999997,2.06,2.03,4.02,3.1599998,2.76,2.22,2.52,4.89,7.5699997,9.28,6.71,5.7999997,5.99,9.3,12.42,13.13,16.4,19.43,18.16,18.13,24.789999,32.57,27.31,24.16,22.529999,23.119999,17.65,19.109999,9.91,9.03,10.45,9.21,4.63,2.56,1.64,1.3,1.12,2.55,1.16,1.27,1.56,4.36,5.2,2.74,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08,0.56,0.82,1.35,0.29999998,1.02,1.4399999,1.28,0.71,0.48999998,1.09,5.0499997,1.79,0.0,0.099999994,0.61,2.32,3.28,2.85,4.85,8.76,36.41,55.489998,24.55,23.35,16.67,7.99,0.87,1.5699999,1.29,0.12,0.22999999,0.0,0.0,0.0,0.22,0.0,0.0,0.0,0.0,0.28,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,3.1499999,4.2,3.1799998,0.89,1.3199999,0.0,0.7,1.5899999,2.8,4.16,4.79,4.45,4.3399997,0.96,0.08,0.0,0.79999995,0.29999998,0.22999999,0.87,0.64,3.1799998,3.99,5.06,2.1599998,1.22,0.79999995,0.11,0.0,0.0,0.0,0.13,1.39,1.8299999,2.8799999,2.61,1.29,0.45,0.0,0.19999999,1.53,2.99,5.42,1.18,0.0,0.16,0.35999998,1.09,3.99,8.29,15.7699995,0.9,1.5699999,2.61,2.56,1.9799999,1.89,1.51,0.94,1.41,2.2,4.13,4.4,3.99,1.3199999,0.9,0.55,0.32,0.19,0.16,0.16,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.099999994,0.089999996,0.02,0.0,0.0,0.0,0.0,0.04,0.14,0.32999998,0.19,0.19999999,0.14999999,0.14,0.14,0.17,0.19,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.34,0.37,0.32,0.39,0.42,0.53,1.54,2.6799998,2.51,1.01,0.35,3.37,9.09,13.61,16.039999,21.359999,35.32,44.16,40.98,35.59,24.01,21.199999,16.26,8.639999,1.9,1.06,1.22,1.3199999,1.49,1.15,2.72,3.23,3.6799998,2.3999999,1.8499999,2.84,6.7599998,5.0899997,5.2999997,6.97,13.179999,17.39,15.45,18.66,20.189999,22.82,27.74,36.399998,49.309998,56.199997,49.73,51.36,34.8,21.189999,19.22,10.0,4.41,13.65,14.32,6.5499997,5.23,5.5899997,2.4099998,1.8199999,2.11,3.21,1.68,0.48999998,0.59999996,0.22,0.14,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.59,0.28,0.77,0.71,0.42,0.0,0.13,0.96999997,0.96999997,0.53999996,0.01,0.0,1.3,1.1,0.0,0.0,0.0,0.049999997,0.0,0.0,0.72999996,5.43,27.05,38.98,22.949999,2.25,16.15,4.21,0.0,4.22,0.0,0.42,11.7699995,1.6999999,0.0,0.0,0.0,0.0,0.0,0.0,0.44,0.37,0.17,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,3.1499999,4.2,8.75,10.4,6.47,4.87,4.2,4.2,4.24,4.89,4.14,4.5899997,4.2799997,1.91,1.05,0.62,1.3199999,1.86,0.71,0.08,1.0799999,4.5299997,3.52,0.55,0.0,0.21,0.17999999,0.0,0.0,0.0,0.01,0.52,2.51,5.21,7.98,10.34,6.49,1.99,0.089999996,0.83,2.49,5.73,7.98,3.8999999,0.98999995,0.0,0.0,0.44,3.8999999,11.36,27.16,2.62,3.4299998,4.79,5.1,5.35,5.02,4.97,3.8999999,3.6699998,3.7099998,3.79,3.6499999,2.97,1.16,0.81,0.57,0.35,0.17999999,0.21,0.22,0.14,0.06,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.049999997,0.42,0.37,0.39,0.32999998,0.22,0.04,0.0,0.0,0.0,0.03,0.089999996,0.06,0.01,0.02,0.02,0.0,0.049999997,0.17999999,0.25,0.19,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14,0.58,1.29,1.8499999,1.43,1.75,1.3299999,1.75,2.81,2.54,1.12,4.13,11.92,22.91,27.23,31.789999,42.95,54.719997,48.21,43.61,31.769999,26.72,21.869999,14.53,6.04,1.92,2.11,2.34,1.1999999,1.0699999,1.39,2.4299998,4.65,4.33,2.46,2.97,3.79,3.75,2.4299998,5.2,15.059999,15.78,13.179999,20.609999,24.59,32.489998,36.989998,38.66,58.32,79.86,62.64,66.439995,49.28,29.41,22.26,10.0,3.99,11.67,13.66,4.13,11.809999,13.28,4.21,2.9399998,3.3999999,4.31,1.9599999,0.08,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14999999,1.36,0.39999998,0.0,0.0,0.0,0.0,0.0,0.0,0.06,0.19999999,0.0,3.1799998,0.61,0.34,0.35,0.28,0.0,0.0,0.04,0.03,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,5.5899997,15.839999,24.25,17.91,6.77,7.1,0.72999996,0.0,1.8299999,1.7199999,0.13,3.9299998,4.1,0.42,0.28,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.26999998,2.1,8.47,14.5199995,12.98,6.98,6.7599998,5.06,5.5899997,6.5499997,7.41,6.8399997,7.1299996,6.29,7.6699996,9.67,9.349999,6.06,2.78,0.0,0.25,1.92,2.59,0.0,0.049999997,0.25,0.29999998,0.19,0.0,0.0,0.0,0.02,0.63,1.61,2.1299999,4.19,7.73,4.99,0.29999998,0.35999998,2.2,4.13,9.349999,5.42,0.75,0.0,0.08,0.71999997,2.69,10.7,25.269999,3.4499998,5.06,6.0299997,6.35,5.79,6.1099997,6.54,6.35,6.42,6.2599998,4.75,3.6799998,2.22,0.90999997,0.85999995,0.53999996,0.38,0.22,0.06,0.11,0.11,0.14999999,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14999999,0.61,0.45999998,0.29,0.34,0.26,0.04,0.0,0.0,0.06,0.14999999,0.12,0.03,0.04,0.089999996,0.08,0.03,0.0,0.0,0.03,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.099999994,0.9,1.8199999,3.4399998,5.04,4.0299997,3.1299999,2.0,2.9199998,3.74,3.37,5.7999997,14.19,31.13,39.82,47.039997,53.05,58.75,59.219997,54.84,43.77,32.85,26.59,17.47,10.0199995,3.3899999,2.56,3.23,2.03,1.36,1.37,1.62,2.57,4.42,1.75,4.12,4.71,4.58,1.38,3.22,12.87,11.12,11.66,20.789999,27.859999,38.95,39.2,34.98,48.78,76.63,61.129997,59.92,48.21,29.369999,20.63,10.12,4.8599997,7.52,10.92,3.58,5.2599998,12.62,8.5,5.62,7.66,7.83,3.48,0.13,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02,1.3399999,0.42999998,0.0,0.0,0.0,0.0,0.0,0.0,0.32999998,0.71999997,0.0,5.74,0.94,0.06,1.0,0.25,0.0,0.049999997,0.04,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13,2.75,9.62,14.21,4.74,6.18,3.24,1.05,0.0,0.0,0.0,0.0,1.28,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.71,9.12,11.49,6.74,5.67,7.71,8.33,9.37,10.2,9.36,8.19,10.09,11.7699995,16.67,20.22,21.76,14.96,0.32999998,0.0,0.0,0.0,0.0,0.17,0.45,0.5,0.32999998,0.0,0.0,0.0,0.0,0.02,0.42,0.0,0.0,0.32999998,1.73,0.66999996,0.97999996,0.90999997,0.45999998,0.06,0.0,0.0,0.0,0.06,0.61,2.03,4.36,10.03,3.98,4.75,5.8199997,6.81,6.83,6.96,6.5299997,6.89,7.25,7.3199997,5.8199997,3.27,1.65,0.98999995,0.69,0.61,0.63,0.65,0.34,0.03,0.03,0.049999997,0.04,0.06,0.07,0.0,0.06,0.049999997,0.0,0.0,0.0,0.0,0.13,0.26999998,0.32999998,0.14,0.04,0.0,0.0,0.01,0.17999999,0.31,0.58,0.55,0.16,0.04,0.11,0.17999999,0.07,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.11,0.29,1.43,3.4299998,6.97,9.75,9.84,7.2799997,5.8799996,4.39,4.2599998,7.69,16.98,41.44,55.86,58.55,68.38,74.369995,55.77,54.949997,31.22,24.66,18.46,13.99,9.08,3.9199998,1.48,1.6899999,1.6999999,1.35,1.5799999,2.28,4.37,2.58,1.74,1.7199999,3.47,2.85,2.07,1.68,8.4,8.4,9.42,16.14,25.1,34.11,36.96,31.22,37.05,51.969997,38.19,37.6,28.97,21.439999,12.94,8.28,4.36,5.3199997,7.0099998,4.88,9.139999,23.81,28.17,14.09,15.28,16.119999,9.29,0.88,0.13,0.03,0.0,0.11,0.099999994,0.04,0.0,0.0,0.03,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.29,0.55,0.0,3.83,0.48999998,0.16,0.14999999,0.0,0.0,0.01,0.03,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.22,0.59999996,0.95,16.529999,30.539999,13.219999,39.05,14.589999,0.21,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.04,0.39999998,4.37,6.49,4.39,3.49,4.44,5.3399997,5.7,10.5,7.94,11.69,13.34,18.56,23.539999,37.21,41.079998,36.62,2.33,0.01,0.0,0.0,0.0,0.049999997,0.19,0.17,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.3,3.85,1.5999999,0.12,0.049999997,0.099999994,0.049999997,0.02,0.25,0.7,1.43,3.72,3.6999998,4.3399997,4.5,5.3199997,6.1099997,7.43,8.41,7.7999997,7.23,7.14,6.74,3.9599998,1.66,1.09,0.66999996,0.32999998,0.21,0.08,0.0,0.099999994,0.19999999,0.089999996,0.04,0.0,0.32999998,0.19999999,0.31,0.39,0.31,0.12,0.03,0.0,0.0,0.0,0.0,0.14999999,0.26,0.16,0.089999996,0.02,0.22,0.82,1.29,1.9799999,1.77,0.47,0.08,0.04,0.17999999,0.19,0.08,0.06,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13,0.39999998,1.1899999,4.52,9.16,17.59,20.22,13.33,6.54,5.38,5.7,16.59,45.649998,63.719997,71.4,71.72,68.65,44.809998,39.629997,23.39,13.78,10.88,8.57,6.93,4.48,2.3899999,1.92,1.8399999,4.37,4.45,2.7,3.98,4.46,2.9399998,1.7199999,4.3199997,5.47,3.85,2.1699998,6.7999997,6.8799996,9.63,14.75,18.96,25.68,31.619999,34.66,37.23,31.22,21.34,17.72,10.849999,10.46,7.08,3.85,2.6699998,4.2799997,4.5099998,5.79,12.0,19.189999,32.309998,25.14,35.57,29.67,11.46,1.3,0.48,0.9,0.17999999,0.42,0.71,0.31,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.04,0.71999997,0.37,1.3399999,0.16,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.55,1.61,0.93,1.35,5.25,35.86,60.94,15.58,67.95,33.61,6.04,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.26999998,0.0,0.089999996,0.63,1.36,3.98,6.91,1.12,0.44,2.6299999,3.6599998,5.0299997,5.67,7.3399997,14.58,19.77,26.289999,29.51,34.09,37.28,31.279999,9.21,5.0,1.14,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.17,0.11,0.01,0.099999994,0.19999999,0.13,0.0,0.0,0.39,4.0099998,2.8799999,2.35,4.02,3.8,4.29,5.52,6.15,7.7599998,8.16,7.14,6.89,6.8199997,5.1,1.64,0.89,0.65,0.39999998,0.21,0.04,0.0,0.01,0.06,0.13,0.13,0.04,0.19999999,0.62,0.51,0.22999999,0.17,0.12,0.0,0.0,0.0,0.0,0.0,0.0,0.02,0.17,0.089999996,0.0,0.02,0.26,1.0,2.6699998,3.26,1.9399999,1.64,0.65999997,0.06,0.11,0.29,0.25,0.099999994,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02,0.07,0.08,0.35999998,0.78,3.9199998,11.37,26.019999,30.34,22.24,8.37,3.6799998,3.61,10.91,37.36,63.02,68.08,73.95,72.68,48.35,29.929998,20.39,11.45,6.8599997,5.62,5.23,4.37,3.8999999,6.73,4.77,7.5899997,13.099999,4.94,1.37,3.85,4.64,3.97,4.98,8.88,7.0,4.66,7.68,9.309999,12.79,19.64,20.43,21.38,22.619999,25.82,29.13,21.41,14.63,10.929999,5.6299996,4.72,4.7599998,2.81,2.45,3.4199998,4.2999997,5.2799997,8.099999,15.73,13.78,31.33,55.75,43.1,49.59,89.56,29.8,2.96,1.29,1.09,1.9799999,1.1,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02,0.0,0.42,0.47,0.29999998,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,3.82,4.19,3.26,4.08,20.46,34.239998,57.61,12.7,17.949999,8.97,4.0699997,0.0,0.32999998,0.45999998,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.19999999,0.24,0.0,0.0,0.17,0.28,0.0,0.61,1.0699999,0.0,0.0,0.19999999,0.59,4.08,7.1499996,0.19,0.089999996,2.84,3.33,2.22,2.3999999,5.0499997,5.24,11.2,16.08,17.82,14.08,12.57,18.38,12.11,8.33,5.0899997,3.54,0.63,0.22,0.099999994,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02,0.19999999,1.06,0.16,0.55,1.53,2.69,8.41,0.78,0.96,2.62,3.32,4.11,4.92,5.42,6.7599998,6.45,6.3599997,6.46,6.19,2.6799998,1.5699999,0.69,0.45,0.28,0.12,0.03,0.0,0.0,0.0,0.0,0.06,0.11,0.0,0.0,0.0,0.07,0.22,0.14999999,0.16,0.049999997,0.01,0.0,0.0,0.0,0.0,0.0,0.02,0.02,0.0,0.0,0.06,0.65999997,1.52,0.41,0.53,1.06,0.55,0.04,0.0,0.099999994,0.049999997,0.0,0.02,0.01,0.03,0.0,0.0,0.0,0.01,0.07,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.04,0.04,0.11,0.17,0.45,0.45,1.3399999,6.5099998,17.34,32.68,35.77,32.079998,16.58,4.5899997,1.03,7.12,19.13,47.44,54.199997,52.01,56.239998,49.39,29.32,16.97,12.21,5.7,3.34,2.77,3.31,3.24,5.3599997,5.69,4.65,8.99,6.8599997,1.18,1.24,3.03,5.12,6.0099998,10.57,13.099999,8.66,7.49,9.3,13.5199995,16.15,20.59,19.359999,15.9,18.88,21.88,19.189999,12.61,7.35,3.27,1.3399999,1.68,1.5,1.79,2.53,3.05,4.18,4.89,7.8799996,9.09,29.449999,63.809998,82.7,129.34,76.58,20.99,2.24,1.06,3.6899998,5.08,2.52,0.07,0.0,0.0,0.0,0.0,0.0,0.0,0.53999996,1.8,0.58,0.47,0.0,0.06,0.04,0.0,0.0,0.0,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.98999995,4.3399997,6.29,2.6399999,15.23,59.579998,32.45,7.2599998,0.69,1.13,2.33,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.089999996,1.23,2.3,2.24,0.90999997,0.72999996,0.16,0.71999997,1.55,1.28,1.4,1.4,0.13,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.21,0.03,0.14999999,0.35,1.9499999,1.75,1.7199999,1.15,1.9,2.4299998,8.16,12.889999,8.929999,8.04,9.099999,5.77,2.36,0.78,0.22999999,0.35,0.04,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.24,2.97,6.7599998,19.31,14.38,3.06,5.0299997,1.2099999,0.66999996,2.09,3.03,2.8799999,2.9399998,3.6699998,4.5,5.2799997,5.2999997,5.5099998,6.3399997,2.8799999,0.95,0.53,0.28,0.11,0.03,0.0,0.0,0.0,0.0,0.02,0.08,0.17999999,0.26999998,0.16,0.08,0.0,0.0,0.0,0.0,0.04,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02,0.0,0.0,0.0,0.0,0.08,0.06,0.11,0.02,0.0,0.0,0.0,0.02,0.04,0.02,0.0,0.14,0.25,0.21,0.06,0.0,0.0,0.0,0.0,0.03,0.07,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07,0.34,0.48,0.63,0.59999996,0.90999997,1.11,3.4199998,11.09,26.199999,32.17,34.809998,29.06,18.23,5.44,0.87,2.09,7.2999997,18.32,33.96,35.559998,42.96,40.989998,25.779999,11.61,7.45,4.85,2.12,0.87,0.83,1.23,1.18,2.25,6.35,7.95,4.48,1.88,1.0799999,3.86,7.6299996,10.4,10.16,17.789999,16.85,12.73,11.65,11.429999,13.759999,17.42,18.529999,12.0,10.0,15.82,16.869999,11.8,5.06,1.81,0.71999997,0.38,0.11,0.21,1.26,1.3399999,2.62,3.3,3.05,4.96,37.57,72.619995,101.77,56.149998,23.279999,7.6,1.0799999,0.89,5.92,9.469999,5.04,0.68,0.22999999,0.0,0.0,0.0,0.0,0.06,1.6999999,3.51,2.03,2.44,0.07,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02,0.29,1.4499999,4.89,8.33,2.87,2.74,37.13,30.64,1.4699999,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.35,3.34,1.91,0.17,0.72999996,1.3299999,0.59999996,0.35999998,0.79999995,1.0799999,0.68,0.79999995,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.16,0.12,0.089999996,0.07,0.04,0.089999996,0.75,3.0,9.099999,11.66,5.2599998,8.3,2.59,1.8,1.8,1.06,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.06,5.48,0.48999998,2.47,4.14,10.05,14.799999,18.8,11.12,0.59,1.6899999,2.32,2.8999999,2.6799998,3.54,4.5299997,5.06,5.0899997,4.38,3.57,2.22,0.94,0.52,0.32999998,0.099999994,0.03,0.28,0.099999994,0.0,0.0,0.0,0.0,0.01,0.089999996,0.24,0.03,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02,0.0,0.0,0.0,0.0,0.04,0.099999994,0.089999996,0.03,0.01,0.049999997,0.08,0.049999997,0.03,0.04,0.04,0.02,0.0,0.0,0.0,0.03,0.04,0.13,0.26,0.45999998,0.45999998,0.35,0.089999996,0.02,0.07,0.14,0.22999999,0.25,0.17,0.03,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.11,0.14,0.42,1.39,2.08,2.72,3.1899998,3.62,3.08,6.8799996,16.16,30.83,31.07,34.809998,24.13,12.0,6.81,4.0299997,5.1,5.2799997,9.7,21.369999,25.269999,22.529999,23.369999,18.17,8.79,3.09,1.7199999,0.72999996,0.58,0.53,0.16,0.65999997,0.71999997,2.81,8.88,7.14,3.6599998,3.6799998,7.3199997,11.849999,13.54,16.94,17.49,23.82,22.779999,18.31,14.2,13.19,16.82,18.029999,15.639999,9.29,7.5099998,9.48,7.7799997,3.7099998,0.96,0.32999998,0.39999998,0.41,0.01,0.099999994,0.5,1.5,2.09,0.56,1.4,27.89,31.23,54.489998,21.359999,15.7699995,4.5299997,0.56,1.09,9.84,16.57,11.809999,2.3899999,0.57,0.0,0.0,0.0,0.0,0.64,2.46,2.24,5.21,4.77,0.41,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02,0.03,0.0,0.0,0.0,0.0,0.0,0.01,0.52,0.82,2.6599998,3.54,1.53,0.0,1.8499999,2.2,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.02,2.9199998,1.91,0.44,0.0,0.0,0.13,0.0,0.03,0.03,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13,0.56,0.75,0.66999996,0.22,0.17,0.44,0.5,0.14999999,0.59999996,0.59999996,0.45999998,1.1999999,0.9,1.06,2.05,1.06,0.12,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.39999998,1.5,5.52,7.77,18.14,1.0699999,1.6899999,1.91,2.8,3.9499998,4.24,4.45,4.95,5.73,5.64,2.75,0.75,0.12,0.07,0.089999996,0.03,0.02,0.099999994,0.03,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.12,0.16,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.14,0.13,0.0,0.0,0.0,0.049999997,0.099999994,0.11,0.11,0.13,0.06,0.11,0.089999996,0.08,0.03,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.12,0.42,0.72999996,0.71,0.79999995,0.53999996,0.41,0.32999998,0.42999998,0.59999996,0.7,0.59,0.19,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.02,0.01,0.01,0.04,0.58,0.94,1.48,3.3899999,5.8199997,7.0099998,8.63,10.0,10.95,6.7999997,9.969999,15.259999,24.359999,29.83,21.109999,10.78,9.5199995,13.0,12.91,10.07,7.48,10.38,14.889999,11.259999,7.98,7.22,5.37,3.08,1.3299999,0.55,0.53999996,1.41,1.16,0.049999997,0.78,1.03,1.56,2.46,2.26,5.79,8.179999,14.799999,18.289999,20.13,18.539999,20.6,27.539999,27.47,18.51,13.67,12.66,17.16,18.93,13.88,5.3399997,1.88,2.36,1.29,0.55,0.62,0.66999996,0.14999999,0.099999994,0.08,0.12,1.3399999,1.5799999,0.08,0.22,0.96999997,5.54,16.789999,11.53,4.43,1.28,0.26999998,1.68,6.8399997,13.84,13.13,3.32,0.79999995,0.82,0.29999998,0.0,0.0,0.90999997,4.25,2.74,10.7699995,5.94,0.58,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.099999994,0.26,0.0,0.0,0.0,0.02,0.0,0.0,0.03,0.04,0.0,0.0,0.24,0.39,0.53,0.31,0.17999999,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.27,0.66999996,0.0,0.0,0.0,0.0,0.0,0.0,0.08,0.08,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.5,0.71999997,0.39,0.089999996,0.0,0.0,0.049999997,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.06,1.41,0.16,0.0,0.0,0.14,0.08,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.4399999,4.0099998,12.139999,5.72,3.58,13.03,0.9,1.9799999,1.99,2.3799999,3.4499998,3.84,3.9299998,3.84,4.85,5.92,3.9299998,0.90999997,0.16,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02,0.12,0.13,0.07,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.16,0.17999999,0.0,0.0,0.06,0.089999996,0.17999999,0.29999998,0.26,0.16,0.099999994,0.049999997,0.0,0.099999994,0.049999997,0.03,0.0,0.0,0.0,0.0,0.0,0.02,0.099999994,0.47,0.74,1.4,2.31,2.6599998,2.36,1.4399999,1.1999999,1.25,1.26,1.18,0.74,0.21,0.02,0.0,0.0,0.0,0.0,0.089999996,0.21,0.31,0.85999995,0.90999997,2.85,3.3999999,6.44,11.98,14.03,16.01,19.529999,21.59,23.66,21.15,16.539999,13.88,20.48,20.89,20.25,14.34,12.96,15.179999,12.469999,6.92,4.42,6.87,6.29,4.45,2.78,3.55,3.31,2.28,1.49,1.48,1.79,3.1699998,2.02,1.5699999,1.36,1.56,2.76,2.85,6.24,9.98,11.429999,13.809999,15.61,19.41,16.529999,20.98,27.869999,24.63,16.529999,11.8,14.54,20.84,18.75,13.59,3.9499998,0.5,1.42,2.31,2.6399999,2.75,0.78999996,0.17,0.53999996,0.74,1.68,1.6999999,0.45,0.03,0.099999994,0.84,4.7799997,4.95,1.48,0.11,0.11,0.29999998,0.94,5.5099998,6.0299997,4.35,1.74,1.49,1.4699999,0.0,0.0,0.35,2.51,4.38,14.349999,5.3399997,0.48999998,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.049999997,0.04,0.0,0.0,0.04,0.049999997,0.0,0.0,0.0,0.0,0.14,0.89,1.9499999,1.09,0.32,0.04,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.04,0.089999996,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.049999997,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.78999996,2.26,12.2699995,16.789999,17.3,11.61,0.049999997,1.2099999,1.29,1.9,3.25,3.1899998,3.22,3.11,3.6899998,5.33,4.0899997,1.4499999,0.65,0.26999998,0.06,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.03,0.089999996,0.19,0.34,0.31,0.45999998,0.26999998,0.13,0.03,0.7,1.64,0.26999998,0.06,0.0,0.07,0.07,0.17999999,0.59999996,0.29,0.71,1.8399999,3.8799999,6.0699997,6.62,6.81,4.22,2.48,2.21,2.07,1.9599999,1.25,0.42,0.04,0.0,0.14,0.01,0.24,0.47,0.96,2.81,2.69,5.62,8.7,12.309999,18.0,22.34,24.699999,32.02,31.73,41.84,36.149998,21.529999,10.889999,10.83,14.88,16.0,18.029999,17.47,22.779999,22.74,12.69,5.43,1.0799999,2.36,2.3,2.04,2.6399999,3.4199998,3.4499998,3.1699998,3.36,3.52,4.3199997,6.1099997,6.45,4.62,1.8199999,2.6699998,3.9599998,6.3199997,11.599999,13.259999,14.63,12.5,13.21,18.119999,15.04,18.89,21.5,17.64,13.71,12.28,21.15,31.22,27.859999,12.45,2.04,3.59,8.36,9.059999,8.83,5.39,0.96,1.23,1.43,1.9,1.3299999,0.14999999,0.0,0.0,0.44,0.58,0.75,0.45,0.26,0.0,0.0,0.0,0.93,3.1599998,2.49,0.77,3.47,1.3199999,0.0,0.0,0.01,0.19,4.25,11.8,3.4199998,0.19999999,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06,0.59999996,1.3199999,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.02,0.049999997,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,5.8199997,10.87,17.1,7.58,0.0,0.03,0.44,0.94,2.19,2.81,2.76,2.87,3.03,3.1299999,2.8899999,1.28,0.64,0.39999998,0.32999998,0.24,0.0,0.0,0.0,0.0,0.0,0.0,0.099999994,0.13,0.089999996,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02,0.07,0.049999997,0.06,0.01,0.16,0.22999999,0.55,0.63,0.41,0.07,0.0,0.0,0.14,0.75,0.58,0.099999994,0.26999998,1.04,3.26,3.57,2.24,3.1599998,3.1699998,5.3599997,7.5499997,8.59,10.03,11.38,7.6699996,4.5,3.23,2.78,2.83,2.27,0.93,0.049999997,0.049999997,0.48,0.95,2.21,3.01,5.3199997,5.6099997,7.85,13.45,16.33,20.449999,27.47,33.34,44.629997,44.43,47.829998,46.329998,28.699999,17.23,5.79,8.51,10.969999,14.69,22.35,22.08,30.97,29.769999,16.359999,4.6,1.3399999,1.5999999,2.57,3.1999998,3.29,4.7599998,6.22,5.79,5.44,5.98,7.8199997,9.49,9.46,4.31,3.04,4.72,4.3399997,9.679999,13.87,14.34,14.049999,10.04,13.25,16.039999,12.23,14.599999,15.82,17.779999,13.73,16.529999,24.65,30.369999,26.57,5.66,3.8799999,12.66,15.759999,14.08,11.759999,4.18,0.71999997,1.5,1.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14999999,0.0,0.0,0.01,0.02,0.0,0.0,0.0,0.0,2.78,6.81,1.8,0.02,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08,0.14,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.049999997,0.08,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.97999996,7.0499997,4.23,1.5999999,0.0,0.0,0.0,0.26,1.3,1.8299999,2.24,2.55,3.22,2.73,1.9799999,0.84,0.44,0.41,0.11,0.22999999,0.24,0.17999999,0.26,0.0,0.0,0.02,0.22,0.29999998,0.22,0.14,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.03,0.089999996,0.099999994,0.06,0.11,0.089999996,0.25,0.72999996,1.77,1.64,0.71999997,0.16,0.02,0.0,0.11,0.52,0.26999998,1.12,3.6699998,6.79,11.28,10.33,8.849999,10.349999,13.86,13.049999,12.69,13.37,15.83,12.54,7.52,5.7599998,4.93,4.25,3.34,2.03,1.0,1.73,4.2,8.5,8.49,8.76,10.32,15.54,18.15,21.32,24.21,35.079998,51.3,59.98,63.3,57.46,58.05,45.629997,25.24,4.7799997,3.22,3.75,5.31,16.58,15.009999,14.7699995,19.42,10.28,4.35,2.21,2.12,3.6499999,5.67,7.41,8.099999,10.51,12.349999,10.26,9.29,10.469999,11.55,12.2699995,6.67,2.31,3.3899999,4.7599998,6.92,11.65,13.849999,11.96,10.34,8.92,10.719999,10.55,11.219999,15.969999,20.199999,19.25,14.16,16.4,18.68,26.939999,19.42,6.74,8.61,17.25,15.74,12.11,8.929999,2.0,0.48,0.42999998,0.0,0.0,2.61,1.8,0.0,0.0,0.0,0.16,0.51,0.12,0.0,0.0,0.0,0.0,0.03,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.81,1.87,0.53999996,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.12,0.17999999,0.29,0.39999998,0.11,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.049999997,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,4.74,1.68,2.22,0.03,0.099999994,0.04,0.049999997,0.63,1.2099999,1.37,2.18,3.27,3.28,2.33,1.0699999,0.78,2.21,1.9699999,0.02,0.11,0.53,0.59999996,0.08,0.03,0.01,0.0,0.04,0.08,0.08,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.22,0.14999999,0.22999999,0.39,0.26,0.32,0.57,0.59,0.47,0.089999996,0.0,0.0,0.0,0.28,0.53,0.72999996,1.5799999,2.7,8.15,9.05,14.23,9.75,15.24,18.939999,18.49,16.69,16.08,14.07,10.2699995,8.01,5.58,5.45,7.3599997,7.06,4.61,9.19,15.809999,22.39,21.06,22.289999,25.269999,27.539999,23.67,29.609999,43.879997,53.44,63.77,76.229996,75.909996,72.4,64.17,26.189999,10.29,1.6899999,0.93,0.65999997,2.57,9.66,7.3199997,5.14,3.1699998,1.9399999,1.02,1.52,4.67,8.34,12.04,14.74,13.49,15.88,17.619999,14.37,15.21,15.809999,15.99,14.21,4.99,2.02,4.0299997,6.18,10.349999,13.95,13.29,9.13,8.86,11.74,14.37,12.67,13.11,15.389999,17.17,13.969999,12.25,12.74,15.57,19.21,13.139999,5.43,8.67,11.53,8.309999,6.7999997,4.0299997,0.68,0.049999997,0.0,0.0,0.0,4.7799997,0.58,0.03,0.0,1.0,2.45,1.67,0.0,0.0,0.0,0.02,0.12,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.04,0.06,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.01,0.08,0.14,0.11,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.9399999,7.33,0.0,0.02,0.68,0.57,0.26,0.55,0.59999996,0.69,0.95,1.89,1.86,1.09,0.48999998,2.25,5.41,4.8199997,1.8199999,2.74,3.56,2.3,0.32,0.22,0.11,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.049999997,0.01,0.01,0.19,0.45999998,0.59999996,0.65999997,0.38,0.089999996,0.32,0.72999996,0.71999997,0.89,0.7,0.08,0.0,0.13,0.71,0.58,0.44,0.71999997,1.14,2.26,6.0699997,7.7799997,8.28,12.36,21.84,29.109999,35.53,31.179998,17.16,12.48,11.44,17.44,21.52,26.71,30.65,42.87,35.62,36.59,49.489998,59.91,60.44,58.62,46.989998,54.76,40.69,35.42,53.21,48.86,38.739998,37.07,14.7699995,6.39,0.34,0.32999998,0.14999999,0.34,2.09,4.9,3.4399998,1.64,0.29,0.82,1.86,3.36,6.56,11.509999,19.38,22.67,21.439999,19.779999,19.22,17.99,17.31,19.52,25.369999,16.24,3.86,3.01,5.48,7.6699996,11.79,15.33,13.849999,10.599999,10.7,13.509999,15.009999,12.88,11.86,13.37,13.509999,11.62,9.3,9.7,7.95,10.13,5.83,5.29,5.2999997,4.33,3.23,2.54,0.78,0.04,0.0,0.0,0.02,0.42,0.69,0.75,0.89,1.23,6.64,17.789999,18.449999,4.7,0.24,0.02,0.07,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.049999997,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06,0.0,0.0,0.0,0.0,0.0,0.47,3.97,0.13,0.39999998,0.47,2.03,1.24,0.98999995,0.12,0.32999998,0.44,0.91999996,0.85999995,0.71,0.53,0.29,0.39,1.68,2.52,2.01,2.37,2.11,0.78999996,1.67,1.8199999,0.14999999,0.099999994,0.08,0.0,0.0,0.0,0.0,0.0,0.01,0.08,0.11,0.0,0.0,0.0,0.0,0.0,0.02,0.07,0.07,0.02,0.08,0.14999999,0.11,0.03,0.22,0.47,0.85999995,1.02,0.74,0.51,0.87,0.39,0.51,0.77,1.78,1.76,0.48,0.24,0.19,0.95,1.13,1.3,1.22,1.11,5.43,5.92,1.81,9.74,34.53,70.04,104.11,130.55,75.08,42.399998,41.379997,48.739998,62.219997,72.08,49.05,61.25,41.66,31.869999,44.329998,69.35,97.92,113.1,71.43,59.329998,25.9,15.74,11.17,10.83,8.71,5.92,1.1,0.31,0.0,0.0,0.0,0.03,0.29999998,0.74,0.5,0.32,0.14,0.03,0.13,1.64,4.49,7.18,11.44,20.029999,26.17,23.73,18.18,15.82,14.15,14.5,21.92,25.13,15.429999,5.0299997,5.42,6.87,9.25,12.03,17.23,18.92,15.259999,11.36,8.98,10.44,11.139999,10.98,11.88,10.65,10.929999,16.08,7.2999997,12.98,12.509999,9.599999,6.0299997,3.24,3.48,2.74,1.88,1.0799999,0.34,0.03,0.0,0.17,0.48,0.64,1.3399999,1.37,4.43,11.86,12.41,11.7699995,12.05,5.5,1.22,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.39,0.93,0.0,0.0,0.0,0.0,0.0,1.5,1.48,1.0,0.03,0.66999996,1.31,2.6699998,0.35,0.03,0.28,2.2,0.35999998,0.19999999,0.34,0.26,0.51,0.19,1.17,1.5899999,1.8199999,0.96,0.79999995,0.84999996,0.65,0.26,0.39,0.29999998,0.28,0.25,0.55,0.82,1.88,3.6899998,3.53,1.53,0.32,0.22999999,0.11,0.14999999,0.11,0.0,0.0,0.0,0.0,0.04,0.02,0.04,0.049999997,0.0,0.0,0.0,0.0,0.01,0.049999997,0.089999996,0.29,0.35999998,0.39,0.52,0.72999996,0.72999996,0.45999998,1.39,1.18,0.91999996,0.65,0.59,1.0799999,0.94,0.89,0.44,0.13,0.39999998,0.56,0.25,0.39,0.52,0.89,1.8299999,3.6599998,4.5099998,6.41,11.929999,13.469999,17.67,34.69,60.399998,70.93,83.03,84.32,79.97,64.659996,69.38,72.53,60.28,50.309998,46.27,33.809998,20.029999,35.69,50.36,57.3,87.4,86.6,35.84,16.89,7.8799996,2.96,2.28,1.3399999,0.26,0.0,0.0,0.19,0.16,0.0,0.0,0.0,0.06,0.049999997,0.01,0.0,0.03,0.28,2.1399999,7.3399997,9.389999,8.7699995,11.09,17.449999,19.63,16.58,13.86,12.75,12.179999,13.82,20.13,22.51,13.29,5.83,6.7599998,9.7699995,14.04,14.54,13.87,17.41,17.34,10.5199995,8.679999,9.41,9.809999,10.44,10.639999,10.8,22.65,13.91,18.619999,30.179998,27.789999,10.24,3.82,1.5799999,1.27,1.53,1.5699999,1.0699999,0.78,2.07,5.1099997,5.45,5.38,8.03,8.95,9.92,12.44,6.2599998,3.98,5.7799997,8.349999,2.45,0.0,0.0,0.049999997,0.25,0.049999997,0.0,0.0,0.0,0.0,0.0,0.0,0.06,0.03,0.04,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.01,0.0,0.0,0.0,0.0,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.38,0.7,0.0,0.0,0.0,0.0,0.84,4.36,7.48,9.55,8.55,10.96,10.349999,10.7699995,3.75,2.44,4.27,9.04,6.3599997,2.62,1.81,0.049999997,0.03,0.089999996,0.19,0.68,0.90999997,1.23,1.05,0.75,1.06,0.32,0.0,0.59,1.39,2.08,1.49,1.25,0.89,0.44,0.83,1.22,0.91999996,0.52,0.32999998,0.19999999,0.32,0.089999996,0.02,0.0,0.0,0.0,0.099999994,0.099999994,0.07,0.0,0.0,0.0,0.0,0.099999994,0.41,0.29,0.16,0.62,1.18,0.90999997,0.93,1.31,1.61,1.67,1.9599999,1.1899999,0.78,0.84,0.59999996,0.37,0.45999998,0.26999998,0.0,0.11,0.61,0.42999998,0.28,0.63,0.98999995,1.8,2.62,3.9599998,7.8399997,15.929999,23.48,36.41,42.57,50.329998,63.46,86.21,114.24,105.649994,78.07,61.6,61.5,60.18,47.44,44.219997,33.87,24.289999,26.289999,41.28,35.739998,55.59,36.53,26.49,6.06,2.02,1.14,0.39999998,0.08,0.0,0.0,0.0,0.16,0.89,0.66999996,0.03,0.0,0.0,0.0,0.0,0.08,0.089999996,0.0,1.02,4.5,9.71,12.889999,10.28,8.38,8.0,12.11,14.24,16.859999,19.279999,15.5,14.2699995,22.949999,20.789999,10.16,5.75,6.95,12.12,17.39,18.47,11.58,11.17,14.71,14.33,12.55,10.37,9.03,10.0,13.82,21.68,16.18,14.24,20.699999,14.299999,6.62,6.0699997,3.1999998,1.3,1.02,0.7,0.26,1.0,4.73,8.48,9.429999,11.559999,11.58,8.97,10.41,11.679999,7.91,6.0099998,4.65,2.3,0.049999997,0.0,0.01,0.44,0.75,0.29999998,0.0,0.0,0.0,0.0,0.0,0.0,0.02,0.38,0.59999996,0.11,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.04,0.02,0.07,0.13,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.37,0.11,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.59999996,1.74,0.96,0.88,2.18,5.66,10.87,22.109999,20.58,21.279999,19.0,21.02,12.719999,13.049999,16.48,19.609999,12.469999,16.369999,7.3399997,0.0,0.0,0.0,0.0,0.07,0.03,0.88,0.47,0.19999999,0.26,0.17,0.049999997,0.21,0.96999997,1.15,0.65,0.47,0.85999995,0.61,0.45999998,0.88,0.48,0.13,0.13,0.28,0.78999996,0.48,0.13,0.099999994,0.04,0.0,0.0,0.0,0.01,0.01,0.0,0.0,0.12,0.24,0.42,0.69,0.74,0.58,0.85999995,1.9399999,1.89,1.28,1.24,1.73,2.27,1.62,0.93,0.66999996,0.75,0.9,0.96999997,0.39999998,0.14999999,0.29999998,1.06,1.86,2.3,2.1399999,1.67,2.07,3.57,7.41,10.7,18.09,36.98,61.39,57.78,50.649998,53.699997,66.909996,89.02,104.88,95.159996,81.42,61.289997,64.729996,52.39,54.489998,50.53,46.42,37.82,20.74,8.54,15.559999,20.58,17.76,4.6,2.1,3.1299999,1.1,0.049999997,0.0,0.0,0.0,0.0,0.049999997,0.08,0.03,0.02,0.01,0.0,0.0,0.04,0.29,0.53,0.32,1.5,4.0899997,8.69,12.639999,11.0199995,9.7,7.2999997,10.179999,15.059999,20.26,17.39,15.929999,16.84,18.26,16.449999,10.08,6.33,6.7,13.0199995,15.339999,13.84,9.92,8.83,12.059999,16.26,17.199999,11.59,8.37,8.74,10.95,10.26,7.68,5.97,3.26,3.79,2.72,5.0499997,5.62,3.79,2.1699998,2.18,2.55,5.18,9.54,13.599999,22.23,14.2,6.5099998,2.9099998,3.78,4.21,3.6699998,4.43,1.8399999,0.44,0.099999994,0.07,0.06,0.13,0.049999997,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.089999996,0.55,0.44,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.03,0.0,0.0,0.53999996,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.089999996,0.13,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.16,1.15,2.24,2.3,1.66,1.03,7.71,12.46,21.689999,32.739998,37.21,43.18,48.53,56.8,38.48,29.599998,32.809998,39.399998,37.0,39.46,24.279999,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.0,0.0,0.01,0.01,0.01,0.0,0.03,0.14,0.17999999,0.29999998,0.55,0.39999998,0.19,0.48999998,0.56,0.58,0.39999998,0.06,0.17999999,0.14999999,0.19999999,0.48,0.25,0.0,0.0,0.0,0.0,0.0,0.07,0.19,0.34,0.45999998,0.26999998,0.39,0.72999996,0.85999995,0.96999997,1.27,2.28,3.4299998,5.12,2.82,2.73,2.48,1.5,0.85999995,1.04,0.74,0.34,0.26,0.28,0.39999998,1.42,2.4199998,2.8799999,3.01,3.5,6.24,7.81,12.86,21.539999,36.95,59.07,68.82,90.78,117.32,134.12999,129.25,135.0,130.73999,104.579994,83.78,80.29,71.89,79.71,63.03,49.52,56.11,32.61,20.76,4.3199997,3.3999999,12.07,4.98,0.68,1.23,0.24,0.25,0.24,0.04,0.0,0.0,0.06,0.0,0.0,0.03,0.22999999,0.25,0.25,0.29999998,0.099999994,0.28,0.53,0.16,0.74,2.36,4.38,6.83,8.79,8.389999,7.96,11.0,18.949999,20.93,14.429999,11.969999,13.5,16.699999,15.38,10.5,7.37,6.19,12.9,12.95,6.48,5.02,5.99,7.91,13.59,17.859999,13.95,7.91,5.42,3.31,5.35,6.7599998,5.19,1.37,0.89,1.18,3.37,5.94,5.7999997,5.96,4.74,4.67,7.5099998,10.48,12.07,5.8199997,3.3,5.22,5.99,0.76,0.07,0.85999995,2.62,3.1399999,2.11,2.07,0.59,0.21,0.0,0.0,0.0,0.02,0.0,0.0,0.0,0.0,0.02,0.02,0.32,0.17,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06,0.07,0.0,0.0,0.59999996,0.64,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.51,2.6,2.6399999,2.36,0.82,0.81,9.54,13.349999,20.31,34.1,36.96,51.35,54.579998,60.12,57.8,50.379997,51.61,71.06,67.38,58.21,42.25,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.42999998,0.66999996,0.29,0.12,0.0,0.0,0.11,0.89,0.78,0.96999997,0.78,0.38,0.5,0.65,0.24,0.26,0.17,0.31,0.35999998,0.22,0.19,0.12,0.17,0.06,0.0,0.0,0.0,0.01,0.08,0.049999997,0.34,0.71999997,0.51,0.75,1.93,2.95,2.81,2.71,3.28,5.72,5.37,3.1499999,4.11,4.2599998,1.79,0.58,0.69,0.55,0.29,0.48999998,0.65,1.13,2.62,5.35,5.0299997,2.3,4.72,10.639999,12.61,17.18,24.84,35.8,46.649998,69.72,120.43,133.23,123.93,104.7,123.04,126.619995,116.369995,127.71999,95.35,100.119995,58.92,56.62,71.71,67.58,38.649998,6.19,1.8399999,6.5899997,2.5,0.47,0.089999996,0.0,0.04,0.96999997,0.65999997,0.65,0.06,0.26999998,0.13,0.01,0.04,0.08,0.17,0.48,0.71,1.0799999,0.28,0.22999999,0.78,0.93,1.18,1.93,2.28,4.15,6.58,8.47,8.86,12.719999,17.539999,20.09,13.509999,10.2,10.92,14.94,14.95,10.78,7.21,5.6,14.19,11.08,4.0499997,2.73,3.1299999,4.87,9.84,18.17,10.17,4.88,3.02,4.7,8.71,9.0199995,7.3599997,4.45,2.37,1.4499999,6.91,11.15,10.46,9.2,4.3399997,3.31,1.75,1.29,1.29,2.95,3.97,1.99,0.37,1.6899999,1.9399999,2.05,1.68,0.52,1.56,4.38,0.19999999,0.0,0.0,0.03,0.11,0.08,0.01,0.0,0.0,0.01,0.0,0.049999997,0.17999999,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.0,0.0,0.0,1.81,0.25,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.83,0.47,0.39,0.42,1.9799999,7.75,11.7,18.529999,30.63,42.8,52.449997,59.27,70.65,60.739998,63.5,58.8,83.009995,68.49,58.14,51.42,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.04,0.44,0.83,1.4599999,1.29,0.01,0.19999999,0.91999996,0.96,0.81,0.69,0.96,0.42,0.14,0.03,0.049999997,0.14999999,0.28,0.07,0.41,0.57,0.11,0.29999998,0.48999998,0.56,1.12,1.66,1.23,0.81,0.12,0.16,0.62,1.79,2.34,4.47,8.98,11.59,13.799999,7.93,5.8599997,6.12,5.9,4.72,5.43,4.35,1.9599999,0.84,1.17,0.78999996,0.47,0.94,1.79,2.8,4.5099998,7.83,8.96,7.5,7.1,8.59,9.67,16.42,26.779999,42.1,46.75,74.119995,104.22,87.479996,64.97,62.12,89.259995,119.28,111.909996,107.24,102.14,72.82,71.43,80.13,79.509995,44.559998,10.16,6.2999997,2.8799999,1.16,0.69,0.0,0.0,0.0,0.75,1.43,2.35,1.49,0.03,0.04,0.16,0.17999999,0.14999999,0.25,0.29,0.53,0.89,0.96999997,0.48999998,0.7,1.77,2.6,2.85,3.22,3.6499999,2.6799998,4.65,5.85,8.059999,9.809999,15.809999,15.49,13.16,11.5,9.36,10.34,13.66,13.389999,7.7999997,6.99,10.09,7.48,3.9499998,2.03,2.53,5.3399997,7.96,5.8799996,5.06,5.94,7.31,11.429999,10.65,7.3999996,5.47,4.37,2.81,2.2,6.37,7.6299996,8.7,6.2799997,2.21,1.3,1.86,2.95,3.1399999,3.3999999,1.01,0.97999996,2.82,4.71,5.6299996,5.17,4.27,3.1699998,2.23,1.6899999,0.59999996,0.74,1.23,1.17,0.51,0.14,0.0,0.0,0.0,0.0,0.0,0.01,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.79,1.31,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.35,2.87,5.66,10.38,16.05,22.189999,32.27,57.62,81.729996,105.54,98.99,76.7,45.739998,52.96,47.0,52.91,46.95,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.64,0.35999998,0.0,0.26999998,0.82,1.9799999,1.18,0.07,0.14999999,0.06,0.14999999,0.0,0.07,0.35999998,0.45999998,0.7,0.83,0.59,0.78,1.79,3.04,4.19,4.45,3.6799998,4.25,4.25,1.27,2.3799999,6.7799997,8.95,7.6099997,20.88,25.24,16.34,14.13,11.05,6.91,5.91,6.37,5.44,7.6299996,9.0199995,8.46,6.0,2.34,0.93,0.78999996,1.63,2.6299999,6.2599998,9.46,9.34,9.13,8.28,8.599999,6.6299996,5.3399997,5.12,8.29,8.46,16.71,33.73,41.21,33.21,36.38,46.57,59.949997,65.58,60.699997,48.23,67.71,105.03,66.63,45.95,29.05,4.69,1.51,1.43,1.5799999,1.54,0.0,0.26999998,0.96,0.32999998,0.91999996,2.37,2.06,0.66999996,0.34,0.12,0.24,0.38,0.41,0.35,0.48999998,1.0,1.18,1.06,0.63,2.33,4.11,5.58,6.08,7.99,4.68,2.11,2.05,3.1799998,5.6099997,9.84,12.19,10.21,6.96,7.68,7.95,6.5,7.06,8.99,7.06,4.12,3.12,3.52,3.36,2.1499999,5.39,5.24,4.75,5.15,7.96,13.66,15.679999,12.5199995,5.79,2.8999999,1.48,1.28,2.73,4.94,9.059999,13.599999,17.69,11.139999,4.24,3.85,5.2,6.47,8.36,4.63,4.24,5.0099998,7.12,9.11,11.01,10.2699995,7.5299997,4.56,2.8999999,2.3999999,2.12,2.34,2.6699998,3.08,0.78,0.0,0.0,0.0,0.0,0.0,0.0,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,6.12,2.26,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.17999999,0.35,1.6999999,4.0299997,8.429999,11.8,14.809999,18.4,43.719997,52.86,75.85,92.299995,66.93,48.579998,70.659996,65.979996,67.17,45.64,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.0,0.0,0.0,0.11,0.52,0.61,0.69,0.53,0.25,0.35,0.17999999,0.14999999,0.06,0.16,0.83,1.5899999,1.55,1.15,1.5799999,2.9099998,5.25,7.3799996,6.15,4.92,3.21,2.6599998,2.84,3.9199998,7.5499997,10.429999,16.21,14.45,17.66,17.31,12.24,9.0199995,9.73,12.259999,10.58,10.87,11.559999,8.28,9.71,7.3199997,3.8899999,3.03,2.8799999,4.14,7.96,11.75,14.78,13.48,11.74,8.24,3.4099998,2.0,0.42999998,0.7,2.75,6.0,9.3,19.14,20.609999,9.34,14.5199995,18.289999,17.82,16.869999,35.93,50.26,37.82,20.41,10.44,0.64,0.0,0.34,0.39,0.94,0.0,0.099999994,1.22,1.4,0.28,0.71999997,0.48999998,0.14999999,0.22,0.48,0.95,1.42,1.13,1.64,1.68,0.94,0.87,0.78999996,0.48999998,0.62,1.99,4.5699997,6.52,6.23,5.85,3.58,2.37,2.62,1.51,2.12,5.43,10.87,9.139999,4.8399997,2.8899999,3.84,4.5499997,3.61,2.8799999,2.78,2.22,1.74,1.37,2.86,4.5299997,6.0899997,7.1499996,6.87,6.37,8.349999,9.809999,8.889999,8.25,3.6699998,1.16,0.48,2.47,1.8299999,3.1,10.96,19.06,11.71,5.41,5.49,8.8,10.429999,11.82,7.9199996,10.389999,14.24,12.429999,13.849999,19.109999,19.289999,13.719999,8.679999,5.0099998,2.72,0.96,0.37,1.27,2.51,0.59999996,0.0,0.0,0.0,0.04,0.08,0.0,0.0,0.0,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.78,3.11,1.9,0.089999996,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06,0.37,0.39,0.06,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.049999997,0.0,0.0,0.42999998,3.26,6.21,6.93,10.86,24.33,33.66,31.939999,43.76,52.98,73.34,63.649998,69.01,52.629997,49.09,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.04,0.13,0.19999999,0.35999998,0.39,0.21,0.51,0.35,0.0,0.0,0.01,0.19,0.22999999,0.35,0.57,1.4,3.6399999,6.47,7.22,6.62,3.4499998,1.8399999,3.33,5.1099997,5.7799997,10.26,14.19,15.719999,13.48,13.59,12.559999,10.91,13.75,13.94,16.14,12.13,8.91,7.5899997,6.7,8.37,10.3,7.3199997,3.3,3.1499999,3.5,5.19,9.15,9.5,8.69,6.24,3.9399998,2.02,1.38,2.58,5.45,9.849999,15.11,21.38,15.99,7.91,5.8399997,5.0099998,3.01,6.1299996,19.13,28.119999,21.449999,2.9399998,0.26,0.0,0.0,0.0,0.0,0.07,0.0,0.0,0.0,0.03,0.02,0.0,0.0,0.0,0.0,0.04,0.5,0.59999996,1.52,1.18,1.5,1.9499999,4.19,6.92,3.75,1.41,1.11,1.29,2.1399999,4.2799997,5.96,4.39,4.04,4.58,3.85,2.85,1.3299999,2.59,7.89,12.08,9.059999,4.72,1.2099999,1.5799999,1.48,0.59,0.42999998,0.75,0.81,1.36,3.6599998,5.74,6.17,6.12,8.96,5.3399997,3.1399999,3.7099998,6.5499997,7.58,3.8999999,2.97,2.28,1.15,1.75,3.51,4.45,3.27,2.54,3.9199998,4.95,5.87,7.3999996,3.8,7.14,18.06,22.59,20.4,20.0,23.99,23.71,16.369999,8.21,2.24,0.11,0.0,0.17,0.26,0.02,0.0,0.0,0.0,0.03,0.04,0.01,0.0,0.0,0.049999997,0.089999996,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.04,0.47,6.68,2.37,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.12,0.84999996,1.13,0.45999998,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02,0.089999996,0.0,0.0,0.78999996,1.43,1.7199999,2.1599998,7.1499996,12.58,25.97,20.76,28.89,52.87,90.159996,93.45,68.909996,53.949997,41.05,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.049999997,0.0,0.01,0.04,0.03,0.099999994,0.11,0.0,0.0,0.0,0.0,0.04,0.37,1.3399999,2.01,2.22,1.99,2.84,3.06,4.93,3.46,2.52,2.24,3.6,8.29,13.99,15.61,13.66,11.3,12.12,11.65,11.07,10.55,12.25,14.839999,11.86,7.85,6.3999996,4.5499997,7.93,9.059999,7.0,4.69,3.6799998,4.5499997,5.2999997,6.2999997,7.5499997,8.71,8.92,5.68,3.4499998,4.8199997,5.91,4.23,5.0,5.24,1.66,0.14999999,0.17,0.38,0.53,2.3999999,5.3399997,7.48,5.8599997,1.77,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.08,0.14999999,0.65,0.0,0.0,0.0,0.0,0.0,0.07,0.51,0.98999995,1.5699999,2.95,3.3999999,4.54,8.4,10.36,7.69,4.5299997,2.29,1.9799999,2.59,4.6,5.5299997,4.9,5.15,5.5299997,5.8199997,6.29,4.22,3.3999999,2.7,1.9699999,1.49,0.53,0.26999998,0.44,0.42,0.45,0.69,0.69,0.74,1.91,4.7599998,6.5899997,7.75,26.91,15.28,4.02,1.92,2.6499999,3.79,3.55,3.33,3.32,2.75,1.9699999,2.1399999,2.59,2.23,1.27,1.4,2.03,3.02,2.24,0.64,1.4699999,4.88,7.8399997,6.62,5.43,5.0899997,5.5499997,4.13,2.07,0.51,0.049999997,0.22999999,0.39999998,0.65,0.12,0.41,0.06,0.0,0.089999996,0.17999999,0.02,0.0,0.0,0.0,0.08,0.13,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.099999994,0.07,0.02,6.37,8.42,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.31,0.53,0.22999999,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.04,0.13,0.26999998,0.29,0.099999994,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.22,0.0,0.08,0.39999998,0.47,0.26,1.05,4.72,10.32,19.56,12.7699995,18.779999,34.77,44.27,91.189995,84.15,63.039997,52.969997,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.17,0.19,0.14,0.17999999,0.22999999,0.25,0.45999998,0.21,0.14999999,0.089999996,0.03,0.52,0.5,0.41,0.39999998,1.05,1.03,0.35,0.21,0.58,0.83,0.65,1.17,1.54,4.73,6.75,8.139999,8.29,10.48,13.54,10.55,7.33,7.3799996,8.8,10.2699995,11.48,11.63,12.099999,9.69,5.35,6.31,9.2699995,14.559999,13.469999,13.63,12.32,10.55,10.809999,11.86,10.809999,10.349999,18.289999,16.17,10.76,9.12,5.4,3.34,0.91999996,0.19,3.79,4.08,9.69,11.84,0.93,0.0,0.049999997,0.0,0.0,0.0,0.0,0.07,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.04,0.63,0.0,0.0,0.0,0.0,0.0,0.12,2.82,9.0199995,9.37,11.01,13.5,12.21,13.11,13.73,10.62,6.79,7.1099997,7.6499996,7.95,6.69,6.71,6.24,5.77,4.16,2.49,1.3,0.45,0.7,0.42,0.049999997,0.22,0.45999998,0.88,1.0,0.52,0.77,0.84,0.88,2.7,4.75,2.81,3.6299999,3.4399998,2.1399999,0.45999998,0.17,1.2099999,2.29,2.32,4.0899997,2.29,1.12,0.77,0.77,1.36,0.66999996,0.39,0.66999996,1.01,1.25,1.89,5.22,8.92,11.3,9.639999,5.37,2.95,1.8299999,0.96,0.29,0.83,2.8899999,1.7199999,0.64,0.32,0.68,9.16,20.58,5.97,1.42,0.28,0.65999997,0.06,0.0,0.0,0.0,0.0,0.01,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07,0.26999998,0.0,6.06,11.469999,0.13,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.42999998,0.74,0.96999997,0.89,0.65999997,0.049999997,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.35,0.66999996,0.0,0.0,0.13,0.19999999,1.0,3.36,7.3399997,8.16,7.31,10.63,12.759999,20.1,26.08,56.12,93.579994,106.78,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.049999997,0.099999994,0.099999994,0.26,0.38,0.65999997,0.78999996,0.58,0.39,0.13,0.01,0.08,0.26,0.47,0.14999999,0.12,0.25,0.13,0.19999999,0.22,0.35999998,0.5,0.88,2.02,3.25,3.6999998,5.2,7.48,9.4,6.8599997,5.08,4.8199997,5.6,5.72,6.3799996,8.66,9.75,11.54,12.75,14.63,20.17,32.329998,37.69,29.779999,23.789999,16.869999,10.91,9.04,10.4,15.54,28.88,25.519999,22.17,21.289999,8.26,4.0899997,2.28,1.17,4.89,8.55,17.34,14.37,2.6799998,0.0,0.0,0.0,0.87,2.0,2.1499999,1.8299999,0.0,0.03,0.0,0.0,0.07,0.32999998,0.65,7.1299996,8.54,0.26,0.12,0.04,0.08,0.53999996,1.22,3.1699998,4.48,6.69,8.23,14.28,16.89,14.5199995,15.0,16.94,13.509999,9.37,7.81,6.48,4.99,6.71,5.6299996,4.0099998,2.9399998,1.5,1.49,0.90999997,0.19999999,0.63,0.45999998,0.16,0.45,0.63,0.57,0.95,0.71999997,0.45,0.48999998,0.81,2.48,3.32,3.11,2.0,1.5999999,0.45999998,0.07,0.62,1.89,1.5899999,2.52,1.53,1.52,1.3,1.06,0.87,0.82,1.14,1.3299999,0.53,0.08,1.18,4.79,8.16,10.58,10.7699995,8.679999,8.139999,6.46,3.74,2.3799999,3.6899998,5.79,1.12,0.0,0.0,0.35,17.84,46.45,17.75,4.69,4.33,0.84,0.59999996,0.0,0.0,0.0,0.0,0.0,0.06,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08,0.0,7.2,13.29,1.51,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.26999998,0.45999998,1.01,0.96,1.13,0.25,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.35,0.59,0.0,0.0,0.089999996,0.19999999,0.81,2.33,5.68,4.46,3.74,6.91,9.7,16.3,20.34,62.91,80.4,90.68,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.049999997,0.089999996,0.17999999,0.41,0.42999998,0.56,0.77,0.28,0.19,0.17,0.21,0.59,0.71999997,0.12,0.03,0.37,0.34,0.099999994,0.13,0.53999996,0.48999998,0.32999998,0.17,0.39,0.62,0.72999996,2.0,2.3999999,3.11,3.32,4.5299997,5.41,4.14,3.34,3.85,4.71,3.8999999,4.38,9.059999,13.62,15.69,17.75,20.949999,33.52,48.44,60.84,67.14,61.64,53.789997,47.129997,38.079998,29.179998,43.82,34.11,28.32,9.42,2.4199998,1.29,2.1299999,3.4199998,8.03,14.04,8.19,3.55,0.22999999,0.0,0.0,0.0,0.02,2.4299998,3.58,2.45,0.0,0.0,0.12,0.04,0.12,0.66999996,2.53,9.41,9.38,0.14,0.07,0.26999998,0.53999996,1.41,3.59,9.99,16.1,15.53,13.15,14.74,15.889999,18.949999,18.56,16.76,16.38,14.33,10.51,5.94,3.57,2.85,3.1999998,2.4099998,0.87,0.35,0.48999998,0.48999998,0.42,0.44,0.39999998,0.34,0.32,0.45,0.84999996,0.84,0.53999996,0.049999997,0.099999994,0.52,0.59,1.61,3.3,2.9099998,1.65,1.3399999,1.9799999,1.24,0.64,0.65,1.15,2.18,2.32,1.68,2.33,0.74,0.37,0.089999996,0.06,0.099999994,1.26,6.0699997,11.48,11.25,8.05,4.3399997,3.74,3.25,2.9199998,3.54,2.84,4.48,4.0699997,2.6,1.5899999,0.45,0.11,6.7799997,17.119999,5.1,1.43,5.6,5.1099997,2.1599998,1.28,0.65,0.13,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,3.06,10.61,7.31,0.12,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.04,0.19999999,0.28,0.62,0.29999998,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02,0.19999999,0.17999999,0.72999996,1.38,1.5999999,2.1699998,8.36,10.5199995,14.92,18.41,42.75,72.15,93.92,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02,0.19,0.049999997,0.07,0.26999998,0.37,0.35999998,0.21,0.19,0.22,0.38,0.04,0.0,0.01,0.19,0.17,0.24,0.48,0.48,0.28,0.24,0.17,0.39999998,0.90999997,1.2099999,2.32,4.44,3.81,3.1399999,2.83,2.8899999,2.8899999,3.74,6.12,8.87,11.23,10.71,11.11,11.099999,11.13,10.92,14.589999,23.1,36.19,45.68,47.71,46.05,48.809998,38.829998,26.97,24.699999,19.81,8.51,0.96999997,1.4699999,1.27,1.05,0.35999998,0.77,1.1,0.17,0.04,0.0,0.0,0.0,0.0,0.0,0.0,0.35999998,1.53,1.11,1.22,2.3899999,1.29,1.65,1.05,1.99,4.15,3.81,0.14,0.0,0.099999994,0.11,0.16,0.48999998,4.81,10.82,18.619999,19.449999,16.49,16.07,14.16,16.47,19.05,19.09,19.05,19.66,11.139999,5.38,1.9,1.42,1.5699999,1.13,0.69,0.02,0.0,0.0,0.099999994,0.7,0.72999996,0.5,0.9,1.56,1.03,1.36,1.13,0.56,0.11,0.07,0.14,0.11,0.5,0.74,0.56,0.42,0.26999998,0.26,0.26999998,1.02,1.5799999,1.13,0.7,0.98999995,1.73,0.35,0.0,0.0,0.32,1.4399999,4.83,9.849999,12.28,10.639999,7.93,4.0,1.51,0.28,0.35,0.97999996,1.55,3.5,10.309999,13.679999,6.7799997,1.51,0.04,0.0,0.0,0.38,1.8199999,2.98,1.17,1.41,2.97,3.1599998,0.71,0.0,0.03,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,8.79,5.5899997,1.17,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.04,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.14999999,0.03,0.0,0.0,0.0,0.0,0.29,0.24,0.0,0.0,0.0,0.0,0.0,0.29,0.76,0.45,0.13,0.0,0.0,0.0,0.37,0.71,0.16,1.35,0.76,2.57,9.51,12.639999,14.299999,13.79,25.34,63.39,78.22,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.089999996,0.22999999,0.22,0.29999998,0.51,0.47,0.32999998,0.28,0.28,0.32999998,0.38,0.62,0.21,0.03,0.24,0.25,0.29999998,0.5,0.25,0.26,0.35,0.41,0.79999995,1.52,2.6299999,3.46,3.8899999,4.7599998,3.6899998,2.84,3.33,3.81,2.06,2.99,5.7999997,9.2,15.299999,18.949999,14.7699995,7.29,4.77,6.92,12.679999,19.76,21.859999,23.59,26.189999,23.199999,14.34,9.08,5.65,4.21,3.9399998,4.62,6.14,4.39,1.4499999,0.48999998,0.0,0.089999996,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.0799999,4.16,7.6099997,4.0,5.42,11.469999,6.08,0.19,0.22,0.34,0.68,0.52,0.0,0.0,0.0,0.0,0.08,2.81,7.14,13.59,20.41,15.549999,14.7699995,12.9,10.17,6.58,6.16,8.08,8.57,6.72,4.5699997,1.75,0.98999995,1.81,1.4499999,1.28,0.58,0.14,0.089999996,0.0,0.03,0.21,0.52,0.45,0.45999998,1.81,1.86,1.63,0.9,0.22,0.17,0.22,0.13,0.01,0.07,0.06,0.04,0.099999994,0.39999998,1.6899999,0.85999995,0.47,0.42,0.42999998,0.39999998,0.68,1.3199999,0.53,0.08,0.049999997,0.06,0.44,0.97999996,1.4399999,1.91,3.3799999,3.61,2.45,0.89,1.06,3.47,0.78,2.04,7.3599997,18.88,14.139999,14.4,5.79,1.0799999,0.03,0.19,1.03,1.03,0.21,0.32999998,2.09,7.14,5.66,1.62,0.42999998,0.099999994,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,3.76,5.1099997,2.47,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.04,0.14999999,0.049999997,0.0,0.04,0.11,0.02,0.0,0.0,0.0,0.0,0.0,0.01,0.099999994,0.56,0.68,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.64,0.78999996,0.59999996,0.53999996,0.04,0.0,0.0,0.049999997,0.12,0.0,0.0,0.0,0.0,0.0,0.62,1.3399999,0.88,0.24,0.75,1.75,2.24,2.71,1.6899999,1.0,0.71,0.94,2.27,7.04,13.32,16.119999,16.39,31.06,68.65,84.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.049999997,0.51,0.90999997,0.65999997,0.78,0.59999996,0.37,0.25,0.14,0.38,0.53,0.59999996,0.55,0.14,0.06,0.39,0.74,0.29,0.48999998,0.55,0.51,1.16,1.6899999,2.11,3.24,3.85,3.77,3.48,3.1899998,2.79,2.3999999,2.6399999,2.18,1.68,3.09,4.29,8.26,8.69,10.94,7.62,2.62,7.43,20.35,27.05,22.949999,16.619999,8.48,4.87,2.9399998,3.6599998,14.5199995,14.86,9.53,19.68,16.15,7.68,4.17,2.37,1.0,0.26999998,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.22999999,8.13,6.47,17.19,12.17,2.9299998,4.49,4.91,0.52,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.28,2.82,6.0099998,9.2,16.789999,19.81,12.17,10.54,6.31,2.8,1.09,1.39,2.36,1.8499999,0.59,1.41,1.8299999,2.1299999,3.53,3.1799998,2.99,2.9299998,0.78999996,0.24,0.11,0.0,0.02,0.21,0.35,0.07,0.0,0.69,0.68,0.24,0.34,1.28,1.91,0.84,0.39,1.5699999,0.95,1.1999999,1.4,2.57,1.1999999,0.44,0.25,0.59,1.1999999,0.96,0.47,0.65999997,0.45999998,0.52,0.51,0.74,1.18,0.9,0.44,0.11,0.32999998,1.29,1.06,4.2799997,9.78,4.0899997,0.0,0.0,2.09,3.87,2.4099998,0.53999996,0.06,0.0,0.0,0.17999999,0.35,0.19,0.45999998,1.16,3.87,7.3599997,3.11,3.1599998,0.62,0.04,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,6.04,1.41,0.0,0.0,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06,0.14,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.099999994,1.8,3.56,2.2,0.42,0.11,0.06,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.48,0.93,0.82,0.62,0.11,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.48,0.91999996,0.48,0.74,2.31,3.83,4.0,2.62,3.28,6.41,9.03,6.96,1.35,6.2,16.77,23.39,34.25,52.059998,74.9,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.26,0.62,0.48,0.38,0.35999998,0.21,0.28,0.17999999,0.29999998,0.39999998,0.32999998,0.28,0.45999998,0.52,0.62,0.78999996,0.37,1.28,1.65,1.14,2.0,2.97,3.9199998,4.93,6.5699997,8.66,10.309999,11.46,11.849999,9.45,4.63,3.8899999,2.75,2.6799998,4.5499997,6.87,6.5699997,4.4,4.42,6.68,15.73,29.849998,32.25,28.8,21.64,16.23,10.37,6.48,2.44,0.59999996,0.52,2.4299998,1.4599999,0.85999995,0.63,0.37,0.37,0.29999998,0.03,0.0,0.0,0.0,0.0,0.16,0.41,0.28,6.1099997,4.69,5.83,10.41,21.06,15.2,5.73,2.81,0.0,0.0,0.0,0.07,0.66999996,0.64,0.47,0.24,0.099999994,0.01,3.6399999,20.0,23.32,20.9,13.809999,10.58,8.73,2.73,0.85999995,0.69,1.61,1.38,1.4699999,1.3299999,0.32,0.48,0.89,2.3999999,7.0,5.12,3.08,2.52,0.96999997,0.089999996,0.06,0.0,0.0,0.03,0.11,0.07,0.01,0.03,0.19,0.19,0.11,0.01,0.0,0.14999999,0.59,0.22999999,0.56,0.5,0.22,0.099999994,0.099999994,0.0,0.19,0.34,0.14,0.0,0.32999998,0.91999996,0.69,0.42999998,0.26,1.0699999,0.94,0.57,0.32,0.06,0.52,1.3199999,1.5799999,1.5899999,0.75,0.08,0.19999999,0.42,1.6999999,0.48999998,0.08,0.0,0.0,0.0,0.0,0.02,0.28,0.83,1.5,2.25,2.8899999,1.62,4.2799997,3.6499999,0.42,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.6999999,1.77,0.0,0.0,0.01,0.07,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.04,5.17,12.84,5.6099997,1.2099999,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.089999996,0.26999998,0.26,0.07,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.099999994,1.3399999,1.9499999,5.5,11.15,15.94,12.639999,7.52,12.88,11.45,20.05,18.46,12.48,8.54,11.639999,13.759999,28.76,48.73,76.72,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.099999994,0.32,0.7,0.65999997,0.39999998,0.049999997,0.0,0.32999998,0.65999997,0.65,0.55,0.45999998,0.39,1.28,1.0799999,0.64,1.06,0.90999997,1.4,1.43,1.55,2.24,2.8,3.4299998,4.91,7.0899997,9.33,10.9,14.67,18.939999,16.539999,11.259999,5.56,3.78,4.8199997,7.98,10.0199995,9.24,8.639999,9.61,11.66,10.99,12.7699995,10.28,8.45,7.18,7.52,4.5,2.09,1.86,0.69,0.099999994,0.0,0.0,0.0,0.14999999,0.13,0.02,0.0,0.68,4.19,5.0299997,8.22,11.08,8.809999,7.44,6.1099997,1.9499999,1.91,0.45,0.59999996,2.78,4.46,1.66,0.16,0.11,0.65999997,1.9499999,2.03,2.74,1.54,0.78,2.6699998,9.04,35.95,47.629997,30.019999,18.779999,11.95,6.44,4.02,3.26,6.39,10.8,16.56,15.08,9.75,4.48,0.97999996,0.14,0.83,3.1599998,4.3199997,5.2799997,2.73,0.42999998,0.07,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.089999996,0.17999999,0.17999999,0.07,0.19,0.32999998,0.07,0.0,0.0,0.55,0.32,0.03,0.25,0.11,0.16,0.26999998,0.83,0.97999996,0.52,0.089999996,0.11,0.29999998,0.41,0.39999998,0.45,0.34,0.59999996,0.35,0.32999998,0.37,0.56,1.22,2.6699998,0.62,0.12,0.32999998,1.15,0.35999998,0.17999999,0.11,0.0,0.0,0.0,0.049999997,0.42999998,1.38,2.57,3.4499998,4.15,3.51,4.2,5.5299997,2.23,0.13,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.049999997,0.0,1.11,0.0,0.0,0.0,0.02,0.049999997,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,3.6299999,13.0,6.95,1.55,0.04,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.099999994,1.1899999,3.73,5.7799997,5.41,5.33,5.44,6.0299997,11.219999,21.3,19.119999,20.01,31.769999,33.16,31.109999,30.25,32.11,54.5,61.48,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02,0.64,1.26,0.76,0.17999999,0.26,0.52,0.65999997,0.76,1.16,1.3199999,0.96,1.5799999,1.36,0.32999998,1.03,1.86,1.18,1.77,1.54,1.4599999,1.12,1.17,1.23,2.46,3.11,3.07,5.83,10.78,16.41,19.23,17.09,11.99,7.49,3.8999999,5.0499997,8.59,10.099999,9.139999,7.3199997,4.74,4.0699997,7.62,8.49,5.66,5.3199997,2.56,1.63,0.17999999,0.089999996,0.0,0.0,0.0,0.0,0.32999998,0.57,0.0,0.0,0.19999999,3.8799999,9.34,11.49,14.549999,14.36,11.74,20.72,6.15,7.47,0.63,0.22999999,0.96999997,3.1499999,2.34,0.48,1.06,2.6499999,3.8,1.11,1.4399999,0.91999996,0.89,5.62,22.31,44.39,33.32,12.05,10.639999,11.259999,5.4,2.53,1.74,7.71,12.54,17.24,9.74,11.92,5.75,0.82,0.22999999,0.84,5.06,1.9799999,2.23,1.7199999,0.66999996,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.07,0.0,0.0,0.03,0.099999994,0.0,0.049999997,0.14999999,1.09,2.1,1.93,0.38,0.049999997,0.21,0.28,0.83,1.7199999,1.9799999,1.09,0.31,1.36,1.6899999,1.67,0.13,0.049999997,0.9,1.1,1.22,2.26,0.42,0.19999999,10.99,15.98,0.03,0.0,0.0,0.0,0.17999999,0.39,0.0,0.0,0.0,0.13,0.68,2.6799998,4.2599998,5.97,7.0899997,7.96,6.0099998,6.5,5.81,0.61,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.0,0.089999996,0.0,0.0,0.0,0.0,0.049999997,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.76,4.74,6.15,1.8499999,0.11,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.04,0.53,1.5899999,3.47,2.98,2.02,1.75,3.55,9.51,18.71,25.47,27.97,26.08,30.779999,40.86,29.939999,42.27,56.219997,55.789997,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02,0.14999999,0.14999999,0.01,0.0,0.0,0.14999999,2.22,1.9499999,1.7199999,2.1499999,3.1399999,2.59,1.49,0.88,1.5,2.82,4.47,5.64,6.48,7.19,5.02,2.6499999,2.11,2.31,1.76,2.87,2.47,1.52,1.18,1.13,1.4,1.76,1.49,1.1,0.77,1.66,5.08,10.87,14.7,14.66,12.87,6.7999997,3.23,2.61,3.72,4.73,6.0099998,3.8799999,3.09,3.4499998,4.06,4.0299997,3.6399999,3.81,2.32,0.42,0.07,0.0,0.0,0.14999999,0.32999998,0.37,0.81,0.26,0.01,0.88,1.92,1.66,1.4699999,2.6599998,3.9299998,2.81,1.64,0.64,1.43,1.79,1.9799999,1.87,3.4499998,2.8899999,1.0799999,0.95,0.94,1.49,0.37,2.23,5.24,5.22,11.83,31.71,55.69,63.94,55.26,18.59,1.9,5.29,7.5499997,4.6,2.03,6.04,8.75,8.38,5.7999997,4.2599998,4.95,4.2999997,1.87,0.89,4.67,3.22,0.48,0.03,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.099999994,0.0,0.04,0.11,0.45999998,0.7,1.09,0.29,0.0,0.0,0.0,0.11,0.59999996,0.64,0.049999997,0.57,0.96,2.04,3.21,3.05,1.17,0.71999997,1.43,1.28,0.17,0.0,0.0,0.03,3.3999999,1.28,0.0,0.0,0.0,0.0,0.12,0.099999994,0.0,0.0,0.0,0.35,3.03,7.89,10.349999,12.599999,12.559999,11.25,7.97,9.32,3.4199998,0.17999999,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.03,0.0,0.0,0.0,0.0,0.01,0.04,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.12,1.8,3.49,1.3199999,0.13,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.089999996,0.0,0.0,0.0,0.26999998,1.18,5.5299997,9.389999,13.9,8.08,15.009999,19.189999,17.83,28.73,44.93,58.78,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06,0.12,0.01,0.0,0.0,0.0,0.0,4.0099998,5.77,3.84,4.29,6.08,6.2,4.94,2.98,4.06,7.12,12.78,18.83,31.21,37.14,22.619999,10.87,5.39,3.6399999,2.23,2.49,4.65,4.0699997,2.52,1.37,0.74,0.52,0.64,0.42,0.32999998,0.26999998,0.66999996,1.8299999,4.99,6.75,6.23,5.95,2.84,1.15,1.06,2.56,3.07,6.37,4.41,2.75,5.98,8.92,6.19,4.0299997,6.73,5.38,0.59999996,0.0,0.02,0.089999996,0.0,0.26999998,0.26,0.0,0.02,1.14,1.25,0.64,0.55,0.39,1.7199999,2.28,2.1,0.13,0.19999999,0.48999998,3.3799999,6.25,2.8799999,9.33,12.95,4.66,1.14,0.19,0.13,1.16,3.6799998,7.33,16.55,22.72,27.48,42.89,60.91,46.64,11.03,8.65,11.07,10.25,10.25,9.74,5.24,1.05,0.78999996,3.34,10.74,8.28,5.6099997,2.0,3.6499999,2.37,0.71999997,0.03,0.0,0.0,0.0,2.58,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.04,0.049999997,0.16,0.03,0.0,0.0,0.0,0.0,0.03,0.13,0.14,0.26,0.22,0.19,2.22,2.1699998,1.8299999,2.56,1.4399999,0.82,0.61,0.52,0.16,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.26999998,0.0,0.0,0.0,0.0,0.0,1.36,10.139999,17.35,20.529999,23.16,22.26,13.34,11.61,9.389999,1.02,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.03,0.0,0.0,0.0,0.0,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.0,0.0,0.48999998,1.8499999,1.0,0.13,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07,0.19999999,0.93,2.19,4.71,4.93,3.6999998,3.85,6.71,15.87,40.809998,31.67,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.28,0.12,0.07,0.0,0.0,0.049999997,0.24,3.4399998,5.92,5.71,7.3599997,10.36,11.5199995,11.94,10.53,12.54,15.46,23.289999,37.39,50.809998,53.61,40.48,27.33,9.83,4.02,2.36,0.55,0.75,3.53,4.66,2.79,1.74,1.06,1.01,0.78999996,0.41,0.14999999,0.17,0.14,0.34,0.84,2.3999999,2.8899999,3.6899998,4.06,3.22,1.65,1.43,6.33,9.7,7.5899997,8.139999,10.75,13.21,9.01,7.3999996,8.15,3.8,0.24,0.02,0.02,0.0,0.13,0.48999998,0.03,0.0,0.0,0.0,0.04,0.21,2.02,5.5699997,3.4499998,0.28,0.099999994,0.07,0.62,4.9,7.21,2.8999999,8.809999,31.109999,24.619999,4.1,1.18,0.81,1.28,3.85,4.0,7.04,13.03,13.389999,14.849999,22.119999,28.91,18.32,18.31,14.38,12.99,11.05,5.29,5.97,4.7599998,2.22,0.16,2.95,1.8,0.0,0.84999996,1.0,0.16,0.29999998,1.64,0.049999997,2.09,0.38,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.35,0.31,0.0,0.0,0.02,0.0,0.91999996,0.32999998,0.28,0.22999999,0.87,0.58,0.14,1.09,1.1999999,0.71,0.03,0.0,0.02,0.08,0.13,0.0,0.08,0.03,0.0,0.0,0.0,0.0,0.03,3.37,16.08,29.25,39.35,41.0,27.4,14.61,14.15,4.14,0.65999997,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.0,0.11,0.65999997,0.71999997,0.11,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.11,0.14,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.22,0.81,1.3299999,0.96999997,0.03,0.0,1.16,4.25,16.14,16.88,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.04,0.099999994,0.02,0.0,0.03,0.58,0.53,0.16,0.03,0.0,0.08,0.44,1.3299999,4.0899997,8.57,9.75,13.24,20.869999,26.43,28.88,28.68,31.34,35.32,41.32,51.34,56.77,52.67,36.989998,17.13,4.44,1.5799999,1.1999999,0.38,0.26,0.64,3.1299999,4.58,2.9199998,1.77,0.75,0.47,0.51,0.9,1.4599999,1.16,0.7,0.42,0.82,1.1,2.9299998,6.0899997,7.62,6.16,3.84,1.51,3.6699998,10.74,8.95,5.06,6.33,5.02,2.96,2.86,2.26,0.57,0.0,0.25,0.5,0.45,0.0,0.0,0.0,0.45999998,0.0,0.0,1.29,12.12,33.89,18.65,0.55,0.17,0.0,0.13,0.58,1.55,0.76,2.1699998,15.92,10.4,3.26,0.59,0.07,1.24,8.12,6.02,4.7999997,9.78,14.99,13.11,15.28,16.779999,16.789999,20.22,26.93,22.06,16.859999,10.11,4.23,0.26999998,0.0,0.0,0.0,0.12,0.16,0.06,0.02,0.0,0.19,1.91,1.3,0.26999998,0.08,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.29,0.14,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.26,0.48999998,0.34,0.17999999,0.03,0.29,2.1699998,7.56,1.22,0.39999998,0.089999996,0.0,0.0,0.0,0.0,0.0,0.06,3.4199998,24.58,55.28,71.369995,45.51,27.05,17.26,7.43,2.8899999,0.42,0.06,0.089999996,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.0,0.0,0.06,0.19999999,0.04,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.26999998,0.45,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.7,0.34,0.01,0.0,0.0,0.45999998,2.1,4.5,8.82,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02,0.13,0.03,0.0,0.0,0.04,0.14,0.0,0.0,0.04,0.5,1.67,3.77,7.6299996,12.929999,17.0,25.869999,34.579998,41.52,45.5,45.23,50.579998,53.35,57.079998,57.64,50.84,36.52,21.51,10.48,8.429999,4.2799997,1.88,1.1899999,0.72999996,0.98999995,1.41,2.48,3.4299998,3.51,2.37,2.08,1.29,1.14,1.38,1.77,2.18,1.65,2.72,2.49,2.3799999,6.24,4.58,4.98,5.5,3.28,1.12,2.34,5.38,3.27,0.64,0.47,0.11,0.35999998,0.28,0.14,0.049999997,0.06,0.06,0.0,0.0,0.0,0.0,0.0,0.0,0.07,2.3899999,9.29,20.96,15.95,0.53999996,0.03,0.14,0.45999998,0.65,1.42,2.22,3.01,6.48,10.29,5.67,2.31,1.68,2.1599998,4.39,8.01,12.86,11.5199995,9.05,9.139999,12.96,14.38,12.75,12.509999,20.63,26.08,13.12,3.36,2.47,1.3299999,0.88,0.06,0.14,0.42,3.55,3.58,0.81,0.12,0.0,0.08,1.4,0.32,0.07,1.4499999,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.31,0.12,0.35,1.04,1.13,0.26999998,0.0,0.0,0.06,0.16,0.0,0.01,0.01,0.29,0.35999998,0.12,0.06,3.27,10.63,22.75,8.599999,0.049999997,0.099999994,0.0,0.0,0.0,0.0,0.0,0.0,0.099999994,4.5099998,34.239998,62.219997,57.629997,41.92,19.73,4.0299997,2.82,2.4099998,2.83,2.47,0.07,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.02,0.0,0.08,0.35,0.03,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.24,0.42,0.049999997,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.049999997,0.96999997,1.01,0.07,0.0,0.0,0.17999999,1.6899999,3.56,4.74,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08,0.26,0.74,1.01,2.2,6.23,10.66,13.61,16.949999,23.67,35.86,44.489998,44.84,43.32,44.23,43.96,41.7,37.149998,23.51,15.03,10.12,8.28,6.1,3.3,3.55,2.74,1.38,1.62,1.61,1.9699999,2.1399999,2.61,2.9299998,2.52,2.4199998,2.35,2.18,1.65,2.6299999,2.96,2.46,3.4399998,2.72,2.12,4.08,3.74,2.07,0.78,0.51,0.08,1.05,0.9,1.73,0.17,0.0,0.0,0.0,0.0,0.59,0.5,0.17,0.84,0.71999997,0.0,0.0,0.64,4.83,0.32,0.39999998,0.39,1.9499999,0.14,0.16,0.0,0.0,0.08,0.08,0.38,1.66,3.84,7.39,19.17,36.19,11.8,6.7599998,10.45,20.4,45.26,68.369995,60.41,36.309998,13.29,7.1099997,8.309999,11.08,13.4,29.21,44.809998,22.789999,7.6699996,5.02,2.3999999,1.03,0.12,0.39,1.2099999,3.01,13.03,9.04,2.22,0.14999999,0.0,0.0,1.9799999,0.07,0.0,0.14,0.06,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02,0.17999999,0.57,0.42999998,0.13,0.39999998,0.099999994,0.0,0.04,0.01,0.02,0.19999999,0.37,0.17999999,0.0,2.1,11.5199995,4.52,0.03,0.11,0.0,0.0,0.0,0.0,0.0,0.0,0.07,0.14,3.62,24.609999,22.779999,25.269999,12.04,2.22,8.7699995,14.2,14.099999,11.57,1.6999999,0.03,0.04,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07,0.03,0.0,0.0,0.0,0.0,0.04,0.04,0.04,0.07,0.9,0.37,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.35999998,1.3,0.29999998,0.02,0.0,0.01,1.5699999,4.49,4.79,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08,0.26,0.7,0.96,1.76,2.96,6.33,11.969999,14.65,21.63,31.01,39.309998,40.57,42.41,37.11,33.54,24.72,22.39,21.15,18.08,7.2999997,2.6399999,2.84,1.0,0.69,1.4,1.3,0.71999997,0.89,1.52,2.6799998,3.27,3.56,3.6999998,3.56,3.58,4.21,3.6999998,2.9199998,2.56,4.8399997,5.77,5.6299996,2.96,0.88,2.26,3.4099998,1.4699999,0.89,0.19,0.04,0.12,0.04,0.049999997,0.07,0.099999994,0.22,0.24,0.38,0.22,0.11,2.09,6.64,6.24,6.44,2.5,2.27,0.11,0.0,0.0,0.08,0.11,0.0,0.0,0.0,0.0,0.0,0.42999998,1.9599999,13.889999,26.91,38.649998,67.58,69.5,55.329998,40.25,27.66,36.23,61.239998,69.45,53.71,31.66,16.38,11.44,6.98,7.2,26.55,34.76,16.07,6.31,2.21,1.99,0.14,0.0,1.0799999,1.73,2.98,6.5699997,20.68,13.45,3.9399998,0.75,0.44,0.17999999,1.53,0.9,0.07,0.19,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.04,0.089999996,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.08,0.049999997,0.21,0.42,0.22,0.39999998,14.049999,24.8,18.81,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.19999999,1.7099999,0.97999996,3.6999998,7.87,3.8899999,2.1299999,5.35,15.7699995,29.029999,29.3,18.93,14.799999,6.06,1.29,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.11,0.11,0.0,0.0,0.0,0.0,0.04,0.02,0.01,0.01,0.7,0.35999998,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.04,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.099999994,1.04,1.1999999,0.099999994,0.0,0.0,0.63,1.9499999,4.91,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07,0.63,0.82,0.78999996,1.4,2.78,5.83,11.63,19.24,29.89,38.78,36.29,40.09,35.2,22.55,18.64,17.619999,15.299999,11.42,5.0899997,3.1699998,4.72,3.37,1.4599999,0.83,0.81,1.14,1.67,2.24,3.1299999,5.17,8.679999,11.849999,9.2699995,8.42,8.11,6.73,5.8799996,5.93,5.2599998,6.52,5.18,3.55,2.85,0.98999995,0.79999995,0.47,0.81,1.5699999,0.88,0.39999998,0.52,0.099999994,0.099999994,0.099999994,0.51,1.5899999,2.61,5.22,3.47,0.82,1.0799999,2.35,0.58,0.0,0.0,0.049999997,0.48999998,2.9299998,4.06,1.1899999,0.0,0.0,0.0,0.0,0.0,0.06,3.3999999,8.97,31.48,75.39,98.369995,113.049995,142.84,126.27,96.31,42.66,23.92,32.25,49.41,51.16,46.57,38.93,9.099999,6.47,21.93,24.789999,11.58,6.77,1.7199999,0.04,0.02,0.06,0.48,1.7099999,5.2,2.98,4.93,7.54,3.34,1.03,2.34,0.62,0.89,0.59,2.11,1.27,0.53999996,0.28,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.099999994,0.47,0.97999996,1.0699999,0.31,0.0,0.0,0.0,0.0,0.0,0.11,0.25,0.099999994,0.099999994,0.099999994,0.0,5.81,38.649998,37.0,0.0,0.0,0.0,0.0,0.02,0.53999996,0.72999996,0.0,0.79999995,3.49,4.64,1.0799999,0.84,0.75,3.99,24.16,47.59,48.36,27.01,15.599999,20.72,13.98,0.37,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07,0.0,0.0,0.22999999,0.42,0.04,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02,0.48,0.16,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.31,1.14,0.47,0.049999997,0.0,0.0,0.01,0.11,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.44,0.88,0.45,0.39999998,1.16,2.35,3.9199998,7.1299996,12.969999,26.039999,37.27,37.34,42.68,34.86,17.47,14.7,13.88,16.18,16.23,13.349999,9.86,6.0899997,3.49,1.99,0.62,0.14,0.39,0.64,1.06,0.81,3.6899998,5.52,7.25,10.91,12.849999,12.099999,11.0199995,11.71,12.5199995,13.44,9.0199995,6.42,3.97,2.9299998,4.74,5.12,1.93,0.32999998,0.24,1.09,1.77,1.9499999,2.18,0.48999998,0.13,0.14999999,1.49,3.1499999,4.08,3.0,1.26,0.9,4.98,3.59,0.5,1.53,2.54,4.12,9.51,8.51,2.62,0.78999996,0.65,0.04,1.1,0.26,0.52,6.8599997,16.3,24.67,31.439999,46.96,81.79,114.52,136.11,116.57,54.469997,36.61,44.739998,64.86,77.54,83.86,69.409996,25.66,11.8,5.16,8.98,4.5099998,1.7099999,0.089999996,0.74,1.65,2.54,3.3799999,3.1,0.82,1.4499999,1.0799999,2.3,2.7,0.25,2.1299999,0.74,0.049999997,0.0,0.88,1.17,1.64,0.29999998,0.03,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.07,0.12,0.02,0.0,0.21,0.45999998,0.26999998,0.0,0.0,0.0,0.0,0.16,0.28,0.099999994,0.0,0.0,0.0,0.14,8.71,0.0,0.0,0.0,0.0,0.52,2.6399999,4.69,1.0,0.04,1.42,3.9499998,3.05,3.6299999,2.4099998,3.52,15.45,37.44,53.059998,46.719997,23.76,21.189999,35.36,3.54,0.0,0.01,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02,0.049999997,0.0,0.049999997,0.39,0.13,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.049999997,0.0,0.0,0.0,0.47,0.44,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.7,1.25,0.089999996,0.03,0.06,0.56,1.51,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14999999,0.28,0.11,0.049999997,0.089999996,1.1,4.54,14.29,22.38,33.3,54.699997,56.39,77.56,56.199997,29.849998,13.2,19.1,31.689999,50.18,23.859999,6.68,3.1999998,1.4499999,2.11,1.38,0.87,0.55,0.45,0.47,0.87,1.91,4.3199997,4.5,4.04,4.24,5.14,5.47,7.5099998,10.28,13.2,15.45,12.05,7.99,4.0099998,5.58,10.67,8.309999,2.3999999,0.94,0.96999997,1.29,1.8299999,2.11,1.87,2.85,0.77,0.02,0.08,1.61,2.7,3.4199998,2.86,2.6299999,2.3899999,1.09,2.23,2.73,3.1899998,9.2,11.48,5.33,2.46,6.08,11.63,7.3199997,0.0,0.0,1.0799999,8.2,12.059999,7.69,9.22,17.02,28.26,35.12,27.88,14.65,8.59,14.69,34.03,72.99,110.92,117.34,63.079998,27.51,3.56,1.4399999,2.52,0.79999995,1.93,1.3,1.23,6.0499997,15.45,5.97,1.23,1.5799999,13.0199995,7.18,2.08,1.86,0.9,4.75,0.0,1.43,4.0899997,3.8,4.74,2.28,1.13,0.26,0.04,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02,0.12,0.0,0.01,0.099999994,0.03,0.0,0.0,0.0,0.0,0.34,0.17,0.02,0.0,1.35,2.09,0.45,0.0,0.0,0.0,0.0,0.0,0.12,0.22999999,0.07,0.0,0.0,0.0,0.93,0.0,0.0,0.0,0.0,0.35,3.27,6.31,7.68,1.36,1.37,6.7799997,11.07,11.45,12.57,2.95,6.29,13.969999,31.24,36.76,39.48,26.71,44.68,25.34,0.13,0.0,0.04,0.03,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.0,0.0,0.07,0.099999994,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.06,0.0,0.0,0.06,0.44,0.29,0.08,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.17999999,0.66999996,0.82,0.51,0.17999999,0.39999998,1.6999999,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08,0.29999998,0.08,0.0,0.14999999,2.3,14.2699995,26.51,35.559998,53.48,69.97,71.27,37.16,21.77,15.25,20.21,32.25,50.53,21.67,11.34,0.93,1.3,1.4399999,0.77,1.48,2.57,0.52,0.12,0.19999999,0.14999999,0.26999998,0.59,1.18,1.79,0.81,0.57,0.78999996,2.83,5.52,7.7,11.07,5.68,4.2,2.46,3.1499999,5.83,3.4299998,0.75,0.17999999,0.39,0.19,0.049999997,0.16,0.03,0.13,0.0,0.0,0.14999999,0.66999996,3.09,4.8199997,2.58,0.87,1.65,3.25,4.19,3.53,3.03,0.69,4.5499997,6.0299997,3.85,7.0899997,6.87,0.0,0.0,0.0,0.0,0.84,0.28,0.049999997,0.0,0.25,3.6699998,6.15,5.24,4.38,2.75,5.52,22.4,57.079998,68.979996,79.659996,21.35,10.26,1.12,2.99,0.39999998,0.76,0.17999999,2.96,0.83,15.37,9.179999,2.34,1.26,1.49,0.0,0.0,1.75,2.75,1.8199999,6.7599998,6.7999997,6.73,8.11,9.17,11.83,6.98,2.73,0.21,0.0,0.0,0.0,0.0,0.0,0.0,0.06,0.0,0.0,0.14,0.96,0.17,0.0,0.22999999,1.0699999,0.19999999,0.0,0.0,0.0,0.0,0.17,0.03,0.02,0.19999999,0.35999998,0.099999994,0.0,0.0,0.0,0.0,0.0,0.0,0.08,0.14,0.02,0.0,0.0,0.51,0.0,0.0,0.0,0.0,0.0,0.82,4.54,3.9399998,1.37,6.5,12.49,17.449999,18.67,28.22,14.21,6.21,10.12,14.91,23.21,15.48,18.71,41.379997,40.239998,2.26,0.0,0.0,0.049999997,0.0,0.04,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02,0.03,0.01,0.0,0.0,0.0,0.0,0.11,0.26,0.22,0.049999997,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.02,0.29999998,0.78,0.79999995,0.47,0.01,0.77,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.11,0.11,0.39999998,0.17,0.81,1.41,4.98,16.1,25.91,32.26,75.92,72.299995,36.95,21.59,16.44,17.41,16.779999,14.48,9.08,7.7799997,4.5699997,4.21,5.8399997,2.52,2.3899999,2.44,0.82,0.17,0.099999994,0.13,0.26,0.32,0.06,0.07,0.44,0.75,0.42999998,0.85999995,1.53,1.5899999,2.4199998,2.58,1.79,0.74,0.48,0.59999996,2.06,0.04,0.0,0.099999994,0.07,0.14,0.099999994,0.29,0.08,0.0,0.0,0.04,4.06,0.24,0.56,0.28,0.06,0.11,0.39999998,1.12,0.69,1.8399999,1.4,0.35,0.0,0.91999996,3.1799998,1.75,0.71,0.56,0.0,0.26,0.089999996,0.0,0.0,0.0,0.049999997,1.22,3.08,3.58,3.79,1.9499999,1.01,1.86,6.8199997,11.389999,20.24,6.12,2.98,0.53999996,2.11,2.05,0.35999998,0.32999998,2.02,0.68,0.71,1.22,1.3399999,0.58,0.11,0.08,0.58,11.13,21.77,3.75,14.54,18.449999,11.99,21.859999,12.559999,13.9,7.37,3.78,0.19999999,0.0,0.0,0.01,0.08,0.14999999,0.26,0.69,0.099999994,1.25,0.11,1.05,0.26999998,0.0,0.16,1.9699999,1.68,0.12,0.03,0.0,0.32,0.26,0.0,0.14,0.35,0.32999998,0.32999998,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.08,0.049999997,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.61,0.79999995,0.22,0.94,18.96,26.789999,26.82,35.5,34.71,23.699999,21.31,12.98,12.07,7.64,5.0899997,31.689999,44.42,7.69,0.94,0.0,0.0,0.0,0.04,0.089999996,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14,0.71999997,0.34,0.0,0.0,0.0,0.0,0.0,0.01,0.099999994,0.21,0.11,0.01,0.0,0.0,0.0,0.0,0.049999997,0.14999999,0.099999994,0.0,0.12,0.62,1.1,1.2099999,0.81,0.48999998,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.53999996,2.62,8.7699995,16.32,6.67,4.39,18.25,29.119999,39.96,75.24,53.93,37.57,22.25,25.16,21.55,20.0,14.33,3.62,2.22,1.29,1.9,5.1,3.4199998,0.59999996,0.61,0.39999998,0.01,0.0,0.02,0.03,0.11,0.14,0.02,0.0,0.16,0.52,1.13,0.64,1.8199999,0.68,1.0699999,0.31,0.04,0.06,0.04,0.51,0.84999996,1.23,0.19999999,0.0,0.71999997,0.96,2.19,2.77,0.0,0.0,0.0,0.17,0.0,0.22999999,1.26,0.89,0.03,0.02,0.0,0.0,2.35,0.25,1.66,0.0,0.12,0.0,0.19999999,0.42,2.04,0.19,1.16,3.29,0.0,0.0,0.0,0.0,0.21,0.76,3.4499998,5.85,0.44,0.58,0.03,1.73,0.0,0.26,0.88,0.24,2.69,1.1999999,0.83,2.23,0.78999996,1.8299999,4.69,2.12,0.0,0.0,1.42,0.62,0.37,0.82,13.2,24.5,2.59,28.75,33.39,22.24,33.43,16.77,15.21,7.99,1.03,0.0,0.0,0.0,0.099999994,1.3,2.97,1.35,0.69,0.06,0.62,0.45999998,0.21,0.049999997,0.29999998,0.07,0.32,0.90999997,1.29,1.8499999,0.74,1.2099999,0.63,0.01,0.39,0.72999996,0.26999998,0.03,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.02,0.089999996,0.11,0.049999997,0.03,0.099999994,0.0,0.0,3.57,30.05,21.6,27.67,40.62,25.98,26.14,21.55,15.48,4.44,4.39,13.599999,37.92,11.3,1.66,0.69,0.0,0.0,0.0,0.14999999,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02,0.34,1.09,1.56,0.04,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.04,0.02,0.0,0.0,0.0,0.0,0.12,0.47,0.29999998,0.0,0.0,0.07,0.53999996,1.15,1.31,1.09,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.25,2.86,14.889999,21.84,6.37,5.19,19.22,43.44,36.37,36.69,24.15,27.01,24.019999,24.76,27.099998,29.23,25.66,12.55,9.01,5.13,2.61,3.33,3.4399998,1.81,0.62,0.9,1.24,0.47,0.14999999,0.25,0.17,0.08,0.78,0.39999998,0.0,0.64,0.51,0.22999999,0.25,0.52,0.03,0.45999998,0.42,0.01,0.01,0.03,1.5999999,3.7099998,1.9499999,0.35,0.0,0.98999995,0.35999998,2.3799999,1.11,0.32999998,0.13,0.07,0.0,0.049999997,1.67,8.7,8.139999,1.16,0.0,0.0,0.55,0.0,2.8999999,2.57,0.049999997,0.26,0.48,0.42999998,1.26,1.24,0.0,0.68,0.26999998,0.84,3.52,4.37,0.28,0.17999999,2.44,0.62,0.04,0.68,2.3899999,1.7199999,1.28,1.41,0.90999997,0.51,2.11,0.04,0.19999999,1.9699999,3.06,6.04,5.52,2.55,9.62,2.09,1.49,1.12,0.06,3.28,12.099999,21.99,2.03,19.439999,27.0,20.289999,22.6,19.99,22.439999,17.279999,2.3,0.0,0.0,0.0,0.04,1.15,3.62,1.68,0.59,0.9,0.74,0.78999996,0.0,0.22,0.34,0.04,0.0,0.19,1.43,5.58,6.52,4.1,1.27,0.22999999,0.35,0.0,0.0,0.0,0.0,0.08,0.22,0.03,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.22999999,0.37,0.66999996,0.83,0.91999996,0.97999996,0.79999995,0.63,5.44,14.679999,21.59,11.9,20.96,26.26,10.94,16.08,7.73,4.62,6.54,22.39,29.539999,9.01,0.45,1.62,0.16,0.0,0.0,0.099999994,0.099999994,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.099999994,0.65,1.52,0.34,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.11,0.75,0.62,0.0,0.0,0.0,0.04,1.29,1.25,1.24,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.75,12.009999,10.51,1.78,6.96,31.49,58.039997,34.6,29.529999,17.16,12.74,15.25,11.96,15.809999,19.22,13.19,7.54,5.93,3.6499999,2.6,4.08,4.25,6.14,5.0899997,2.4199998,0.71,0.91999996,1.14,0.45999998,0.83,0.59,0.39,0.0,0.0,0.0,0.0,0.06,0.68,2.54,1.26,0.75,2.73,0.47,0.11,0.0,1.15,3.26,5.49,2.61,0.0,0.08,0.06,0.03,0.32,0.0,1.16,0.48,0.11,0.0,0.35999998,3.3999999,11.0,9.13,0.14,0.0,0.0,0.0,0.65,2.9299998,0.07,1.06,0.35,0.0,0.38,1.56,0.65,4.16,3.6799998,7.1299996,7.95,3.73,1.3,0.0,0.37,0.84999996,1.16,2.52,3.1,0.0,1.1899999,6.71,2.0,2.3799999,0.82,1.4,0.0,1.36,3.11,1.54,1.3399999,1.8199999,5.7599998,7.17,7.73,1.16,1.78,10.309999,2.8999999,4.19,6.3599997,12.429999,46.02,35.76,32.75,28.73,30.25,27.72,3.87,0.0,0.0,0.0,0.28,0.89,3.36,4.3199997,1.51,0.35,0.11,0.099999994,0.13,0.14,0.08,0.01,0.19,0.41,1.24,7.1099997,8.97,6.12,1.99,0.22,0.26,0.08,0.0,0.0,0.0,0.14999999,0.26999998,0.17,0.0,0.0,0.02,0.03,0.0,0.25,0.0,0.06,0.21,0.0,0.04,0.31,0.71999997,1.4699999,1.88,2.55,3.04,2.9199998,3.31,15.599999,23.96,13.469999,10.179999,16.33,9.469999,5.96,6.58,1.12,3.08,7.64,25.9,9.73,0.37,0.7,0.099999994,0.22,0.0,0.03,0.13,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.12,0.35,0.29999998,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.84,1.04,0.31,0.0,0.0,0.0,0.29999998,0.02,0.57,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.11,9.5,3.9499998,2.4299998,6.2599998,27.39,43.11,28.609999,13.59,9.76,6.5099998,6.33,6.69,7.48,12.889999,2.77,0.82,1.3399999,3.3,2.97,3.48,4.3399997,5.91,3.6599998,3.1799998,2.6799998,1.02,1.3399999,0.65999997,0.69,0.9,1.1999999,0.72999996,0.11,0.0,0.089999996,2.19,3.3,4.5699997,6.12,1.3199999,3.4399998,1.78,1.9799999,0.03,1.06,2.9199998,4.95,5.33,0.45999998,2.34,1.02,0.0,0.0,0.0,0.65999997,2.4199998,0.68,0.0,0.0,0.78,6.37,8.87,2.11,0.35999998,0.0,0.0,0.01,0.06,0.0,0.0,0.0,0.0,0.0,0.0,0.19999999,1.0799999,3.01,6.45,9.22,3.1699998,3.78,0.59,3.1399999,0.16,0.21,1.26,0.90999997,0.04,0.88,5.64,5.43,5.8799996,5.8399997,1.03,0.31,0.58,0.12,0.02,0.65999997,0.45,3.72,5.48,3.81,10.63,14.33,10.75,2.3899999,29.449999,49.899998,24.46,43.25,33.05,28.5,25.88,35.62,21.449999,3.98,0.0,0.099999994,0.17999999,0.45999998,0.81,1.81,4.46,6.06,0.22999999,0.02,0.02,0.39999998,1.0,0.049999997,0.35999998,0.68,3.25,4.1,4.52,6.46,11.059999,4.8399997,0.31,0.32,0.12,0.0,0.0,0.0,0.0,0.19999999,0.19999999,0.0,0.0,0.03,0.29,0.28,1.26,1.3399999,0.099999994,0.59999996,0.0,0.12,0.35,1.11,1.62,3.03,3.9399998,4.73,5.68,6.0299997,6.87,13.61,10.639999,11.13,13.299999,10.7,6.8199997,3.9499998,3.35,0.91999996,1.22,14.29,10.25,0.39999998,0.13,0.089999996,0.24,0.0,0.02,0.049999997,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.03,0.06,0.11,0.01,0.0,0.0,0.0,0.0,0.0,0.01,0.04,0.04,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02,0.0,0.0,0.0,0.0,0.44,1.39,1.01,0.07,0.0,0.0,0.0,0.0,1.26,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.28,2.5,0.78,2.47,6.5099998,37.7,48.92,39.25,19.699999,11.16,8.5199995,8.92,9.38,3.49,1.2099999,1.05,2.22,5.08,5.7,6.48,7.6499996,5.72,4.2,6.6099997,3.6699998,2.29,1.37,0.94,0.37,0.06,0.26999998,2.29,2.96,1.4,0.21,0.0,0.58,3.51,5.24,6.5699997,3.9099998,1.3,1.12,3.36,0.42,7.39,3.57,4.45,6.0699997,3.1399999,1.1,0.31,0.0,0.0,0.0,0.32999998,1.04,0.74,1.54,0.0,0.0,0.22,1.06,0.06,2.01,0.37,0.04,0.01,0.45999998,1.54,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.32999998,3.03,4.9,0.68,0.0,0.34,0.0,0.11,0.64,4.31,7.87,6.02,4.0699997,6.1099997,4.39,3.4199998,5.99,0.0,6.67,8.5199995,0.04,0.0,0.089999996,0.78,0.85999995,1.0,9.75,27.05,8.5,0.02,11.0199995,40.57,38.129997,49.23,33.95,32.2,28.289999,29.619999,13.95,4.37,0.0,0.04,0.04,1.27,3.47,1.0799999,5.1,9.08,2.6399999,1.54,1.67,1.8,1.2099999,0.38,0.26999998,1.15,2.52,3.53,1.7099999,3.73,11.179999,8.88,0.29999998,0.12,0.049999997,0.0,0.0,0.0,0.0,0.0,0.03,0.0,0.0,0.01,0.29999998,0.94,2.31,11.059999,3.07,1.4,0.03,0.06,0.47,1.7199999,2.8899999,3.74,5.04,6.23,7.5299997,8.71,9.65,10.7,14.889999,17.56,18.89,16.99,12.29,7.85,7.3399997,7.1499996,7.8599997,13.88,4.21,2.69,1.8399999,1.4499999,1.09,0.96,0.06,0.06,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.29,0.35,0.41,0.17999999,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.14,0.22999999,0.049999997,0.0,0.0,0.0,1.48,1.9799999,0.85999995,0.17,0.24,1.3299999,1.61,2.05,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.19999999,7.7799997,2.1499999,0.52,2.96,29.0,44.36,43.98,49.69,34.27,22.24,11.849999,7.46,3.78,0.55,1.49,1.79,2.35,2.69,3.54,3.22,3.72,1.5899999,2.08,3.85,4.89,2.4099998,0.35,0.13,0.0,0.0,1.43,3.1499999,2.1699998,1.01,0.28,0.0,2.51,2.6799998,1.68,2.21,1.43,0.71,1.2099999,1.2099999,12.74,3.25,1.53,3.79,4.36,0.02,0.0,0.02,0.0,0.0,0.28,0.72999996,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.34,0.29,0.22999999,1.3299999,1.6899999,0.5,0.0,0.0,0.0,0.0,0.0,0.04,2.49,5.24,4.74,2.12,0.12,0.0,0.0,0.0,2.9399998,8.45,10.33,5.0,9.059999,7.04,0.28,0.71,5.33,2.84,7.7,19.34,0.94,0.44,0.0,0.0,0.0,3.61,2.62,3.1399999,11.059999,3.6999998,7.7,17.21,40.25,43.989998,42.219997,32.809998,44.73,35.86,13.139999,3.8899999,0.0,0.0,0.0,0.77,2.1599998,1.3,4.16,5.64,4.5299997,7.64,17.01,2.98,1.49,2.1699998,2.24,0.84999996,0.97999996,1.93,1.14,0.62,1.88,5.68,0.38,0.08,0.26,0.049999997,0.0,0.0,0.0,0.0,0.29,0.099999994,0.0,0.0,0.02,0.76,3.0,20.75,23.91,2.71,0.06,2.01,1.8299999,1.16,2.6699998,4.48,6.19,7.7999997,9.63,11.4,12.46,17.199999,21.76,23.75,20.85,20.699999,16.529999,15.179999,17.71,21.46,32.53,42.899998,20.1,8.2,8.37,6.42,4.49,3.9499998,0.84,0.01,0.089999996,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.37,0.47,0.41,0.21,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.099999994,0.14999999,0.06,0.0,0.0,0.45999998,1.25,0.94,0.08,0.29,1.02,2.3899999,2.95,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,3.51,20.949999,3.97,0.19999999,2.12,24.66,54.149998,63.73,46.309998,37.21,25.98,18.72,11.11,4.99,1.35,0.53999996,0.58,0.53999996,1.01,1.5699999,1.28,2.1399999,1.1,0.19,0.96,2.1399999,1.4399999,0.0,0.01,0.0,0.0,0.37,1.22,1.0,0.79999995,1.64,0.72999996,0.08,0.35,0.099999994,0.03,0.9,1.3399999,0.19999999,1.63,4.49,1.26,0.78999996,1.03,1.06,1.37,0.42,0.02,0.02,0.0,0.0,0.35,0.07,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02,0.03,0.14,0.0,0.37,4.0,1.76,0.0,0.0,0.0,0.02,0.0,0.08,1.05,4.8399997,3.9599998,1.88,0.55,0.0,0.0,0.03,2.4299998,2.9099998,0.03,4.25,2.24,0.47,0.78,1.6999999,2.8,2.03,3.02,10.809999,10.71,5.97,0.0,0.0,0.0,0.35,0.29999998,0.07,1.0799999,2.73,4.24,14.049999,36.39,61.5,62.829998,44.75,113.759995,140.56,75.78,4.17,0.089999996,0.0,0.0,0.26,0.84999996,1.3399999,3.49,5.37,7.0099998,21.039999,26.4,9.94,6.8599997,3.9399998,3.31,0.42,0.72999996,1.17,0.65999997,0.08,1.12,2.85,0.84999996,0.19,0.02,0.03,0.0,0.0,0.0,0.02,0.85999995,0.91999996,0.0,0.0,0.0,0.049999997,1.9,11.5,33.309998,21.32,1.8399999,0.45,7.35,3.57,1.3,2.82,6.0099998,8.889999,11.94,20.13,22.279999,25.9,32.18,36.23,28.279999,21.55,21.14,26.789999,24.93,43.1,66.979996,86.299995,70.36,27.859999,11.54,11.82,10.5,6.37,1.9599999,0.0,0.04,0.13,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07,0.29,0.16,0.08,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.02,0.0,0.0,0.14,0.35,0.26999998,0.53999996,2.03,4.5099998,3.77,2.83,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.8399999,8.26,4.35,0.39999998,0.82,10.599999,23.59,34.23,31.019999,27.019999,19.369999,13.73,6.0699997,0.85999995,1.24,0.88,0.22,0.71,0.82,1.12,0.11,0.75,0.96,0.17,0.29999998,0.38,0.0,0.0,0.0,0.0,0.0,0.0,6.71,10.49,19.1,17.42,6.43,1.05,1.18,0.84,0.79999995,3.04,2.3899999,0.58,2.23,3.87,3.87,0.39,3.4299998,6.0899997,3.62,1.92,0.19,0.07,0.0,0.0,0.07,0.14,0.13,0.0,0.03,0.0,0.0,0.0,0.0,0.0,1.9699999,0.42,0.0,0.0,0.22999999,0.06,0.0,0.11,0.07,1.17,0.31,0.0,0.0,0.95,0.06,0.0,0.0,0.0,0.0,0.099999994,0.19999999,0.0,0.17999999,6.6099997,12.44,7.9199996,7.06,6.96,1.0799999,2.44,7.35,14.34,19.8,3.97,0.01,0.0,0.07,0.0,0.95,3.35,3.57,2.26,3.4399998,8.69,37.36,65.52,54.17,53.789997,80.009995,127.229996,75.979996,7.75,0.58,0.0,0.0,0.0,0.06,0.56,2.09,4.0499997,7.02,15.36,19.09,22.07,30.08,8.86,1.9799999,0.65999997,0.56,0.51,0.41,0.28,0.02,3.28,2.87,1.15,0.04,0.06,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,4.68,21.09,19.96,12.57,2.36,1.35,7.64,0.59,0.29,1.81,5.79,9.849999,23.35,47.76,56.059998,54.879997,55.82,41.51,31.98,24.33,31.32,37.23,34.579998,75.59,118.63,127.649994,73.9,14.929999,3.1,4.0699997,3.36,1.67,0.78999996,0.0,0.16,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.17,0.03,0.03,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08,0.57,1.01,2.3899999,6.54,9.42,8.309999,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.22999999,0.61,0.37,0.98999995,0.94,1.05,4.99,28.189999,27.14,21.369999,17.15,15.57,9.86,2.45,1.03,0.35999998,0.59999996,1.68,0.48999998,0.53,0.03,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.56,4.8599997,7.23,1.53,1.1999999,1.12,5.31,12.62,25.14,22.88,5.45,3.04,8.05,9.13,5.68,1.4499999,3.59,5.81,3.1299999,0.64,0.0,0.0,0.0,0.45999998,0.0,0.03,1.4499999,0.049999997,2.08,0.93,0.0,0.089999996,0.07,0.0,3.8799999,2.22,0.0,0.0,0.0,0.0,0.11,1.06,0.98999995,0.14999999,0.44,0.38,0.02,0.07,0.0,0.0,0.0,0.0,0.0,0.0,0.56,2.22,2.1599998,3.78,9.8,11.2,10.96,11.7699995,4.8599997,5.33,5.7599998,14.309999,9.45,2.3799999,0.0,0.06,1.54,1.53,3.9199998,17.06,7.19,3.09,4.8399997,4.14,8.22,17.199999,35.93,80.29,61.85,33.71,72.74,20.4,0.13,0.0,0.0,0.0,0.0,0.08,1.76,4.58,8.4,6.96,16.94,47.559998,53.149998,13.509999,3.1999998,1.1,0.22,0.53999996,3.84,0.51,2.4299998,1.22,9.5199995,3.4199998,0.32,5.75,3.87,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,7.44,16.529999,13.259999,15.74,11.66,5.0499997,0.22999999,0.42,0.56,1.01,5.0899997,11.11,39.219997,85.509995,108.13,76.09,56.89,44.35,38.85,31.26,51.629997,65.67,58.62,115.74,147.79,120.63,38.18,0.79999995,0.03,0.14,0.93,0.06,0.0,0.12,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.37,0.62,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.26,0.95,2.32,7.35,17.23,0.07,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08,0.39999998,0.26999998,0.17,0.06,0.82,4.65,15.7699995,13.41,20.8,31.74,24.99,10.73,3.8,0.29999998,0.03,0.03,0.0,0.0,0.0,0.0,0.07,0.91999996,4.37,9.679999,3.12,0.0,0.0,0.0,0.03,0.02,0.03,0.31,0.65999997,0.69,3.97,1.1999999,2.1499999,10.42,41.489998,65.42,47.45,35.84,22.13,13.099999,2.82,2.4199998,0.47,0.04,0.099999994,0.02,0.0,0.0,0.0,0.0,0.17,0.0,0.07,0.17,0.87,54.03,28.09,4.3399997,0.0,0.31,0.0,0.0,0.25,0.0,0.0,0.0,0.0,0.0,0.29,0.0,0.0,0.59,1.28,0.64,0.39,0.0,0.0,0.0,0.0,0.0,0.0,1.61,6.39,4.72,1.4399999,4.52,4.75,1.13,3.49,4.27,6.0699997,7.85,4.61,1.39,1.62,0.06,0.08,3.51,5.21,7.6499996,31.08,10.88,1.8499999,2.9099998,0.42,1.37,8.139999,16.19,43.29,53.289997,17.32,35.13,10.7699995,0.0,0.0,0.0,0.0,0.0,0.0,0.89,5.02,7.56,5.41,5.22,4.49,13.11,5.58,3.4399998,1.42,1.09,0.22,1.13,0.29,2.04,0.83,6.2799997,3.1899998,0.32,13.299999,9.4,1.4699999,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.76,9.09,9.62,11.53,30.96,32.59,11.86,1.4699999,6.12,22.949999,26.08,13.719999,17.73,49.84,117.7,93.49,51.059998,50.37,43.399998,21.21,37.969997,58.96,93.47,67.89,32.44,105.36,32.01,1.5699999,0.0,0.099999994,0.06,0.0,0.0,0.11,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.88,0.65999997,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.0,0.0,0.0,0.07,1.18,3.1899998,13.62,7.6,3.6699998,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14999999,0.0,0.91999996,5.92,39.09,41.43,35.899998,33.29,18.48,6.8599997,2.6,0.14999999,0.26,0.0,0.0,0.0,0.0,0.0,0.35,2.6299999,6.27,5.62,1.3399999,0.0,0.96,0.77,0.0,0.29,0.48,0.34,1.15,1.31,6.2999997,15.79,15.049999,10.9,18.93,30.269999,23.539999,32.469997,27.21,23.73,7.08,0.45999998,2.6299999,0.14,0.03,0.03,0.0,0.90999997,0.53999996,0.19,0.099999994,1.63,10.5199995,2.29,0.69,54.62,59.079998,10.559999,0.22,0.11,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.22999999,0.0,0.0,0.26,0.049999997,0.049999997,0.02,0.0,0.0,0.16,0.22,0.0,0.0,1.4,0.26999998,4.41,5.9,4.16,2.6799998,2.22,0.17,0.61,2.26,0.45999998,0.7,2.35,0.77,0.94,3.02,8.139999,6.66,28.84,9.98,0.81,1.01,1.9799999,5.02,11.61,9.969999,18.699999,49.059998,20.65,36.55,11.88,0.0,0.0,0.0,0.0,0.0,0.0,0.48999998,2.56,5.54,6.81,5.99,6.66,4.94,3.6499999,3.1499999,1.9499999,1.61,0.47,0.12,0.55,0.38,16.65,31.82,3.47,1.53,26.75,31.47,36.45,19.17,0.06,2.72,1.2099999,0.0,0.0,0.0,0.0,0.47,3.7099998,2.71,4.48,7.6299996,3.26,10.48,21.68,26.8,14.049999,6.22,27.22,35.55,35.79,26.939999,21.17,68.06,76.13,51.71,41.93,40.579998,24.609999,18.02,30.4,56.02,42.21,9.07,17.21,4.4,1.31,0.0,0.07,0.03,0.03,0.01,0.099999994,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.32999998,1.13,0.41,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02,0.24,0.099999994,0.0,0.0,0.0,0.78999996,1.5,4.89,32.239998,3.05,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.049999997,0.04,0.37,0.29999998,0.08,0.08,0.01,0.07,0.0,3.21,0.19999999,1.64,2.03,0.68,1.64,2.99,22.93,27.019999,17.16,11.03,5.23,3.35,1.22,0.24,0.17,0.0,0.11,0.48,0.03,0.0,0.06,0.0,0.04,0.0,0.0,0.93,1.48,1.86,2.96,4.72,6.2999997,3.83,3.24,5.6299996,9.01,10.48,8.2,6.6299996,23.3,37.79,32.11,24.3,38.69,36.329998,18.5,3.9599998,3.55,1.64,0.08,0.45,6.04,7.0699997,4.98,2.33,2.36,1.8199999,13.509999,3.7099998,0.32999998,3.21,5.8799996,2.1699998,4.5,1.4,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.049999997,0.0,0.14999999,0.0,0.0,0.02,0.48,0.07,0.76,1.3199999,0.0,0.0,0.0,1.74,3.8,5.69,2.1499999,4.5699997,1.5899999,0.0,0.0,0.0,0.79999995,3.8899999,7.0899997,1.86,2.4199998,1.3399999,2.07,4.36,6.0299997,1.5799999,0.0,0.19999999,5.83,10.94,5.5699997,2.78,2.8,6.98,15.849999,9.67,3.29,0.0,0.0,0.59,2.71,0.39999998,0.0,0.16,1.27,2.96,6.18,20.99,28.51,14.599999,8.679999,6.5299997,2.0,1.78,0.78999996,0.14,0.0,0.34,27.3,67.84,3.1799998,0.55,14.0199995,36.41,58.89,14.929999,1.16,5.0899997,4.11,1.48,0.64,0.0,0.0,0.37,5.0099998,13.139999,15.53,4.77,6.56,5.65,5.31,11.86,19.89,16.359999,21.949999,31.359999,24.6,15.639999,12.45,25.189999,34.149998,35.87,43.12,43.53,18.34,3.4299998,13.03,33.489998,48.289997,6.18,0.95,0.31,2.6399999,0.0,0.07,0.03,0.03,0.04,0.07,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.02,0.45,1.23,1.15,0.45,0.0,0.08,0.08,0.25,0.06,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02,0.19,0.72999996,0.34,0.0,0.0,0.0,0.56,1.55,2.98,0.0,0.03,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.65999997,1.31,2.57,3.1,4.18,3.6799998,6.33,18.91,9.36,19.4,4.63,0.0,0.35,10.04,15.17,5.64,29.99,11.24,1.92,4.15,3.85,0.53,0.04,0.0,0.31,0.0,0.0,0.0,0.0,1.37,1.36,0.84,0.089999996,0.0,0.0,0.0,0.14,0.52,3.04,3.08,8.15,15.75,15.44,9.4,6.58,11.42,9.07,1.89,0.77,3.5,16.07,47.579998,33.16,33.43,27.83,13.29,6.99,0.88,1.27,0.0,0.03,3.4299998,7.81,3.1999998,1.15,1.13,3.1799998,0.0,0.26,0.11,0.0,1.0799999,10.29,4.67,7.56,1.1899999,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.19,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.5,0.71999997,1.03,0.79999995,0.26,0.71,0.0,0.0,0.0,0.0,0.0,1.6999999,7.3599997,1.92,2.82,3.32,0.75,4.98,3.4099998,0.48,0.21,0.62,5.85,7.35,2.33,3.52,2.3799999,0.0,0.0,0.51,0.45,1.14,0.17,0.0,5.1,3.46,0.0,0.0,0.06,2.46,15.7699995,36.02,60.0,37.78,23.199999,9.92,3.0,0.85999995,1.03,0.97999996,1.31,3.4399998,14.969999,33.16,1.62,0.26999998,12.2,16.52,19.939999,9.19,4.8399997,11.2,17.199999,4.5699997,1.53,0.02,0.0,1.63,6.96,18.41,42.309998,23.359999,6.14,10.889999,25.369999,11.04,7.3399997,11.469999,22.109999,22.49,11.849999,4.13,7.6299996,12.79,11.98,17.72,23.51,22.519999,9.139999,4.31,1.78,14.17,22.25,5.0699997,1.7199999,6.3399997,8.34,6.2,0.04,0.01,0.48,0.049999997,0.06,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.19,0.63,2.51,2.1,1.67,0.89,0.39999998,0.38,0.57,0.55,0.06,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07,0.14,0.65999997,1.06,0.59999996,0.03,0.0,0.0,0.26,1.03,1.38,1.1999999,1.1899999,0.12,0.11,0.79999995,2.07,2.22,2.86,4.77,4.58,14.7,23.75,45.129997,31.51,12.38,9.469999,24.25,22.59,23.109999,47.18,13.5,1.5899999,6.1,40.579998,34.87,29.789999,49.629997,25.09,9.99,4.45,5.44,0.17,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.48,1.68,2.6599998,8.74,10.04,4.2799997,0.57,0.21,2.47,8.349999,16.31,12.79,13.179999,9.61,5.5299997,2.74,4.0499997,2.36,0.71999997,0.31,0.37,2.86,14.13,16.96,12.04,4.91,2.4099998,6.33,14.19,12.42,4.47,6.06,6.5899997,2.29,1.0799999,8.99,23.57,15.03,6.5499997,1.22,0.0,0.0,1.7199999,1.4599999,12.08,2.78,1.15,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.07,0.0,0.0,0.0,0.0,0.29999998,0.0,0.0,0.01,0.049999997,0.24,0.07,0.0,0.0,0.0,0.14,0.19,0.0,0.0,0.0,0.48999998,0.13,0.19999999,0.099999994,0.0,0.0,0.0,1.49,1.87,1.31,2.87,1.3299999,6.04,6.6499996,3.4299998,1.7099999,1.88,6.17,4.69,1.78,1.66,0.099999994,0.0,0.12,6.92,17.21,50.559998,4.9,0.0,1.03,13.42,17.94,9.2699995,4.0,17.3,28.21,50.64,60.48,48.84,34.27,12.679999,4.1,1.66,2.52,4.25,13.73,19.57,11.0,5.22,0.48,1.8499999,10.17,10.76,14.07,16.91,15.889999,30.39,50.09,16.789999,4.75,1.78,0.41,1.29,11.98,16.58,36.71,56.28,41.95,21.85,13.429999,23.56,28.029999,15.469999,14.429999,21.98,14.309999,7.5699997,11.3,16.699999,27.88,16.69,12.25,8.73,6.1299996,18.88,6.46,2.4199998,5.0099998,3.82,10.0,18.039999,19.31,16.09,13.57,4.08,2.24,1.67,0.06,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.42999998,1.48,3.46,3.12,2.02,1.7199999,0.79999995,0.31,0.28,0.95,4.5299997,6.08,3.22,2.22,1.56,1.01,0.96999997,0.85999995,0.28,0.06,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.04,0.04,0.049999997,0.16,0.26999998,0.9,1.1899999,0.94,0.38,0.01,0.0,1.3299999,0.32999998,0.22,0.28,0.82,0.22999999,5.16,15.23,20.75,14.91,20.619999,25.33,40.17,48.28,88.36,94.509995,39.43,17.46,8.33,24.13,21.01,25.57,26.74,4.7999997,3.6999998,24.5,61.129997,42.82,33.91,40.309998,29.529999,10.05,2.34,1.11,0.0,0.01,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14,0.32999998,2.09,1.67,1.55,2.6,3.47,6.97,21.46,18.83,19.07,11.74,6.6499996,4.36,9.309999,5.04,3.08,1.0,0.07,1.92,9.0,13.65,12.33,3.6899998,0.68,0.75,0.0,0.0,8.26,9.33,4.99,9.95,9.8,19.699999,25.32,24.68,8.09,2.47,0.0,0.0,5.14,0.47,1.52,2.46,4.65,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.78,0.0,0.0,0.0,0.04,0.88,0.29999998,0.0,0.28,1.03,0.59999996,0.21,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.22999999,0.13,0.0,0.0,0.0,0.0,1.6899999,0.87,1.67,1.5899999,5.17,7.25,7.71,3.6299999,1.81,3.1699998,1.79,1.9599999,9.04,1.7099999,0.17,0.06,0.65999997,25.67,99.909996,11.349999,0.0,0.19999999,7.17,8.7699995,4.35,16.109999,38.09,39.6,56.62,58.85,46.079998,23.15,10.96,4.95,2.57,2.07,5.87,30.789999,45.77,21.99,4.8399997,0.0,3.9599998,15.389999,15.23,20.91,24.65,31.519999,45.61,82.54,43.41,22.519999,6.0,1.68,1.67,8.19,22.619999,36.719997,53.449997,69.58,78.09,40.2,23.22,21.279999,33.11,21.439999,16.91,14.53,13.17,17.67,27.539999,35.059998,34.84,17.46,6.1,6.8599997,27.5,19.779999,4.98,12.5199995,16.96,32.899998,39.28,29.769999,27.23,30.84,13.17,2.9299998,2.96,0.06,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.96999997,3.84,9.179999,11.45,10.0,9.78,7.94,5.56,2.7,2.08,5.52,10.24,7.18,3.58,4.9,6.0299997,4.44,2.57,1.25,0.65999997,0.07,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.19,0.19999999,0.29999998,0.53,0.89,1.31,1.29,1.55,0.65,0.12,0.14999999,0.0,0.0,0.0,0.14999999,2.8799999,15.44,47.559998,48.629997,31.019999,55.11,75.57,116.579994,90.2,71.299995,65.689995,23.83,15.679999,7.95,21.27,22.46,26.81,15.04,3.4199998,6.95,17.72,30.539999,29.57,24.25,22.769999,24.07,19.99,6.21,1.28,0.5,0.26999998,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07,0.02,0.95,3.1999998,5.48,8.67,6.35,3.8799999,2.08,2.4099998,8.7699995,9.059999,7.77,9.8,9.34,6.92,3.78,4.1,4.49,7.91,9.2,10.7,10.04,4.12,0.01,0.0,0.0,0.04,3.4199998,3.73,0.22,1.11,2.4199998,11.809999,9.3,9.42,1.02,0.17999999,0.06,0.0,0.03,2.51,5.1,0.0,10.98,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.19,0.0,0.11,0.83,0.22999999,0.0,0.049999997,0.0,0.0,0.099999994,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.98999995,1.4399999,1.04,1.0799999,1.04,5.3599997,3.46,6.5099998,2.3,0.049999997,0.0,2.72,8.72,3.33,1.65,0.39,0.0,2.85,13.139999,5.72,1.6899999,0.0,0.19999999,3.31,6.91,12.0,25.599998,40.84,45.489998,47.3,35.66,19.699999,7.2,1.8199999,1.78,8.37,4.71,9.99,17.5,15.53,8.12,2.8999999,6.17,30.67,28.06,27.09,46.26,77.119995,87.22,82.04,53.39,41.86,26.859999,12.4,5.44,6.37,19.64,43.29,58.05,74.93,90.27,85.06,45.719997,20.47,9.679999,12.73,26.76,24.939999,21.109999,26.539999,38.42,54.02,70.229996,40.18,13.469999,10.29,34.93,59.37,29.66,6.19,23.289999,37.86,42.44,28.65,15.639999,7.5099998,0.95,0.59999996,0.78,0.03,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.39999998,1.48,2.96,3.76,4.0699997,4.42,4.79,4.46,4.19,4.7,5.85,14.49,14.74,8.309999,6.73,12.559999,12.9,5.42,3.26,1.74,0.78,0.14999999,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13,0.39999998,0.51,0.71,0.90999997,1.17,1.5799999,2.76,2.28,2.34,0.88,0.65,0.19,0.0,0.0,4.7599998,13.429999,54.53,46.53,27.16,55.26,76.96,136.23999,95.579994,56.27,53.42,32.91,12.799999,8.32,17.529999,17.1,10.889999,0.53,0.76,2.61,6.3199997,14.759999,19.64,12.0,11.889999,15.42,6.92,2.22,0.06,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.17,1.24,3.05,4.15,3.8999999,5.31,4.5499997,2.45,3.6699998,4.83,2.34,1.43,4.3399997,3.57,4.5499997,2.48,1.8199999,8.139999,9.37,9.28,6.17,2.72,0.099999994,0.53,0.5,0.02,0.0,0.089999996,0.7,0.06,0.0,0.06,0.02,0.0,0.0,2.82,2.28,0.0,0.0,0.099999994,0.44,0.0,0.84,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.95,0.19999999,0.06,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.04,0.22,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.34,0.0,0.56,1.16,0.21,0.29,0.78,2.49,4.5699997,0.79999995,0.0,0.0,0.19999999,0.68,0.85999995,0.84,0.089999996,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.16,2.02,7.44,21.9,32.93,40.41,42.53,25.25,11.719999,3.24,1.28,1.6999999,11.679999,2.01,2.76,8.74,12.87,8.599999,9.599999,35.37,43.2,35.57,53.649998,101.67,121.56,129.26,86.67,55.8,55.0,72.2,56.449997,22.32,16.09,16.89,37.69,70.11,93.479996,93.6,80.83,64.75,51.25,20.609999,7.56,9.45,17.18,23.5,37.26,52.66,72.72,120.409996,95.67,34.32,21.47,39.04,49.34,49.78,10.48,19.64,27.08,45.629997,42.5,11.42,1.16,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.16,0.53999996,0.59999996,0.61,0.89,0.94,1.0699999,1.3,3.1499999,6.73,17.77,17.02,10.2699995,12.07,14.889999,8.75,4.2,3.01,1.6899999,0.53,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02,0.35,0.87,0.98999995,1.0799999,1.17,1.0,1.17,1.4599999,5.0899997,3.35,2.6399999,1.38,0.0,0.01,4.0899997,11.639999,33.13,32.68,31.55,45.68,57.539997,82.2,53.61,50.67,52.16,32.969997,13.41,14.49,19.67,5.31,1.5899999,0.71999997,1.43,4.25,3.74,5.64,11.559999,13.219999,8.88,5.6,3.1499999,0.52,0.21,0.04,0.02,0.0,0.0,0.0,0.0,0.01,0.089999996,0.29,0.37,0.44,0.53,0.91999996,1.3,1.8199999,2.6499999,2.28,5.87,10.07,7.5699997,4.5699997,1.9699999,0.5,0.42999998,0.55,2.01,2.1699998,3.07,5.58,8.0,7.77,4.5699997,3.26,1.8199999,1.04,0.59,0.26999998,0.089999996,0.0,0.0,0.13,0.089999996,0.0,0.0,0.0,0.0,0.0,1.1999999,1.04,0.31,0.19999999,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.28,1.99,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.14999999,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.87,0.29999998,0.03,0.87,0.41,0.0,0.0,0.089999996,0.32999998,0.0,0.0,0.0,0.0,0.0,0.17999999,0.13,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.25,2.72,8.08,16.25,26.99,24.66,11.69,2.02,0.19999999,0.45,0.06,0.22999999,0.9,4.17,17.58,33.82,20.58,14.17,17.949999,12.95,13.48,48.34,83.0,105.42,112.32,85.09,61.329998,69.25,114.18,110.96,51.469997,57.94,52.23,36.12,61.699997,115.13,94.21,70.27,48.96,43.25,55.219997,39.93,8.61,11.62,29.519999,51.0,78.45,105.729996,146.25,143.55,80.09,35.94,36.76,28.41,18.84,4.66,16.24,29.08,50.95,67.67,20.01,0.56,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.089999996,0.11,0.29999998,1.5,4.6,15.299999,12.719999,9.349999,10.03,8.24,3.82,4.31,4.1,2.1299999,0.52,0.13,0.06,0.0,0.0,0.0,0.0,0.0,0.0,0.099999994,0.78999996,1.27,1.55,1.4399999,1.25,1.03,1.15,1.89,2.82,2.53,2.31,0.02,0.17,3.23,22.029999,21.15,30.17,51.62,37.04,35.63,36.059998,19.35,24.08,31.49,27.439999,20.279999,19.66,21.98,4.27,1.88,2.1499999,4.04,1.87,0.25,0.69,2.58,3.4299998,2.09,0.21,0.44,0.03,0.03,0.0,0.64,0.47,0.0,0.0,0.13,0.96999997,2.05,3.22,3.49,2.21,1.93,4.0099998,3.3899999,4.31,4.2799997,4.41,5.2599998,5.17,3.6,2.21,1.01,0.12,0.0,0.17,7.3599997,4.31,4.2799997,2.59,1.9,2.12,3.12,4.36,2.4099998,1.36,0.7,0.12,0.0,0.0,0.44,3.3799999,7.3599997,0.88,0.0,0.0,0.0,0.0,3.74,5.54,0.9,0.78,0.74,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.17,0.84,0.29,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.53999996,0.04,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.58,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.24,8.96,16.619999,9.639999,1.22,0.0,0.07,0.0,0.0,0.26999998,0.53999996,5.8199997,18.89,18.33,6.31,7.49,13.96,11.349999,7.89,3.9099998,5.62,15.5,39.96,56.85,47.05,42.07,63.489998,77.03,54.8,69.15,69.35,38.6,51.82,87.229996,103.18,65.97,40.899998,27.92,30.859999,19.49,37.57,30.109999,59.98,79.29,112.34,114.39,121.329994,137.45,119.909996,62.68,68.159996,59.19,34.68,10.25,45.39,45.46,24.96,28.949999,3.55,0.089999996,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.81,2.62,8.49,9.42,7.46,6.79,4.13,4.06,5.54,4.93,3.04,1.0,0.65,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.29999998,1.7199999,2.03,1.79,1.67,1.15,0.62,0.9,1.38,1.81,1.67,0.78999996,1.13,2.23,31.26,26.48,35.2,40.28,14.0,9.41,9.49,4.04,12.83,16.09,18.23,26.98,24.26,24.4,6.12,1.1,1.49,1.18,0.26999998,0.01,0.0,0.0,0.03,0.07,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.31,0.75,1.09,1.76,2.0,3.74,7.06,10.54,9.96,3.1799998,2.12,1.39,1.42,0.84,0.79999995,0.28,0.0,0.0,0.0,0.17999999,1.9699999,2.18,6.77,7.5099998,9.599999,5.7599998,4.5,2.51,3.1499999,5.64,6.7799997,5.06,2.6,0.62,3.1399999,3.56,0.45999998,0.56,0.0,0.0,0.01,1.62,6.75,5.25,1.22,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.03,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.37,5.5499997,17.24,8.26,0.35999998,0.14,0.53,0.08,0.03,0.19999999,2.22,4.64,3.52,2.44,1.8,24.029999,25.66,4.5699997,1.7099999,1.6999999,3.12,31.8,57.16,46.82,46.17,37.62,24.48,32.219997,30.369999,18.97,19.15,28.359999,75.4,110.79,119.159996,67.729996,27.189999,7.7999997,13.67,14.75,23.14,28.63,55.77,83.65,107.85,106.119995,106.22,106.579994,101.939995,70.58,94.1,74.15,48.02,18.55,49.94,86.75,33.079998,2.1299999,0.56,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08,0.79999995,1.51,7.9199996,7.5299997,6.0499997,3.57,3.4399998,4.9,5.92,6.79,3.8899999,2.1299999,1.06,0.0,0.0,0.0,0.0,0.0,0.0,0.04,1.3,1.9799999,1.9399999,1.89,1.3,0.16,0.31,1.05,1.4399999,1.1999999,2.8899999,3.36,17.6,27.42,2.6,4.75,2.84,0.55,0.89,1.43,0.24,0.51,2.02,3.86,9.849999,15.849999,13.92,4.97,1.06,0.47,0.01,0.29999998,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08,0.01,0.0,0.02,0.32,1.3299999,5.02,11.87,9.32,2.1,0.93,0.26,0.61,0.71,0.83,1.52,1.13,0.11,0.29999998,6.47,8.13,10.71,10.98,9.099999,9.59,6.98,4.35,2.97,2.4199998,0.98999995,0.71,0.44,0.25,1.5699999,10.17,9.63,4.0099998,4.3399997,1.68,0.19999999,0.06,2.3999999,14.28,10.37,3.84,0.28,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.17,1.1999999,2.61,0.24,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.16,1.0799999,0.14999999,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.5699999,11.13,7.83,2.72,0.56,0.0,0.089999996,0.03,0.02,6.1,13.58,10.7699995,5.91,1.4699999,8.28,9.639999,0.95,1.4399999,8.9,17.99,42.44,54.649998,36.87,27.64,14.75,8.36,5.1099997,1.81,6.14,11.969999,42.82,91.71,125.96,116.439995,64.07,42.02,7.95,43.68,31.72,30.96,66.189995,50.07,77.689995,107.79,126.63,86.159996,63.719997,62.92,82.17,104.149994,39.18,45.32,26.189999,20.619999,64.049995,15.17,0.82,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.099999994,0.56,1.51,6.6099997,5.49,2.1699998,1.76,3.31,4.8399997,5.75,9.679999,6.5899997,2.31,0.65,0.0,0.0,0.0,0.0,0.0,0.0,0.65,1.9399999,2.04,1.93,1.5799999,0.14,0.0,0.13,0.11,0.16,4.99,4.72,5.96,2.4199998,0.11,0.0,0.0,0.0,0.0,0.0,2.1399999,3.49,5.6099997,3.3899999,3.9399998,7.5299997,10.53,7.14,1.7099999,0.14999999,0.19999999,0.71,0.71,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.34,0.55,0.17,0.48999998,1.1,0.48,0.44,0.63,0.34,0.03,0.29,0.22,0.14999999,0.07,0.0,0.03,0.03,0.37,0.51,3.74,7.8599997,12.44,12.509999,8.37,9.61,9.69,6.1299996,6.49,4.5699997,2.78,1.29,0.03,0.0,0.75,1.27,1.02,2.95,2.18,0.48,3.26,3.46,2.03,0.32,0.66999996,4.62,3.01,1.04,0.14,0.0,0.06,0.19,0.13,0.0,0.02,0.53,0.29,0.03,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.32999998,1.22,3.82,1.63,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.41,2.85,0.83,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.19999999,3.55,4.77,0.97999996,0.17999999,0.0,1.65,0.7,0.01,11.16,30.0,5.5,4.18,5.39,9.21,8.0,0.74,1.3299999,15.2,19.39,9.2699995,10.59,29.019999,46.219997,5.14,0.19999999,0.51,6.7999997,22.68,38.69,76.85,152.34,174.4,119.17,53.17,65.799995,31.76,21.689999,29.82,34.969997,64.979996,62.25,77.009995,113.31,111.38,55.11,39.27,36.53,54.0,62.55,34.62,52.219997,28.599998,10.99,1.5799999,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.41,0.88,3.87,1.9799999,1.02,1.17,2.28,3.76,6.44,9.54,3.58,1.78,0.38,0.01,0.0,0.0,0.0,0.0,0.22,1.64,2.03,1.8299999,1.53,0.45,0.0,0.0,0.0,0.0,2.86,2.96,2.21,0.0,0.0,0.0,0.0,0.0,0.0,1.17,17.58,27.22,18.15,6.71,4.95,5.71,2.48,1.05,0.68,0.099999994,0.42999998,0.9,1.3,0.0,0.0,0.0,0.0,0.0,0.0,0.04,0.13,0.19,0.099999994,0.02,0.19999999,0.53999996,0.19,3.02,5.75,0.84999996,0.87,1.92,2.08,2.71,0.57,0.01,0.0,0.03,0.26,0.89,0.19,0.089999996,0.75,2.1299999,3.1799998,2.78,3.35,5.74,11.86,14.559999,15.78,11.98,5.58,1.89,0.32999998,0.049999997,0.45999998,2.62,2.23,0.56,1.3199999,0.68,0.0,0.0,1.6999999,1.48,0.099999994,0.099999994,0.74,0.45999998,0.19999999,0.01,0.0,0.14,0.22,0.06,3.31,7.3599997,9.59,7.2,2.51,0.049999997,0.0,0.0,0.0,0.0,0.0,0.04,0.29999998,0.64,4.5899997,2.52,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.099999994,0.08,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06,0.04,0.22999999,0.14,0.01,4.7,8.87,9.9,0.90999997,14.95,48.09,3.6899998,12.74,8.36,4.35,0.42,2.77,4.5899997,11.639999,5.7,4.0099998,11.84,5.0299997,6.27,13.429999,16.119999,11.179999,22.269999,61.079998,55.07,71.88,70.439995,91.57,40.43,20.539999,90.29,71.72,57.28,89.79,86.159996,52.18,58.34,70.38,81.84,55.379997,29.65,30.099998,29.369999,28.67,48.77,72.78,31.09,8.26,1.06,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.03,0.03,0.03,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.29999998,0.61,1.0799999,0.7,0.77,0.94,1.4599999,4.0499997,5.73,6.81,3.47,1.38,0.22999999,0.01,0.0,0.0,0.0,0.0,1.1,1.5799999,1.5699999,1.26,0.71,0.0,0.0,0.0,0.0,0.35,0.13,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.35,10.95,20.46,23.699999,16.039999,8.099999,3.9299998,0.97999996,0.06,0.0,0.06,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13,0.58,1.27,1.75,0.84,0.11,0.0,0.21,0.64,0.42,1.42,0.44,0.12,0.14,0.099999994,0.14,0.17,0.02,0.0,0.07,0.55,0.63,0.31,1.66,1.65,1.9599999,3.98,2.1599998,0.55,6.0499997,8.29,6.8599997,7.04,5.95,3.97,2.1,1.22,0.31,0.01,0.26999998,0.61,0.78999996,0.79999995,0.07,0.0,0.0,1.91,3.9099998,0.66999996,0.03,2.77,2.1699998,2.07,0.14999999,4.0499997,2.87,0.06,0.0,16.449999,32.36,24.05,21.539999,9.26,2.19,3.04,0.38,0.03,0.14999999,0.0,0.0,0.0,0.0,0.22999999,0.089999996,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.32999998,0.08,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.9,0.9,0.0,4.8199997,12.92,29.89,13.67,0.03,5.45,2.37,15.839999,12.849999,0.64,0.02,1.31,24.07,29.82,20.789999,11.19,1.63,4.4,18.41,66.47,86.009995,34.66,39.67,36.51,10.87,19.05,37.61,11.469999,3.34,8.66,55.77,48.34,116.52,138.48999,132.26,47.16,34.53,41.64,63.629997,38.84,43.92,45.899998,30.869999,27.05,33.69,31.46,51.26,12.389999,0.08,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.03,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02,0.099999994,0.02,0.28,0.35999998,0.45,0.39999998,0.69,2.85,2.48,5.5,2.48,1.1899999,0.099999994,0.02,0.0,0.0,0.0,0.47,1.1,1.2099999,1.15,0.85999995,0.04,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.28,9.28,18.41,22.58,20.67,10.13,2.6,0.32999998,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.35,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.25,1.1999999,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.049999997,0.5,0.97999996,1.1999999,2.61,4.5,7.54,7.7799997,3.21,0.13,0.03,0.099999994,0.77,0.72999996,0.38,0.48999998,0.42999998,0.88,0.88,0.44,2.46,2.86,5.87,2.09,0.91999996,0.02,0.0,0.17,1.68,3.6999998,5.83,4.52,4.85,4.0099998,0.02,0.07,0.0,0.0,3.26,11.36,37.649998,36.219997,38.92,26.14,21.23,12.38,15.54,9.23,5.31,4.42,1.75,0.06,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.04,0.76,1.16,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14,1.79,29.22,27.56,56.899998,110.39,4.45,3.05,12.84,21.67,10.309999,0.47,1.1999999,29.73,58.539997,38.61,17.27,9.389999,24.14,8.809999,19.289999,24.42,46.28,26.05,42.93,53.89,22.67,2.56,31.13,17.51,0.79999995,0.51,5.16,43.02,98.159996,83.61,69.689995,38.26,23.35,31.84,32.98,51.899998,71.52,66.77,41.239998,20.949999,34.94,37.8,10.87,3.08,0.38,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02,0.04,0.03,0.01,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.19,0.22999999,0.14,0.099999994,0.7,1.66,2.18,2.6699998,1.76,0.44,0.02,0.0,0.0,0.0,0.03,0.35,0.29999998,0.91999996,0.9,0.13,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08,2.32,8.059999,12.19,14.2,10.48,5.8599997,1.87,0.62,1.5699999,0.47,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.099999994,0.72999996,0.32,0.01,0.0,0.51,1.3299999,4.3399997,5.15,8.66,10.7,14.61,17.19,10.219999,5.35,2.3999999,0.39999998,0.0,0.0,0.0,0.22999999,1.51,1.05,1.81,6.3399997,7.22,5.14,2.71,1.51,0.13,0.0,0.0,0.83,2.9299998,5.44,3.08,0.17999999,0.32,0.35,0.0,0.0,2.29,4.11,12.219999,42.149998,49.469997,49.469997,31.779999,26.92,14.12,20.16,20.48,10.389999,9.09,5.37,1.09,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.59,1.5999999,3.32,0.47,0.0,0.0,0.0,0.0,0.0,0.44,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,23.32,24.019999,39.1,60.16,27.47,31.689999,39.379997,39.719997,9.69,0.42999998,0.29,26.32,32.219997,17.93,21.23,1.4699999,4.3199997,2.31,4.71,46.92,68.63,38.57,19.27,41.7,43.43,8.99,14.25,18.199999,13.4,9.0,12.7699995,27.48,85.159996,68.32,60.039997,22.199999,8.45,11.57,32.899998,66.36,56.699997,35.239998,9.74,2.4299998,12.41,15.71,0.01,0.16,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.55,0.57,0.099999994,0.39999998,0.58,1.12,1.16,0.82,0.22,0.0,0.0,0.0,0.0,0.02,0.03,0.47,0.48,0.26999998,0.0,0.0,0.0,0.0,0.0,0.0,0.08,0.52,0.52,0.44,0.08,2.1699998,2.8799999,9.0,6.04,3.6499999,3.12,2.6699998,0.96,0.07,0.71,0.41,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.06,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.38,0.53,0.02,0.0,0.04,0.22999999,0.21,0.16,0.02,0.16,0.39,1.01,1.23,5.6299996,4.4,1.8299999,0.65999997,0.17999999,0.02,0.0,0.0,0.049999997,2.84,5.83,6.83,3.49,0.17,0.0,0.0,0.0,0.0,0.0,0.06,1.4699999,0.7,0.77,5.25,18.35,2.53,0.17999999,4.36,0.32,2.52,13.94,29.189999,31.929998,28.23,9.23,6.23,16.699999,22.51,23.17,13.94,8.34,3.74,0.41,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.5,10.55,13.809999,26.73,11.55,2.6299999,0.52,0.0,0.0,0.03,0.06,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.05,3.51,0.0,0.07,41.129997,18.0,3.8,18.71,0.61,2.06,12.13,7.17,15.41,13.45,0.34,0.26,0.32,4.7999997,73.53,29.82,8.55,14.78,24.26,32.37,8.08,10.42,13.92,16.34,24.73,58.149998,86.52,69.93,31.33,23.789999,24.859999,17.109999,35.61,34.53,38.51,24.98,11.13,3.3899999,0.22,0.12,0.31,0.59,0.57,0.14,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02,0.55,0.53,0.11,0.06,0.42999998,0.59,0.51,0.19999999,0.03,0.0,0.0,0.0,0.0,0.0,0.04,0.16,0.04,0.0,0.0,0.0,0.52,0.0,0.0,0.0,0.08,0.12,0.0,0.0,0.0,0.41,4.43,2.95,1.93,1.77,0.45999998,0.0,0.0,2.48,3.54,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.04,0.049999997,0.0,0.0,0.0,0.0,0.0,0.04,0.16,0.13,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.29999998,0.79999995,0.03,0.52,1.56,2.58,2.8899999,0.48999998,0.049999997,0.19,0.84999996,2.6799998,3.21,2.75,1.24,0.53,0.22999999,0.08,0.95,2.28,5.46,7.1499996,1.65,0.29,0.0,0.0,0.0,0.0,0.0,0.57,1.56,1.4399999,0.89,4.46,9.099999,9.26,1.65,0.26,0.0,0.17999999,0.12,0.79999995,12.9,25.55,21.71,10.63,2.6299999,10.139999,22.859999,22.5,20.71,14.69,5.0699997,1.1999999,0.07,0.0,0.14,0.14,0.01,0.14,0.47,0.84,1.4599999,1.35,2.05,2.04,0.97999996,0.089999996,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.65,0.37,1.6999999,7.62,0.52,0.0,0.53,1.6899999,1.04,0.049999997,0.0,0.14999999,0.48999998,2.1,10.95,6.98,2.08,0.25,1.7099999,1.3299999,0.0,1.7199999,4.77,12.88,32.09,61.21,114.47,52.84,10.12,3.9199998,14.78,30.779999,47.7,39.079998,28.43,15.53,3.03,0.75,0.88,4.6,16.72,5.5099998,0.72999996,0.59,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.17,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.25,0.42,0.91999996,0.71999997,0.17999999,0.11,0.0,0.08,0.049999997,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14,0.0,0.0,0.39999998,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.29999998,0.42999998,0.0,0.17999999,0.71999997,0.26999998,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08,0.26999998,0.049999997,0.0,0.0,0.0,0.0,0.01,0.07,0.48999998,0.64,0.71999997,0.91999996,0.5,0.13,0.0,0.25,0.32999998,0.0,0.0,0.0,0.0,0.0,0.07,0.48,1.5999999,1.64,0.39,0.07,0.35999998,1.09,0.76,0.52,0.16,0.06,0.14,0.19999999,0.14,0.01,0.0,0.24,0.64,2.08,1.56,0.0,0.22,0.71,1.93,0.64,2.83,4.7,2.76,0.26,0.0,0.51,3.0,0.95,0.22999999,0.0,0.0,0.0,1.62,5.0,5.2599998,7.56,6.64,6.21,3.59,3.12,7.5099998,9.15,8.82,5.9,2.8899999,0.52,0.02,0.38,0.76,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.68,1.28,1.15,0.97999996,0.07,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.47,0.81,0.0,0.97999996,11.28,7.54,7.5099998,0.22999999,0.39,1.05,0.22999999,0.14,0.78,2.44,8.49,2.3999999,0.04,2.03,1.4699999,2.28,0.12,0.97999996,2.3999999,12.009999,30.72,28.51,34.719997,43.8,18.369999,5.85,23.779999,48.48,43.53,57.48,53.219997,14.29,0.83,0.0,1.09,7.2,13.74,16.199999,6.33,0.13,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.08,0.03,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.04,2.69,7.46,1.68,0.0,0.0,0.0,0.11,0.08,0.0,0.0,0.0,0.0,0.0,0.0,0.19999999,1.39,0.39,0.0,0.0,0.0,0.82,0.51,0.71,0.34,0.0,0.77,0.77,0.0,0.0,0.59999996,0.0,0.39999998,0.0,0.76,0.58,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08,0.53,1.14,4.5099998,4.31,1.62,0.75,1.16,0.65,0.35999998,0.16,0.099999994,0.02,0.0,0.0,0.0,0.0,0.03,0.0,0.04,0.01,0.12,0.35,0.26999998,0.32,0.22,0.06,0.04,0.049999997,0.0,0.0,0.0,0.089999996,0.95,0.9,0.47,0.21,1.37,5.3199997,4.21,2.04,3.56,0.98999995,0.17999999,0.08,0.64,0.47,0.08,0.06,0.32,0.049999997,0.7,1.79,4.0099998,5.7799997,3.9299998,1.79,0.21,0.0,0.32999998,0.78,1.4399999,1.64,1.05,0.44,0.14,0.01,0.0,0.0,0.14,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.48999998,0.78,4.36,18.33,16.91,2.96,1.25,1.8499999,4.72,1.11,0.0,0.16,0.14999999,0.0,0.0,1.9699999,4.5699997,0.089999996,0.32999998,0.0,0.0,1.39,6.2599998,19.46,27.689999,35.309998,69.74,58.18,21.199999,18.69,33.719997,27.65,48.469997,45.829998,21.99,1.3399999,0.94,11.7699995,18.939999,4.19,9.309999,1.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.26,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.11,0.049999997,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.17999999,5.43,7.5699997,1.4599999,0.08,0.0,0.0,0.06,0.099999994,0.0,0.0,0.0,0.0,0.0,0.07,1.04,1.39,0.0,0.0,0.0,0.0,0.79999995,0.81,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.94,0.9,0.83,0.39,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.95,1.56,3.4099998,0.29999998,0.35999998,0.53,0.12,1.14,1.4399999,1.1899999,1.24,0.84999996,0.65,0.53,0.38,0.099999994,0.099999994,0.02,0.0,0.0,0.13,0.48,0.5,0.26999998,0.0,0.0,0.0,0.0,0.0,0.02,0.06,0.04,0.0,0.41,0.71,2.7,1.63,2.56,4.64,2.48,3.77,5.8399997,6.24,5.8199997,10.9,9.63,5.38,0.29999998,0.45999998,0.64,0.0,0.0,0.0,0.0,0.0,1.4399999,2.3,1.7099999,2.35,1.3199999,0.57,0.14,1.75,5.74,9.44,4.7799997,0.28,0.0,0.0,0.04,0.02,0.0,0.24,0.14,0.81,0.19999999,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.19999999,0.06,0.0,0.0,0.39,0.13,4.5499997,5.0299997,1.36,0.0,0.0,0.9,3.28,0.89,8.03,5.5299997,3.1699998,0.17,0.0,0.0,3.3899999,3.08,2.03,8.94,38.32,26.939999,16.77,21.279999,8.83,13.62,1.48,6.75,42.899998,64.93,53.61,4.74,0.12,1.1899999,3.6999998,0.0,0.0,0.0,0.06,0.04,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.5,0.79999995,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.21,1.24,1.52,0.96999997,0.0,0.0,0.0,0.0,0.08,0.0,0.0,0.0,0.0,0.0,0.0,0.07,0.0,1.1899999,0.39999998,0.39999998,0.0,0.31,0.0,0.9,0.0,0.19999999,0.0,0.0,0.0,0.0,0.13,0.55,0.45,0.13,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.11,0.45,0.0,0.0,0.0,0.04,0.19999999,0.07,0.04,0.28,0.08,0.02,0.06,0.17999999,0.32,0.58,1.06,1.27,0.90999997,0.88,0.34,0.04,0.01,0.01,0.0,0.0,0.17,0.83,2.6599998,0.28,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.04,0.32,0.35999998,0.03,0.64,1.12,4.7999997,9.96,8.23,5.8599997,10.61,15.2699995,18.23,18.0,5.75,1.8399999,0.71999997,0.11,0.0,0.51,0.55,2.3,2.22,3.11,1.0699999,0.26,2.53,3.03,4.27,7.62,7.0099998,2.0,0.41,0.06,0.0,0.06,0.06,0.0,0.0,0.17,1.1999999,0.25,0.04,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.32,0.37,0.0,0.0,0.0,0.02,0.0,0.02,0.0,0.0,0.0,0.0,0.0,0.02,0.0,0.76,2.4199998,2.78,1.31,4.8399997,25.57,11.58,5.98,10.679999,4.22,1.92,0.0,2.73,2.51,0.66999996,2.54,25.869999,5.49,0.74,2.57,0.14999999,0.48999998,0.41,0.32,8.4,12.23,4.16,0.69,0.0,0.0,0.0,0.0,0.45999998,3.3799999,0.14999999,0.17999999,0.34,0.44,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.35,0.07,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.5,0.0,0.0,0.0,0.0,0.03,0.0,0.0,0.0,0.0,0.0,0.08,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.06,0.29999998,0.22999999,0.0,0.0,2.6699998,4.38,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.19,0.22,0.87,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.6999999,1.17,0.03,0.0,0.06,0.48999998,0.79999995,0.29,0.0,0.0,0.0,0.0,0.0,0.04,0.049999997,0.16,0.55,0.78,0.55,0.74,0.44,0.22999999,0.19,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.049999997,1.4,4.2999997,6.33,11.11,5.85,4.04,5.81,5.6099997,5.7999997,5.73,1.76,1.1,1.3,0.65999997,0.13,0.0,0.0,0.66999996,3.01,1.53,1.02,1.01,0.29999998,0.19999999,0.0,0.0,0.48999998,0.71999997,0.57,0.13,0.14999999,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.32999998,0.9,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.51,1.02,1.3399999,1.48,17.73,48.3,15.46,0.29,0.26,1.9,9.58,2.81,0.08,1.22,2.9299998,0.48,0.39999998,1.7099999,0.38,0.71999997,0.0,0.32,0.38,4.08,7.44,6.08,3.1699998,0.0,0.0,0.0,0.0,0.0,0.42,5.79,15.66,6.8599997,6.5699997,0.02,4.7999997,0.37,0.19999999,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07,0.25,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.04,0.07,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.5,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,3.34,5.18,1.54,0.79999995,0.0,0.62,0.5,1.8299999,1.9499999,0.62,0.21,0.0,0.0,0.0,0.0,0.0,0.0,0.22999999,0.35999998,0.16,1.0,0.78999996,0.17,0.01,0.03,0.26,0.57,0.71999997,0.78,0.049999997,0.17999999,0.48999998,0.74,1.3399999,1.12,0.59999996,0.32999998,0.44,0.26999998,0.13,0.12,0.099999994,0.07,0.0,0.0,0.0,0.0,0.0,0.049999997,0.089999996,0.07,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.28,1.05,1.3399999,2.9299998,5.17,4.9,2.46,1.11,0.52,0.83,0.24,0.63,0.34,0.07,0.0,0.0,0.0,0.11,0.35999998,0.39999998,0.089999996,0.17,1.5899999,2.1399999,0.56,1.4,3.51,5.5499997,5.38,4.0,2.56,1.24,0.52,0.32,0.13,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.35999998,1.4,2.9399998,2.9299998,4.49,0.88,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.59,0.32,0.0,0.0,0.22999999,2.03,0.25,0.0,0.0,0.0,0.0,0.0,0.0,0.42,1.89,7.3799996,3.9599998,3.3799999,6.93,0.0,0.0,1.8199999,4.9,2.51,3.84,1.6999999,0.0,0.02,0.0,0.0,0.02,0.96999997,3.28,3.1799998,2.18,17.34,94.189995,86.24,51.23,19.8,0.45,0.0,0.0,0.0,0.0,13.86,20.15,32.46,42.32,21.439999,0.0,0.52,0.0,0.06,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.25,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.17999999,0.19999999,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.53999996,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.49,1.53,0.0,0.48999998,1.11,0.66999996,0.47,0.0,0.26999998,1.6899999,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14,0.11,0.0,0.17999999,0.5,0.47,0.39999998,0.22,0.25,0.17,0.14999999,0.0,0.31,0.17,0.28,0.45999998,0.31,0.17999999,0.099999994,0.14999999,0.02,0.04,0.29,0.38,0.08,0.32,0.38,0.21,0.19,0.16,0.22,0.17999999,0.29999998,0.35999998,0.22999999,0.049999997,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.65999997,0.39,0.0,0.0,0.089999996,0.12,0.7,1.03,1.43,0.42999998,0.01,0.0,0.0,0.0,0.12,0.08,0.0,0.0,0.07,0.84,0.93,0.0,0.0,0.79999995,0.78999996,1.55,2.05,4.37,11.82,11.99,9.74,8.71,3.51,1.13,1.4699999,0.17,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08,0.34,0.71999997,2.12,4.58,1.67,0.68,0.78999996,0.22,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.31,2.03,0.0,0.0,0.0,0.07,0.56,0.0,0.0,0.0,0.0,0.0,0.0,0.26999998,6.1299996,11.349999,7.8199997,9.96,2.36,0.39999998,0.0,2.1,14.2699995,4.5899997,0.38,0.02,0.0,0.0,0.0,0.0,0.0,0.19999999,0.26999998,0.17,0.13,15.03,68.4,56.23,7.45,6.7999997,0.0,0.0,1.26,6.16,13.75,19.039999,8.46,36.5,42.489998,18.18,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02,0.57,0.42999998,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.31,0.34,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08,0.53999996,0.26999998,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.62,0.47,1.79,2.6499999,1.14,0.0,0.0,0.91999996,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.39,0.48,0.0,0.28,0.56,0.13,0.099999994,0.14999999,0.14999999,0.22999999,0.61,0.91999996,2.3899999,2.6499999,1.81,0.93,0.42,0.099999994,0.0,0.11,0.099999994,0.03,0.0,0.06,0.45,0.31,0.32,0.62,1.0,2.04,1.53,0.58,0.22999999,0.01,0.0,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.19,1.66,6.31,9.05,2.04,0.0,0.0,0.0,0.0,0.02,0.02,0.08,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.29999998,0.91999996,2.22,0.75,0.0,0.0,0.08,0.63,1.9499999,3.24,3.4399998,2.06,1.9599999,4.45,1.63,3.75,9.59,2.5,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.51,1.87,3.6699998,1.93,0.45999998,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.41,0.82,0.0,0.0,0.0,0.0,0.049999997,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,3.1,5.99,3.8999999,6.8199997,0.17,0.88,8.09,0.69,0.06,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13,0.45,0.26999998,0.0,2.5,4.35,0.48,0.0,0.0,0.0,2.7,9.7699995,11.969999,6.62,0.59999996,33.48,0.0,0.0,0.0,3.97,0.13,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.07,0.0,0.0,0.0,0.0,0.25,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.29999998,0.26999998,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.22999999,0.74,1.04,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.22999999,0.26999998,1.15,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.25,0.83,0.19999999,0.0,0.17,1.29,1.29,0.77,0.38,0.16,0.01,0.44,1.05,2.05,2.8799999,1.78,1.18,1.3199999,2.36,1.93,1.1999999,1.17,1.77,1.78,1.5799999,1.39,0.85999995,0.5,0.69,0.37,0.41,1.3,2.46,1.8499999,1.68,1.37,0.78,0.17999999,0.099999994,0.11,0.04,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.05,2.79,1.23,0.35,1.24,1.24,0.48,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.38,1.49,2.51,0.35999998,0.03,0.0,0.03,0.31,0.71,1.12,0.84999996,0.55,0.98999995,3.1799998,8.17,7.8999996,8.55,12.12,5.8199997,0.0,0.0,0.0,0.0,0.0,0.0,0.17999999,0.57,0.58,0.35999998,0.13,0.04,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.25,2.3999999,0.32,0.97999996,0.90999997,0.11,0.13,0.17999999,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.37,22.38,0.0,0.0,0.0,0.0,1.74,3.77,0.89,0.0,0.02,1.15,15.7699995,30.369999,28.599998,3.4199998,7.6499996,0.049999997,0.12,0.29999998,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.04,0.0,0.01,0.17999999,0.35999998,0.25,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.089999996,0.07,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.19999999,0.0,0.08,0.53999996,0.44,0.03,0.03,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.24,0.0,0.0,0.0,0.0,2.05,0.0,0.0,0.84,0.21,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.16,0.53,0.0,0.0,0.16,0.0,0.0,0.0,0.0,0.0,0.11,0.17999999,0.35,0.56,0.45,1.06,1.48,1.4499999,3.06,4.2599998,3.6599998,3.73,3.59,2.62,2.44,2.9099998,4.5499997,5.0699997,5.17,4.45,3.36,2.1699998,1.4699999,0.57,0.14999999,0.38,0.53,0.74,1.99,2.74,3.05,1.31,0.17999999,0.32,0.37,0.14,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.52,2.07,6.3399997,6.25,4.0,0.29999998,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.39,0.26,0.03,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.65999997,0.87,2.9099998,3.9299998,2.1399999,1.3,0.14999999,0.17999999,0.65,0.32,0.17999999,0.32,0.22,0.35,0.28,0.11,0.01,0.0,0.0,0.0,0.0,0.26,0.08,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.48,0.48999998,0.26999998,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.099999994,0.7,2.8999999,0.08,0.0,0.78,1.61,5.44,19.17,26.75,26.41,16.44,0.099999994,0.04,0.19,0.0,0.0,0.0,0.0,0.0,0.0,0.16,0.64,0.21,0.099999994,0.099999994,0.14999999,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.17,0.11,0.17999999,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.17999999,1.93,0.75,0.0,0.0,0.0,1.4499999,1.1999999,0.0,0.64,0.16,0.0,0.0,0.0,0.0,0.0,0.08,0.02,0.34,1.79,2.97,0.98999995,0.13,0.0,0.0,0.0,0.0,0.0,0.14999999,0.48,1.5699999,2.3899999,1.0,0.64,0.64,0.61,0.099999994,0.62,0.65,1.06,2.04,3.06,3.6299999,3.84,5.3599997,7.1099997,6.5699997,6.47,6.47,6.43,3.8999999,2.22,1.26,1.99,2.45,2.19,3.49,2.52,2.98,2.01,1.3199999,0.66999996,0.22,0.03,0.0,0.0,0.12,0.37,0.17999999,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.11,0.21,0.37,0.48,0.19,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.03,0.0,0.0,0.01,0.049999997,0.0,0.0,0.11,0.79999995,1.61,2.75,2.74,1.9,2.35,3.02,4.49,3.1799998,2.01,3.8999999,4.13,4.3199997,3.52,2.05,0.79999995,0.14,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.61,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.45999998,0.11,0.0,0.0,0.0,0.0,4.97,2.83,2.44,3.1499999,1.4499999,0.17,0.01,0.049999997,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.049999997,0.06,0.03,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13,0.35,0.81,0.32,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.1999999,2.6499999,1.25,0.0,0.0,0.39999998,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.099999994,0.48,2.46,4.0,6.66,2.19,0.049999997,0.0,0.0,0.0,0.0,0.17999999,1.53,3.74,2.2,1.35,1.14,1.15,0.31,0.07,0.04,0.39999998,0.53999996,0.5,1.1,1.55,2.1399999,3.1599998,3.51,4.56,4.91,6.12,6.8799996,6.37,3.99,3.27,2.52,3.27,3.98,4.1,4.2599998,3.99,3.29,2.6699998,3.7099998,6.5,2.82,0.65999997,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08,1.23,0.84,0.19999999,0.03,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.04,0.04,0.19999999,0.42999998,1.03,0.83,0.37,0.38,0.06,0.29,2.26,4.94,8.28,9.36,10.2699995,12.099999,12.03,15.799999,13.299999,7.97,4.21,1.63,0.35,0.089999996,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.22,0.45,0.08,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.04,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06,0.0,0.53999996,0.38,0.08,0.0,0.0,0.0,0.0,0.0,1.56,0.0,0.17999999,0.0,0.0,0.45999998,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.22999999,1.4,0.0,0.0,0.59999996,1.3399999,2.35,9.92,4.7,1.18,0.0,0.28,0.38,0.26,0.93,2.19,3.1599998,1.5799999,0.65,0.95,1.48,1.4699999,1.02,0.81,0.64,0.48,0.45999998,0.42,0.29999998,0.64,1.5,2.83,3.73,4.0499997,4.65,5.71,5.99,4.74,3.27,1.76,1.43,2.76,4.88,6.41,6.66,6.5499997,4.91,4.43,4.35,3.46,0.87,0.26999998,0.06,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.049999997,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.089999996,0.32,0.90999997,1.39,1.7099999,0.96,1.29,1.63,3.87,7.1,4.64,4.91,6.96,9.73,11.759999,13.49,19.39,14.599999,9.58,5.04,2.79,1.05,0.26,0.37,1.8299999,2.49,2.06,2.3899999,1.9,0.97999996,0.38,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.19,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07,0.049999997,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.099999994,0.07,0.089999996,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.04,0.04,0.11,0.11,0.0,0.0,0.0,0.0,0.52,0.0,0.39999998,0.42999998,0.29999998,0.96999997,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.31,2.77,2.8,4.0,1.22,0.0,0.0,0.0,0.0,0.42999998,0.58,0.39999998,0.48999998,0.94,0.65999997,0.48999998,0.53999996,0.68,1.0699999,1.2099999,1.0699999,1.3399999,1.5799999,0.79999995,1.23,2.02,1.9699999,2.12,2.71,2.77,2.83,3.76,4.79,4.63,3.3899999,1.8399999,0.96999997,0.42999998,0.44,2.46,4.29,4.7999997,3.3999999,2.56,1.5699999,1.0,0.65999997,0.62,0.21,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.089999996,0.45,1.12,1.01,0.39,0.47,1.78,2.6,3.79,6.6099997,10.9,11.13,8.57,6.5699997,7.91,9.309999,10.98,7.89,4.5099998,2.8999999,0.83,0.45,3.1899998,4.81,4.5,4.42,4.39,2.3899999,1.26,0.07,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02,0.12,0.32,0.099999994,0.099999994,0.0,0.0,0.16,0.22999999,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.04,0.04,0.17,0.0,0.0,0.0,0.59999996,0.7,0.0,0.26999998,1.9599999,3.1899998,0.0,0.0,0.0,0.0,0.0,4.67,0.0,0.0,0.0,0.0,0.099999994,1.74,1.9,0.82,2.6499999,0.71999997,0.08,0.0,0.0,0.0,0.41,0.089999996,0.0,0.0,0.12,0.06,0.01,0.12,0.19999999,0.48999998,0.98999995,1.8,2.9199998,2.33,0.59,0.47,0.96999997,2.1699998,2.22,2.85,2.6599998,1.8199999,1.81,2.9199998,3.83,4.46,4.2,2.6799998,1.35,0.89,0.17,0.34,1.3199999,1.29,1.35,0.82,0.53,1.4,1.81,2.05,0.099999994,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.29999998,1.4,1.8,1.05,1.49,1.79,1.53,2.85,5.12,6.31,5.8599997,4.65,3.77,5.91,8.87,8.5,5.7799997,4.3199997,4.0299997,1.9599999,0.71999997,3.3899999,3.52,3.28,3.72,2.78,1.3399999,0.37,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.55,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.28,0.84999996,0.17999999,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13,0.17999999,0.0,0.0,0.0,0.0,0.07,0.0,0.08,0.099999994,0.17,0.07,0.099999994,0.07,0.28,1.0699999,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13,0.76,0.0,0.0,0.0,0.0,0.35,0.0,0.94,3.1599998,0.0,0.0,0.0,0.0,7.77,0.71,0.0,0.0,0.0,0.0,0.64,0.32999998,1.1899999,2.6399999,3.1,1.5999999,0.65,0.07,0.0,0.03,0.17,0.24,0.26999998,0.5,0.68,0.56,0.22,0.35999998,0.65,0.44,0.56,0.58,0.95,0.61,0.52,2.37,3.37,4.5299997,5.0499997,3.33,2.8999999,2.6399999,2.6499999,2.75,3.06,3.55,3.85,3.83,2.87,2.03,1.4399999,1.09,0.29999998,0.78999996,1.5699999,2.9399998,3.07,2.35,0.91999996,0.45,0.14,0.11,0.03,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02,0.06,0.14,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.04,0.45999998,0.29999998,1.0699999,1.99,2.51,1.74,2.46,3.12,2.76,2.8899999,2.8899999,3.4099998,4.94,8.17,7.2599998,5.6099997,5.7799997,4.33,3.01,2.77,2.35,2.9099998,2.8799999,2.7,2.33,1.39,0.78,0.25,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.099999994,0.42,0.32,0.089999996,0.0,0.0,0.06,0.32,0.14999999,0.13,0.22999999,0.16,0.04,0.049999997,0.47,0.95,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.22,2.1499999,2.31,2.31,0.47,0.0,0.0,0.22999999,0.0,0.45,4.08,4.97,2.1699998,3.3999999,1.8199999,1.24,0.0,0.62,0.53999996,0.0,0.04,0.88,5.0499997,2.84,6.25,5.5,1.26,0.14,0.04,0.0,0.5,0.66999996,1.25,2.24,2.29,3.4099998,3.54,2.62,1.17,0.38,0.19999999,0.77,1.1999999,0.81,1.0799999,2.0,5.8199997,5.62,3.1799998,5.2999997,4.83,3.74,4.97,5.64,5.93,6.22,5.72,4.88,3.97,3.06,1.88,0.57,0.06,0.03,0.56,2.54,1.9499999,1.5899999,1.38,0.53,0.53999996,0.64,1.17,0.28,0.0,0.0,0.0,0.0,0.03,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.42,0.59,1.51,1.16,1.23,1.39,1.86,3.33,3.3999999,4.62,9.45,10.73,10.87,10.46,8.71,6.02,5.43,3.8799999,2.7,3.1399999,3.9199998,3.6699998,3.73,3.1399999,1.7099999,1.03,0.21,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07,0.049999997,0.0,0.0,0.0,0.0,0.0,0.03,0.28,0.52,0.45,0.22,0.5,1.09,0.91999996,0.48999998,0.17999999,0.08,0.03,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.81,3.22,2.87,0.65,0.48,2.45,0.22,0.85999995,1.09,0.39999998,0.84,0.41,0.78999996,0.35999998,2.02,1.75,1.17,2.29,0.95,0.0,0.0,0.0,0.0,0.94,2.18,3.51,3.1599998,0.22,0.02,0.01,0.19,0.35,0.42999998,0.44,0.21,0.17999999,0.29999998,0.42,0.62,2.06,2.3799999,1.02,0.14999999,0.19999999,0.32999998,0.38,0.75,2.0,4.23,5.72,4.93,2.9299998,3.54,5.0699997,6.73,9.26,9.849999,8.61,7.45,7.64,5.02,4.6,3.03,2.08,1.4499999,0.84,0.5,0.62,0.37,0.19999999,0.28,0.65,1.66,1.53,1.17,0.58,0.16,0.049999997,0.099999994,0.099999994,0.03,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02,0.099999994,0.11,0.099999994,0.06,0.099999994,0.35999998,1.22,0.81,1.74,1.89,2.69,2.57,2.07,2.74,4.17,5.68,8.309999,8.679999,10.63,10.88,8.599999,8.53,9.92,10.099999,9.139999,8.26,6.02,3.1499999,1.63,0.39999998,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.049999997,2.34,4.13,1.6999999,2.6,0.84,0.79999995,0.29,0.01,0.0,0.0,0.01,0.14,0.21,0.29999998,0.22999999,0.26999998,0.07,0.03,0.08,0.06,0.38,0.97999996,1.03,0.81,0.45,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.11,0.16,0.12,3.37,5.7999997,4.42,2.1399999,3.87,9.08,3.28,3.4399998,2.73,2.62,0.0,0.0,0.0,0.0,1.09,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.29999998,0.0,0.32999998,0.34,0.59,2.49,2.47,0.59999996,1.48,1.73,1.67,2.8799999,3.4499998,4.04,2.57,2.27,1.5,0.45999998,0.65,0.04,0.11,0.089999996,0.5,1.53,2.23,1.8499999,2.09,3.1799998,3.32,4.4,5.04,6.27,7.2799997,8.059999,7.9199996,7.83,8.0199995,6.2999997,5.38,3.97,2.52,1.27,0.17,0.0,0.0,0.0,0.03,0.51,1.06,0.98999995,0.34,0.9,0.39,0.14,0.11,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.04,0.01,0.0,0.03,0.34,0.35999998,0.64,0.94,1.17,0.91999996,0.93,1.31,2.31,3.76,6.08,8.82,12.78,13.929999,14.929999,18.23,18.69,16.97,14.37,11.32,6.77,3.28,1.4599999,0.31,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.19999999,3.6299999,5.44,5.74,28.0,34.55,43.02,33.86,4.21,0.32999998,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.35,0.59,2.47,4.2999997,5.81,9.309999,7.7999997,1.8499999,0.5,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.98999995,0.0,0.0,0.03,0.0,0.19,1.28,0.089999996,0.08,2.7,0.0,0.04,1.37,0.22999999,0.04,0.48,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,4.17,0.01,0.03,0.22999999,3.62,8.22,7.5299997,7.66,8.929999,7.5699997,10.929999,11.25,7.35,4.63,2.8899999,1.64,0.98999995,0.39999998,0.28,0.089999996,0.0,0.21,0.22999999,0.82,1.03,0.29,0.26,1.64,5.7599998,10.71,10.29,9.349999,7.31,6.2999997,6.71,7.54,7.6099997,7.16,5.8799996,4.65,3.37,2.0,1.09,0.37,0.13,0.06,0.01,0.14,0.55,0.39999998,0.21,0.56,0.48,0.35,0.089999996,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.29999998,0.53,0.19,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08,0.71999997,1.52,1.27,0.9,0.5,0.32999998,0.57,0.64,0.90999997,1.9799999,3.1999998,5.47,11.349999,16.5,18.99,19.789999,16.109999,11.849999,7.6499996,4.0899997,2.11,1.18,0.51,0.14,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.19999999,1.05,1.76,10.66,27.15,41.95,53.01,60.18,30.76,8.25,2.02,0.16,0.0,0.0,0.0,0.0,0.089999996,2.19,7.64,8.9,6.8399997,10.66,14.78,14.429999,11.059999,5.21,1.4,0.06,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.049999997,0.04,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,13.13,0.42999998,0.0,0.0,0.0,0.0,0.0,0.0,0.02,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08,0.17,0.48,0.0,0.0,0.0,0.0,0.0,6.27,0.75,0.08,1.03,1.4,3.4499998,6.67,5.99,14.559999,12.36,16.039999,15.549999,12.5199995,7.0299997,5.99,4.3399997,2.76,1.75,1.01,0.29,0.35,0.55,0.16,0.04,0.0,0.0,0.0,0.22999999,2.4099998,8.48,11.36,14.0199995,12.13,7.02,4.44,4.36,3.86,5.45,6.7999997,5.92,4.5,3.35,2.6,2.1499999,1.36,0.83,0.58,0.35,0.29,0.06,0.12,0.62,0.66999996,0.39999998,0.22,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.049999997,0.31,0.16,0.28,0.39,0.19,0.16,0.22,0.22,0.42,0.47,0.63,1.5699999,3.4399998,4.88,5.8399997,5.0,2.6799998,2.12,1.48,0.96,0.58,0.29,0.099999994,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.41,1.3,10.62,23.68,37.0,35.73,45.219997,35.71,19.26,10.28,2.73,0.69,0.03,0.0,0.0,0.17,1.3299999,4.8599997,10.559999,6.6,4.0099998,4.18,5.7799997,7.98,8.87,3.61,0.29,0.04,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.48,2.78,1.9399999,1.91,1.3,1.63,1.5799999,1.26,0.84,1.3399999,1.35,0.53,0.22999999,2.01,4.87,0.0,0.0,0.0,0.0,0.0,0.089999996,0.71,0.90999997,0.59999996,0.39,2.97,7.98,2.35,3.35,7.99,7.16,8.33,9.08,7.64,7.8199997,6.45,5.14,3.1699998,1.7099999,0.74,1.01,0.62,0.099999994,0.0,0.0,0.0,0.0,0.0,0.0,1.1999999,2.73,7.18,10.639999,10.099999,7.74,5.37,4.22,5.06,6.77,4.21,2.8899999,2.8899999,3.1999998,2.7,2.9299998,2.8999999,2.3899999,1.4499999,1.6899999,2.3999999,2.6,0.48999998,0.19,0.13,0.049999997,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07,0.28,0.45,0.44,0.29,0.13,0.14,0.25,0.47,0.71999997,0.66999996,1.28,1.67,0.84999996,0.14999999,0.17,0.31,0.5,0.93,1.03,0.75,0.22999999,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.48,6.1,13.65,30.65,36.26,39.71,40.03,30.23,19.23,10.96,8.0,2.74,0.089999996,0.0,0.06,0.01,0.84,1.5899999,2.33,2.1399999,1.18,1.2099999,1.43,1.55,1.7099999,1.49,1.31,0.66999996,0.24,0.06,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.0,3.46,4.11,3.27,4.23,6.72,7.22,7.02,9.73,14.23,16.24,17.34,15.19,11.469999,6.6099997,3.05,1.3199999,0.48,0.5,0.17,0.13,0.06,0.29,0.66999996,0.94,0.66999996,0.47,0.53,2.04,3.6699998,4.45,3.61,3.33,6.7799997,7.71,9.05,8.17,6.3399997,4.9,4.31,2.54,1.23,0.45999998,0.16,0.06,0.01,0.0,0.0,0.0,0.01,0.41,0.78999996,0.42,1.63,3.37,4.47,4.65,3.57,3.0,3.01,2.71,2.74,3.73,4.95,2.87,2.54,2.34,2.28,3.02,3.24,4.3199997,5.25,2.11,0.78999996,0.25,0.22999999,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.16,0.32999998,0.71,1.38,1.9399999,2.24,1.81,1.02,0.75,0.59999996,0.77,0.97999996,0.84999996,0.32,0.0,0.0,0.04,0.17999999,0.41,0.53999996,0.45,0.22999999,0.089999996,0.06,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.81,4.71,15.349999,26.279999,47.36,59.859997,45.59,31.769999,16.449999,9.58,4.77,3.3999999,0.82,0.08,0.01,0.0,0.26,0.94,2.27,3.09,3.3999999,1.93,0.45999998,0.45999998,1.4499999,3.9499998,5.5699997,6.27,5.8799996,6.3399997,9.86,10.42,3.37,0.77,0.03,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.31,0.79999995,0.55,1.0799999,2.1499999,2.58,2.32,3.5,6.1,8.11,11.96,8.48,4.02,3.74,2.0,1.6899999,0.9,2.31,3.1799998,2.98,1.1999999,0.35,0.099999994,0.13,0.02,0.02,0.07,1.11,3.79,10.49,17.59,13.12,6.8199997,4.2799997,3.82,2.72,3.1399999,4.24,2.79,2.61,2.2,1.8499999,1.0799999,0.62,0.29999998,0.08,0.02,0.19,0.14,0.37,1.0,1.28,1.9599999,2.04,2.2,1.29,1.01,1.55,1.9799999,1.56,1.91,5.06,5.97,6.8399997,5.29,3.26,1.88,1.29,1.76,2.31,3.77,7.06,4.98,3.29,1.7199999,1.4699999,1.14,0.57,0.26,0.11,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.12,0.55,1.1899999,0.98999995,1.52,1.54,1.3399999,1.16,1.01,1.61,2.21,1.18,0.42,0.07,0.0,0.03,0.29999998,0.56,0.48999998,0.26999998,0.12,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.22999999,1.0,3.04,10.44,29.01,40.079998,30.64,21.91,11.509999,5.7599998,4.06,4.02,5.79,2.99,1.67,1.17,0.39,0.08,0.78,2.76,4.42,3.6499999,2.1399999,0.87,0.41,0.69,2.0,4.46,11.5,23.58,39.64,46.48,36.54,28.57,10.54,2.54,0.63,0.16,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.03,1.56,1.5799999,0.08,0.0,0.17999999,0.0,0.0,0.0,0.0,0.03,1.89,0.12,0.049999997,0.0,0.06,0.35999998,1.06,3.31,5.0699997,3.86,0.63,0.08,1.05,3.51,5.97,6.2599998,4.25,2.0,0.78999996,0.22,0.07,0.37,0.93,1.8299999,4.3399997,9.98,9.469999,7.6699996,5.12,2.22,1.05,0.51,0.94,1.81,2.1399999,1.16,1.6999999,1.9599999,2.09,1.42,0.64,0.51,0.42999998,0.32,0.08,0.14999999,0.13,1.1999999,2.9099998,2.79,1.64,1.37,0.95,0.35999998,0.79999995,0.69,1.0699999,1.9,2.21,2.56,2.73,2.76,2.9199998,2.47,2.04,1.6899999,1.09,1.89,2.1299999,3.97,3.6,4.49,4.56,4.06,2.47,1.41,0.74,0.29,0.08,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.03,0.22999999,0.32999998,0.61,1.11,1.29,1.5899999,1.51,1.4399999,1.27,1.3199999,1.5799999,1.5,1.03,0.53999996,0.32,0.13,0.03,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.19,1.89,10.66,21.75,23.72,20.31,15.349999,10.389999,6.47,3.9499998,6.95,6.39,3.78,3.1499999,2.56,1.11,0.35999998,0.19999999,0.14,0.11,0.29,0.07,0.12,0.37,0.32,0.22,2.11,7.8399997,17.789999,31.849998,42.59,40.239998,22.33,10.809999,5.56,2.04,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.0,0.0,0.0,0.0,0.12,1.3199999,1.88,1.04,0.34,0.0,0.07,1.0,0.0,0.07,0.44,0.14,0.32,3.83,3.9399998,6.5499997,8.07,1.1,0.59999996,0.0,0.96,1.0,0.53,0.9,1.1899999,0.97999996,0.29999998,0.12,0.06,0.17,0.37,1.5999999,4.16,7.68,7.5299997,4.04,2.3799999,2.18,1.0799999,0.98999995,3.05,4.5699997,3.12,1.79,1.77,2.6,3.34,4.0099998,3.9399998,2.3,0.71999997,0.19,0.02,0.07,0.01,0.26999998,0.5,0.41,0.83,0.52,0.22,0.12,0.089999996,0.17999999,0.32,0.59,0.95,1.41,1.26,1.25,1.06,0.74,0.56,0.48,0.45999998,0.45999998,0.59,1.01,1.63,2.27,2.69,3.26,3.02,1.91,0.95,0.45999998,0.14999999,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02,0.81,2.6799998,2.3999999,1.9399999,1.06,0.87,0.77,0.07,0.29,0.45999998,0.45999998,0.35,0.21,0.07,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07,4.87,8.139999,9.86,10.41,10.57,9.09,6.2599998,4.2799997,2.6399999,2.2,3.9099998,6.16,6.35,3.62,2.0,1.3299999,1.09,0.77,0.12,0.0,0.0,0.0,0.02,0.06,0.78,3.83,5.5299997,10.17,11.84,11.84,10.889999,8.72,4.27,1.3299999,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.17999999,0.13,0.17999999,0.45999998,0.63,2.5,3.01,2.02,0.69,0.24,0.87,0.0,0.22999999,0.61,0.96,0.25,0.12,0.0,1.76,20.279999,6.39,0.68,1.26,1.5799999,0.76,0.089999996,0.03,0.08,0.06,0.0,0.0,0.0,0.0,0.0,0.089999996,0.42999998,2.31,2.04,2.81,1.8499999,3.09,4.49,5.5299997,6.1099997,8.95,6.85,5.2799997,3.6999998,1.6999999,1.4599999,3.33,5.6299996,6.8799996,5.97,2.6699998,0.14,0.04,0.01,0.03,0.01,0.19,0.44,1.0,1.1899999,1.9,3.3899999,6.39,4.5699997,1.4499999,0.32999998,0.22,0.44,0.41,0.48999998,0.45,0.38,0.17999999,0.12,0.03,0.03,0.07,0.31,0.65,0.34,0.11,0.03,0.14,0.19999999,0.25,0.13,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.049999997,0.22999999,1.16,1.5999999,1.3,1.39,1.4499999,1.7199999,0.32999998,0.04,0.049999997,0.08,0.049999997,0.03,0.03,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.48,1.8399999,4.38,9.25,6.0299997,9.76,7.5699997,10.389999,7.81,4.29,2.84,2.55,5.7599998,7.9199996,6.0699997,3.46,2.96,3.09,5.0299997,7.2599998,6.67,3.25,0.79999995,0.17,0.08,0.22999999,2.45,3.6499999,5.19,5.12,2.75,0.52,0.02,0.03,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14999999,0.78,0.59999996,1.3199999,2.8899999,5.21,3.97,4.0899997,3.9299998,0.42,3.1599998,1.3399999,2.3899999,1.13,1.5799999,1.9499999,2.44,2.69,1.5799999,2.3,2.71,0.78999996,0.75,2.85,0.56,0.69,0.26999998,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.089999996,0.39999998,0.71,0.28,0.32,0.099999994,2.1,2.78,5.98,8.29,10.36,10.639999,8.71,3.8999999,1.88,1.62,2.36,3.82,5.15,7.37,8.25,6.98,2.26,0.91999996,0.68,0.65,0.96999997,0.53,1.17,3.01,2.61,2.57,2.4199998,1.64,0.7,0.29999998,0.24,0.089999996,0.06,0.049999997,0.08,0.08,0.07,0.0,0.0,0.0,0.0,0.089999996,0.06,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07,0.44,1.12,1.5699999,1.5999999,1.36,0.7,0.65,1.0799999,1.24,1.22,1.0699999,0.88,0.59,0.39,0.24,0.07,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.39,1.06,1.2099999,8.29,12.38,13.719999,9.13,6.3599997,4.46,4.8599997,1.81,1.8399999,1.78,1.42,3.1899998,0.90999997,1.06,1.3399999,1.53,1.52,1.62,0.91999996,0.19999999,0.099999994,0.75,2.46,2.1399999,2.55,2.9399998,1.3299999,0.42999998,0.089999996,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13,0.59,0.93,0.82,0.39999998,0.17999999,0.41,0.52,0.37,0.22999999,0.06,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02,0.39999998,0.96999997,0.48999998,0.32,0.35,0.0,0.0,0.0,0.68,0.0,0.0,0.38,2.12,0.58,1.53,1.8199999,1.8,1.56,1.5799999,1.5799999,1.4,0.0,0.0,2.23,0.24,0.0,0.0,0.0,0.03,0.24,0.58,0.47,0.42,0.72999996,0.26999998,0.59,2.0,1.9,1.41,1.35,0.96,0.75,1.01,2.05,3.0,5.5299997,7.1499996,8.86,9.49,8.389999,8.62,9.94,9.809999,10.309999,10.79,9.7,7.19,5.92,3.53,1.7199999,1.55,1.29,1.54,1.7199999,1.05,0.55,0.22,0.02,0.42999998,1.65,2.3999999,2.54,2.74,2.26,0.97999996,0.35999998,0.099999994,0.17,0.19999999,0.29,0.21,0.06,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.03,0.16,0.41,0.74,0.82,0.53999996,0.48999998,0.41,0.42999998,0.32999998,0.25,0.19,0.14,0.089999996,0.04,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.57,0.0,0.03,0.07,0.01,0.0,0.03,0.26999998,0.71,0.79999995,1.27,1.74,1.06,1.23,1.01,0.53,0.42999998,0.44,0.32999998,0.16,0.01,0.34,2.28,3.6699998,7.73,5.02,4.45,3.6999998,2.99,2.09,0.98999995,0.82,0.96,0.59,0.53999996,0.53999996,0.56,0.93,1.3399999,1.15,0.66999996,0.42,0.24,0.29999998,0.5,0.62,0.19999999,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.11,0.089999996,0.0,0.0,0.089999996,0.22999999,0.06,0.0,0.22,0.29999998,0.089999996,0.0,0.04,0.19999999,0.03,0.0,0.0,0.0,0.03,0.22,0.13,0.03,2.58,1.73,1.28,0.53999996,4.14,2.75,0.82,0.0,0.41,0.17999999,0.11,1.4399999,1.5,1.28,2.3,3.01,0.71999997,0.5,0.62,1.3199999,3.84,7.45,14.74,13.7,10.24,9.61,8.91,7.5499997,7.93,5.04,3.31,3.79,3.72,5.0699997,6.42,5.13,4.65,3.31,1.4399999,0.41,0.099999994,0.03,0.44,1.38,2.6599998,4.74,4.5899997,4.64,2.57,1.91,2.03,2.2,1.48,1.27,0.65999997,0.39,0.22999999,0.03,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07,0.0,0.0,0.14999999,0.099999994,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.049999997,0.08,0.03,0.0,0.0,0.12,0.42,0.93,1.53,2.03,2.22,1.78,1.06,0.44,0.14999999,0.049999997,0.06,0.08,0.13,0.84,3.52,10.69,14.54,20.039999,15.19,10.07,6.69,4.52,3.49,3.61,4.42,5.33,4.72,3.22,1.92,1.66,1.4699999,1.1999999,1.06,0.98999995,0.81,0.37,0.11,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06,0.41,0.45,0.04,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.11,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.04,0.01,0.0,3.87,9.75,7.1,8.7699995,6.72,1.86,0.9,0.19999999,0.0,0.62,2.9299998,4.68,4.8199997,4.1,2.59,0.17999999,1.17,2.71,1.1999999,0.75,0.75,1.67,7.33,10.67,10.639999,10.469999,15.339999,16.07,12.2,9.54,9.0199995,5.39,5.52,5.2599998,5.02,6.25,6.33,3.87,1.79,0.85999995,0.5,0.22999999,0.16,0.45999998,0.96,2.07,4.64,5.06,4.39,3.8799999,3.07,3.6499999,2.86,2.85,1.74,1.16,0.94,0.35999998,0.11,0.02,0.0,0.0,0.22999999,0.39999998,0.12,0.16,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02,0.04,0.0,0.0,0.0,0.0,0.0,0.01,0.02,0.14,0.17999999,0.11,0.07,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.19999999,0.47,0.82,0.25,0.13,0.45999998,1.0799999,1.8499999,2.8999999,3.46,3.73,3.29,2.35,0.97999996,0.45999998,0.29,0.34,0.39,0.45999998,3.1299999,10.639999,24.539999,19.91,26.97,24.74,18.869999,13.41,9.75,9.179999,9.21,9.44,11.15,11.92,10.05,8.79,7.71,6.79,5.64,4.62,3.85,2.83,1.74,0.96999997,0.45999998,0.48,0.56,0.37,0.07,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07,0.47,0.96,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.11,0.02,0.0,0.0,0.0,0.0,0.0,0.14,0.69,0.12,0.0,0.0,1.5699999,10.74,12.0199995,3.32,1.5,0.37,1.5999999,4.2,7.41,6.73,8.59,7.58,4.83,1.6999999,0.17999999,0.0,0.0,0.03,0.26999998,0.099999994,1.91,2.45,3.37,1.91,2.84,2.8899999,5.47,6.04,9.429999,11.13,9.25,7.04,5.33,4.75,4.5299997,4.0,2.73,1.41,1.14,0.96999997,0.88,0.59,0.34,0.16,0.07,0.22,1.13,1.5699999,1.53,1.4599999,1.67,2.05,2.2,2.53,2.1699998,2.1399999,1.31,1.12,0.19999999,0.03,0.14999999,0.45,0.74,0.68,0.32,0.17999999,0.01,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.39,1.29,1.9399999,1.3,0.39999998,0.11,0.06,0.0,0.0,0.0,0.01,0.08,0.14,0.19999999,0.21,0.14999999,0.12,0.08,0.049999997,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.04,0.24,0.77,0.26,0.07,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.099999994,1.28,4.56,7.95,8.16,5.33,4.5299997,11.16,11.66,6.12,3.6,4.15,6.2799997,7.3999996,7.0099998,5.41,3.26,1.67,1.01,1.13,1.9399999,6.29,19.16,37.69,30.64,31.519999,34.12,29.82,21.76,15.889999,13.03,11.04,9.969999,10.7,10.98,10.179999,9.05,8.0,7.08,5.95,4.89,4.0,2.95,2.09,1.3,0.63,0.59,0.68,0.5,0.25,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.22999999,1.6899999,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.22999999,0.0,0.87,1.5999999,3.0,4.72,3.85,2.36,1.4,0.13,0.0,0.0,0.0,0.02,0.25,0.04,0.12,0.13,0.17999999,0.099999994,0.0,0.22,0.68,0.88,1.23,1.5999999,2.9199998,3.72,4.5299997,4.87,4.5,3.25,2.69,1.89,1.4599999,0.59999996,0.74,0.48999998,0.35999998,0.37,0.22999999,0.21,0.31,0.26999998,0.39999998,0.14,0.28,0.59999996,1.68,3.03,3.1899998,3.4299998,2.1299999,1.4,1.67,0.74,0.59,0.32999998,0.29999998,0.35,0.14,0.13,0.12,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02,0.34,1.8199999,3.6599998,6.74,9.96,7.54,1.9,0.48,0.03,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.02,0.06,0.099999994,0.06,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.26,0.74,0.19,0.03,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.04,0.02,0.0,0.61,5.7599998,16.84,24.64,20.17,19.949999,26.33,31.349998,25.939999,16.9,8.889999,5.0499997,5.79,7.5099998,8.55,7.8199997,6.5,4.7799997,3.34,4.31,8.309999,18.74,36.59,34.64,31.439999,37.809998,38.55,34.92,30.97,25.88,19.33,14.509999,11.96,10.17,8.79,7.2999997,6.49,5.44,4.49,3.6,2.7,1.9399999,1.15,0.59999996,0.29999998,0.32999998,0.51,0.59,0.31,0.04,0.03,0.02,0.02,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.32,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.07,0.21,1.05,0.19999999,0.0,0.0,0.0,0.02,0.08,0.0,0.0,0.0,0.099999994,0.14999999,0.13,0.39999998,0.04,0.03,0.0,0.11,0.48,0.88,2.57,2.86,1.54,2.22,3.02,4.19,4.67,4.14,3.48,2.27,1.53,0.82,0.44,0.099999994,0.089999996,0.32,0.71999997,1.03,1.3399999,0.90999997,1.0,1.4399999,2.3899999,3.3,2.1299999,1.6999999,2.18,1.3,0.47,0.02,0.0,0.0,0.02,0.04,0.03,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.59999996,3.9199998,8.36,10.94,13.259999,10.61,6.49,4.2799997,3.31,1.8499999,1.2099999,0.53999996,0.29999998,0.099999994,0.049999997,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.31,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.6399999,11.45,23.92,29.369999,27.5,24.56,26.71,27.98,25.13,19.57,13.46,8.17,5.62,5.0099998,5.99,6.15,5.56,4.6,3.98,5.45,8.389999,11.73,15.78,22.02,31.23,37.42,45.3,46.1,38.91,28.91,19.51,15.799999,14.13,13.5,12.71,11.46,9.92,8.65,7.35,5.47,3.98,3.07,2.1699998,1.5899999,1.26,1.15,1.06,0.64,0.37,0.32,0.25,0.17999999,0.16,0.099999994,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.45999998,0.79999995,1.6899999,1.4499999,2.54,2.1499999,0.82,0.77,0.14999999,0.099999994,0.03,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.089999996,0.42,0.97999996,1.4599999,1.9,2.3799999,2.3,2.24,1.93,1.4,0.87,0.48999998,0.11,0.03,0.01,0.0,0.0,0.11,0.29999998,0.96999997,1.04,0.53,0.42999998,1.27,1.79,0.72999996,0.17,0.19,0.11,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.28,3.9199998,5.98,5.2999997,5.6299996,4.11,3.4099998,2.8899999,3.09,2.57,2.32,1.92,1.35,0.63,0.31,0.11,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02,0.78,5.12,11.07,16.46,20.32,22.82,23.99,23.939999,21.51,17.72,14.009999,9.51,6.47,4.88,4.91,5.0299997,4.48,3.1399999,2.84,2.99,3.1599998,3.9099998,5.64,7.31,10.3,15.759999,26.23,34.239998,32.38,26.49,20.18,16.199999,14.12,13.08,11.849999,10.889999,9.75,8.46,7.29,6.08,4.67,3.31,2.48,1.81,1.31,0.76,0.19,0.02,0.12,0.34,0.21,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.52,0.17999999,0.099999994,0.31,0.24,0.11,0.24,1.25,1.67,2.54,4.0499997,4.38,2.6499999,2.34,1.0699999,3.1899998,1.81,0.25,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.04,0.11,0.28,0.42,0.61,0.48,0.55,0.51,0.38,0.19,0.06,0.01,0.0,0.0,0.0,0.0,0.04,0.07,0.049999997,0.12,0.39999998,0.56,1.04,0.98999995,0.65999997,0.34,0.51,0.38,0.0,0.07,0.17,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.28,0.81,0.71999997,0.55,0.58,0.59999996,0.97999996,0.76,0.61,0.45,0.48,0.47,0.32999998,0.17,0.06,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06,1.1,3.8799999,6.2799997,9.44,12.94,17.4,18.24,17.9,15.36,12.17,8.33,5.8599997,4.04,4.04,4.5499997,4.6,4.47,3.35,3.35,4.0699997,3.8899999,3.85,5.0899997,6.1,5.54,5.33,11.88,18.74,20.35,18.18,16.039999,14.45,13.17,11.32,10.01,9.19,7.8799996,6.7799997,6.04,4.79,3.98,3.3,2.26,1.86,1.74,0.65999997,0.17999999,0.01,0.17,0.35999998,0.14999999,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.22999999,3.4099998,2.54,2.04,3.6599998,4.04,2.09,0.04,0.38,0.26,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.06,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13,0.29999998,0.19999999,0.12,0.01,0.0,0.0,0.0,0.0,0.0,1.24,0.51,0.42999998,0.65999997,0.41,0.76,0.39,0.22,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.04,0.28,0.31,0.0,0.0,0.0,0.0,0.0,0.02,0.049999997,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.01,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.19,1.3199999,1.9799999,2.3799999,3.5,6.5499997,9.559999,12.44,12.53,9.96,7.08,4.25,2.4199998,1.86,2.79,3.4499998,3.3799999,3.33,2.52,1.9499999,2.12,2.22,2.36,1.9599999,1.42,1.62,3.99,7.98,10.8,11.34,10.36,11.0199995,12.24,11.36,11.759999,13.7699995,15.179999,16.16,17.5,18.71,20.279999,22.99,27.48,33.94,25.38,12.87,3.29,1.53,0.95,0.39999998,0.31,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.7,1.38,0.32,1.88,5.6099997,5.23,6.77,17.64,10.53,0.68,0.29,0.64,0.59999996,0.22999999,0.19,0.69,0.17999999,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.04,0.04,0.04,0.02,0.0,0.0,0.089999996,0.16,0.57,2.6399999,5.35,6.85,4.8199997,3.82,2.04,1.3399999,1.1999999,0.59999996,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.35999998,0.93,0.26,0.12,0.0,0.0,0.0,0.0,0.0,0.0,0.049999997,0.02,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.31,0.72999996,0.34,0.48999998,2.24,4.04,6.49,7.8399997,7.47,6.41,4.61,2.4099998,1.0799999,0.57,0.95,1.16,1.64,1.67,0.78,0.52,1.0699999,1.67,1.68,0.95,0.7,0.87,1.26,1.9399999,3.26,3.8999999,4.14,4.2799997,4.18,7.04,11.2,14.67,17.34,19.96,22.65,25.439999,28.63,38.95,49.61,42.46,25.63,13.9,13.0199995,9.349999,2.71,0.84999996,0.089999996,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.099999994,0.53,0.74,1.79,0.28,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.26,0.0,0.0,1.65,1.68,1.43,1.3,1.63,1.35,3.35,3.1599998,2.8,2.24,0.84999996,1.8,1.93,1.76,4.71,12.5,8.2699995,0.93,0.099999994,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.049999997,0.04,0.24,2.1299999,2.61,3.1499999,4.77,4.33,3.03,0.5,0.25,0.07,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.17999999,0.16,0.16,0.03,0.0,0.0,0.0,0.0,0.01,0.22,0.85999995,2.18,2.83,2.8899999,3.12,3.9399998,2.97,1.3299999,0.42999998,0.03,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02,0.099999994,0.26,0.58,1.87,3.6599998,3.78,3.4099998,3.1799998,2.53,1.89,1.15,0.63,0.45,0.19999999,0.16,0.12,0.04,0.01,0.07,0.099999994,0.03,0.07,1.36,3.99,3.98,4.0899997,4.0,2.75,3.04,3.6299999,4.5899997,5.43,5.6099997,7.52,9.389999,11.139999,13.83,14.929999,17.32,23.5,23.939999,21.31,18.039999,19.76,17.91,5.85,1.14,0.099999994,0.04,0.04,0.04,0.049999997,0.06,0.03,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13,2.1699998,2.6399999,0.35,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.11,5.5,17.98,13.799999,3.4199998,7.37,2.34,0.57,0.16,0.0,0.07,1.8399999,3.6599998,0.19,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.32,0.42,2.1299999,5.27,6.15,6.2599998,4.83,3.12,0.81,0.25,0.04,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.04,0.32,1.8499999,2.4199998,3.4199998,4.5899997,4.68,4.58,3.6299999,2.27,0.9,0.12,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.17999999,0.71999997,1.0699999,1.15,1.15,1.66,1.66,1.53,1.1,0.9,0.69,0.22,0.12,0.03,0.07,0.099999994,0.07,0.11,0.31,0.53,0.34,0.35999998,2.32,4.41,4.15,5.0099998,6.96,9.2699995,12.29,15.94,12.55,6.67,3.6,4.38,7.3399997,7.83,6.66,6.7799997,6.8599997,7.6499996,10.09,12.69,12.799999,11.21,6.21,1.5699999,0.17999999,0.03,0.03,0.08,0.12,0.22999999,0.13,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13,1.1,0.65999997,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.39999998,2.51,11.36,9.559999,8.25,5.46,4.92,0.14999999,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.099999994,0.59999996,1.49,2.6699998,2.55,4.7999997,6.69,5.79,4.0,1.1,0.08,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.08,0.03,0.04,0.37,1.13,1.9599999,2.6599998,2.84,2.09,1.0699999,0.42,0.089999996,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08,1.01,0.38,0.089999996,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14,0.58,1.16,1.24,1.0,0.87,0.75,1.06,1.23,0.74,0.34,0.12,0.099999994,0.01,0.03,0.089999996,0.21,0.59999996,1.31,1.5899999,1.36,0.97999996,1.42,2.97,4.1,5.72,7.0499997,10.11,12.48,10.88,6.06,3.59,2.35,3.54,5.97,7.74,9.389999,9.7699995,9.33,8.34,6.8599997,5.5299997,4.22,1.61,0.35,0.03,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.099999994,0.099999994,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.26,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.06,3.49,9.37,6.98,3.47,0.61,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.089999996,0.41,1.18,1.68,1.39,0.82,0.31,0.04,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.9,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08,0.28,0.57,0.64,0.29,0.25,0.16,0.099999994,0.29999998,0.37,0.28,0.22,0.17,0.049999997,0.07,0.38,0.61,0.93,2.24,4.02,3.8,3.29,3.23,4.46,6.25,6.52,5.33,3.1699998,1.78,1.56,2.18,3.26,3.9299998,4.23,5.1,4.99,3.76,2.6599998,1.67,0.48,0.19999999,0.24,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,6.3599997,12.37,5.58,0.0,0.0,0.19,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.19,1.03,0.37,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.26,1.8299999,4.0899997,5.0,4.95,2.83,0.32999998,0.24,0.04,0.04,0.06,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.049999997,0.28,0.53,0.32999998,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.12,0.28,0.52,0.44,0.21,0.04,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13,2.77,1.48,0.24,0.34,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.11,0.07,0.03,0.08,0.12,0.089999996,0.089999996,0.39999998,1.0699999,1.31,0.95,0.42,0.22999999,0.19,0.03,0.13,0.59,1.28,1.43,1.49,1.55,1.81,2.6399999,2.23,1.77,1.3199999,1.75,2.05,2.77,2.6599998,1.53,1.64,2.44,1.9599999,1.43,0.93,0.12,0.07,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,9.4,26.07,25.58,4.42,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06,0.61,2.29,5.54,7.97,10.54,12.15,8.809999,4.0099998,1.13,0.51,0.08,0.08,0.07,0.03,0.01,0.0,0.0,0.0,0.0,0.0,0.11,1.3299999,3.31,3.3999999,1.68,0.34,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.61,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.32,0.74,0.48,0.12,0.02,0.03,0.099999994,0.14999999,0.07,0.0,0.19999999,0.62,0.74,0.71,0.76,0.84,0.79999995,0.29,0.089999996,0.08,0.19,0.45,0.61,0.45,0.17999999,0.31,0.90999997,1.9599999,1.8199999,1.87,1.8199999,0.82,1.05,1.4699999,0.94,0.14,0.099999994,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.04,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02,0.0,0.12,0.34,0.38,0.53999996,0.93,1.49,2.1399999,2.96,3.7099998,7.22,11.63,11.05,3.9099998,1.87,14.2699995,7.71,0.0,0.0,0.0,0.0,0.0,0.0,0.93,1.26,7.29,29.98,6.69,0.77,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.11,0.29,0.56,0.9,2.2,4.0299997,7.85,12.73,15.0,12.13,5.9,1.56,0.29,0.06,0.06,0.08,0.06,0.0,0.0,0.58,1.4,0.79999995,0.26999998,1.24,4.0699997,6.73,5.4,2.54,0.55,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.32999998,0.59,0.35,0.08,0.089999996,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13,0.44,0.75,0.81,0.38,0.24,0.34,0.35,0.39999998,0.45,0.45999998,0.41,0.31,0.65999997,1.25,1.0799999,1.63,1.39,0.71,0.22,0.07,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.07,0.16,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.58,2.01,4.5899997,6.93,11.86,12.429999,14.16,12.5199995,13.4,15.28,15.15,11.01,9.71,3.8899999,3.36,12.54,26.189999,23.8,1.17,0.0,0.0,0.0,0.0,8.54,19.5,15.2699995,2.33,2.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02,0.02,0.0,0.0,0.07,0.41,1.3,3.26,6.37,8.309999,7.98,5.44,2.04,0.65,0.14,0.02,0.0,0.099999994,1.12,3.11,5.25,5.69,4.75,2.62,1.63,3.1899998,4.49,4.8599997,3.6699998,1.91,0.96,0.31,0.03,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06,0.76,9.83,2.1499999,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.049999997,0.11,0.17,0.29999998,0.35,0.089999996,0.0,0.0,0.0,0.099999994,0.14999999,0.21,0.35999998,0.45,0.47,0.55,0.66999996,0.77,0.82,0.78999996,0.75,0.59999996,0.53,0.39999998,0.68,0.89,0.64,0.32,0.13,0.03,0.03,0.01,0.0,0.0,0.0,0.01,0.03,0.17999999,0.56,0.66999996,0.61,0.39999998,0.19,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.26999998,0.29,0.32999998,0.88,1.01,1.61,4.49,2.9399998,2.55,4.35,4.19,0.0,0.0,0.0,0.0,0.0,0.79999995,2.76,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.11,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.049999997,0.38,1.79,0.11,0.049999997,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02,0.13,0.31,0.39,0.84,1.8,3.9099998,5.69,6.2799997,4.83,2.96,1.24,0.24,0.93,2.4199998,4.0099998,6.2,8.389999,9.5199995,11.469999,10.87,7.33,3.1799998,1.73,1.4499999,3.02,4.0699997,3.78,2.35,1.1,0.29999998,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.07,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.12,5.24,2.48,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02,0.42,0.53999996,0.17,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06,0.099999994,0.04,0.089999996,0.22,0.32,0.39,0.84999996,1.16,1.22,1.39,1.36,1.05,1.05,0.42,0.0,0.04,0.12,0.19,0.13,0.089999996,0.03,0.0,0.0,0.0,0.0,0.24,0.79999995,1.52,1.54,0.88,0.22,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.61,1.7099999,1.5799999,2.8,2.56,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.45,0.19,0.22999999,0.45999998,0.06,0.64,0.06,0.0,0.0,0.0,0.0,0.0,0.06,0.03,0.0,0.22999999,1.4599999,1.88,4.58,17.58,10.82,1.54,0.06,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.17,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.04,0.29,0.68,0.37,0.42,0.59,1.12,2.24,3.07,4.2799997,4.38,3.54,2.6699998,3.9399998,6.08,7.5299997,8.87,10.05,11.36,14.11,15.33,16.67,15.78,11.17,6.37,2.51,4.61,8.69,10.3,7.19,1.62,0.42,0.089999996,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02,0.08,0.08,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02,0.12,0.41,0.84999996,0.45,0.06,0.0,0.0,0.0,0.13,0.22999999,0.11,0.14999999,0.17999999,0.14,0.13,0.099999994,0.07,0.06,0.14,0.35999998,0.68,1.14,1.65,1.79,1.67,1.03,0.65999997,0.26,0.19999999,0.26999998,0.08,0.0,0.06,0.06,0.0,0.0,0.0,0.0,0.22999999,0.69,0.96999997,0.59,0.099999994,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.97999996,0.53999996,0.17999999,0.63,0.53999996,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.24,0.0,0.0,0.0,0.0,0.11,0.0,0.11,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.66999996,2.87,4.18,4.54,11.34,13.049999,2.75,0.45,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.21,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.17,0.59,1.3,3.0,5.72,8.28,6.71,5.8199997,7.98,12.13,14.309999,18.23,20.35,18.26,18.46,21.43,24.34,23.96,19.22,9.179999,8.73,12.69,13.61,6.97,2.6799998,1.25,0.39,0.099999994,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.04,0.14999999,0.29999998,0.29,0.03,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.03,0.0,0.0,0.0,0.06,0.34,0.56,0.24,0.04,0.099999994,0.089999996,0.049999997,0.049999997,0.08,0.08,0.11,0.089999996,0.11,0.29999998,0.95,1.23,0.96,0.85999995,0.79999995,0.39,0.31,0.17,0.07,0.39,0.19999999,0.07,0.0,0.0,0.0,0.02,0.19999999,0.34,0.29999998,0.07,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.45,0.81,0.0,0.0,0.0,0.0,0.0,0.0,0.08,0.44,0.61,0.68,0.78999996,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.09,0.14999999,0.01,0.0,0.16,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.22999999,1.09,2.35,2.6699998,4.69,6.43,6.3199997,6.99,9.349999,12.45,16.47,19.13,20.609999,20.449999,21.66,23.939999,27.019999,26.21,24.67,21.92,14.83,14.48,11.4,6.1,2.81,1.24,0.93,0.34,0.14999999,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06,0.42,0.75,0.90999997,1.7099999,2.8899999,3.9599998,7.08,2.59,0.049999997,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08,0.37,0.57,0.57,0.53,0.45999998,0.31,0.099999994,0.049999997,0.07,0.08,0.21,0.29999998,0.32,0.52,0.93,1.1999999,1.05,0.78,0.45,0.11,0.089999996,0.089999996,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.19,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.099999994,1.1999999,5.3399997,3.58,4.75,0.28,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.45,22.51,7.25,1.68,1.09,0.71,0.90999997,0.71,0.06,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.22999999,1.41,2.59,2.34,3.35,2.97,2.98,2.84,5.52,9.08,10.8,15.099999,17.9,18.9,20.23,23.57,26.71,28.34,27.43,21.699999,16.44,13.99,9.95,5.23,2.1399999,1.37,0.42,0.22,0.16,0.089999996,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.17999999,0.94,2.01,6.52,6.54,0.34,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.11,0.21,0.22,0.21,0.22999999,0.35,0.59,0.51,0.24,0.04,0.089999996,0.22999999,0.41,0.68,1.0,1.15,1.04,0.71,0.089999996,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07,0.71999997,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.9499999,10.349999,13.58,12.49,7.0299997,2.22,0.44,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,3.25,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.17999999,0.42999998,0.91999996,9.3,15.23,2.18,9.639999,28.46,20.84,1.26,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.17,0.08,0.17,0.13,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.099999994,0.65999997,1.56,3.25,4.24,3.57,1.99,1.9399999,2.34,4.1,6.7999997,11.349999,17.39,20.55,21.039999,16.56,15.549999,18.93,24.189999,23.9,23.449999,19.21,15.12,11.17,5.0699997,1.7199999,0.89,0.55,0.38,0.22,0.11,0.03,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.19999999,0.22,0.26,0.26,0.31,0.16,0.38,0.88,1.0799999,1.78,1.5699999,0.93,0.29,0.02,0.0,0.0,0.0,0.03,0.049999997,0.08,0.14999999,0.53,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.38,1.9699999,1.36,0.84,0.82,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.31,5.87,10.05,0.0,0.0,0.0,0.59999996,0.66999996,0.0,0.0,0.0,0.32999998,0.45999998,1.1999999,0.66999996,0.7,2.78,0.25,5.8799996,2.18,0.57,0.0,0.0,0.0,0.0,0.06,1.11,2.6,0.47,0.69,0.68,2.21,0.44,0.07,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06,0.22,1.01,2.8,3.34,3.12,2.72,2.6799998,2.69,2.73,5.96,13.78,22.06,30.449999,31.76,26.93,23.189999,24.33,26.46,25.83,23.74,19.88,16.59,11.2699995,5.08,2.34,0.90999997,0.48999998,0.35999998,0.32999998,0.25,0.17,0.099999994,0.03,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.04,0.12,0.17,0.17999999,0.17999999,0.12,0.06,0.099999994,0.08,0.049999997,0.03,0.01,0.0,0.16,0.41,0.7,0.81,0.51,0.31,0.07,0.02,0.0,0.03,0.089999996,0.16,0.29999998,0.68,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.19,0.7,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.90999997,8.94,7.3999996,0.75,0.03,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.53,5.08,0.0,0.0,0.0,0.0,1.5699999,2.56,0.0,0.0,0.32,0.45999998,1.16,0.53,0.26999998,0.55,0.17999999,0.16,0.0,0.0,0.0,0.0,0.0,0.0,0.13,0.089999996,0.19999999,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.04,0.35999998,0.19,0.13,0.04,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.04,0.03,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.19,0.52,0.63,1.24,2.3,3.05,3.28,4.68,4.7999997,3.9499998,3.08,5.72,11.34,21.0,30.849998,32.25,33.07,34.62,37.69,36.96,34.76,29.789999,21.449999,16.71,15.049999,10.099999,5.47,3.22,1.8199999,0.97999996,0.38,0.25,0.28,0.24,0.16,0.06,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.65999997,0.93,0.45,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.049999997,0.14,0.17999999,0.17,0.14,0.099999994,0.14,0.12,0.16,0.17,0.049999997,0.07,0.06,0.0,0.0,0.0,0.049999997,0.07,0.06,0.02,0.0,0.03,0.06,0.14999999,0.34,0.66999996,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.049999997,0.13,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,2.11,7.2799997,12.87,9.12,1.22,0.049999997,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13,0.38,0.04,0.35999998,0.19999999,0.35999998,0.65999997,0.45,0.0,0.0,0.0,1.93,9.36,4.97,0.04,0.0,0.0,0.0,0.0,0.0,0.0,0.049999997,0.82,0.56,0.35999998,0.48999998,0.84,3.27,4.22,1.6899999,0.96,0.03,0.0,0.049999997,0.0,0.0,0.0,0.0,0.0,0.0,0.049999997,0.099999994,0.03,0.0,0.0,0.0,0.0,0.0,0.0,0.02,0.39,1.1999999,1.28,1.5799999,2.34,3.21,4.68,5.93,6.6,5.83,5.56,5.66,8.55,15.799999,30.279999,43.17,48.079998,52.21,49.43,46.51,44.95,37.71,32.28,27.439999,21.01,15.61,12.7699995,9.16,6.0699997,3.79,2.01,1.05,0.48999998,0.22999999,0.21,0.14999999,0.089999996,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13,1.43,2.8799999,2.98,1.55,0.26,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.03,0.06,0.089999996,0.11,0.08,0.16,0.41,0.77,0.55,0.39,0.25,0.08,0.0,0.0,0.03,0.08,0.19999999,0.45999998,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.55,0.39999998,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.11,0.28,0.13,3.9499998,0.35,0.04,0.39,6.68,19.5,23.51,11.91,1.27,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.16,0.93,0.29999998,0.90999997,0.89,1.35,1.52,1.49,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.13,1.31,2.09,2.31,3.53,4.77,5.75,6.45,7.5899997,8.33,8.32,7.5,7.94,12.83,23.019999,40.14,50.3,57.96,56.48,55.12,48.079998,40.89,34.739998,30.73,25.699999,20.9,16.34,10.71,8.22,6.97,4.83,2.61,1.41,0.69,0.24,0.089999996,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14999999,0.89,1.4499999,0.47,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.26,0.51,0.63,0.61,0.71,0.65,0.65,0.35,0.12,0.06,0.14,0.32999998,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,4.22,9.679999,0.77,0.26999998,0.14,0.21,0.0,0.24,0.87,0.13,3.35,6.2799997,4.9,0.97999996,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08,0.38,1.81,1.0699999,0.89,0.13,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.59999996,1.36,2.08,2.5,5.23,6.04,6.29,7.46,9.83,12.24,12.57,12.849999,13.889999,18.69,28.18,41.55,51.239998,56.75,57.71,56.969997,49.379997,44.0,36.69,28.3,22.26,16.32,11.83,9.22,7.69,5.72,4.0299997,2.51,1.48,0.84999996,0.47,0.22,0.07,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02,0.02,0.03,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.04,0.26,0.53999996,0.55,0.24,0.06,0.28,0.35999998,0.47,0.65,0.79999995,0.0,0.0,0.0,0.02,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07,0.099999994,0.04,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,6.17,0.06,0.089999996,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.089999996,0.14999999,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.26999998,1.11,4.36,3.9299998,3.23,3.6499999,5.94,8.57,12.509999,15.73,17.539999,19.9,29.56,45.219997,56.149998,55.379997,50.48,46.62,48.17,48.879997,44.789997,38.5,29.56,21.46,14.259999,10.179999,8.13,6.08,3.8799999,2.7,1.8299999,1.36,0.84,0.39999998,0.099999994,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.049999997,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06,0.22,0.19999999,1.5,0.0,0.0,0.0,0.0,0.0,0.089999996,0.53,0.31,0.04,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02,0.0,0.35,0.53999996,0.61,0.78999996,1.0799999,0.0,0.0,0.0,0.19,0.55,0.25,0.0,0.0,0.0,0.03,0.049999997,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.48,0.64,0.14999999,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02,0.16,0.93,0.25,0.0,0.0,1.36,0.45,0.0,0.0,0.5,0.049999997,0.0,0.0,0.01,0.02,0.0,0.0,0.0,0.0,0.0,0.13,0.049999997,1.39,0.31,0.089999996,0.0,0.0,0.0,0.0,0.41,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.22999999,0.29999998,0.22999999,0.0,0.0,0.0,0.01,0.32999998,0.14,0.0,0.01,0.07,0.08,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.03,0.0,0.0,0.049999997,0.21,0.28,0.22999999,0.19999999,0.02,0.0,0.11,0.78,0.7,0.16,0.08,0.28,1.5,2.9099998,4.33,4.37,3.1499999,2.45,3.55,5.99,8.79,12.309999,16.44,27.08,40.78,51.55,52.239998,46.309998,42.07,47.14,50.219997,47.8,45.18,39.27,28.34,17.72,12.69,10.16,7.21,4.81,2.97,1.8499999,1.16,0.74,0.29,0.04,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08,0.11,0.04,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.16,0.0,0.0,0.08,0.84999996,1.03,0.41,0.12,0.0,0.0,0.0,0.0,0.0,0.01,0.03,0.03,0.02,0.07,0.089999996,0.14999999,0.099999994,0.089999996,0.13,0.19999999,0.17,0.14999999,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.02,0.04,0.14999999,0.29999998,0.52,0.76,0.0,0.0,0.0,0.11,1.12,0.98999995,0.29,0.0,0.0,0.0,0.099999994,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.04,0.03,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.04,0.03,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.32,0.32,0.08,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.17999999,0.24,0.0,0.0,0.03,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.09,9.34,9.7699995,0.37,0.0,0.0,0.0,0.82,2.71,0.06,0.0,0.0,0.0,0.0,0.0,0.0,0.13,0.39999998,0.17,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.099999994,0.04,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.07,0.04,0.0,0.11,0.45,0.53,0.5,0.41,0.19,0.19999999,1.04,2.26,2.86,1.8,0.44,0.0,0.5,1.1,1.22,1.4599999,1.8199999,3.62,4.2599998,4.49,4.8599997,7.08,10.37,15.74,29.019999,40.51,50.84,55.149998,48.16,45.309998,46.2,51.07,50.84,41.399998,28.939999,21.789999,16.869999,12.61,8.22,4.98,3.08,1.78,1.03,0.59,0.14999999,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08,0.32,0.16,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13,0.32999998,0.45999998,0.48999998,1.22,0.13,0.0,0.22999999,0.0,0.07,0.35999998,0.66999996,0.35999998,0.42,0.07,0.14999999,0.63,0.35,0.02,0.0,0.089999996,0.42999998,0.58,0.17,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.02,0.01,0.01,0.02,0.02,0.049999997,0.24,0.26999998,0.0,0.0,0.0,0.02,0.45,1.5799999,1.27,0.38,0.0,0.0,0.07,0.07,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.049999997,0.17,0.13,0.0,0.0,0.29,0.22,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.11,0.79999995,1.01,0.099999994,0.03,0.04,2.1499999,1.37,0.0,0.0,0.0,0.0,1.5999999,0.14,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14,0.31,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.22,0.89,0.61,0.78999996,0.55,0.12,0.0,0.0,0.0,0.17,0.19999999,0.13,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.14,0.25,0.32999998,0.29999998,0.26,0.65999997,1.8,3.6799998,5.71,6.7,4.63,0.71999997,0.01,0.04,0.06,0.71,2.26,5.25,6.21,4.77,3.98,5.81,7.99,13.07,24.35,36.98,48.559998,51.02,46.26,44.989998,49.309998,49.71,46.01,37.01,27.55,19.779999,15.33,12.04,8.19,4.14,2.49,1.49,1.22,0.64,0.19,0.03,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02,0.17,0.26,0.099999994,2.74,4.56,3.1499999,1.28,4.69,1.26,0.84,3.3899999,3.47,1.23,1.01,1.05,1.15,1.0699999,0.76,0.64,0.11,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.02,0.01,0.01,0.02,0.01,0.03,0.03,0.08,0.0,0.0,0.0,0.0,0.03,1.0,3.07,1.64,0.19,0.0,0.02,0.12,0.07,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.049999997,0.14999999,0.28,0.14999999,0.0,0.08,0.35999998,0.35,0.08,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.71,0.5,0.25,0.24,0.089999996,0.049999997,0.03,0.0,0.0,0.0,0.0,0.22999999,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02,0.26,1.36,2.05,2.51,3.03,0.88,1.36,1.56,0.26,0.0,0.0,0.26999998,1.13,1.53,1.6899999,1.5799999,0.72999996,0.11,0.0,0.0,0.78,1.5999999,4.63,5.2799997,2.72,0.95,0.39999998,0.26999998,0.34,0.28,0.08,0.16,0.16,0.089999996,0.099999994,0.11,0.38,1.6899999,2.75,3.97,6.1,8.11,8.82,5.8399997,1.4499999,0.16,0.22,0.25,0.90999997,2.54,3.3999999,3.79,3.6899998,4.7599998,5.95,9.59,19.0,29.07,36.13,41.28,40.28,42.51,43.34,42.809998,37.559998,32.059998,25.63,17.699999,13.42,10.19,6.48,3.5,1.8,1.05,0.7,0.44,0.19,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02,1.04,3.55,3.11,6.15,14.58,12.38,6.18,4.42,4.68,6.94,10.69,8.05,3.6699998,2.53,1.38,1.0,0.48999998,0.84,1.14,0.17,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.03,0.03,0.03,0.03,0.02,0.03,0.04,0.0,0.0,0.0,0.0,0.0,0.08,1.8199999,3.9099998,2.46,0.42999998,0.0,0.0,0.12,0.22999999,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.11,0.06,0.26999998,0.29999998,0.08,0.02,0.48999998,0.69,0.58,0.51,0.34,0.21,0.13,0.03,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.29999998,0.03,0.0,0.0,0.0,0.07,0.07,0.24,0.93,1.37,1.18,2.12,2.78,5.2999997,3.9599998,1.99,3.06,2.6499999,5.49,3.6299999,3.56,3.3799999,1.53,1.17,1.4499999,2.22,2.3899999,0.55,0.0,0.0,0.0,0.34,1.39,1.7099999,0.81,0.91999996,0.71,0.85999995,0.90999997,0.28,0.19999999,0.13,0.12,0.08,0.11,0.24,1.5999999,3.27,3.75,3.8899999,4.5499997,7.8399997,8.559999,7.89,3.87,0.45,0.35999998,0.099999994,0.26999998,1.66,3.55,5.54,6.97,4.65,4.7599998,6.5299997,11.54,18.97,28.609999,32.5,33.69,34.36,39.52,39.25,34.89,27.49,21.38,17.02,13.599999,10.099999,7.2,4.6,2.53,1.54,0.84,0.35999998,0.14999999,0.02,0.13,0.17,0.04,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13,0.21,0.62,0.76,0.47,2.51,4.66,4.17,5.45,4.35,5.6099997,5.45,7.37,6.7,4.5299997,3.03,1.09,0.32,0.22,0.08,0.049999997,0.13,0.24,0.089999996,0.19999999,0.39999998,0.0,0.0,0.0,0.13,0.29,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.02,0.0,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.11,2.21,4.66,4.5099998,1.87,0.099999994,0.0,0.13,0.14999999,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02,0.17,0.17999999,0.48999998,0.66999996,0.26999998,0.0,0.71999997,1.39,1.5,2.52,2.52,2.24,1.9799999,1.37,1.01,1.05,0.84999996,0.63,0.45999998,0.25,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.099999994,0.17999999,0.17,0.34,0.06,0.0,0.06,0.07,0.089999996,0.35999998,0.72999996,1.81,4.02,1.5999999,0.32999998,0.78,1.5799999,2.8,0.78999996,1.36,2.01,6.33,9.19,10.139999,9.09,5.1,3.78,4.15,2.72,1.76,2.47,0.58,0.14,0.0,0.0,0.08,0.75,0.89,0.96999997,1.41,1.3299999,1.3399999,0.48,0.04,0.07,0.11,0.13,0.24,1.17,2.0,3.6299999,5.19,6.98,6.92,6.33,5.5899997,4.7599998,3.79,2.8899999,2.11,1.29,0.45,0.17999999,0.66999996,2.54,4.45,5.45,5.19,5.3399997,6.2999997,9.01,13.33,18.529999,22.23,28.769999,31.65,36.18,38.03,34.32,26.81,20.71,17.0,14.559999,11.679999,9.04,7.19,4.8199997,2.47,1.09,0.32,0.049999997,0.01,0.08,0.16,0.03,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.39999998,1.14,0.089999996,0.0,0.13,2.35,4.44,4.2,2.45,3.59,3.6599998,3.55,3.8899999,2.84,3.4499998,2.37,0.82,0.32999998,0.19,0.0,0.0,0.0,0.0,0.29999998,1.0699999,1.1899999,0.68,0.19,0.099999994,0.04,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.049999997,1.1,4.0499997,3.56,1.56,0.089999996,0.11,0.14999999,0.07,0.47,0.06,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.089999996,0.42999998,0.42999998,1.4599999,1.43,0.0,0.0,2.26,2.96,3.3999999,5.56,5.5499997,5.7999997,5.2999997,3.98,3.99,3.7099998,3.1399999,2.57,2.21,0.96,0.32,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.53,0.97999996,0.02,0.17999999,0.089999996,0.71,1.31,1.26,0.66999996,0.79999995,1.4,3.8,2.8799999,0.5,0.14999999,0.0,0.0,3.1299999,6.16,7.7599998,11.65,11.83,10.04,6.98,3.4199998,4.77,6.42,6.39,4.88,5.0099998,4.4,1.5899999,0.25,0.0,0.04,0.71,2.8799999,2.3999999,2.28,2.1,2.59,1.4,1.3299999,0.83,0.42999998,0.01,0.099999994,0.48,2.48,5.68,7.74,8.15,10.17,9.66,10.13,7.0899997,2.48,1.3,2.46,4.31,5.06,1.31,0.32999998,0.29,0.88,2.7,3.53,4.31,5.21,7.12,8.95,10.03,12.15,19.97,25.75,30.269999,32.27,29.98,27.849998,25.46,20.14,15.69,12.83,10.219999,8.42,5.8199997,3.4299998,1.87,0.59999996,0.049999997,0.19999999,0.07,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.03,0.04,0.06,0.17999999,0.13,0.17,0.35,0.12,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.089999996,0.56,0.25,0.78,0.59,0.53999996,0.35999998,0.65999997,0.76,0.11,0.02,0.12,0.22,0.26,0.44,0.42999998,0.28,0.21,0.42999998,0.39999998,0.32999998,0.19,0.049999997,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.099999994,0.96,2.3899999,3.09,2.3799999,1.49,0.94,0.08,0.79999995,0.9,0.13,0.0,0.0,0.0,0.0,0.03,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.12,0.59,0.66999996,2.29,2.08,0.0,0.0,3.4099998,4.58,5.56,7.9199996,7.5499997,8.13,6.87,5.47,6.16,5.68,5.15,5.06,3.56,1.48,1.06,0.69,0.31,0.14999999,0.049999997,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02,0.04,0.0,0.29999998,0.44,0.9,0.099999994,0.57,2.11,2.71,3.4399998,3.83,3.6599998,2.8,0.95,0.63,0.44,0.56,1.77,2.6799998,3.4099998,8.82,15.089999,21.42,24.18,20.91,15.049999,7.0,5.17,5.9,6.8399997,7.6699996,8.139999,5.98,2.49,1.25,0.71999997,0.78,0.56,1.01,2.21,6.1299996,6.68,6.02,6.52,5.91,7.8599997,8.41,2.4199998,1.68,2.22,5.45,11.73,13.88,13.139999,14.44,14.009999,11.21,11.259999,7.19,3.8,3.3999999,5.69,6.85,5.67,2.1299999,0.45999998,0.03,0.26,1.3199999,1.8199999,3.35,5.48,5.14,9.179999,11.969999,13.719999,17.42,20.67,27.59,28.47,25.289999,21.41,18.55,15.799999,12.21,9.82,8.28,5.74,3.84,3.1,2.36,1.17,0.77,0.47,0.12,0.0,0.0,0.0,0.0,0.04,0.049999997,0.099999994,0.12,0.29,0.29999998,0.41,0.66999996,0.17,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.03,0.06,0.099999994,0.13,0.08,0.07,0.53,0.35,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.17,0.85999995,1.88,5.6,3.9499998,2.05,0.72999996,0.13,0.59,0.94,0.22999999,0.0,0.0,0.0,0.099999994,0.41,0.06,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.17999999,0.79999995,0.90999997,3.51,3.1699998,0.0,0.0,4.56,6.06,7.33,9.51,9.66,10.19,7.7799997,7.2999997,7.98,6.85,6.73,6.47,3.9099998,2.61,3.04,2.84,2.18,1.55,0.84,0.42,0.13,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.089999996,0.11,0.42999998,0.37,0.35,0.48,0.0,0.0,0.53999996,0.89,0.91999996,2.75,3.35,3.48,4.62,3.02,2.35,2.44,3.01,4.0899997,9.04,11.179999,13.23,17.63,21.289999,21.859999,23.64,22.83,21.41,18.47,20.029999,21.21,13.049999,5.56,1.25,0.59999996,2.19,3.51,2.48,3.06,3.75,3.9399998,5.12,4.94,4.75,6.79,10.33,14.21,13.679999,8.46,6.8599997,8.98,9.48,8.01,6.12,5.37,12.7,19.859999,13.349999,10.75,6.46,4.72,8.23,10.2699995,10.73,5.58,1.66,0.57,0.39999998,0.26999998,0.38,1.75,4.14,3.82,3.6699998,8.69,15.99,16.75,15.62,16.0,21.89,27.289999,29.63,25.18,19.59,13.5,8.95,6.5499997,4.94,4.54,4.75,4.5,3.8799999,2.69,1.79,0.9,0.25,0.0,0.099999994,0.11,0.22999999,0.26999998,0.17999999,0.19,0.26999998,0.21,0.17999999,0.22999999,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.12,0.42,0.66999996,0.81,1.53,1.8399999,1.55,2.1699998,2.2,0.24,0.08,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.52,3.04,6.3799996,3.4299998,1.87,1.26,0.28,0.53999996,0.53999996,0.0,0.08,0.02,0.049999997,0.5,0.71999997,0.03,0.0,0.0,0.0,0.0,0.0,0.089999996,0.68,0.48,0.14999999,0.03,0.0,0.0,0.0,0.21,0.90999997,0.93,3.7099998,3.25,0.11,0.03,4.63,6.19,7.5899997,10.78,11.599999,11.55,9.15,9.58,9.5,8.42,8.349999,7.18,4.04,3.75,3.1799998,3.11,3.27,2.18,1.41,1.0799999,0.78,0.38,0.32999998,0.48999998,0.64,0.81,0.59,0.94,0.87,0.91999996,0.65,0.34,0.13,0.0,0.0,0.0,0.0,0.0,0.02,0.42999998,0.37,0.52,0.13,0.0,0.0,0.0,0.0,0.0,0.12,0.39999998,1.1899999,1.77,2.31,4.22,6.89,7.94,9.69,11.28,10.17,8.0199995,10.01,11.07,18.17,26.56,33.5,37.219997,36.71,35.48,32.82,26.31,12.91,2.8899999,4.6,5.43,7.29,8.48,8.889999,10.48,12.469999,13.259999,14.11,17.369999,16.19,13.849999,12.059999,10.76,7.54,6.74,9.5199995,10.45,9.5199995,8.4,6.54,5.3199997,7.0099998,12.889999,14.299999,11.809999,8.2699995,9.7699995,12.73,13.0199995,10.41,5.69,3.3899999,3.35,3.6,1.88,1.05,1.51,0.77,0.78999996,2.77,8.349999,14.53,17.16,13.5,13.15,14.69,19.74,26.25,29.51,29.289999,20.91,13.88,9.3,6.54,4.8199997,3.8899999,3.21,2.56,2.74,2.97,1.75,0.9,0.77,0.55,0.04,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02,0.03,0.07,0.08,0.13,0.11,0.29999998,1.1,2.02,0.32999998,0.14,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13,1.36,1.7199999,1.23,2.77,1.36,0.08,0.04,0.0,0.07,0.13,0.099999994,0.5,0.96999997,0.19999999,0.089999996,0.61,0.0,0.0,0.0,0.14999999,0.52,1.15,0.96,0.26999998,0.24,0.07,0.099999994,0.12,0.58,0.71999997,2.8899999,2.46,0.42999998,0.0,2.83,4.41,6.2,10.099999,11.53,9.86,9.48,11.179999,9.78,9.469999,9.61,6.18,3.6799998,3.4199998,3.23,3.25,1.9399999,1.53,1.02,1.04,0.78999996,0.78999996,2.06,3.29,3.9499998,4.08,3.99,4.5099998,4.4,4.36,3.86,3.4299998,2.01,0.81,0.17,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.11,0.03,0.55,0.16,0.01,0.11,1.5799999,2.6299999,5.91,9.78,10.5199995,11.46,12.45,10.809999,5.97,3.81,5.74,5.73,11.599999,14.49,21.01,28.58,31.05,32.5,28.81,31.98,18.699999,12.57,12.259999,13.099999,14.219999,12.98,11.04,12.44,14.46,17.529999,22.029999,22.08,18.23,12.36,6.7799997,2.9199998,2.11,2.96,5.81,7.49,7.79,7.0,6.41,4.92,4.54,6.6499996,13.13,18.82,16.71,15.49,14.33,13.929999,8.82,5.42,5.15,9.2699995,10.58,6.0299997,1.48,0.35,0.56,1.42,3.1399999,6.46,12.32,15.599999,11.42,9.48,10.01,12.08,20.34,23.74,29.939999,30.21,23.22,15.7699995,9.73,6.6099997,3.74,2.62,2.3,2.6499999,3.32,3.23,2.73,1.6899999,0.22,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.9799999,0.95,2.69,1.78,0.81,0.0,0.0,0.03,0.06,0.19,0.19,0.42,0.13,0.0,1.9799999,0.29,0.0,0.0,0.0,0.099999994,1.52,3.6,1.14,0.72999996,2.24,0.7,0.06,0.22,1.9799999,2.37,4.73,0.85999995,0.79999995,3.8899999,5.3599997,5.33,8.679999,9.12,6.17,6.97,8.11,8.63,8.2699995,7.99,4.35,4.42,3.47,4.71,2.9199998,1.1999999,0.35999998,0.78999996,0.68,0.56,1.4,2.6799998,3.24,3.9099998,4.08,4.23,4.56,4.31,4.41,4.87,4.29,3.34,2.55,1.92,1.11,0.65,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02,0.02,0.0,0.25,1.0799999,1.1,1.06,3.11,4.23,6.93,10.07,8.559999,9.92,14.65,12.19,5.6299996,4.36,4.92,3.3899999,5.7799997,8.84,13.889999,23.82,28.57,21.67,27.13,34.96,33.78,17.369999,9.099999,7.95,8.36,8.36,9.24,11.07,20.74,30.96,33.739998,27.99,22.029999,17.029999,11.36,5.27,1.9399999,1.38,3.73,6.49,6.85,7.21,7.5699997,6.77,4.88,3.76,4.15,11.37,22.41,25.06,20.279999,15.219999,12.7,12.0,9.48,9.19,13.21,14.61,9.9,1.9,0.78999996,0.65999997,0.35999998,1.36,2.8999999,5.5699997,9.78,11.469999,10.58,9.099999,9.139999,14.839999,19.97,22.369999,24.939999,24.88,20.609999,13.24,9.05,4.91,2.6299999,1.91,2.2,1.6999999,2.1,1.61,1.0799999,2.34,1.89,0.7,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.04,0.0,0.07,0.12,0.0,0.0,0.0,0.08,0.35999998,0.14,0.03,0.08,0.39,1.5,1.15,0.71999997,0.089999996,0.0,0.21,0.48999998,0.17999999,0.13,0.12,0.68,1.53,2.46,0.79999995,0.0,0.0,0.0,0.32,0.71,0.34,0.089999996,3.08,11.37,1.38,0.0,0.25,3.9099998,4.83,4.96,2.57,9.66,15.7699995,19.199999,12.7699995,8.809999,9.4,8.33,8.54,9.5,9.4,7.8799996,4.2999997,4.73,3.9499998,5.64,3.74,1.38,0.39,1.13,0.84999996,0.65,1.51,2.6799998,3.75,4.7599998,4.1,4.31,3.8899999,3.6399999,3.1799998,2.59,2.22,2.23,1.81,1.1999999,1.56,1.87,2.2,1.02,0.28,0.0,0.0,0.0,0.0,0.14,0.17,0.04,0.0,0.0,0.42999998,1.0,1.79,4.75,5.74,6.1,6.22,7.2599998,8.809999,13.69,14.48,10.809999,8.55,3.4399998,0.82,4.5,9.719999,14.509999,19.84,21.97,17.59,16.449999,26.73,27.16,21.16,12.25,8.72,7.45,8.07,9.95,12.59,16.21,22.33,30.779999,31.25,26.31,20.33,16.58,11.759999,6.0299997,2.87,2.35,3.1499999,3.54,4.94,7.75,7.83,5.5899997,4.3399997,4.68,6.31,8.71,14.0199995,19.32,19.25,18.84,18.68,17.359999,19.539999,20.699999,18.24,15.45,10.349999,4.6,1.11,0.29,0.14999999,0.41,2.02,3.9499998,9.5,14.61,15.549999,11.88,8.2699995,8.75,12.059999,16.449999,20.42,20.39,17.06,13.13,8.59,4.8399997,2.73,1.4399999,1.3399999,1.26,0.47,0.53,1.02,2.02,2.32,1.9599999,1.51,0.90999997,0.42999998,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08,0.0,0.0,0.0,0.17,0.34,0.62,0.25,0.0,0.0,0.17999999,1.1999999,3.4499998,2.74,0.13,0.06,0.59999996,1.02,0.37,0.03,0.02,0.01,1.4499999,1.91,0.53999996,0.61,1.9,3.1499999,2.4099998,0.12,0.0,0.0,0.0,0.16,0.37,0.19999999,0.11,3.83,13.37,0.82,0.0,0.11,1.52,5.6,2.82,3.97,11.469999,19.039999,30.13,23.689999,15.509999,11.62,10.73,13.24,12.09,10.95,12.889999,11.559999,11.34,7.95,6.14,3.4399998,1.36,1.75,1.26,0.65,1.68,3.1299999,4.15,4.6,3.29,4.2599998,4.5,4.5699997,3.6299999,2.6399999,2.22,2.37,2.22,1.8199999,1.8499999,1.14,0.55,0.52,1.1,1.22,0.41,0.049999997,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.22999999,2.06,4.87,11.15,11.0199995,8.46,6.99,9.75,9.929999,7.3199997,6.7799997,2.84,3.06,4.47,3.82,7.69,13.2699995,11.13,10.48,7.1499996,6.8399997,10.03,8.22,8.01,8.47,8.42,7.52,8.349999,11.83,12.15,13.799999,14.66,15.61,18.09,15.7,11.62,11.09,9.7,7.2799997,4.0699997,3.32,3.4199998,4.16,5.3399997,6.15,5.41,4.38,4.49,6.62,9.83,8.8,6.0099998,9.13,15.49,23.23,25.779999,20.42,20.34,24.8,25.46,19.35,15.33,8.29,2.9199998,0.89,0.03,0.21,1.4399999,3.01,8.72,12.45,18.09,16.58,9.75,7.69,9.0,15.799999,16.16,14.44,10.84,9.34,7.31,6.1099997,3.9599998,2.57,0.7,0.03,0.0,0.089999996,0.41,0.78999996,1.16,1.22,1.29,1.61,1.49,0.98999995,0.91999996,0.66999996,0.17,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.099999994,0.0,0.0,0.0,0.42999998,0.12,0.07,0.0,0.07,0.089999996,0.7,1.15,0.14999999,0.0,0.0,0.17,4.5299997,7.6,0.85999995,0.77,0.28,0.32999998,0.66999996,0.17,0.19,0.17999999,1.56,4.7999997,1.3199999,0.56,2.62,3.1699998,2.9099998,0.08,0.0,0.0,0.0,0.0,0.0,0.14999999,0.78999996,2.6499999,5.73,0.52,0.01,0.0,1.4699999,3.58,2.29,1.39,8.63,11.259999,12.53,13.49,11.96,7.47,6.8999996,9.82,11.49,12.21,14.98,18.25,15.78,12.54,7.39,4.62,3.9199998,4.54,3.36,3.83,4.2599998,4.68,5.4,4.48,5.24,3.72,1.88,1.3,0.48,0.24,0.77,2.02,1.5999999,1.75,2.1699998,1.8499999,1.86,0.59,0.9,1.4399999,1.22,0.89,1.2099999,0.84999996,0.72999996,0.52,0.52,0.16,0.14,0.0,0.0,0.0,0.38,1.36,3.7099998,5.37,4.37,7.72,9.75,8.32,3.6999998,2.09,0.06,0.13,1.56,3.1699998,2.22,6.7799997,10.24,9.389999,6.81,3.4399998,2.52,5.2799997,7.06,7.18,8.91,8.22,5.8199997,5.69,6.56,6.22,5.48,5.12,6.19,5.71,5.41,7.2799997,7.43,7.31,5.43,4.83,5.89,6.58,6.19,4.71,4.92,4.56,3.81,4.5299997,6.22,9.41,8.25,4.94,4.58,9.53,16.94,20.4,17.84,15.69,17.65,22.13,22.48,24.31,16.56,8.53,1.9799999,0.26999998,0.0,0.65999997,1.67,3.74,9.26,16.68,19.35,17.05,15.73,17.41,16.77,18.119999,14.63,10.88,8.88,7.6699996,6.0099998,4.08,1.75,0.41,0.04,0.01,0.0,0.049999997,0.11,0.24,0.35999998,0.5,0.51,0.39,0.32,0.22999999,0.089999996,0.06,0.049999997,0.04,0.11,0.07,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.25,0.29,0.21,0.0,0.04,0.04,0.07,0.08,0.19,0.38,1.77,1.63,0.87,0.17999999,0.02,0.13,0.0,0.0,0.0,0.17,2.1599998,1.3299999,0.03,0.0,0.0,0.76,4.0,0.98999995,0.96,0.25,0.0,0.51,0.35999998,0.94,1.1899999,2.05,3.99,2.49,0.61,3.37,2.81,1.4599999,0.0,0.0,0.0,0.0,0.0,0.0,0.29999998,2.23,1.49,2.6,0.35,0.0,0.22999999,2.01,1.3399999,0.37,1.35,3.1,4.67,3.25,3.84,4.48,3.62,2.71,4.0299997,5.17,6.35,8.559999,14.799999,11.059999,7.37,4.71,2.49,3.53,7.98,10.639999,9.559999,6.06,3.55,2.28,4.33,1.87,0.5,0.35999998,0.7,1.65,2.47,4.5699997,6.18,5.87,5.8799996,6.52,5.83,4.56,2.75,1.99,1.29,1.61,1.31,1.74,1.8,1.56,1.7099999,2.46,1.78,1.3299999,0.42,0.22,0.03,0.0,0.0,0.06,0.57,1.37,1.03,4.6,3.6699998,2.81,1.23,1.9799999,5.0699997,5.43,4.71,5.2999997,6.49,9.04,10.639999,12.7699995,13.0199995,9.78,9.639999,12.2,11.889999,12.79,16.029999,13.92,7.7,5.22,2.9199998,2.0,1.03,1.27,1.49,2.26,5.3599997,4.89,5.5,6.66,7.79,11.429999,10.69,9.07,7.79,7.0899997,7.04,7.4199996,6.08,3.97,3.58,3.9499998,4.37,4.46,4.0699997,6.95,9.23,12.65,12.4,11.86,14.28,15.7699995,21.66,27.3,24.939999,13.759999,5.27,0.53,0.03,0.01,0.66999996,1.48,5.37,12.82,21.109999,27.09,24.34,26.539999,24.58,19.66,15.16,10.75,9.23,7.3399997,5.24,3.48,2.25,1.31,0.91999996,0.55,0.21,0.01,0.0,0.0,0.02,0.07,0.089999996,0.11,0.099999994,0.02,0.0,0.04,0.14,0.21,0.39,0.32,0.28,0.12,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.16,0.08,0.0,0.25,2.37,3.79,1.03,0.01,0.01,0.01,0.01,0.01,0.04,0.41,0.35999998,0.16,0.0,0.0,0.0,0.0,0.0,0.0,0.07,0.83,1.24,0.0,0.0,0.0,0.11,0.57,0.19,0.089999996,0.39,0.16,0.57,1.05,2.79,1.68,1.37,4.49,1.48,0.39,0.52,0.39,0.29,0.0,0.0,0.0,0.0,0.0,0.0,0.32999998,1.3299999,1.01,3.26,1.15,0.55,0.71999997,3.54,2.4299998,0.84,1.8199999,7.1499996,9.67,8.55,5.96,5.3599997,5.29,7.1099997,7.6499996,10.58,7.14,10.4,16.19,10.62,8.78,4.49,4.75,5.98,5.45,5.31,3.59,1.01,2.6,2.83,1.27,0.58,1.5799999,3.23,4.1,5.45,6.66,8.07,11.219999,11.139999,9.179999,6.58,5.72,4.47,4.3199997,1.8,1.35,1.15,0.78999996,1.1899999,1.35,0.97999996,1.54,1.42,1.23,1.22,0.77,0.14999999,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.96999997,3.22,4.71,5.89,5.66,8.78,10.15,11.13,9.03,9.889999,9.21,9.28,12.54,14.19,13.2699995,11.83,12.179999,14.34,16.89,19.029999,20.64,20.109999,15.24,9.349999,5.44,3.7099998,3.8,4.54,5.35,2.57,2.57,4.5899997,5.89,7.77,10.34,11.259999,11.8,11.11,9.12,10.679999,11.37,11.849999,10.37,6.2,3.6499999,4.2,4.72,5.64,5.52,7.1099997,7.19,7.6099997,8.92,10.08,11.75,13.179999,16.91,19.91,21.84,15.429999,7.8199997,1.24,0.11,0.06,0.24,1.26,4.14,11.61,22.43,30.179998,31.73,27.01,19.08,12.04,8.83,9.679999,11.349999,12.4,10.41,7.87,5.71,4.42,2.99,2.27,1.9,1.66,1.03,0.35,0.07,0.0,0.03,0.06,0.12,0.12,0.08,0.01,0.0,0.0,0.0,0.0,0.0,0.01,0.02,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.11,0.12,0.14999999,0.59,1.99,6.81,9.11,2.21,0.84999996,1.14,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.099999994,0.0,0.0,0.0,0.0,0.0,0.0,0.16,0.04,0.0,0.0,0.02,0.57,0.96999997,1.17,0.04,0.26,0.5,0.57,0.38,2.56,3.04,0.85999995,3.1699998,1.4399999,0.41,0.34,0.62,0.13,0.0,0.0,0.0,0.0,0.0,0.0,0.42,0.53999996,0.58,3.82,1.81,1.74,2.72,4.0299997,0.52,0.77,1.9599999,2.79,6.98,10.61,3.4099998,2.3999999,8.09,10.679999,6.25,6.2999997,7.7999997,11.03,8.8,4.72,8.349999,13.32,12.059999,6.6299996,2.6,0.78,0.48,4.36,7.68,9.599999,8.84,7.2,7.91,6.67,5.5899997,8.389999,11.34,12.45,11.179999,8.86,4.58,2.03,1.49,1.16,1.14,0.37,1.68,0.39,0.29,0.16,0.07,0.26999998,0.16,0.25,0.089999996,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.22999999,1.1,1.27,2.57,4.56,8.33,9.41,9.4,9.23,7.1499996,8.99,12.65,13.78,12.73,10.639999,10.63,12.86,14.87,15.63,16.38,16.39,13.049999,9.46,7.16,6.6,6.5699997,7.39,3.75,2.9399998,2.02,2.8,4.0099998,5.06,4.97,7.1,9.9,12.15,12.45,15.17,16.869999,15.66,12.61,8.41,7.0499997,8.44,6.72,6.49,4.85,4.92,6.37,6.54,5.98,6.46,6.99,7.9199996,10.5199995,12.75,16.199999,16.76,10.429999,4.85,1.24,0.83,1.77,3.1499999,6.2,12.09,21.06,25.33,25.92,20.16,12.559999,10.33,13.11,15.73,16.539999,15.57,14.49,14.82,15.639999,15.0199995,11.92,8.679999,4.93,4.46,2.61,1.4699999,0.22,0.07,0.0,0.02,0.07,0.19999999,0.28,0.47,0.7,0.77,0.26999998,0.0,0.01,0.08,0.25,0.31,0.14999999,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.53999996,6.87,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.29,0.55,0.75,0.89,1.12,1.4,7.17,11.74,1.42,10.04,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.049999997,0.03,0.07,0.0,0.0,0.0,0.0,0.0,0.02,0.22,0.089999996,0.17999999,0.74,2.01,2.69,1.35,0.68,0.58,0.79999995,0.03,0.61,0.68,0.39999998,0.81,0.31,0.53999996,0.41,1.06,0.28,0.089999996,0.099999994,0.0,0.0,0.089999996,0.17999999,0.19,0.38,0.84999996,3.22,1.09,2.36,7.1,2.71,0.32999998,2.08,1.8399999,0.19,4.42,10.44,1.49,8.32,10.42,4.97,2.24,3.06,7.8199997,8.82,2.98,8.349999,11.78,10.59,9.34,6.0499997,2.76,2.53,11.13,13.25,13.92,15.179999,15.28,15.69,13.73,9.44,7.12,8.96,9.09,7.74,3.53,1.68,0.98999995,0.19999999,0.11,0.049999997,0.06,0.0,0.94,0.32999998,0.45,0.04,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.79999995,0.48,2.02,2.61,2.56,3.6499999,5.13,5.13,5.21,6.69,7.0,6.69,6.79,7.25,7.12,8.389999,10.08,11.15,10.42,8.92,9.69,8.0,5.8599997,6.62,5.21,2.8899999,1.9699999,2.54,3.36,2.32,2.23,3.73,6.18,10.38,14.049999,15.32,17.77,22.76,21.41,16.67,14.7,14.389999,12.3,9.09,5.74,4.49,6.0899997,5.0699997,4.62,3.9199998,2.8899999,3.23,5.6099997,9.7699995,15.429999,17.55,18.21,17.18,13.0,7.2999997,3.4199998,3.27,4.5499997,7.35,11.37,14.2699995,14.299999,13.23,10.2699995,9.12,12.19,14.57,14.86,14.23,15.219999,18.16,20.32,20.97,21.43,21.5,21.46,19.18,12.969999,7.68,2.09,0.39999998,0.089999996,0.06,0.06,0.049999997,0.08,0.089999996,0.11,0.099999994,0.0,0.0,0.0,0.03,0.12,0.03,0.099999994,0.07,0.13,0.22,0.31,0.19,0.04,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,8.2,12.809999,0.089999996,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.12,0.11,0.099999994,0.17,0.14,2.51,4.98,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.01,0.0,0.26,0.94,0.96999997,0.75,0.93,2.1499999,3.75,6.64,7.75,2.73,0.56,0.57,0.74,0.48,1.62,0.37,0.85999995,0.14999999,0.29,0.07,1.37,1.22,0.04,0.0,0.08,0.25,0.22999999,1.0,1.66,2.73,0.42999998,0.59999996,1.7099999,0.53,0.049999997,1.48,0.94,0.04,0.91999996,1.89,1.27,7.14,6.7799997,2.22,0.74,3.02,3.9099998,3.46,3.58,4.0699997,5.6,5.69,4.41,4.04,4.39,11.15,18.949999,21.369999,20.369999,19.38,17.449999,15.67,14.21,9.389999,7.2,6.0699997,2.96,1.41,0.96999997,0.17999999,0.0,0.0,0.01,0.56,0.47,0.089999996,0.11,0.22999999,0.07,0.049999997,0.16,0.22999999,0.56,0.71999997,0.32,0.08,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.049999997,0.26,0.59999996,1.81,1.61,1.92,3.1999998,4.38,5.58,7.06,8.099999,8.639999,7.3199997,7.98,8.0199995,6.5,7.37,8.74,7.3199997,4.7,4.61,4.25,3.25,3.25,3.37,5.04,4.45,2.58,4.2599998,7.1499996,9.94,12.48,14.32,15.889999,18.09,22.76,23.279999,23.289999,20.4,18.08,13.719999,9.28,5.3399997,3.51,3.46,2.3799999,1.8499999,2.1499999,3.86,3.98,6.98,12.259999,17.88,20.82,22.529999,22.6,22.67,18.27,11.83,8.9,7.48,7.44,7.22,6.81,6.27,5.96,7.0,8.73,9.24,7.96,6.7,9.639999,14.2,17.92,20.67,23.199999,24.98,24.89,23.25,19.289999,17.14,7.6299996,2.78,1.09,0.53,0.42999998,0.39,0.24,0.35,0.5,0.63,0.78,0.62,0.19999999,0.0,0.04,0.16,0.089999996,0.03,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.68,5.4,4.25,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08,1.35,1.9399999,0.58,0.089999996,0.14,0.17,0.19,0.84999996,0.45,4.12,3.24,0.55,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.11,0.41,0.02,0.7,1.43,3.06,2.9099998,2.12,3.6799998,8.4,10.59,10.929999,7.7799997,1.14,0.76,1.13,0.66999996,0.89,0.77,0.71999997,0.17999999,0.0,0.0,2.21,4.0899997,0.57,0.0,0.0,1.14,0.17999999,2.4299998,2.1,0.98999995,0.77,0.78999996,0.48999998,0.0,0.0,0.42,0.32999998,0.22999999,0.0,0.01,1.64,1.09,6.7,0.91999996,1.43,2.31,3.34,4.44,1.4399999,2.4299998,2.76,2.53,2.12,5.41,10.01,11.63,10.42,14.09,15.91,20.65,21.22,11.429999,8.559999,6.6099997,5.47,2.47,1.1,1.38,1.54,0.90999997,0.81,0.74,0.71,0.35999998,0.61,0.52,0.72999996,0.68,0.59999996,0.65999997,1.62,3.01,3.3799999,2.53,1.3299999,0.61,0.22,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.04,0.089999996,0.84,3.1799998,4.35,5.71,8.4,10.71,12.07,10.48,9.099999,7.81,6.68,6.8999996,8.51,6.46,4.5699997,3.47,3.83,6.2,7.3599997,6.8399997,6.2,5.42,6.5899997,8.21,9.95,13.849999,18.49,20.689999,18.02,17.44,20.0,23.01,23.85,20.51,16.3,12.45,7.8999996,4.44,2.3799999,3.5,5.14,5.49,5.91,6.6099997,7.27,8.94,11.469999,15.0199995,19.619999,23.83,26.71,34.67,38.75,38.149998,29.099998,15.83,10.29,11.509999,11.099999,9.179999,7.98,6.69,5.58,5.04,3.3,4.81,6.52,9.3,11.41,14.44,16.77,19.08,17.55,16.5,13.95,8.429999,4.73,2.79,1.48,1.3199999,1.0699999,0.66999996,0.38,0.03,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.04,0.14,0.22999999,0.34,0.48,0.53,2.58,6.5699997,2.29,1.5899999,1.4399999,0.04,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.22999999,0.32999998,0.0,0.0,0.32999998,0.17999999,0.65,2.4199998,3.77,6.96,6.3999996,5.73,9.7699995,9.599999,5.58,4.37,2.6299999,0.96999997,1.18,0.31,0.17999999,0.22999999,0.08,0.0,0.0,0.0,0.48999998,3.12,0.87,0.01,0.06,2.9299998,0.24,1.56,0.91999996,1.18,1.66,1.4499999,0.42,0.0,0.049999997,0.76,0.83,0.29999998,0.0,0.26,1.3199999,3.1799998,2.62,0.26,1.01,0.63,2.25,2.8899999,1.0699999,4.46,4.35,3.07,3.1,6.75,6.95,7.45,10.809999,12.75,14.98,14.299999,8.98,5.99,5.6299996,3.52,2.1499999,1.28,2.01,3.11,4.41,5.66,7.5499997,7.46,8.309999,8.58,6.56,6.15,4.3399997,2.82,1.1999999,0.45,1.0,1.16,0.93,0.79999995,0.93,1.0,0.71999997,0.74,0.76,0.58,0.32999998,0.68,0.22999999,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.16,1.1999999,2.24,5.39,8.24,10.599999,13.059999,12.17,10.69,9.139999,6.89,8.21,9.03,5.73,3.7099998,1.9799999,3.25,4.75,4.0899997,4.36,4.11,5.38,6.6099997,10.16,13.69,18.52,22.859999,22.63,20.82,17.21,17.789999,20.49,22.05,19.83,14.95,8.639999,5.23,3.9099998,5.8199997,7.74,11.73,11.0199995,10.16,9.76,7.35,8.59,8.42,10.87,15.61,22.34,26.99,33.23,35.14,42.719997,41.55,35.29,32.98,25.519999,21.1,23.82,24.73,17.93,10.25,6.5299997,6.6299996,4.5699997,3.47,5.3599997,8.599999,11.08,11.32,11.57,10.0199995,8.72,8.21,7.39,6.5299997,5.5299997,4.27,2.6599998,1.39,0.41,0.049999997,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06,0.13,0.17999999,0.24,0.29999998,0.52,0.52,0.76,1.09,0.51,0.59,0.39999998,0.07,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.11,0.84,0.44,0.17999999,0.04,0.76,0.32999998,0.32999998,0.93,1.5899999,2.58,2.9099998,4.08,3.85,4.5099998,1.8,0.96999997,1.55,2.1399999,1.93,0.29999998,0.0,0.0,0.0,0.0,0.0,0.0,0.13,0.69,0.19999999,0.01,0.04,1.51,0.13,0.65,0.75,0.45999998,0.85999995,0.84,0.0,0.0,0.04,0.61,0.59999996,0.0,0.0,0.78999996,1.17,1.91,0.44,0.11,0.32,0.61,0.96,1.7199999,0.85999995,5.69,6.58,2.2,1.22,2.86,3.35,8.62,11.0199995,8.639999,9.639999,8.41,5.46,2.32,1.0799999,1.26,2.23,2.69,4.31,6.3599997,6.42,5.3599997,5.54,7.0699997,6.49,5.5899997,5.48,6.48,4.94,2.8,0.94,0.56,0.29,0.38,0.39,0.42999998,0.32,0.51,0.32,0.12,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.17,1.75,3.99,6.29,9.719999,11.48,11.09,10.66,8.67,5.8599997,5.95,4.91,6.1099997,5.27,1.9799999,1.76,4.25,4.68,4.5299997,4.41,5.38,8.97,14.83,17.949999,19.89,21.99,22.63,21.99,20.22,17.83,16.55,15.16,12.809999,9.929999,6.92,7.1299996,7.8999996,12.349999,12.98,14.32,13.41,10.04,7.25,4.13,4.89,6.6,8.0199995,14.13,21.15,24.23,26.9,33.48,41.579998,48.39,45.75,38.219997,33.059998,27.269999,30.97,35.29,24.22,20.34,21.32,11.11,4.74,3.9299998,4.13,5.29,6.8399997,6.79,6.8399997,6.0499997,7.49,9.66,11.63,12.08,11.74,8.389999,4.5099998,1.52,0.29,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.04,0.07,0.049999997,0.17999999,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.22,2.06,1.37,0.07,0.0,0.65,1.13,1.8299999,2.22,3.9599998,1.74,0.65,1.53,2.6699998,4.98,2.6599998,0.32,1.31,3.56,2.44,0.52,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.049999997,0.0,0.0,0.01,0.58,0.02,0.11,0.13,0.04,0.44,0.42,0.0,0.0,0.21,0.26999998,0.06,0.0,0.17,0.52,0.21,0.57,0.01,0.06,0.14999999,0.48,0.45999998,0.52,1.5899999,2.6699998,3.4099998,3.7099998,3.3799999,3.11,3.6499999,11.05,26.039999,17.3,8.389999,6.24,4.62,5.04,6.24,5.81,5.2,5.0499997,4.02,2.6799998,1.5699999,1.65,1.1,1.1999999,0.14999999,0.9,1.01,0.59,0.22,0.19,0.049999997,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.17,0.29,2.98,9.849999,12.94,16.22,14.099999,9.63,8.0,6.49,5.42,4.8599997,5.66,4.83,3.1599998,3.51,4.9,5.18,3.25,3.24,6.83,13.309999,15.679999,16.17,17.539999,18.91,18.93,20.06,19.3,16.5,13.809999,11.139999,8.17,7.0299997,8.41,8.29,9.3,12.59,11.92,13.69,13.32,9.559999,6.3799996,3.59,2.8999999,4.2,7.3799996,9.92,14.889999,19.289999,22.24,26.64,33.68,42.899998,50.98,47.129997,42.129997,38.52,40.14,41.059998,41.37,37.26,27.08,17.039999,9.12,5.12,3.9199998,3.1499999,2.83,2.31,2.49,3.53,6.5099998,9.71,11.66,10.67,7.3999996,4.1,1.8199999,0.26999998,0.0,0.01,0.06,0.099999994,0.16,0.17,0.13,0.19999999,0.21,0.21,0.35,0.17,0.13,0.12,0.0,0.0,0.02,0.049999997,0.03,0.08,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,1.1,1.87,0.77,0.35,0.16,0.08,1.13,2.58,6.85,4.75,0.25,1.24,5.3199997,8.08,2.48,0.31,0.61,3.25,2.19,0.42999998,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.44,0.0,0.0,0.0,0.0,0.32,0.0,0.0,0.0,0.02,0.0,0.0,0.08,0.59,0.14,0.0,0.0,0.03,0.19999999,0.04,0.11,0.38,0.69,2.1499999,2.32,2.48,2.75,6.91,4.65,5.18,11.92,15.78,9.99,9.469999,14.969999,14.009999,10.37,7.8999996,4.39,2.86,1.09,0.41,0.45999998,1.13,0.88,0.0,0.94,0.53,0.35999998,0.13,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.21,1.87,8.059999,11.36,8.0199995,7.5,6.79,7.35,6.6099997,5.87,6.27,8.53,6.71,4.61,4.79,4.7,2.08,1.9499999,3.79,7.2999997,8.95,10.08,12.96,16.17,16.699999,16.13,17.63,17.92,18.76,17.27,12.559999,9.0199995,9.01,9.21,7.77,7.02,7.91,10.0,11.65,11.71,9.429999,6.42,3.1,2.9199998,3.6899998,6.64,8.09,10.59,13.32,16.07,18.279999,21.699999,29.429998,37.059998,40.17,39.69,38.91,43.329998,51.91,50.6,48.079998,38.18,25.92,18.06,7.97,6.41,4.0099998,2.79,1.86,2.06,2.69,2.8,3.21,3.27,2.81,2.06,0.16,0.0,0.0,0.0,0.03,0.07,0.099999994,0.08,0.0,0.099999994,0.17,0.099999994,0.07,0.13,0.03,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13,1.1899999,1.99,1.04,1.13,0.14,0.45999998,0.81,2.48,2.76,0.22,1.63,3.9499998,4.0699997,1.9799999,0.61,0.14999999,2.04,0.96,0.13,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.39999998,0.0,0.0,0.0,0.0,0.16,0.0,0.0,0.0,0.0,0.0,0.0,0.14999999,0.26,0.099999994,0.11,0.0,0.08,0.19,0.0,0.0,0.14,0.47,0.47,1.64,1.9799999,3.47,6.29,6.24,10.88,19.22,20.289999,18.97,14.41,13.49,9.45,4.69,1.68,0.42999998,0.02,0.0,0.04,0.14999999,0.19999999,0.13,0.53999996,0.21,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.02,0.29,2.57,3.26,2.47,4.5099998,5.1099997,5.14,5.71,6.19,6.5899997,7.18,5.95,5.71,5.33,2.97,0.85999995,1.48,3.1799998,4.5099998,5.54,8.45,12.83,15.61,17.07,18.31,17.51,18.029999,21.539999,18.98,15.04,13.2,11.95,9.429999,7.1,5.31,6.48,6.7599998,7.6699996,9.11,8.46,6.71,4.3199997,2.9399998,3.4499998,4.46,7.48,8.0199995,9.33,10.79,12.69,13.639999,17.47,22.93,31.32,30.09,34.719997,41.7,51.52,52.71,45.02,38.54,24.93,12.46,7.71,5.23,5.17,3.73,2.74,1.9399999,1.91,1.86,1.22,0.63,0.26,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02,0.089999996,0.13,0.089999996,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.19,0.31,0.41,0.45999998,1.14,0.9,1.15,0.41,0.66999996,0.89,0.03,1.3399999,3.24,2.26,0.55,0.22999999,0.01,0.76,0.42,0.04,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13,0.38,0.0,0.0,0.0,0.0,0.14,0.0,0.0,0.0,0.0,0.0,0.28,0.28,0.0,0.04,0.29999998,0.0,0.03,0.0,0.0,0.0,0.29999998,0.51,0.17,0.7,1.11,5.58,8.26,11.21,18.64,27.8,34.13,30.449999,18.33,7.2599998,1.66,0.29999998,0.04,0.0,0.0,0.0,0.0,0.38,0.03,0.08,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.089999996,0.13,0.41,1.9699999,3.05,3.6,3.73,5.73,6.64,7.33,6.5099998,6.06,6.1099997,3.76,2.47,2.6,3.86,4.68,6.85,11.57,14.09,16.77,18.93,20.58,20.83,24.18,24.98,21.84,18.42,16.83,15.96,12.24,7.3199997,4.7599998,4.5499997,5.04,5.5899997,6.43,8.97,10.44,9.38,6.6299996,5.27,4.92,6.31,7.14,6.18,6.74,8.09,10.37,13.71,15.139999,17.49,18.27,21.449999,30.14,36.23,38.399998,35.059998,26.49,15.759999,7.47,4.0299997,2.97,2.49,2.6399999,2.79,2.71,2.27,1.49,0.89,0.29999998,0.11,0.099999994,0.12,0.07,0.29,0.48,0.52,0.29999998,0.099999994,0.0,0.03,0.04,0.07,0.04,0.0,0.0,0.0,0.0,0.01,0.049999997,0.07,0.03,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.11,0.83,0.77,0.65,0.35,0.0,0.59,4.17,5.2799997,1.05,0.26,0.07,0.0,0.59999996,1.28,0.35999998,0.08,0.089999996,0.0,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07,0.0,0.0,0.0,0.0,0.0,0.049999997,0.0,0.0,0.0,0.0,0.04,0.03,0.049999997,0.0,0.06,0.19,0.0,0.0,0.0,0.0,0.02,0.47,0.19999999,0.11,0.04,0.5,6.0299997,8.98,11.099999,14.349999,20.619999,27.0,20.22,11.01,2.44,0.22999999,0.0,0.0,0.0,0.0,0.0,0.02,0.07,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.11,0.04,0.04,0.72999996,1.09,0.9,3.47,7.97,7.4199996,6.6499996,6.0699997,6.0099998,7.6099997,6.45,4.7799997,3.7099998,5.15,7.37,9.34,10.59,12.599999,15.5199995,18.55,19.6,21.46,24.039999,24.119999,21.34,18.32,17.16,14.24,11.429999,7.0899997,3.62,3.23,3.87,4.61,4.68,6.2999997,7.79,8.26,8.79,5.64,4.7,5.0,6.97,5.0899997,4.27,4.97,7.06,8.809999,9.29,9.0199995,10.09,12.66,15.38,17.32,19.63,17.9,16.18,10.7,7.16,6.25,6.0699997,3.8899999,3.11,3.1299999,3.47,2.59,2.1599998,1.26,0.84999996,0.53,0.29,0.57,0.74,0.5,0.38,0.26999998,0.07,0.0,0.0,0.0,0.0,0.099999994,0.099999994,0.099999994,0.13,0.089999996,0.14,0.17,0.22,0.19999999,0.19999999,0.049999997,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.35999998,1.48,1.15,0.28,0.32999998,0.38,0.84999996,2.08,3.99,0.96999997,0.28,0.14999999,0.0,0.21,0.37,0.02,0.0,0.01,0.0,0.31,0.35,0.16,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13,0.14,0.0,0.0,0.0,0.0,0.0,0.04,0.0,0.0,0.0,0.0,0.07,0.099999994,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02,0.11,0.0,0.0,0.06,2.84,10.4,13.49,9.45,8.429999,14.799999,16.869999,9.99,5.08,1.04,0.31,0.14,0.12,0.16,0.06,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.049999997,0.19,0.22,0.01,0.0,0.0,0.0,0.0,0.19,0.32,0.26,1.91,6.2799997,7.16,7.23,6.92,7.85,8.9,7.71,7.62,7.44,7.75,9.11,10.69,11.57,13.009999,15.2,16.92,17.359999,19.199999,19.75,19.72,19.46,17.359999,15.29,15.559999,11.86,9.09,7.0299997,6.15,5.43,3.99,2.45,3.01,4.0099998,4.95,5.33,4.18,3.09,2.71,2.74,2.81,2.69,2.4299998,3.25,3.76,4.38,4.22,3.46,5.31,9.0,11.7699995,12.88,10.37,8.45,8.55,8.2699995,7.3799996,5.27,3.6999998,3.58,3.6,4.8599997,5.73,5.71,4.0699997,3.03,1.63,1.01,0.71999997,0.45,0.38,0.31,0.07,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.91999996,1.5799999,0.69,0.12,0.90999997,1.03,0.56,1.0,0.5,0.21,0.12,0.0,0.03,0.04,0.0,0.0,0.0,0.0,0.53999996,0.48,0.22999999,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.04,0.099999994,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.11,0.48999998,1.15,2.84,3.1699998,3.02,9.82,15.089999,12.509999,6.43,2.62,0.89,0.95,0.62,0.59999996,0.63,0.44,0.17,0.0,0.099999994,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07,0.04,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08,0.14999999,0.13,0.25,0.14,0.099999994,0.08,0.08,0.14,0.14999999,0.03,1.31,4.7,6.1099997,6.99,9.08,10.66,9.5199995,9.719999,11.2,9.44,5.58,6.45,8.48,11.349999,14.009999,13.84,16.5,16.97,17.23,16.13,15.139999,16.47,15.219999,14.25,13.61,11.809999,11.74,10.469999,9.2699995,5.83,4.5,3.9399998,3.6499999,3.6599998,4.5499997,5.46,5.25,3.47,1.17,0.52,1.01,1.39,1.26,1.77,2.04,2.3899999,2.4299998,2.25,1.79,3.24,4.68,6.44,5.38,4.1,4.49,5.37,6.17,5.25,4.22,3.58,3.31,2.95,2.57,2.85,3.23,4.0,3.9499998,3.33,2.3899999,1.49,0.55,0.0,0.04,0.17,0.24,0.22,0.08,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.04,0.17,0.26999998,0.08,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.35999998,0.42,1.24,1.1899999,0.13,0.099999994,0.41,0.13,0.049999997,0.07,0.03,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.42,0.47,0.26,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.19,1.55,2.31,3.6899998,2.82,3.28,10.3,11.9,7.3599997,2.79,1.67,1.2099999,1.51,1.87,1.3,0.78999996,0.24,0.02,0.28,0.53999996,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.0,0.28,0.25,0.12,0.03,0.01,0.28,0.32,0.02,0.0,0.0,0.0,0.0,0.02,0.19,2.33,1.38,0.45,0.53999996,0.59,0.71,0.74,0.22999999,0.38,1.3299999,3.1999998,6.77,8.07,11.05,10.91,9.809999,10.59,11.19,8.099999,7.3399997,8.139999,9.88,12.139999,14.09,13.969999,14.67,16.25,16.23,16.83,15.24,13.65,12.3,11.46,12.389999,12.04,12.46,11.54,10.29,8.61,7.6499996,6.8799996,6.29,5.22,4.93,5.0699997,5.35,4.88,2.9199998,1.29,0.72999996,0.72999996,0.96999997,1.5799999,2.11,1.9499999,1.76,1.51,1.23,1.64,1.64,1.75,1.41,0.90999997,0.71999997,0.84999996,1.43,2.0,2.45,2.3899999,2.33,2.32,2.3,2.8799999,4.36,3.9099998,3.98,3.7099998,2.85,2.12,2.3,2.1299999,1.8299999,1.43,0.7,0.5,0.16,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.04,0.07,0.03,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.26,0.53,0.76,0.78999996,0.66999996,0.77,0.68,0.5,0.39999998,0.28,0.24,0.11,0.07,0.04,0.0,0.07,1.1899999,1.39,0.90999997,0.56,0.03,0.01,0.049999997,0.0,0.0,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.26999998,0.22999999,0.04,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.55,1.03,1.91,1.48,2.78,7.6099997,11.429999,13.21,9.17,2.24,1.0699999,1.75,2.01,3.06,3.1499999,3.54,4.02,0.88,0.66999996,0.79999995,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02,0.29,1.4499999,1.27,1.31,0.65,0.28,0.0,0.01,0.53,0.58,0.0,0.0,0.01,0.03,0.03,0.02,0.19999999,0.42,0.13,0.37,0.63,0.96,1.5,2.09,1.93,0.93,1.5999999,1.61,1.6899999,3.98,4.61,4.19,6.08,6.8999996,7.96,8.95,8.099999,6.99,7.73,9.29,10.139999,11.13,13.179999,13.849999,14.19,14.73,15.19,14.589999,12.59,11.389999,11.0,12.2699995,13.5,14.07,13.259999,11.44,9.5,8.36,8.45,6.5299997,5.45,3.98,3.23,3.28,4.0499997,3.31,1.53,0.69,0.32,0.68,1.3399999,1.66,1.4699999,0.88,0.47,0.22,0.07,0.0,0.089999996,0.26,0.29999998,0.14999999,0.01,0.01,0.17999999,0.22999999,0.65,1.4399999,2.1399999,3.33,3.51,1.91,0.41,0.22999999,0.28,0.29999998,1.3,0.79999995,0.37,0.24,0.089999996,0.04,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02,0.19,0.39,0.42,0.57,0.66999996,0.22,0.11,0.0,0.13,0.04,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.089999996,0.17,0.0,0.0,0.0,0.0,0.38,0.45,0.22999999,0.17999999,0.35999998,0.26999998,0.28,0.84,1.39,1.64,2.0,2.25,2.45,2.04,2.1299999,2.4199998,2.1499999,1.5699999,1.26,0.89,0.59999996,0.47,0.26,0.14,0.17,1.05,2.18,1.09,0.62,0.099999994,0.0,0.0,0.0,0.0,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.44,0.51,0.71999997,1.26,1.52,3.9099998,5.7999997,7.3799996,7.68,3.03,1.14,1.51,2.51,3.75,3.77,2.9299998,2.9299998,1.8399999,0.35999998,1.25,0.65999997,0.12,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.12,0.42,2.62,3.9199998,3.3799999,1.42,0.61,0.08,0.32,1.05,0.17999999,0.0,0.0,0.17,0.45999998,0.42999998,0.37,0.32999998,0.72999996,0.82,0.82,0.65,0.78,1.53,2.05,2.51,1.9799999,1.5899999,2.2,1.76,0.93,2.53,3.6599998,4.81,5.98,6.6499996,7.3799996,7.8399997,7.5,7.27,7.93,9.309999,9.809999,11.53,14.349999,13.0,11.61,11.23,12.11,11.71,11.01,9.33,9.28,10.5,12.92,13.53,13.679999,12.62,12.429999,10.7,10.08,8.87,7.8799996,6.3999996,5.7,4.85,4.14,2.6499999,1.18,0.32999998,0.61,0.90999997,1.11,1.04,0.81,0.69,0.68,0.62,0.19999999,0.0,0.01,0.04,0.28,0.34,0.22999999,0.04,0.03,0.12,0.26999998,0.35999998,0.53999996,0.85999995,0.39999998,0.26,0.12,0.04,0.01,0.08,0.049999997,0.0,0.01,0.03,0.0,0.0,0.0,0.049999997,0.12,0.08,0.04,0.07,0.08,0.03,0.06,0.13,0.089999996,0.049999997,0.17,0.19999999,0.099999994,0.22999999,0.31,0.44,0.52,0.74,0.72999996,0.45999998,0.32999998,0.42999998,0.04,0.02,0.01,0.0,0.0,0.0,0.14999999,0.38,0.47,0.25,0.12,0.14999999,0.55,0.85999995,1.23,0.89,0.61,0.7,1.61,2.0,2.02,1.8399999,2.48,2.47,2.4099998,2.6599998,2.78,3.6299999,3.4199998,3.1799998,2.7,2.3799999,2.1299999,2.1299999,2.36,1.7099999,1.4499999,0.96999997,0.59999996,0.32,0.11,0.08,0.0,0.47,1.39,0.24,0.089999996,0.0,0.0,0.0,0.0,0.0,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.099999994,0.13,0.42,0.65,2.07,5.98,11.849999,10.17,4.23,0.11,0.93,3.24,3.78,3.3799999,3.56,4.2999997,3.81,0.83,0.85999995,0.95,0.14999999,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.31,0.65,2.25,3.8999999,5.83,4.87,3.21,0.83,2.78,2.56,0.26999998,0.0,0.0,0.74,1.17,0.97999996,0.83,1.1899999,1.28,2.01,2.58,2.33,2.26,2.6499999,2.6699998,2.52,2.4099998,2.22,1.78,1.9399999,0.94,0.39,1.76,4.72,6.89,8.34,8.139999,8.62,7.95,7.21,6.7599998,8.309999,8.45,9.21,10.61,11.07,12.44,11.7699995,10.26,10.719999,11.09,11.05,10.3,9.98,10.32,12.2699995,13.96,15.809999,16.89,16.05,13.87,13.21,13.11,12.2699995,11.07,10.78,7.71,5.39,2.6799998,2.23,0.56,0.32,0.19999999,0.41,0.59,0.66999996,1.1899999,1.3399999,1.41,0.90999997,0.14,0.07,0.0,0.08,0.21,0.22,0.11,0.089999996,0.21,0.26,0.16,0.0,0.0,0.0,0.0,0.29999998,0.21,0.089999996,0.08,0.0,0.0,0.0,0.0,0.0,0.0,0.32999998,0.52,0.45,0.32999998,0.34,0.58,0.59,0.22,0.03,0.02,0.39999998,0.88,0.71999997,0.90999997,1.02,1.09,1.18,1.01,0.89,0.72999996,0.35999998,0.68,0.53999996,0.48,0.51,0.29999998,0.17,0.28,0.84999996,1.31,1.67,1.1899999,1.3199999,1.73,1.6899999,1.8299999,2.75,4.22,4.21,2.99,1.73,2.72,3.6399999,2.8899999,2.3999999,2.96,3.6399999,3.6599998,3.98,3.6699998,3.58,3.46,3.11,2.09,1.31,0.97999996,0.61,1.3199999,2.28,1.62,0.5,0.48,0.48,0.41,0.37,0.0,0.29999998,0.88,0.03,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.099999994,0.22999999,0.13,1.09,0.39,1.3299999,4.06,6.5099998,5.1099997,1.73,0.29,1.9599999,3.37,3.5,2.34,2.51,4.27,2.81,0.85999995,1.3399999,0.71999997,0.07,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.29999998,0.57,1.56,4.35,5.93,5.39,5.25,4.04,4.49,1.8299999,0.07,0.0,0.0,1.25,1.79,1.64,0.7,2.09,1.25,0.88,2.78,4.13,3.47,4.06,3.72,3.25,3.6899998,2.6,1.56,1.05,1.05,1.2099999,1.13,3.1399999,6.92,8.3,8.33,8.599999,6.79,6.04,5.98,6.19,6.31,6.8199997,7.31,9.4,8.41,10.94,11.469999,12.25,11.95,12.19,13.41,13.21,12.639999,14.929999,15.95,15.799999,18.039999,19.52,18.07,17.06,15.96,14.67,14.139999,15.61,14.349999,12.639999,9.38,5.33,4.18,2.11,0.89,1.05,0.89,0.65,0.84999996,0.84,0.93,1.53,1.89,1.0699999,0.53999996,0.22999999,0.049999997,0.099999994,0.07,0.0,0.0,0.099999994,0.089999996,0.03,0.0,0.0,0.02,0.28,0.62,0.51,0.41,0.48,0.32999998,0.19999999,0.07,0.29999998,0.53,0.56,0.19999999,0.19,0.21,0.45,1.12,0.98999995,0.53999996,0.95,1.25,1.37,1.43,1.49,1.39,1.93,2.44,2.28,1.9599999,1.64,1.77,2.28,3.85,5.71,4.5699997,3.09,2.0,1.87,2.07,1.64,1.8199999,2.1599998,2.53,4.0499997,4.96,4.41,4.0099998,5.8199997,8.0199995,6.5,4.89,3.23,3.1699998,4.08,4.21,3.3999999,2.37,2.3799999,2.46,2.34,2.75,1.9799999,1.5899999,1.02,0.7,0.53999996,0.84999996,1.22,1.56,2.3999999,2.5,2.09,1.86,1.7099999,1.3,1.0,0.37,0.24,0.69,0.11,0.19,0.04,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.53,1.2099999,0.22,1.3299999,0.91999996,1.4499999,2.51,1.1899999,0.39999998,0.099999994,1.22,1.8499999,1.39,1.64,1.3199999,1.39,0.41,0.35999998,0.97999996,0.93,0.14999999,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03,0.41,0.21,0.63,0.88,1.8199999,3.84,4.08,6.0099998,8.059999,6.8199997,4.48,0.38,0.08,1.92,3.49,3.9299998,4.8599997,3.9199998,1.5699999,4.21,4.0899997,3.05,3.6599998,4.15,5.72,4.2599998,3.83,3.32,2.96,2.27,1.3299999,1.05,1.4499999,1.86,2.71,3.36,4.27,8.82,10.3,9.22,7.71,5.69,4.87,4.63,4.7999997,4.61,4.3399997,5.93,8.11,8.5,9.57,10.34,12.54,13.92,14.929999,15.07,17.77,20.31,21.67,20.85,20.39,22.16,21.89,20.42,19.18,17.84,17.72,18.71,21.3,20.93,19.779999,18.91,14.25,8.7699995,4.19,2.6399999,3.23,2.74,2.54,2.01,1.2099999,1.3299999,2.19,3.56,3.9299998,2.72,1.4,1.04,0.68,0.26,0.03,0.049999997,0.0,0.0,0.02,0.03,0.28,0.51,0.71999997,0.78999996,0.90999997,0.90999997,0.9,0.45999998,0.88,1.3,1.41,0.53999996,0.26999998,0.55,0.59999996,0.44,0.59999996,0.64,0.51,0.47,0.48999998,0.48,0.39,0.42999998,0.5,0.84,0.9,1.1899999,1.65,2.82,4.17,6.83,9.71,9.5199995,6.43,3.9599998,4.52,5.08,6.0699997,7.12,7.49,7.2,6.3599997,6.1299996,6.3999996,6.0499997,5.54,5.13,6.0299997,5.47,4.88,4.71,4.2999997,4.5099998,4.2,3.1999998,2.04,1.41,0.72999996,0.65999997,0.64,0.75,1.05,1.5999999,2.33,2.7,2.6699998,2.54,2.29,2.06,1.7199999,1.41,0.96999997,0.78999996,0.5,0.26999998,0.24,0.14,0.35999998,0.08,0.21,0.07,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.17,0.42,0.44,1.7199999,1.7099999,3.6399999,3.6699998,1.3199999,0.26999998,1.38,1.5,1.5,1.4699999,0.22,0.24,0.12,0.0,0.13,0.58,0.28,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06,0.47,0.099999994,0.26999998,0.96,2.11,2.51,5.6299996,5.8199997,6.93,6.7999997,5.92,4.95,3.02,13.08,11.08,6.37,11.2699995,10.639999,8.2699995,4.43,4.79,4.2799997,6.74,3.77,2.74,2.74,4.1,3.84,3.55,2.74,2.4099998,1.01,0.96,2.4099998,1.55,1.4599999,3.6899998,5.04,3.82,3.47,6.73,7.3799996,6.99,6.04,4.2,3.06,2.51,2.51,2.8799999,2.19,2.1299999,4.85,8.639999,10.88,10.4,11.19,11.15,13.799999,13.19,14.88,18.21,23.41,24.65,25.39,23.71,20.31,18.939999,18.02,17.02,18.55,22.16,26.359999,26.359999,24.8,20.58,17.22,11.719999,8.5,4.0499997,3.21,3.55,4.1,4.58,3.1399999,2.74,2.98,3.9099998,4.39,3.3,1.73,1.4,1.39,0.88,0.29,0.02,0.0,0.0,0.0,0.03,0.22,0.39,0.66999996,1.01,1.26,1.7199999,1.8299999,2.03,2.32,2.32,2.4099998,2.31,2.3899999,1.53,1.37,1.5699999,2.32,2.26,2.1399999,1.8299999,1.88,2.56,3.9099998,5.8399997,7.16,7.0699997,7.6699996,7.47,7.5699997,9.0199995,10.09,8.17,5.4,3.23,3.9399998,3.9499998,3.75,4.15,5.08,6.2799997,7.04,5.46,4.3399997,3.4299998,2.53,2.71,3.33,3.1899998,3.23,3.58,3.97,3.35,1.77,2.24,2.4099998,2.18,2.19,2.1,2.6299999,3.1799998,3.4499998,3.73,3.4299998,2.82,1.86,1.13,0.62,0.42999998,0.29,0.13,0.03,0.0,0.0,0.0,0.0,0.08,0.08,0.14999999,0.01,0.049999997,0.02,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.7,1.6899999,1.88,2.23,1.13,0.59,0.59,1.38,1.51,1.38,0.35999998,0.0,0.0,0.0,0.0,0.13,0.22,0.049999997,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06,0.31,0.0,0.0,1.41,2.2,3.99,7.9199996,6.5299997,9.32,9.929999,7.19,4.04,1.37,3.3799999,3.98,0.96999997,0.68,0.32999998,1.4,2.9199998,9.74,15.089999,16.67,8.63,2.6499999,2.2,2.6499999,2.11,2.02,1.6999999,1.1899999,0.74,0.19,0.82,1.36,1.4399999,1.76,2.8,2.97,2.07,1.62,2.12,3.23,2.81,2.19,1.86,1.48,1.0699999,0.87,1.17,0.91999996,0.45999998,1.13,4.44,7.8599997,8.73,7.89,5.6299996,6.6499996,7.0299997,8.46,8.5199995,12.99,17.949999,20.0,17.1,15.98,16.92,14.9,13.91,18.119999,20.859999,24.01,28.46,24.539999,18.42,14.12,9.83,7.72,5.95,5.1099997,3.8799999,3.4299998,2.6299999,2.23,2.22,2.35,2.87,2.36,1.4,0.93,0.51,0.47,0.26,0.26999998,0.26,0.0,0.13,0.29999998,0.22,0.08,0.13,0.37,0.44,0.48,0.59999996,0.62,1.15,2.1699998,3.9199998,3.62,3.81,2.74,1.66,1.24,2.9099998,2.33,2.18,2.22,2.26,2.35,2.78,3.1,3.59,3.4199998,4.1,4.2999997,5.8599997,7.9199996,7.3199997,5.43,3.74,3.61,3.29,2.44,1.35,0.81,0.7,0.71,0.72999996,0.64,0.74,0.82,1.18,1.5699999,1.4699999,1.4,1.3,1.14,0.64,0.39999998,0.35,0.45999998,0.65999997,0.78,0.87,0.88,0.84999996,0.84999996,0.79999995,0.77,0.32,0.35,0.17,0.13,0.01,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0;
 } 
