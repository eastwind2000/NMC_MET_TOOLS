netcdf ecmwf_r24_2018062500_f096 {
dimensions: 
 lat = 601; 
 lon = 701; 
variables:  
float lat(lat) ; 
   lat:long_name = "latitude" ;
   lat:units = "degrees_north" ;
   lat:standard_name = "latitude" ;
float lon(lon) ;
   lon:long_name = "longitude" ;
   lon:units = "degrees_east" ;
   lon:standard_name = "longitude" ;
float APCP_24(lat, lon) ;
   APCP_24:name = "APCP_24" ;
   APCP_24:long_name = "Total Precipitation" ;
   APCP_24:level = "A24" ;
   APCP_24:units = "kg/m^2" ;
   APCP_24:_FillValue = -9999.f ;
   APCP_24:init_time = "20180625_000000" ;
   APCP_24:init_time_ut = "1529884800.0" ;
   APCP_24:valid_time = "20180629_000000" ;
   APCP_24:valid_time_ut = "1530230400.0" ;
   APCP_24:accum_time = "240000" ;
   APCP_24:_FillValue = 65535 ;
   APCP_24:accum_time_sec = 86400 ;
 // global attributes: 
 :_NCProperties = "version=1|netcdflibversion=4.4.1.1" ;
	:FileOrigins = "ECMWF_HR_APCP24" ; 
	:MET_version = "V7.0" ;
	:Projection = "LatLon" ;
	:lat_ll = "0.0 degrees_north" ; 
	:lon_ll = "70.0 degrees_east" ; 
	:delta_lat = "0.10 degrees" ;
	:delta_lon = "0.10 degrees" ;
	:Nlat = "601 grid_points" ; 
	:Nlon = "701 grid_points" ; 
data:
lat = 0.0,0.1,0.2,0.3,0.4,0.5,0.6,0.7,0.8,0.90000004,1.0,1.1,1.2,1.3000001,1.4,1.5,1.6,1.7,1.8000001,1.9,2.0,2.1000001,2.2,2.3,2.4,2.5,2.6000001,2.7,2.8,2.9,3.0,3.1000001,3.2,3.3,3.4,3.5,3.6000001,3.7,3.8,3.9,4.0,4.1,4.2000003,4.3,4.4,4.5,4.6,4.7000003,4.8,4.9,5.0,5.1,5.2000003,5.3,5.4,5.5,5.6,5.7000003,5.8,5.9,6.0,6.1,6.2000003,6.3,6.4,6.5,6.6,6.7000003,6.8,6.9,7.0,7.1,7.2000003,7.3,7.4,7.5,7.6,7.7000003,7.8,7.9,8.0,8.1,8.2,8.3,8.400001,8.5,8.6,8.7,8.8,8.900001,9.0,9.1,9.2,9.3,9.400001,9.5,9.6,9.7,9.8,9.900001,10.0,10.1,10.2,10.3,10.400001,10.5,10.6,10.7,10.8,10.900001,11.0,11.1,11.2,11.3,11.400001,11.5,11.6,11.7,11.8,11.900001,12.0,12.1,12.2,12.3,12.400001,12.5,12.6,12.7,12.8,12.900001,13.0,13.1,13.2,13.3,13.400001,13.5,13.6,13.7,13.8,13.900001,14.0,14.1,14.2,14.3,14.400001,14.5,14.6,14.7,14.8,14.900001,15.0,15.1,15.2,15.3,15.400001,15.5,15.6,15.7,15.8,15.900001,16.0,16.1,16.2,16.300001,16.4,16.5,16.6,16.7,16.800001,16.9,17.0,17.1,17.2,17.300001,17.4,17.5,17.6,17.7,17.800001,17.9,18.0,18.1,18.2,18.300001,18.4,18.5,18.6,18.7,18.800001,18.9,19.0,19.1,19.2,19.300001,19.4,19.5,19.6,19.7,19.800001,19.9,20.0,20.1,20.2,20.300001,20.4,20.5,20.6,20.7,20.800001,20.9,21.0,21.1,21.2,21.300001,21.4,21.5,21.6,21.7,21.800001,21.9,22.0,22.1,22.2,22.300001,22.4,22.5,22.6,22.7,22.800001,22.9,23.0,23.1,23.2,23.300001,23.4,23.5,23.6,23.7,23.800001,23.9,24.0,24.1,24.2,24.300001,24.4,24.5,24.6,24.7,24.800001,24.9,25.0,25.1,25.2,25.300001,25.4,25.5,25.6,25.7,25.800001,25.9,26.0,26.1,26.2,26.300001,26.4,26.5,26.6,26.7,26.800001,26.9,27.0,27.1,27.2,27.300001,27.4,27.5,27.6,27.7,27.800001,27.9,28.0,28.1,28.2,28.300001,28.4,28.5,28.6,28.7,28.800001,28.9,29.0,29.1,29.2,29.300001,29.4,29.5,29.6,29.7,29.800001,29.9,30.0,30.1,30.2,30.300001,30.4,30.5,30.6,30.7,30.800001,30.9,31.0,31.1,31.2,31.300001,31.4,31.5,31.6,31.7,31.800001,31.9,32.0,32.100002,32.2,32.3,32.4,32.5,32.600002,32.7,32.8,32.9,33.0,33.100002,33.2,33.3,33.4,33.5,33.600002,33.7,33.8,33.9,34.0,34.100002,34.2,34.3,34.4,34.5,34.600002,34.7,34.8,34.9,35.0,35.100002,35.2,35.3,35.4,35.5,35.600002,35.7,35.8,35.9,36.0,36.100002,36.2,36.3,36.4,36.5,36.600002,36.7,36.8,36.9,37.0,37.100002,37.2,37.3,37.4,37.5,37.600002,37.7,37.8,37.9,38.0,38.100002,38.2,38.3,38.4,38.5,38.600002,38.7,38.8,38.9,39.0,39.100002,39.2,39.3,39.4,39.5,39.600002,39.7,39.8,39.9,40.0,40.100002,40.2,40.3,40.4,40.5,40.600002,40.7,40.8,40.9,41.0,41.100002,41.2,41.3,41.4,41.5,41.600002,41.7,41.8,41.9,42.0,42.100002,42.2,42.3,42.4,42.5,42.600002,42.7,42.8,42.9,43.0,43.100002,43.2,43.3,43.4,43.5,43.600002,43.7,43.8,43.9,44.0,44.100002,44.2,44.3,44.4,44.5,44.600002,44.7,44.8,44.9,45.0,45.100002,45.2,45.3,45.4,45.5,45.600002,45.7,45.8,45.9,46.0,46.100002,46.2,46.3,46.4,46.5,46.600002,46.7,46.8,46.9,47.0,47.100002,47.2,47.3,47.4,47.5,47.600002,47.7,47.8,47.9,48.0,48.100002,48.2,48.3,48.4,48.5,48.600002,48.7,48.8,48.9,49.0,49.100002,49.2,49.3,49.4,49.5,49.600002,49.7,49.8,49.9,50.0,50.100002,50.2,50.3,50.4,50.5,50.600002,50.7,50.8,50.9,51.0,51.100002,51.2,51.3,51.4,51.5,51.600002,51.7,51.8,51.9,52.0,52.100002,52.2,52.3,52.4,52.5,52.600002,52.7,52.8,52.9,53.0,53.100002,53.2,53.3,53.4,53.5,53.600002,53.7,53.8,53.9,54.0,54.100002,54.2,54.3,54.4,54.5,54.600002,54.7,54.8,54.9,55.0,55.100002,55.2,55.3,55.4,55.5,55.600002,55.7,55.8,55.9,56.0,56.100002,56.2,56.3,56.4,56.5,56.600002,56.7,56.8,56.9,57.0,57.100002,57.2,57.3,57.4,57.5,57.600002,57.7,57.8,57.9,58.0,58.100002,58.2,58.3,58.4,58.5,58.600002,58.7,58.8,58.9,59.0,59.100002,59.2,59.3,59.4,59.5,59.600002,59.7,59.8,59.9,60.0;
lon = 70.0,70.1,70.2,70.3,70.4,70.5,70.6,70.7,70.8,70.9,71.0,71.1,71.2,71.3,71.4,71.5,71.6,71.7,71.8,71.9,72.0,72.1,72.2,72.3,72.4,72.5,72.6,72.7,72.8,72.9,73.0,73.1,73.2,73.3,73.4,73.5,73.6,73.7,73.8,73.9,74.0,74.1,74.2,74.3,74.4,74.5,74.6,74.7,74.8,74.9,75.0,75.1,75.2,75.3,75.4,75.5,75.6,75.7,75.8,75.9,76.0,76.1,76.2,76.3,76.4,76.5,76.6,76.7,76.8,76.9,77.0,77.1,77.2,77.3,77.4,77.5,77.6,77.7,77.8,77.9,78.0,78.1,78.2,78.3,78.4,78.5,78.6,78.7,78.8,78.9,79.0,79.1,79.2,79.3,79.4,79.5,79.6,79.7,79.8,79.9,80.0,80.1,80.2,80.3,80.4,80.5,80.6,80.7,80.8,80.9,81.0,81.1,81.2,81.3,81.4,81.5,81.6,81.7,81.8,81.9,82.0,82.1,82.2,82.3,82.4,82.5,82.6,82.7,82.8,82.9,83.0,83.1,83.2,83.3,83.4,83.5,83.6,83.7,83.8,83.9,84.0,84.1,84.2,84.3,84.4,84.5,84.6,84.7,84.8,84.9,85.0,85.1,85.2,85.3,85.4,85.5,85.6,85.7,85.8,85.9,86.0,86.1,86.2,86.3,86.4,86.5,86.6,86.7,86.8,86.9,87.0,87.1,87.2,87.3,87.4,87.5,87.6,87.7,87.8,87.9,88.0,88.1,88.2,88.3,88.4,88.5,88.6,88.7,88.8,88.9,89.0,89.1,89.2,89.3,89.4,89.5,89.6,89.7,89.8,89.9,90.0,90.1,90.2,90.3,90.4,90.5,90.6,90.7,90.8,90.9,91.0,91.1,91.2,91.3,91.4,91.5,91.6,91.7,91.8,91.9,92.0,92.1,92.2,92.3,92.4,92.5,92.6,92.7,92.8,92.9,93.0,93.1,93.2,93.3,93.4,93.5,93.6,93.7,93.8,93.9,94.0,94.1,94.2,94.3,94.4,94.5,94.6,94.7,94.8,94.9,95.0,95.1,95.2,95.3,95.4,95.5,95.6,95.7,95.8,95.9,96.0,96.1,96.2,96.3,96.4,96.5,96.6,96.7,96.8,96.9,97.0,97.1,97.2,97.3,97.4,97.5,97.6,97.7,97.8,97.9,98.0,98.1,98.2,98.3,98.4,98.5,98.6,98.7,98.8,98.9,99.0,99.1,99.2,99.3,99.4,99.5,99.6,99.7,99.8,99.9,100.0,100.1,100.2,100.3,100.4,100.5,100.6,100.7,100.8,100.9,101.0,101.1,101.2,101.3,101.4,101.5,101.6,101.7,101.8,101.9,102.0,102.100006,102.2,102.3,102.4,102.5,102.600006,102.7,102.8,102.9,103.0,103.100006,103.2,103.3,103.4,103.5,103.600006,103.7,103.8,103.9,104.0,104.100006,104.2,104.3,104.4,104.5,104.600006,104.7,104.8,104.9,105.0,105.100006,105.2,105.3,105.4,105.5,105.600006,105.7,105.8,105.9,106.0,106.100006,106.2,106.3,106.4,106.5,106.600006,106.7,106.8,106.9,107.0,107.100006,107.2,107.3,107.4,107.5,107.600006,107.7,107.8,107.9,108.0,108.100006,108.2,108.3,108.4,108.5,108.600006,108.7,108.8,108.9,109.0,109.100006,109.2,109.3,109.4,109.5,109.600006,109.7,109.8,109.9,110.0,110.100006,110.2,110.3,110.4,110.5,110.600006,110.7,110.8,110.9,111.0,111.100006,111.2,111.3,111.4,111.5,111.600006,111.7,111.8,111.9,112.0,112.100006,112.2,112.3,112.4,112.5,112.600006,112.7,112.8,112.9,113.0,113.100006,113.2,113.3,113.4,113.5,113.600006,113.7,113.8,113.9,114.0,114.100006,114.2,114.3,114.4,114.5,114.600006,114.7,114.8,114.9,115.0,115.100006,115.2,115.3,115.4,115.5,115.600006,115.7,115.8,115.9,116.0,116.100006,116.2,116.3,116.4,116.5,116.600006,116.7,116.8,116.9,117.0,117.100006,117.2,117.3,117.4,117.5,117.600006,117.7,117.8,117.9,118.0,118.100006,118.2,118.3,118.4,118.5,118.600006,118.7,118.8,118.9,119.0,119.100006,119.2,119.3,119.4,119.5,119.600006,119.7,119.8,119.9,120.0,120.100006,120.2,120.3,120.4,120.5,120.600006,120.7,120.8,120.9,121.0,121.100006,121.2,121.3,121.4,121.5,121.600006,121.7,121.8,121.9,122.0,122.100006,122.2,122.3,122.4,122.5,122.600006,122.7,122.8,122.9,123.0,123.100006,123.2,123.3,123.4,123.5,123.600006,123.7,123.8,123.9,124.0,124.100006,124.2,124.3,124.4,124.5,124.600006,124.7,124.8,124.9,125.0,125.100006,125.2,125.3,125.4,125.5,125.600006,125.7,125.8,125.9,126.0,126.100006,126.2,126.3,126.4,126.5,126.600006,126.7,126.8,126.9,127.0,127.100006,127.2,127.3,127.4,127.5,127.600006,127.7,127.8,127.9,128.0,128.1,128.2,128.3,128.4,128.5,128.6,128.7,128.8,128.9,129.0,129.1,129.2,129.3,129.4,129.5,129.6,129.7,129.8,129.9,130.0,130.1,130.2,130.3,130.4,130.5,130.6,130.7,130.8,130.9,131.0,131.1,131.2,131.3,131.4,131.5,131.6,131.7,131.8,131.9,132.0,132.1,132.2,132.3,132.4,132.5,132.6,132.7,132.8,132.9,133.0,133.1,133.2,133.3,133.4,133.5,133.6,133.7,133.8,133.9,134.0,134.1,134.20001,134.3,134.4,134.5,134.6,134.70001,134.8,134.9,135.0,135.1,135.20001,135.3,135.4,135.5,135.6,135.70001,135.8,135.9,136.0,136.1,136.20001,136.3,136.4,136.5,136.6,136.70001,136.8,136.9,137.0,137.1,137.20001,137.3,137.4,137.5,137.6,137.70001,137.8,137.9,138.0,138.1,138.20001,138.3,138.4,138.5,138.6,138.70001,138.8,138.9,139.0,139.1,139.20001,139.3,139.4,139.5,139.6,139.70001,139.8,139.9,140.0;
APCP_24 = 0.65641034,0.67938465,0.64000005,0.6235898,0.67282057,0.79425645,0.8041026,0.7089231,0.56123084,0.48246157,0.64000005,0.6892308,0.574359,0.46933338,0.46276927,0.5481026,0.53825647,0.42338464,0.3511795,0.36102566,0.39712822,0.5907693,0.61374366,0.571077,0.50543594,0.39712822,0.4201026,0.49230772,0.571077,0.6826667,0.9156924,1.086359,1.1191796,1.3587693,1.6410258,1.3128207,1.8740515,2.1530259,2.3466668,2.484513,2.412308,3.4855387,4.092718,3.8596926,3.2853336,3.7218463,4.394667,4.4898467,4.06318,3.4724104,3.387077,3.889231,3.7382567,3.639795,3.9647183,4.7458467,4.562052,4.699898,5.2381544,5.61559,4.637539,4.4077954,4.568616,5.031385,5.61559,6.042257,5.979898,6.0849237,6.439385,6.9054365,7.125334,7.8473854,7.962257,7.4141545,6.5903597,6.3474874,6.7150774,6.8233852,7.2336416,7.8539495,7.965539,8.2215395,8.165744,7.9163084,7.778462,8.254359,7.8769236,7.817847,7.640616,7.325539,7.2631803,8.080411,8.897642,9.229129,8.832001,7.719385,6.695385,5.789539,5.543385,5.87159,6.042257,5.979898,5.3431797,4.5456414,3.7842054,3.0523078,3.0030773,3.1638978,3.2984617,3.1409233,2.3958976,2.1398976,2.0217438,2.100513,2.2646155,2.228513,2.3729234,2.802872,3.249231,3.5741541,3.767795,4.013949,4.322462,4.7425647,5.297231,5.979898,7.056411,7.762052,8.086975,7.939283,7.171283,6.9776416,6.9382567,7.3649235,8.339693,9.7214365,9.511385,9.662359,9.997129,10.400822,10.804514,11.388719,10.939077,10.029949,9.353847,9.718155,9.196308,8.523488,7.6209235,6.672411,6.1341543,7.39118,8.12636,7.6077952,6.413129,6.422975,6.803693,6.3212314,5.910975,5.681231,4.9132314,4.585026,4.4734364,4.3027697,3.8564105,2.989949,3.761231,4.023795,3.879385,3.498667,3.1442053,2.484513,2.228513,2.1530259,2.1103592,1.9987694,2.097231,2.156308,2.2744617,2.4057438,2.3794873,1.9396925,1.6672822,1.2635899,1.014154,1.7690258,1.782154,1.6114873,1.7591796,2.1103592,1.9364104,1.9495386,2.2088206,2.1234872,1.6410258,1.2504616,2.2153847,2.5665643,2.7241027,2.8192823,2.6847181,3.6004105,3.7940516,3.761231,3.754667,3.754667,3.876103,3.6496413,3.698872,4.0533338,4.1517954,3.892513,3.7382567,3.7940516,3.889231,3.570872,3.9614363,3.9220517,3.761231,3.7218463,3.9680004,3.501949,3.1573336,3.121231,3.4166157,3.9056413,3.7120004,3.6890259,3.8498464,4.3027697,5.280821,5.1954875,4.1485133,3.367385,3.2853336,3.5544617,3.3476925,3.058872,3.1737437,3.6627696,3.9680004,4.0533338,3.9286156,3.56759,3.062154,2.609231,2.92759,2.6847181,2.5271797,2.6387694,2.7602053,2.5796926,2.231795,2.5435898,3.2164104,2.8389745,2.6190772,2.2711797,2.2350771,2.3991797,2.1070771,1.7263591,1.4966155,1.4276924,1.3915899,1.0994873,1.024,0.9517949,0.90256417,0.88615394,0.88615394,2.2153847,3.0523078,3.2820516,3.0851285,2.9144619,2.7798977,2.097231,1.5097437,1.3522053,1.6311796,1.3883078,1.0896411,0.7975385,0.5940513,0.5940513,0.6301539,0.5415385,0.6071795,0.83035904,0.9156924,1.4900514,1.4211283,0.97805136,0.8336411,2.0906668,2.3696413,3.8432825,4.8016415,4.7392826,4.348718,4.923077,4.588308,3.9056413,3.3542566,3.3411283,5.0642056,4.020513,2.097231,0.6235898,0.36758977,0.4266667,0.27897438,0.20348719,0.29538465,0.44307697,0.8467693,1.2570257,1.3981539,1.1224617,0.4266667,0.4266667,0.318359,0.23958977,0.21333335,0.15097436,0.190359,0.41025645,0.69579494,1.0436924,1.5556924,2.0676925,3.0129232,4.4110775,5.8978467,6.7282057,9.452309,13.272616,14.431181,12.763899,11.687386,11.98277,12.786873,12.097642,9.042052,3.892513,6.038975,7.3353853,8.329846,9.393231,10.712616,10.663385,11.090053,11.523283,11.579078,10.955488,12.921437,14.647796,15.0088215,13.952001,12.511181,12.681848,11.234463,9.708308,8.897642,8.835282,8.602257,7.8408213,7.351795,7.529026,8.346257,7.6635904,6.3934364,6.419693,7.8014364,8.789334,10.584617,10.436924,9.143796,7.3714876,5.661539,8.602257,11.122872,11.936821,11.687386,12.970668,7.000616,4.023795,2.7437952,2.0709746,1.1454359,0.5218462,1.6311796,2.6190772,3.2886157,5.097026,3.7415388,5.353026,5.671385,4.056616,3.495385,3.5183592,4.4045134,7.204103,10.912822,12.452104,5.907693,3.7218463,2.7634873,2.8914874,6.941539,3.9023592,4.1517954,6.0980515,8.254359,9.232411,6.2884107,5.6352825,5.398975,4.3585644,1.9528207,5.8486156,4.3290257,6.0324106,10.299078,7.1876926,3.9154875,5.917539,9.206155,10.722463,8.329846,11.431385,9.7903595,7.5487185,6.498462,6.058667,3.5183592,6.0783596,6.2129235,3.2820516,3.5249233,4.20759,4.900103,9.301334,16.466053,20.81149,14.158771,12.068104,10.450052,9.796924,15.16636,9.636104,10.341744,11.250873,10.049642,8.132924,7.6701546,9.291488,10.555078,10.518975,9.750975,7.7981544,8.372514,8.579283,7.318975,5.280821,6.51159,8.149334,8.838565,8.861539,10.131693,7.506052,6.4032826,6.482052,6.741334,5.5072823,7.450257,7.8080006,8.720411,10.059488,9.399796,9.826463,9.941334,9.235693,8.369231,9.186462,9.747693,9.501539,9.91836,10.952206,11.063796,11.795693,11.88759,10.788103,9.462154,10.390975,10.489437,7.88677,6.298257,8.001641,13.824001,11.113027,9.019077,8.346257,8.3364105,6.6527185,6.8594875,6.436103,6.8397956,8.044309,8.546462,9.265231,10.039796,10.981745,11.831796,11.979488,13.919181,13.039591,11.313231,10.397539,11.641437,13.423591,14.49354,14.628103,14.87754,17.562258,15.744001,15.58318,16.026258,15.908104,13.932309,16.006565,18.146463,19.495386,19.551182,18.17272,16.745028,14.933334,14.10954,13.774771,11.565949,11.408411,11.74318,11.280411,10.463181,11.490462,9.80677,10.125129,10.857026,11.067078,10.466462,10.906258,12.27159,12.491488,11.37559,10.620719,10.8767185,10.748719,10.722463,11.247591,12.724514,11.053949,11.61518,11.188514,9.4916935,9.186462,8.625232,8.530052,9.43918,10.725744,10.604308,11.897437,15.363283,19.695591,21.792822,16.738462,18.632206,30.28349,37.172516,37.80267,43.684105,46.50667,48.656414,51.055595,54.64944,60.42585,66.41888,72.84185,76.32739,78.90052,87.98196,110.798775,118.0554,122.50585,129.62791,137.66237,141.27591,133.51057,108.205956,71.643906,42.528824,34.1399,32.354465,31.858873,29.892925,26.230156,27.818668,29.971695,31.202463,33.506466,42.35816,34.45826,35.075283,35.393642,32.758156,30.67077,34.12677,36.040207,35.813747,34.274464,33.67713,32.58749,32.49231,31.678362,30.398361,30.838156,29.984823,27.464207,25.577028,25.00595,24.81231,24.018053,25.787079,28.399591,29.341541,25.314463,25.337439,26.945642,26.98831,24.986258,23.131899,23.768618,25.163488,26.74872,27.83508,27.602053,25.465437,24.208412,23.122053,22.596926,24.12308,23.256617,22.885746,22.836515,22.87918,22.721643,24.22154,26.033234,27.053951,27.349335,28.166567,28.862362,27.480618,26.079182,25.924925,27.510157,26.82749,29.5319,31.130259,30.503387,29.892925,30.099695,29.528618,29.912617,30.368822,27.38872,25.888823,24.507078,24.566156,25.475285,24.720411,23.729233,23.483078,23.519182,23.24677,21.943796,20.978874,21.543386,22.212925,22.354053,22.111181,26.90954,26.194054,25.570463,26.476309,26.184208,22.642874,21.336617,19.88595,18.110361,18.034874,0.69251287,0.58092314,0.54482055,0.57764107,0.6629744,0.7450257,0.69907695,0.60061544,0.47917953,0.4004103,0.48246157,0.47261542,0.42338464,0.39712822,0.40369233,0.40369233,0.34133336,0.3052308,0.27897438,0.2855385,0.3708718,0.41025645,0.42338464,0.4201026,0.42994875,0.50543594,0.6662565,0.5973334,0.5874872,0.7187693,0.8533334,0.85005134,1.020718,1.142154,1.3423591,2.1070771,2.03159,2.034872,2.1858463,2.5074873,2.9735386,3.56759,3.6824617,3.6496413,3.751385,4.210872,3.6430771,3.9253337,4.0992823,3.8596926,3.570872,3.8367183,3.8104618,3.9056413,4.276513,4.844308,5.605744,5.622154,5.504,5.3792825,4.8705645,4.6867695,5.0215387,5.3891287,5.467898,5.10359,5.7042055,6.042257,6.3606157,6.672411,6.73477,7.5520005,7.9130263,7.8145647,7.5454364,7.702975,7.6110773,7.8834877,8.4053335,8.756514,8.2215395,7.5487185,7.565129,7.8506675,8.188719,8.546462,8.395488,8.392206,7.8736415,7.138462,7.460103,8.247795,8.772923,8.871386,8.569437,8.064001,7.328821,6.665847,6.2588725,6.166975,6.298257,6.3245134,5.8486156,5.2315903,4.5423594,3.564308,3.2623591,3.5216413,3.751385,3.6036925,2.9571285,2.9144619,2.9243078,2.9735386,3.0162053,2.9604106,3.2328207,4.06318,4.857436,5.405539,5.85518,6.226052,6.698667,7.1056414,7.3714876,7.5191803,8.018052,8.392206,8.523488,8.323282,7.719385,7.5946674,7.936001,8.395488,8.881231,9.596719,10.541949,11.237744,11.841642,12.619488,13.938873,14.194873,13.3251295,11.963078,10.709334,10.148104,9.875693,9.393231,8.65477,7.8834877,7.5487185,7.860513,8.438154,8.470975,7.8408213,7.131898,6.875898,6.616616,6.4689236,6.304821,5.730462,5.1856413,4.8114877,4.5456414,4.312616,3.9909747,4.2141542,3.82359,3.446154,3.318154,3.2656412,3.1048207,2.9801028,2.8882053,2.809436,2.7175386,2.356513,2.412308,2.5009232,2.4648206,2.3926156,1.6607181,1.6344616,1.5360001,1.2406155,1.2931283,1.394872,1.7066668,1.9265642,1.9528207,1.8904617,2.0086155,2.3302567,2.3401027,1.9856411,1.7033848,2.2580514,2.6157951,3.0030773,3.2951798,3.0162053,3.570872,3.8465643,3.945026,3.8564105,3.4855387,4.076308,4.3552823,4.4964104,4.5095387,4.2371287,3.754667,3.43959,3.3641028,3.4166157,3.314872,3.6758976,3.8400004,3.895795,4.0008206,4.381539,4.4373336,4.46359,4.352,4.2469745,4.5423594,4.0041027,3.6758976,3.7809234,4.164923,4.2896414,4.8016415,4.1452312,3.5052311,3.373949,3.5544617,3.8465643,3.6496413,3.5511796,3.7842054,4.2371287,3.7448208,3.446154,3.3608208,3.3247182,2.9997952,2.5271797,2.681436,2.8488207,2.878359,3.0785644,2.484513,2.2777438,2.4418464,2.7733335,2.8750772,2.7044106,2.7634873,2.9669745,2.9735386,2.1924105,1.9692309,1.4966155,1.4211283,1.7001027,1.6246156,1.6180514,1.723077,1.7920002,1.8379488,2.044718,2.7700515,2.6715899,2.6584618,2.8947694,2.793026,1.8970258,1.5491283,1.3587693,1.1651284,1.0469744,1.2406155,1.0371283,0.88287187,0.764718,0.2297436,0.51856416,0.5415385,0.6892308,0.9485129,0.9156924,1.1782565,0.9288206,1.1191796,1.4933335,0.60061544,2.1530259,3.8728209,6.2884107,7.450257,2.9571285,2.2121027,5.76,5.976616,3.9581542,9.540924,5.034667,2.6584618,1.2340513,0.318359,0.20676924,0.14112821,0.14441027,0.22646156,0.35774362,0.45620516,0.48574364,0.67282057,0.61374366,0.3314872,0.28225642,0.40697438,0.26256412,0.15097436,0.16082053,0.17723078,0.3117949,0.5907693,0.88943595,1.2307693,1.8116925,2.412308,2.9965131,4.893539,7.0432825,6.009436,7.6767187,9.872411,11.283693,11.631591,11.651283,13.312001,14.050463,13.11836,10.650257,7.637334,8.986258,10.125129,10.912822,11.1983595,10.84718,11.030975,11.057232,11.565949,12.3076935,12.114052,13.016617,14.043899,14.651078,14.283488,12.402873,11.040821,9.990565,9.114257,8.36595,7.7981544,7.906462,7.634052,7.6077952,7.765334,7.3321033,6.2884107,5.6385646,6.0750775,7.3682055,8.385642,8.4512825,8.533334,8.411898,7.7292314,5.989744,7.253334,9.353847,11.641437,12.905026,11.382154,6.2720003,4.141949,3.255795,2.422154,0.99774367,0.79425645,3.639795,4.6112823,3.3903592,4.279795,3.508513,4.8804107,5.211898,4.4964104,5.8880005,3.751385,4.082872,5.142975,6.2030773,7.5552826,5.028103,6.1440005,6.3540516,5.031385,5.4908724,5.2644105,3.9417439,3.9384618,4.9460516,3.9581542,7.1483083,6.6067696,5.2512827,4.568616,4.6145644,7.1614366,4.919795,4.716308,7.24677,7.066257,11.556104,16.68595,17.060104,12.668719,8.881231,12.488206,13.617231,12.84595,9.7673855,2.9833848,9.242257,12.455385,9.45559,3.0687182,2.1202054,3.0687182,5.2414365,10.33518,15.471591,13.197129,6.7183595,8.470975,12.137027,14.536206,15.632411,11.264001,9.872411,9.800206,9.8592825,9.32759,9.412924,10.732308,10.249847,8.185436,8.041026,9.760821,8.021334,9.278359,12.36677,8.500513,10.79795,10.115283,8.789334,8.605539,10.804514,5.8847184,4.667077,5.474462,6.6034875,6.3376417,6.9809237,7.752206,8.375795,9.061745,10.509129,9.688616,10.157949,10.811078,11.073642,10.893129,10.8307705,10.686359,10.873437,11.195078,10.8537445,10.758565,11.388719,10.962052,9.494975,8.792616,8.392206,6.7117953,9.833026,15.012104,10.699488,8.818872,9.209436,10.361437,10.804514,9.081436,9.035488,8.956718,9.396514,9.961026,9.337437,9.393231,10.20718,11.0375395,11.451077,11.34277,11.877745,12.596514,13.144616,13.351386,13.22995,11.18195,11.88759,13.863386,16.000002,17.562258,17.80513,18.179283,17.785437,17.014154,17.555695,17.85436,17.339079,17.378464,17.929848,17.526155,17.132309,17.02072,16.292105,14.76595,13.00677,12.534155,12.3766165,11.424822,10.20718,10.880001,9.488411,9.31118,9.393231,9.5146675,10.174359,10.427077,10.896411,11.585642,11.733335,9.813334,9.954462,9.862565,10.571488,11.949949,12.714667,10.699488,12.580104,13.105232,11.45436,11.237744,10.627283,10.541949,11.132719,11.782565,11.1064625,13.659899,15.891693,17.348925,18.054565,18.507488,20.46031,34.563286,43.47077,42.673233,40.500515,45.604107,47.573338,50.832413,56.01149,59.9598,67.508514,75.98277,82.92432,91.726776,111.64883,147.74811,155.97293,154.28596,150.10135,140.31427,127.481445,112.41354,94.26708,74.863594,58.637135,51.081852,40.900925,32.256004,28.714668,33.237335,34.84226,35.245953,34.1399,33.14544,35.8039,34.87836,38.262157,40.81231,40.39549,37.894566,35.219696,34.113644,33.13231,31.917952,31.222157,30.585438,31.222157,31.064617,30.25395,31.143387,31.205746,29.728823,28.343798,27.825233,28.071386,28.137028,28.632618,28.55713,27.454361,25.4359,25.14708,25.288208,24.832003,24.027899,24.388926,24.615387,25.225847,25.977438,26.423798,25.918362,24.388926,24.103386,24.33313,24.546463,24.392206,23.273027,23.509335,23.840822,23.768618,23.561848,24.566156,26.072617,26.548515,26.328617,27.605335,31.08431,30.33272,28.87549,27.969643,26.597746,27.26072,28.347078,29.925745,31.40595,31.527388,30.864412,30.116104,29.751797,29.59754,28.816412,27.2279,24.87795,23.78831,24.208412,24.635078,21.838772,21.316925,21.622156,22.272001,23.748924,20.841026,21.622156,22.889027,22.711796,20.437334,24.297028,26.161232,26.935797,26.978464,26.098873,24.18872,23.18113,21.346462,18.740515,17.18154,0.7187693,0.63343596,0.6170257,0.60389745,0.56123084,0.5021539,0.45620516,0.380718,0.32164106,0.2986667,0.2855385,0.29210258,0.30851284,0.3314872,0.33805132,0.28225642,0.23958977,0.2231795,0.22646156,0.25928208,0.35774362,0.35774362,0.41682056,0.42994875,0.39384618,0.40697438,0.6301539,0.574359,0.53825647,0.6432821,0.8467693,0.90912825,0.90912825,0.9353847,1.211077,2.0939488,2.2711797,2.097231,2.1891284,2.6420515,3.0490258,4.0303593,4.1682053,4.1846156,4.3060517,4.2863593,3.5610259,3.9417439,4.352,4.4734364,4.7228723,4.6178465,4.2863593,3.9975388,4.07959,4.923077,5.687795,5.874872,5.4613338,4.713026,4.1682053,4.1517954,4.3749747,4.7360005,5.0510774,5.0609236,5.792821,6.0717955,6.3376417,6.6527185,6.7183595,7.466667,7.8539495,7.821129,7.515898,7.282872,7.683283,8.208411,8.789334,9.107693,8.5891285,7.64718,7.197539,7.1548724,7.453539,8.018052,8.021334,7.8408213,7.351795,6.872616,7.141744,7.702975,7.75877,7.6143594,7.4929237,7.525744,7.387898,7.565129,7.6143594,7.328821,6.7577443,6.9152827,6.6560006,6.245744,5.7042055,4.7917953,4.345436,4.3716927,4.4832826,4.4373336,4.1517954,4.096,3.9220517,3.7809234,3.764513,3.892513,4.3684106,5.146257,5.865026,6.439385,7.0465646,7.463385,7.9983597,8.4972315,8.805744,8.746667,8.346257,8.41518,8.825437,9.219283,8.992821,9.570462,10.184206,10.571488,10.761847,11.067078,12.002462,12.425847,13.078976,14.01436,14.605129,14.601848,14.10954,13.298873,12.347078,11.444513,11.149129,10.673231,9.905231,9.176616,9.268514,8.910769,8.572719,8.408616,8.43159,8.500513,7.79159,7.53559,7.4699492,7.315693,6.76759,6.265436,5.4941545,4.8804107,4.5489235,4.352,4.394667,3.9253337,3.6036925,3.5511796,3.3772311,3.6135387,3.7973337,3.8104618,3.5872824,3.1277952,2.681436,2.6486156,2.7076926,2.6486156,2.3958976,1.8674873,1.8379488,1.7920002,1.5360001,1.2012309,1.7493335,2.0644104,2.0578463,1.8937438,1.9954873,2.172718,2.428718,2.5928206,2.5895386,2.4549747,2.4024618,2.6157951,3.058872,3.4756925,3.370667,3.6758976,4.092718,4.4077954,4.322462,3.4625645,4.017231,4.384821,4.568616,4.562052,4.3585644,3.9089234,3.636513,3.5347695,3.4888208,3.2853336,3.6627696,4.2863593,4.647385,4.6933336,4.8049235,5.100308,5.159385,4.906667,4.5029745,4.352,4.138667,3.9384618,3.9417439,4.092718,4.07959,4.630975,4.4767184,4.013949,3.5807183,3.4822567,3.82359,3.6135387,3.4166157,3.5840003,4.2469745,4.0369234,3.7743592,3.620103,3.5840003,3.508513,2.9407182,2.8947694,3.249231,3.6594875,3.570872,2.9111798,2.7142565,2.6518977,2.665026,2.9571285,2.8291285,2.733949,2.7798977,2.6978464,1.847795,1.7788719,1.6738462,1.847795,2.2219489,2.3236926,2.284308,2.28759,2.2646155,2.1825643,2.0512822,2.28759,2.4418464,2.6289232,2.7963078,2.733949,1.9200002,1.5688206,1.4309745,1.3817437,1.4408206,1.1749744,1.0043077,0.7417436,0.37743592,0.101743594,0.36758977,0.9288206,1.1060513,0.88287187,0.9156924,1.3259488,0.8369231,0.6859488,1.1323078,1.4539489,4.069744,4.588308,4.519385,4.4832826,4.201026,2.8291285,6.1997952,7.1876926,5.1265645,5.83877,2.802872,1.5195899,0.7778462,0.17394873,0.08533334,0.06235898,0.12471796,0.20676924,0.26584616,0.29210258,0.24615386,0.25928208,0.19692309,0.108307704,0.22646156,0.28225642,0.18051283,0.09189744,0.0951795,0.18379489,0.42338464,0.6826667,1.0108719,1.4375386,1.9790771,2.540308,3.1638978,5.7665644,8.904206,7.762052,7.765334,9.819899,11.762873,13.131488,15.16636,15.573335,14.976001,13.656616,12.018872,10.587898,11.730052,12.412719,12.504617,12.120616,11.631591,12.724514,12.150155,11.867898,12.084514,11.250873,11.418258,12.304411,13.016617,12.872206,11.385437,10.180923,9.747693,9.419488,8.743385,7.4929237,7.762052,7.5552826,7.4010262,7.325539,6.8594875,5.543385,5.4514875,5.8847184,6.488616,7.27959,7.8637953,7.8834877,7.640616,7.181129,6.2916927,5.986462,8.165744,11.579078,13.712411,10.804514,6.2884107,4.5128207,3.5774362,2.4188719,0.82379496,1.9626669,5.733744,6.0192823,2.930872,2.8192823,3.1113849,5.041231,5.2053337,3.8531284,4.8836927,3.058872,3.876103,5.3070774,6.180103,6.166975,4.9788723,5.540103,5.83877,5.4482055,5.5204105,3.3969233,3.3641028,3.3017437,2.5961027,2.1464617,4.1452312,4.0434875,4.132103,4.565334,3.3575387,4.6572313,6.0192823,7.5618467,9.324308,11.237744,16.006565,17.900309,15.251694,10.148104,8.4053335,7.9294367,12.081232,12.816411,8.231385,2.550154,14.592001,13.400617,7.890052,3.6036925,2.6945643,3.9712822,5.986462,8.667898,10.610872,9.068309,5.07077,8.802463,12.386462,12.570257,10.712616,10.295795,11.040821,12.25518,12.068104,7.430565,8.28718,10.269539,10.033232,7.634052,6.5345645,8.4972315,7.0957956,9.488411,14.795488,14.076719,13.778052,11.480617,8.917334,7.768616,9.662359,6.1308722,5.146257,5.986462,6.892308,5.080616,5.668103,7.427283,8.231385,8.51036,11.227899,10.33518,10.177642,10.496001,10.985026,11.303386,12.475078,11.818667,11.277129,11.579078,12.242052,10.450052,10.453334,10.276103,9.3078985,8.2904625,7.5191803,5.330052,8.136206,13.338258,9.324308,7.817847,7.7456417,8.723693,9.15036,6.2030773,7.3747697,7.460103,7.6635904,8.267488,8.63836,7.6964107,8.283898,9.222565,10.04636,11.011283,10.322052,9.734565,10.463181,11.877745,11.503591,11.32636,12.839386,14.480412,15.675078,16.840206,18.057848,18.468103,18.487797,18.533745,19.029335,15.904821,15.192616,17.076513,19.104822,16.183796,15.996719,15.711181,14.336001,12.750771,13.696001,12.76718,11.707078,10.650257,9.757539,9.206155,9.777231,9.997129,9.662359,9.393231,10.633847,10.305642,10.70277,11.841642,12.458668,10.016821,10.637129,10.43036,10.752001,11.992617,13.590976,12.104206,13.115078,13.269335,12.278154,12.901745,12.301129,13.141335,13.945437,13.988104,13.308719,16.259283,17.007591,18.710976,21.59918,22.961233,23.14831,37.79939,50.865234,52.77867,40.454567,46.39508,47.9639,50.510773,54.839798,57.22585,65.7198,75.536415,87.14175,102.28513,124.03201,134.29498,130.1596,121.41293,112.04924,100.29293,89.252106,81.450676,74.76842,68.21416,61.89949,51.012928,42.167797,38.324516,39.322258,41.892105,36.325745,33.7198,31.744003,30.529644,32.672825,35.77436,39.341953,40.61867,39.171284,36.89354,35.521645,35.501953,34.884926,33.358772,32.2199,33.02072,33.191387,32.436516,31.232002,30.788925,29.522053,28.85908,28.609644,28.435694,27.858053,27.46749,27.828514,27.972925,27.224617,25.219284,23.394463,22.183386,21.970053,22.833233,24.549746,25.124104,25.383387,25.938053,26.456617,25.662361,24.339695,24.001642,23.958977,23.903181,23.899899,24.021336,23.706259,22.94154,22.268719,22.774155,23.939283,24.933746,25.521233,26.023386,27.319798,31.071182,31.031797,29.59754,28.071386,26.679796,27.85477,28.672003,29.866669,31.021952,30.57231,30.614977,30.276926,29.741951,28.90831,27.37231,26.17108,24.323284,22.826668,22.071796,21.848618,19.580719,19.80718,20.368412,20.965746,23.138464,21.940514,22.107899,22.390156,21.832207,19.780924,22.38031,26.259695,27.641438,25.80677,23.082668,20.79836,20.306053,20.023796,19.285336,18.330257,0.71548724,0.5907693,0.54482055,0.508718,0.44964105,0.38728207,0.38400003,0.34133336,0.2986667,0.26584616,0.190359,0.20348719,0.24615386,0.27569234,0.26256412,0.20348719,0.17394873,0.16738462,0.18379489,0.2297436,0.31507695,0.38400003,0.47917953,0.5021539,0.47917953,0.56451285,0.6629744,0.5874872,0.571077,0.6859488,0.8172308,0.88287187,0.78769237,0.8598975,1.2340513,1.8445129,2.4746668,2.5271797,2.553436,2.789744,3.1343591,4.2469745,4.585026,4.6834874,4.6769233,4.2863593,3.757949,4.0500517,4.535795,4.9526157,5.3825645,4.903385,4.1452312,3.6135387,3.6857438,4.588308,5.2020516,5.481026,5.225026,4.516103,3.692308,3.7349746,3.8662567,4.2338467,4.8049235,5.3760004,5.924103,6.3179493,6.5772314,6.744616,6.885744,7.269744,7.4929237,7.453539,7.2303596,7.0793853,7.6603084,8.152616,8.710565,9.189744,9.143796,8.316719,7.351795,6.744616,6.8004107,7.634052,7.768616,7.4174366,6.918565,6.5050263,6.3343596,6.7216415,6.672411,6.5280004,6.488616,6.6100516,6.957949,7.683283,8.100103,7.8145647,6.7150774,6.9710774,6.8955903,6.616616,6.180103,5.5597954,5.2709746,5.175795,5.179077,5.1889234,5.110154,5.07077,5.0904617,5.1232824,5.1167183,5.0182567,5.2512827,5.8486156,6.439385,6.931693,7.50277,7.9130263,8.434873,9.140513,9.783795,9.7903595,9.120821,9.127385,9.659078,10.440206,11.050668,12.445539,12.970668,12.796719,12.3076935,12.117334,12.642463,13.010053,13.666463,14.516514,14.9398985,14.667488,14.36554,14.17518,14.083283,13.938873,13.39077,12.632616,11.648001,10.86359,11.158976,11.021129,9.987283,9.284924,9.373539,9.944616,9.07159,8.635077,8.379078,8.04759,7.3714876,6.7905645,6.0750775,5.5072823,5.1954875,5.07077,5.07077,4.460308,4.1124105,4.1517954,3.9712822,4.066462,4.135385,4.164923,4.06318,3.623385,3.1573336,3.006359,2.930872,2.7602053,2.3893335,2.03159,1.9692309,1.9495386,1.8445129,1.6180514,2.1891284,2.428718,2.3466668,2.2022567,2.4910772,2.681436,2.6518977,2.6453335,2.6847181,2.6026669,2.4484105,2.6223593,3.0391798,3.5249233,3.82359,4.0533338,4.4242053,4.673641,4.525949,3.7021542,3.9154875,4.1124105,4.273231,4.384821,4.4373336,4.1550775,4.059898,4.0336413,3.9351797,3.5905645,3.9056413,5.0084105,5.5532312,5.225026,4.7622566,5.2381544,5.5138464,5.2348723,4.588308,4.2896414,4.279795,4.3290257,4.2962055,4.20759,4.263385,4.5095387,4.4832826,4.1156926,3.639795,3.5905645,3.7874875,3.6660516,3.5052311,3.5872824,4.210872,4.5128207,4.2568207,3.8859491,3.6758976,3.7284105,3.4494362,3.1934361,3.4888208,4.056616,3.820308,3.2295387,3.006359,2.7864618,2.6420515,3.0720003,3.2032824,3.062154,2.878359,2.5600002,1.7132308,1.5589745,1.8149745,2.2022567,2.5140514,2.6026669,2.6026669,2.5796926,2.556718,2.4024618,1.8313848,1.9462565,2.4320002,2.6551797,2.605949,2.8914874,2.477949,2.1956925,1.8904617,1.6377437,1.7690258,1.2438976,0.9878975,0.5973334,0.16738462,0.30194873,0.35446155,0.92225647,1.0338463,0.76800007,1.2570257,1.2996924,0.69579494,0.30194873,0.69579494,2.176,3.69559,4.6178465,3.4034874,1.5983591,3.8104618,3.6430771,5.5926156,6.1013336,4.7458467,4.2502565,3.2262566,1.7723079,0.67282057,0.190359,0.049230773,0.24287182,0.21333335,0.18707694,0.23302566,0.24287182,0.17394873,0.09189744,0.06564103,0.108307704,0.19692309,0.16410258,0.10502565,0.06564103,0.08205129,0.190359,0.4397949,0.67938465,1.0371283,1.5163078,1.9954873,2.7306669,3.5052311,5.651693,8.36595,8.707283,8.920616,10.633847,13.13477,15.753847,17.828104,16.137848,14.900514,13.922462,13.15118,12.681848,13.50236,13.545027,13.236514,12.865642,12.593232,13.61395,12.832822,12.137027,11.789129,10.433641,9.905231,10.735591,11.483898,11.480617,10.8307705,9.833026,9.409642,9.173334,8.700719,7.522462,7.77518,7.5421543,7.3616414,7.384616,7.3682055,6.0783596,6.0947695,6.232616,6.2162056,6.675693,7.6603084,7.6603084,6.9710774,6.0849237,5.6943593,5.2512827,6.8430777,9.708308,12.419283,12.895181,7.394462,4.6802053,3.0194874,1.654154,0.7811283,2.3302567,5.277539,5.6385646,3.4527183,2.7963078,2.6551797,3.879385,3.9253337,2.9013336,3.5938463,2.8849232,3.826872,5.0477953,5.4941545,4.417641,4.345436,4.516103,4.2601027,3.7776413,4.1222568,2.1366155,2.4615386,2.4943593,1.8838975,2.5600002,2.3860514,2.281026,3.4658465,5.0051284,3.8006158,4.7228723,7.6176414,9.488411,10.082462,11.897437,12.140308,11.477334,8.933744,6.0947695,7.0859494,6.76759,10.456616,10.568206,6.957949,6.928411,16.229744,11.936821,6.012718,3.895795,4.4701543,6.6592827,7.4240007,6.8299494,5.861744,6.416411,5.10359,8.772923,10.312206,8.333129,7.1548724,9.921641,11.490462,12.041847,10.564924,4.850872,6.669129,9.691898,10.049642,7.581539,5.832206,7.4141545,6.9645133,8.776206,12.757335,14.401642,13.35795,11.841642,9.714872,7.9163084,8.461129,6.2916927,5.579488,6.557539,7.259898,3.5446157,4.903385,7.017026,8.090257,8.323282,9.93477,10.148104,10.259693,10.496001,10.824206,10.939077,12.232206,12.074668,11.605334,11.61518,12.547283,9.91836,9.127385,8.920616,8.648206,8.260923,7.1548724,4.5587697,5.664821,10.81436,15.510976,8.845129,5.98318,6.2063594,7.456821,6.298257,7.75877,8.553026,8.65477,8.4283085,8.631796,7.0498466,6.9349747,7.5618467,8.461129,9.429334,7.958975,7.1220517,8.438154,10.801231,10.469745,11.339488,12.599796,13.515489,14.368821,16.456207,18.287592,17.992207,17.99549,18.54359,17.69354,14.221129,14.811898,16.512001,16.502155,12.114052,20.33559,18.451694,13.377642,10.043077,11.408411,11.273847,10.272821,9.521232,9.160206,8.352821,9.120821,9.911796,9.8363085,9.373539,10.371283,10.551796,10.70277,11.575796,12.212514,9.980719,10.962052,11.244308,11.313231,11.910565,14.034052,13.929027,13.919181,13.584412,13.177437,13.6237955,13.348104,14.434463,14.953027,14.578873,14.585437,17.14872,16.54154,18.386053,22.209642,21.441643,23.04,38.327797,47.71118,44.655594,35.725132,39.1319,40.56616,43.936825,49.046978,51.587288,56.572723,64.03939,75.12616,88.50708,100.41109,91.75303,81.06011,71.34196,64.08862,59.277134,54.767593,54.849644,56.352825,57.110977,55.972107,47.169643,44.061543,44.100925,44.468517,42.0759,33.3719,30.401644,29.830566,30.34913,32.68267,37.26113,40.64821,40.39549,37.32349,35.501953,36.03036,36.532516,35.69559,33.73949,32.41026,34.162876,34.454975,34.070976,33.33908,32.15754,29.863386,29.305439,29.518772,29.38749,27.657848,27.024412,27.155695,27.011284,25.872412,23.345232,21.35631,20.962463,22.186668,24.218258,25.38995,25.380104,25.944618,26.696207,26.971899,25.819899,24.799181,24.136208,23.83754,23.91631,24.408617,25.268515,24.297028,22.757746,21.865026,22.78072,23.778463,24.224823,24.943592,26.006977,26.696207,29.206976,29.764925,29.18072,28.228926,27.654566,27.4839,28.435694,29.67631,30.61826,30.900515,30.519796,29.824003,29.161028,28.432413,27.090054,26.138258,24.97313,23.299284,21.31036,19.705437,18.192411,18.770052,19.603693,20.250257,21.638565,22.419695,21.861746,21.22831,20.73272,19.551182,20.768822,25.380104,27.441233,25.412926,22.150566,19.748104,19.22954,19.698874,20.20431,19.721848,0.61374366,0.41025645,0.318359,0.30851284,0.35446155,0.4135385,0.446359,0.42994875,0.36758977,0.27897438,0.19364104,0.20348719,0.2231795,0.2231795,0.20020515,0.16410258,0.13128206,0.128,0.15753847,0.20676924,0.28225642,0.43323082,0.5349744,0.5874872,0.65969235,0.86646163,0.7515898,0.64000005,0.69251287,0.83035904,0.72861546,0.72861546,0.75487185,0.98461545,1.3981539,1.7920002,2.6223593,3.0949745,3.1245131,3.0030773,3.436308,4.1846156,4.6080003,4.8049235,4.781949,4.4832826,4.1517954,4.1846156,4.519385,4.95918,5.179077,4.6112823,3.636513,3.131077,3.3476925,3.9351797,4.4307694,4.6276927,4.824616,4.850872,4.069744,3.9089234,3.9253337,4.1911798,4.7327185,5.5171285,5.901129,6.49518,6.8299494,6.8266673,6.806975,6.885744,7.072821,7.194257,7.3091288,7.702975,7.8802056,8.04759,8.480822,9.110975,9.524513,8.976411,7.955693,7.1548724,7.02359,7.768616,7.939283,7.5487185,6.9645133,6.380308,5.8092313,6.2063594,6.3967185,6.3868723,6.2490263,6.11118,6.560821,7.2205133,7.6570263,7.506052,6.4689236,6.616616,6.5345645,6.2490263,5.901129,5.7435904,5.87159,5.8256416,5.7468724,5.687795,5.618872,5.6418467,6.0980515,6.550975,6.6494365,6.124308,5.970052,6.439385,6.8594875,7.0498466,7.328821,7.830975,8.5661545,9.6754875,10.811078,11.1294365,10.801231,10.761847,11.083488,11.831796,13.072412,14.8709755,15.179488,14.467283,13.354668,12.612924,12.806565,13.420309,14.070155,14.772514,15.927796,15.66195,14.887385,14.575591,15.228719,16.856617,16.272411,14.959591,13.692719,12.918155,12.78359,13.50236,12.409437,11.319796,11.044104,11.408411,10.400822,9.777231,9.31118,8.786052,7.9917955,7.1154876,6.7872825,6.6560006,6.550975,6.488616,6.452513,5.5597954,5.0051284,5.0576415,5.0609236,4.699898,4.33559,4.2568207,4.3716927,4.2240005,3.6529233,3.373949,3.1015387,2.7602053,2.487795,2.1825643,2.1366155,2.169436,2.2219489,2.3368206,2.425436,2.681436,2.8127182,2.861949,3.1967182,3.3444104,3.0227695,2.6223593,2.3696413,2.3401027,2.6157951,2.8717952,3.2000003,3.6791797,4.3716927,4.578462,4.706462,4.634257,4.3552823,3.9844105,3.7809234,3.8301542,4.0402055,4.2929235,4.4800005,4.309334,4.3618464,4.417641,4.3290257,4.017231,4.2994876,5.7731285,6.373744,5.5958977,4.522667,5.1167183,5.717334,5.5204105,4.71959,4.5128207,4.417641,4.516103,4.5456414,4.4800005,4.529231,4.388103,4.2994876,4.0369234,3.751385,3.9778464,4.069744,4.1091285,3.9942567,3.889231,4.240411,4.893539,4.699898,4.1485133,3.6758976,3.6758976,3.692308,3.4231799,3.5183592,3.9680004,4.128821,3.570872,3.2295387,2.917744,2.7536411,3.1540515,3.6463592,3.764513,3.515077,2.9472823,2.1464617,1.5819489,1.8937438,2.3630772,2.5961027,2.5009232,2.6289232,2.7044106,2.8521028,2.8127182,1.9331284,2.1956925,2.7536411,2.8324106,2.6223593,3.2918978,2.986667,2.937436,2.428718,1.6016412,1.4572309,1.1848207,0.86317956,0.5415385,0.36430773,0.58420515,0.44964105,0.47917953,0.508718,0.7056411,1.5885129,0.9714873,0.761436,0.5546667,0.6629744,2.1333334,1.1848207,3.5872824,3.5840003,1.0633847,1.5622566,3.2065644,4.388103,4.0008206,3.570872,7.2172313,5.6352825,2.681436,0.7450257,0.34133336,0.108307704,0.5218462,0.3446154,0.21989745,0.30851284,0.318359,0.20348719,0.12471796,0.1148718,0.15753847,0.17394873,0.101743594,0.06564103,0.068923086,0.118153855,0.19692309,0.36758977,0.64000005,1.0436924,1.5195899,1.9429746,2.9046156,3.7218463,4.6178465,5.835488,7.6176414,9.728001,11.191795,14.276924,17.93313,17.808413,15.067899,14.247386,14.001232,13.75836,13.7386675,13.8075905,13.459693,13.282462,13.298873,12.983796,12.977232,12.484924,12.156719,11.844924,10.624001,9.554052,10.197334,10.840616,10.86359,10.742155,9.567181,8.694155,8.251078,8.064001,7.6668725,7.88677,7.6931286,7.77518,8.224821,8.556309,7.5487185,7.2369237,6.9382567,6.5280004,6.4557953,6.9054365,7.0531287,6.363898,5.179077,4.71959,5.35959,6.0291286,7.4830775,10.400822,15.386257,8.03118,4.1550775,1.8707694,0.7056411,1.6147693,2.3466668,3.0096412,3.8990772,4.716308,4.565334,2.484513,1.8871796,2.0906668,2.5731285,2.9801028,3.43959,3.7809234,3.69559,3.1376412,2.3138463,3.1081028,3.6168208,2.8750772,1.467077,1.529436,2.359795,1.6902566,1.3883078,2.1070771,3.2918978,3.3608208,3.0884104,3.9975388,5.72718,6.0258465,7.351795,8.786052,8.664616,7.4896417,7.906462,4.4242053,4.2240005,4.2601027,4.2535386,6.685539,10.125129,10.866873,8.766359,7.0957956,12.527591,14.998976,10.538668,5.5762057,3.620103,5.2611284,9.665642,9.488411,6.6560006,3.9089234,4.788513,5.225026,7.259898,7.565129,6.3343596,7.282872,10.656821,10.20718,8.418462,6.304821,3.4034874,5.98318,9.347282,9.544206,6.957949,6.3212314,8.438154,8.132924,7.7292314,8.165744,8.986258,9.760821,10.755282,10.597744,9.222565,7.8703594,5.661539,5.1987696,6.4590774,7.2336416,3.114667,4.818052,6.488616,7.9983597,8.809027,7.9786673,8.966565,10.010257,10.84718,11.1294365,10.420513,10.374565,11.280411,11.720206,11.493745,11.638155,9.176616,7.955693,7.578257,7.762052,8.329846,6.9743595,4.9427695,5.2053337,10.620719,23.926155,12.278154,6.157129,4.6211286,6.2555904,9.160206,9.094564,10.771693,11.16554,9.747693,8.493949,6.925129,6.173539,6.2785645,6.87918,7.200821,5.182359,5.7501545,7.9983597,10.361437,10.59118,9.915077,10.312206,11.1294365,12.534155,15.510976,17.562258,16.997746,16.997746,17.45395,14.966155,14.12595,18.468103,18.661745,13.958565,12.166565,30.756105,24.897642,14.421334,9.16677,8.976411,11.306667,11.250873,10.276103,9.248821,8.418462,8.342975,8.930462,9.202872,9.051898,9.252103,10.476309,10.328616,10.640411,11.283693,10.174359,10.548513,11.69395,12.258463,12.42913,13.945437,15.156514,14.739694,14.237539,14.057027,13.456411,13.656616,14.070155,13.873232,13.430155,14.280207,15.862155,14.572309,15.481437,17.723078,14.506668,21.707489,35.941746,35.84985,24.070566,27.224617,26.601028,28.61949,34.14318,41.176617,44.90175,43.959797,46.273643,51.475697,56.277336,54.449234,48.24944,41.951183,37.40554,35.918774,38.268723,38.1998,40.717133,44.242054,46.84144,46.21785,44.419285,46.260517,45.525337,40.884518,35.895798,30.31631,29.223387,30.710155,32.997746,34.43857,38.7118,41.793644,41.133953,37.79939,36.466873,36.80821,36.31262,34.65518,32.462772,31.300926,32.8599,34.04144,34.95713,35.33785,34.517338,32.515285,31.415798,31.10072,30.660925,28.399591,27.72349,26.981745,25.527798,23.35508,21.087181,20.617847,22.127592,24.513643,26.397541,26.138258,25.363695,26.532104,27.431387,27.050669,25.586874,25.032207,24.605541,24.70072,25.19631,25.455591,26.010258,24.81231,23.40759,22.78072,23.371489,23.955694,24.224823,24.838566,25.580309,25.370258,26.696207,27.562668,28.137028,28.41272,28.182976,26.01354,27.178669,28.868925,30.119387,31.822771,29.906054,28.376617,27.470772,27.264002,27.684105,26.742155,25.770668,24.021336,21.586054,19.38708,17.96595,17.772308,18.546873,19.652925,20.086155,21.421951,20.512821,19.75795,19.80718,19.5479,19.797335,23.5159,25.747694,24.894361,22.711796,21.26113,20.663797,20.834463,21.064207,19.994259,0.32164106,0.23630771,0.2231795,0.2297436,0.24287182,0.3052308,0.26912823,0.23958977,0.2231795,0.20348719,0.16738462,0.2297436,0.20676924,0.190359,0.190359,0.15097436,0.128,0.12143591,0.15753847,0.24287182,0.36758977,0.45292312,0.5284103,0.67282057,0.79425645,0.6104616,0.52512825,0.60389745,0.7450257,0.8041026,0.5940513,0.7417436,0.97805136,1.2898463,1.6935385,2.2416413,2.7798977,3.190154,3.370667,3.4724104,3.876103,4.388103,4.571898,4.6211286,4.7261543,5.080616,4.9821544,4.70318,4.325744,4.1780515,4.8377438,4.886975,4.2830772,3.6004105,3.2623591,3.5544617,3.5446157,3.6594875,4.1780515,4.9493337,5.402257,4.6802053,4.1714873,4.066462,4.381539,4.9427695,5.6385646,5.8945646,6.36718,6.7610264,5.8453336,6.4656415,7.3550773,7.9950776,8.251078,8.362667,8.277334,8.198565,8.41518,8.815591,8.92718,8.681026,8.592411,8.562873,8.477539,8.208411,8.136206,7.8145647,7.456821,7.1909747,7.0793853,7.6898465,7.896616,7.683283,7.273026,7.125334,7.125334,7.4010262,7.6767187,7.716103,7.325539,6.885744,6.370462,5.943795,5.8157954,6.2555904,6.7938466,6.6527185,6.2851286,6.0324106,6.117744,6.045539,6.2194877,6.5805135,6.9054365,6.820103,7.2237954,7.6635904,7.509334,6.8627696,6.547693,7.5454364,9.271795,11.155693,12.727796,13.594257,13.216822,12.501334,12.547283,13.269335,13.367796,14.634667,15.274668,15.474873,15.225437,14.296617,14.431181,14.729847,15.281232,16.147694,17.378464,18.064411,16.183796,14.36554,14.611693,18.310566,18.75036,16.771284,15.379693,14.979283,13.380924,14.480412,13.820719,13.075693,12.980514,13.334975,11.628308,11.136001,11.024411,10.774975,10.177642,8.969847,8.556309,8.556309,8.585847,8.27077,8.195283,7.381334,6.5837955,6.183385,6.196513,5.901129,5.6451287,5.4449234,5.175795,4.578462,3.820308,3.3936412,3.0326157,2.7667694,2.9144619,2.9013336,2.8717952,2.8488207,2.8389745,2.8389745,2.5435898,2.8291285,3.2754874,3.5741541,3.5249233,3.5380516,3.43959,3.0194874,2.5862565,2.9768207,3.5741541,3.7776413,3.9318976,4.273231,4.9427695,4.857436,4.781949,4.568616,4.2174363,3.876103,3.436308,3.764513,4.3651285,4.772103,4.578462,4.210872,4.1189747,4.059898,3.9811285,4.027077,4.663795,6.3507695,7.0957956,6.36718,5.097026,5.5236926,5.8880005,5.661539,4.9296412,4.378257,4.391385,3.9745643,4.1189747,4.7360005,4.637539,4.332308,4.8607183,4.9821544,4.565334,4.578462,4.8344617,4.8049235,4.4898467,4.1550775,4.3651285,5.034667,5.35959,4.84759,3.892513,3.7842054,3.6758976,3.4264617,3.4756925,4.1156926,5.5072823,4.824616,4.066462,3.5610259,3.3247182,3.0654361,3.5807183,3.9745643,4.0041027,3.6726158,3.2196925,2.0118976,2.0644104,2.5895386,2.9538465,2.6847181,2.8816411,2.9210258,3.2754874,3.5544617,2.5173335,2.7602053,3.564308,3.882667,3.6594875,3.8301542,2.6453335,2.7700515,2.2777438,0.9714873,0.39712822,0.39712822,0.37743592,0.51856416,0.6695385,0.3511795,0.42338464,0.31507695,0.42338464,0.74830776,0.86974365,0.69907695,2.0020514,2.0151796,1.0601027,2.546872,1.2800001,2.1070771,2.428718,1.6738462,1.2832822,1.7460514,3.7940516,4.896821,5.21518,7.584821,3.82359,1.591795,0.702359,0.571077,0.2297436,0.49887183,0.41025645,0.36102566,0.40369233,0.24287182,0.15753847,0.18379489,0.23958977,0.25928208,0.19692309,0.08861539,0.068923086,0.0951795,0.13784617,0.19692309,0.30851284,0.69251287,1.211077,1.7132308,2.028308,2.6387694,3.2131286,4.1846156,5.2381544,5.3103595,8.14277,11.753027,15.645539,18.038155,15.855591,15.097437,14.523078,13.846975,13.262771,13.459693,12.432411,12.662155,12.84595,12.461949,11.766154,11.483898,11.414975,11.792411,12.22236,11.674257,10.71918,11.08677,11.300103,10.765129,9.764103,8.825437,8.152616,7.834257,7.8112826,7.8736415,8.3364105,8.280616,8.585847,9.252103,9.399796,8.605539,7.968821,7.24677,6.3212314,5.172513,4.893539,5.2414365,5.579488,5.5893335,5.293949,6.47877,7.716103,9.865847,12.12718,12.0549755,4.716308,2.4451284,1.394872,1.1388719,4.6539493,4.604718,3.0358977,2.8717952,4.699898,6.774154,3.2098465,2.0086155,2.8750772,3.9581542,1.847795,3.6890259,3.3805132,2.5764105,2.4582565,3.754667,2.6551797,1.3193847,1.148718,1.785436,1.1126155,1.9922053,1.8904617,1.4276924,1.1946667,1.7558975,4.9296412,5.658257,5.792821,5.756718,4.5456414,6.157129,7.6701546,6.5345645,3.9417439,4.8082056,6.918565,7.8408213,8.395488,9.176616,10.541949,11.227899,12.278154,9.645949,5.861744,10.026668,15.9343605,11.139283,5.5893335,3.1245131,1.463795,10.30236,11.762873,9.301334,6.1440005,5.2644105,6.373744,6.314667,8.329846,11.149129,9.002667,10.358154,7.5552826,6.5017443,7.3091288,4.31918,6.7216415,8.139488,6.8463597,4.903385,8.162462,12.022155,10.230155,7.939283,6.701949,4.457026,5.5072823,7.719385,9.885539,10.44677,7.4929237,4.7950773,4.716308,5.7042055,6.229334,4.775385,4.2994876,5.58277,8.274052,10.666668,9.688616,8.077128,8.39877,9.412924,10.262975,10.482873,9.895386,9.924924,10.870154,12.07795,11.933539,9.186462,7.958975,7.4207187,7.4010262,8.375795,7.0334363,6.7544622,7.893334,11.254155,18.067694,18.12677,11.395283,4.7983594,2.5337439,6.0717955,3.3017437,4.594872,5.805949,5.3792825,4.378257,3.3772311,3.3378465,3.7973337,4.8344617,7.0793853,4.066462,4.9329233,5.8289237,6.196513,8.759795,6.951385,8.999385,10.597744,10.627283,11.139283,12.225642,14.437745,17.001026,17.992207,14.342566,14.198155,27.579079,31.566772,25.714874,32.08862,41.488415,26.902977,14.372104,12.872206,14.313026,20.197744,20.450462,16.823795,11.631591,7.7357955,10.666668,9.091283,8.155898,8.946873,8.484103,8.690872,9.403078,10.420513,11.592206,12.786873,10.601027,11.766154,13.538463,14.470565,14.434463,15.107284,14.358975,13.686155,13.492514,13.075693,13.308719,13.275898,13.072412,13.033027,13.718975,14.011078,13.423591,13.620514,14.043899,11.933539,25.957747,31.862156,30.631388,26.026669,24.612104,24.12308,27.894156,33.35549,38.429543,41.517952,40.139492,39.27303,39.263184,39.456825,38.226055,38.724926,38.912003,38.767593,38.304825,37.599182,39.696415,41.028927,42.24985,42.55508,39.67344,39.233643,40.20513,40.434875,39.299286,37.687798,34.710976,33.05026,33.204514,34.56,35.41662,38.76103,39.67016,39.207386,38.2359,37.428516,36.98872,36.72616,35.35098,33.194668,32.180515,32.548103,33.929848,34.825848,34.71426,34.04144,33.10277,31.422361,30.260515,29.669746,28.471798,26.361439,24.25108,22.86277,22.357334,22.308104,23.076105,23.361643,23.204103,22.98749,23.45354,24.953438,26.089027,26.43036,25.816618,24.352823,24.119797,25.37354,26.164515,25.711592,24.369232,24.454565,23.476515,22.50831,21.979898,21.697643,22.770874,23.909746,24.264208,23.781746,23.207386,25.554052,26.312206,26.581335,26.584618,25.682053,24.313438,26.095592,27.749746,28.100925,28.077951,26.246567,25.347284,24.310156,23.460104,24.520206,23.77518,22.465643,21.018257,19.961437,19.912207,18.264616,16.150976,15.796514,17.302977,18.645334,19.121233,18.44513,18.162872,18.82913,19.987694,20.548925,21.753437,21.632002,20.027079,18.586258,18.51077,19.508514,20.5719,20.555489,18.189129,0.3314872,0.3249231,0.28225642,0.23958977,0.21661541,0.21989745,0.19364104,0.20348719,0.2100513,0.19692309,0.18051283,0.2297436,0.2297436,0.20676924,0.18051283,0.15097436,0.14769232,0.15425642,0.20348719,0.3052308,0.4266667,0.5316923,0.512,0.5316923,0.61374366,0.6465641,0.6695385,0.6498462,0.72861546,0.9288206,1.1815386,1.142154,1.1651284,1.3587693,1.8379488,2.7175386,2.8947694,3.0752823,3.4034874,3.7743592,3.826872,3.948308,4.4964104,5.2053337,5.8157954,6.0816417,5.917539,5.2512827,4.7917953,4.781949,5.031385,4.8672824,4.709744,4.1714873,3.43959,3.2754874,3.4494362,3.889231,4.4406157,4.965744,5.32677,5.21518,4.781949,4.450462,4.5390773,5.284103,5.6287184,6.114462,6.7872825,7.250052,6.636308,7.076103,8.480822,9.527796,9.731283,9.458873,8.858257,8.740103,8.756514,8.700719,8.500513,8.78277,9.02236,8.953437,8.598975,8.283898,8.36595,8.4283085,8.385642,8.3364105,8.569437,8.937026,8.802463,8.667898,8.585847,8.1755905,7.7357955,7.762052,7.6767187,7.2960005,6.8365135,6.2588725,6.226052,6.1997952,6.157129,6.5969234,7.194257,7.2861543,6.9743595,6.554257,6.5345645,6.518154,6.8332314,6.9677954,6.882462,6.99077,7.637334,8.0377445,7.90318,7.3550773,6.9120007,6.9645133,7.765334,8.792616,9.915077,11.385437,12.051693,12.235488,12.156719,12.2157955,12.977232,15.192616,17.09949,17.634462,16.554668,14.457437,14.775796,15.386257,16.154257,17.174976,18.760206,19.324718,17.08636,15.195899,15.478155,18.44513,19.938463,18.714258,17.207796,16.531694,16.49559,15.8654375,15.829334,15.287796,14.116103,13.154463,11.592206,12.343796,12.750771,12.327386,12.763899,10.9915905,10.509129,9.764103,8.749949,9.025641,8.681026,8.162462,7.6767187,7.253334,6.76759,6.2916927,6.2227697,5.989744,5.467898,4.969026,4.2896414,4.0369234,3.8465643,3.6496413,3.6594875,3.3247182,3.4330258,3.4724104,3.31159,3.2032824,3.3214362,3.4592824,3.7284105,3.9778464,3.7809234,3.754667,3.8071797,3.5872824,3.0818465,2.6223593,3.6496413,4.585026,5.0149746,5.1200004,5.664821,5.3234878,4.900103,4.6867695,4.6802053,4.571898,4.3651285,3.5446157,3.2065644,3.7316926,4.785231,4.8672824,4.706462,4.4438977,4.1780515,3.9417439,4.332308,5.543385,6.7183595,7.0957956,6.012718,5.5696416,5.648411,5.3760004,4.7983594,4.903385,5.0642056,4.4110775,4.1452312,4.4996924,4.7228723,4.4865646,5.2676926,5.691077,5.3234878,4.663795,4.4996924,4.4701543,4.519385,4.594872,4.6572313,5.0838976,5.1856413,4.8836927,4.325744,3.892513,4.1550775,4.394667,4.571898,4.768821,5.2020516,5.428513,4.9854364,4.522667,4.1452312,3.4198978,3.387077,3.6430771,3.9876926,4.164923,3.879385,2.6715899,2.806154,3.2098465,3.3641028,3.3214362,3.6726158,3.7054362,3.4855387,3.186872,3.114667,3.0490258,3.4855387,3.8662567,4.0500517,4.31918,3.2918978,2.3204105,1.4966155,0.8467693,0.3117949,0.41025645,0.48246157,0.4955898,0.46276927,0.44964105,0.7187693,0.5973334,0.508718,0.6826667,1.1881026,1.5622566,1.3620514,0.80738467,1.086359,4.342154,4.673641,4.6867695,3.6036925,1.8412309,1.0010257,2.1202054,3.2328207,4.096,4.332308,3.4100516,2.6945643,1.591795,0.88287187,0.67610264,0.4135385,0.35774362,0.39384618,0.56123084,0.6859488,0.39056414,0.31507695,0.2986667,0.27569234,0.21333335,0.11158975,0.052512825,0.04594872,0.08533334,0.14112821,0.17394873,0.36102566,0.77456415,1.2077949,1.657436,2.297436,3.2000003,3.2262566,3.4691284,4.713026,7.4207187,9.783795,13.98154,16.968206,17.207796,14.680616,15.018668,14.900514,14.516514,14.276924,14.811898,13.4859495,12.504617,12.265027,12.517745,12.337232,11.490462,9.908514,9.350565,10.213744,11.539693,11.533129,11.608616,11.32636,10.377847,8.605539,8.621949,8.408616,7.9195905,7.565129,8.192,8.03118,8.385642,8.979693,9.668923,10.459898,9.95118,9.127385,7.8703594,6.380308,5.1856413,5.159385,4.9362054,5.0477953,5.5729237,6.1505647,7.1680007,8.385642,11.053949,13.63036,11.808822,4.2962055,1.9003079,1.2012309,1.8379488,6.498462,5.3924108,4.5128207,4.1156926,4.3651285,5.346462,4.1550775,5.2742567,6.422975,5.756718,1.8576412,3.3509746,2.294154,1.2012309,1.3357949,2.7175386,2.028308,1.8116925,1.7033848,1.5622566,1.467077,2.5140514,2.3729234,1.9396925,1.9889232,3.1967182,5.4908724,5.58277,5.5302567,5.8092313,5.3037953,5.431795,5.970052,5.3924108,4.1025643,4.453744,5.1987696,6.5378466,7.200821,6.304821,3.367385,5.182359,6.8529234,6.229334,4.6211286,6.803693,10.9915905,11.569232,9.009232,4.844308,1.6607181,3.9844105,4.673641,4.325744,3.5347695,2.858667,10.827488,11.247591,12.274873,14.424617,10.5780525,12.73436,8.805744,8.113232,10.627283,6.99077,6.0849237,6.1538467,5.8125134,5.865026,9.298052,10.33518,8.516924,7.253334,7.1614366,6.0652313,6.8529234,7.6077952,9.130668,10.085744,7.017026,6.6822567,5.9995904,5.9634876,6.2227697,5.093744,5.097026,5.7074876,6.987488,8.3823595,8.713847,8.897642,9.068309,9.3768215,9.895386,10.604308,10.633847,10.082462,10.066052,10.70277,11.10318,8.835282,7.88677,7.8145647,8.4512825,9.915077,8.201847,8.868103,8.661334,8.241231,12.182976,27.77272,19.367386,9.088,7.6570263,14.408206,10.584617,15.195899,17.204514,13.745232,10.115283,11.802258,9.340718,7.4174366,7.6110773,8.421744,8.923898,8.054154,8.864821,11.506873,13.249642,11.178667,14.368821,15.655386,12.724514,8.113232,11.67754,16.042667,17.43754,15.737437,14.441027,17.48677,28.110771,28.865643,19.771078,18.320412,23.561848,19.203283,14.437745,14.575591,21.074053,18.520617,20.289642,23.909746,23.364925,9.091283,8.201847,9.048616,9.219283,8.51036,8.937026,9.905231,9.209436,8.539898,8.989539,11.053949,9.865847,10.06277,11.168821,12.750771,14.421334,14.293334,12.780309,11.85477,12.084514,12.626052,13.610668,13.991385,13.853539,13.643488,14.181745,13.193847,13.203693,14.290052,16.57436,20.233849,39.171284,34.740517,26.10872,23.315695,27.26072,25.426054,25.744411,27.930258,30.516516,30.851284,33.53272,35.22954,35.83016,35.925335,36.78195,37.264412,36.90667,35.324722,33.13231,31.947489,33.29313,34.349953,36.63426,39.33539,39.30585,37.930668,38.006157,38.47877,38.52472,37.56636,35.27221,33.841232,32.557953,32.20677,35.075283,38.05867,37.75672,36.138668,34.189133,31.90154,33.17826,36.000824,36.470158,34.55672,34.110363,34.153027,34.86195,36.32903,37.54667,36.397953,34.1399,32.531696,31.527388,30.500105,28.228926,25.842875,24.73354,24.083694,23.7719,24.359386,24.628515,24.336412,23.794874,23.302567,23.122053,22.242464,23.007181,24.365952,25.291489,24.805746,24.631796,25.458874,25.439182,24.503798,24.33313,24.97313,23.522463,21.989746,21.336617,21.464617,21.710772,21.704206,22.20308,23.125336,23.538874,24.467693,24.562874,24.81231,24.976412,23.59467,25.281643,25.75754,25.51467,25.311182,26.134975,25.074873,25.849438,26.584618,25.938053,23.105642,21.520412,20.319181,19.43631,19.24595,20.585028,19.364103,17.703386,17.122463,17.690258,17.99877,18.376207,18.438566,18.428719,18.806156,20.22072,21.602463,21.471182,20.194464,18.425438,17.11918,16.636719,17.85436,18.208822,16.876308,14.769232,0.28882053,0.26584616,0.25928208,0.26912823,0.29538465,0.3249231,0.30851284,0.28225642,0.26256412,0.24943592,0.23958977,0.23630771,0.24943592,0.26256412,0.26584616,0.22646156,0.21989745,0.2297436,0.26912823,0.33805132,0.45292312,0.508718,0.446359,0.508718,0.6662565,0.62030774,0.69907695,0.7450257,0.8533334,1.024,1.1618463,0.9517949,1.1716924,1.5589745,2.1825643,3.4330258,2.5961027,2.9768207,3.3969233,3.498667,3.7415388,4.023795,4.713026,5.474462,5.9470773,5.72718,5.8814363,5.8880005,5.609026,5.2512827,5.346462,5.293949,5.402257,4.9920006,4.161641,3.7710772,4.138667,4.266667,4.2535386,4.315898,4.788513,5.2348723,5.1167183,4.95918,4.9788723,5.113436,5.4514875,5.9634876,6.547693,7.000616,7.020308,7.4830775,8.480822,9.5606165,10.246565,10.056206,9.176616,9.045334,8.969847,8.766359,8.749949,9.163487,9.137232,8.825437,8.474257,8.402052,8.55959,8.953437,9.019077,8.897642,9.426052,9.498257,9.147078,9.097847,9.334154,9.078155,8.713847,8.024616,7.4765134,7.1483083,6.7314878,6.3277955,6.5083084,6.547693,6.370462,6.554257,7.259898,7.5618467,7.6012316,7.4765134,7.250052,7.030154,6.9776416,6.882462,6.7249236,6.685539,7.1680007,7.381334,7.315693,6.961231,6.3179493,5.901129,6.0783596,6.810257,8.182155,10.420513,11.592206,11.72677,11.237744,11.067078,12.714667,15.67836,17.736206,17.719797,16.15754,15.264822,15.770258,16.344616,16.52513,16.928822,19.222977,19.892515,17.903591,15.740719,15.123693,17.014154,18.7799,18.822565,18.340103,17.959387,17.749334,17.30954,16.39713,15.14995,13.761642,12.465232,12.22236,12.809847,13.049437,12.750771,12.744206,12.232206,11.451077,10.482873,9.672206,9.609847,9.209436,8.736821,8.083693,7.4207187,7.204103,6.0225644,6.180103,6.2720003,5.8223596,5.293949,4.824616,4.1747694,3.8137438,3.8137438,3.817026,3.511795,3.8695388,4.0992823,4.0369234,4.138667,4.1452312,4.0500517,4.0402055,4.210872,4.5489235,4.3290257,4.2174363,3.95159,3.5511796,3.31159,4.197744,4.9821544,5.3070774,5.290667,5.533539,5.8847184,5.533539,5.3005133,5.4449234,5.651693,4.955898,4.1682053,3.8498464,4.092718,4.5062566,4.6966157,5.0182567,5.4875903,5.6352825,4.516103,4.2896414,4.9493337,6.0652313,6.8365135,6.0750775,5.3727183,5.8256416,5.7107697,4.9296412,5.0084105,5.431795,4.9854364,4.4996924,4.391385,4.644103,3.9778464,4.565334,5.2676926,5.504,5.2611284,5.1232824,5.093744,4.962462,4.6933336,4.417641,4.9985647,5.5236926,5.664821,5.3070774,4.5522056,4.598154,4.6276927,4.565334,4.571898,5.044513,5.8125134,5.648411,5.425231,5.2578464,4.4800005,4.1911798,4.391385,4.713026,4.7655387,4.125539,3.387077,3.764513,4.1911798,4.197744,3.9089234,4.453744,4.092718,3.5052311,3.170462,3.3476925,3.0030773,3.2754874,3.9876926,4.670359,4.5587697,3.820308,2.484513,1.4145643,0.84348726,0.35446155,0.27897438,0.4397949,0.58092314,0.6301539,0.69251287,1.273436,0.9321026,0.69579494,0.8467693,0.90912825,1.4966155,1.1881026,1.1520001,2.1366155,4.4800005,3.446154,4.0402055,4.0992823,3.4198978,3.7415388,3.1113849,2.802872,3.1081028,3.6890259,3.5905645,2.353231,1.3456411,0.78769237,0.65312827,0.69579494,0.33476925,0.35446155,0.5218462,0.6301539,0.51856416,0.4004103,0.25271797,0.16082053,0.12471796,0.072205134,0.052512825,0.052512825,0.0951795,0.17723078,0.26912823,0.56451285,0.8763078,1.142154,1.4769232,2.1825643,3.6430771,3.6726158,3.820308,5.0576415,7.77518,12.921437,16.23631,17.618053,17.375181,16.219898,15.520822,13.722258,13.692719,15.090873,14.375385,13.702565,12.435693,11.802258,11.930258,11.867898,11.392001,10.112,9.622975,10.35159,11.523283,11.572514,11.434668,11.2672825,10.65354,8.598975,8.52677,8.454565,7.9983597,7.522462,8.113232,7.5191803,8.155898,8.982975,9.7903595,11.211488,11.122872,9.947898,8.395488,6.7085133,4.6572313,4.2601027,3.820308,4.2568207,5.58277,6.9021544,7.768616,8.444718,10.660104,13.334975,12.58995,4.6900516,1.8904617,1.1881026,2.2055387,7.177847,4.7622566,3.7054362,4.9493337,7.0104623,5.970052,4.20759,3.373949,3.1474874,3.0884104,2.6289232,3.7349746,3.4231799,2.2547693,1.2176411,1.7066668,2.231795,1.9987694,1.7066668,1.7001027,1.9692309,1.7362052,1.4211283,1.1355898,1.2668719,2.4943593,4.0992823,4.781949,6.5312824,8.323282,6.1341543,6.491898,4.598154,3.9417439,5.1265645,5.874872,6.1440005,5.2512827,4.824616,4.7917953,3.383795,5.2644105,8.549745,8.845129,6.806975,8.149334,7.702975,9.03877,9.45559,7.453539,2.7175386,3.170462,3.7349746,3.7448208,3.1015387,2.294154,8.247795,12.635899,14.769232,14.362258,11.546257,12.343796,8.89436,8.684308,11.920411,11.523283,6.163693,4.4964104,4.893539,6.5936418,9.691898,6.449231,5.2381544,5.6254363,6.547693,6.304821,6.987488,7.748924,8.172308,7.7718983,5.989744,6.5772314,5.353026,4.850872,5.1889234,4.066462,5.1626673,4.6834874,5.805949,8.467693,9.373539,8.661334,9.284924,9.796924,9.846154,10.187488,10.656821,9.724719,9.45559,9.987283,9.521232,9.665642,9.554052,8.648206,8.01477,10.31877,7.5881033,7.9983597,8.132924,7.0498466,6.2916927,18.041437,18.139898,15.596309,15.980309,21.418669,16.57436,25.317745,29.741951,24.477541,16.68595,15.474873,11.0375395,7.0859494,6.521436,11.431385,12.511181,9.90195,9.097847,11.339488,13.6237955,10.601027,11.053949,10.433641,8.297027,8.297027,9.672206,11.667693,13.02318,14.086565,16.827078,18.064411,22.127592,21.139694,14.933334,11.050668,10.079181,10.729027,14.020925,18.287592,19.206566,12.521027,15.37313,25.370258,31.678362,15.015386,7.3321033,9.892103,11.218052,8.710565,8.644924,7.899898,7.958975,8.43159,9.133949,10.098872,10.587898,10.948924,10.886565,10.9456415,12.524308,12.209231,11.313231,10.837335,11.224616,12.36677,12.498053,13.128206,13.292309,13.111795,13.804309,12.78359,13.814155,14.854566,15.156514,15.27795,31.40267,29.525335,23.988514,22.87918,28.025438,24.546463,25.51467,29.072412,32.8238,33.795284,35.045746,34.79303,34.668312,35.712,38.38031,38.806976,37.333336,35.27221,33.40472,31.996721,32.43323,33.056824,34.258053,35.797337,36.77867,35.636517,35.623386,35.784206,35.712,35.541336,35.564312,34.753643,32.24944,29.646772,30.979284,34.166157,35.022774,34.871796,34.23836,32.853336,31.8359,33.201233,33.782158,33.030567,33.027283,32.308514,32.05908,33.237335,35.186874,35.633232,34.87508,33.447388,31.658669,29.440002,26.338463,24.71713,24.726976,25.27836,25.600002,25.209438,24.470976,23.689848,22.767591,21.897848,21.54995,20.466873,20.923079,21.779694,22.354053,22.409847,22.419695,23.561848,24.2839,24.070566,23.417439,23.43713,22.754463,21.953642,21.609028,22.288412,21.504002,21.366156,22.022566,23.161438,24.031181,24.116514,24.832003,24.999386,24.500515,24.280617,27.67754,26.79795,24.65149,23.22708,23.489643,22.931694,24.01477,25.222567,24.960001,21.559797,19.971283,18.756924,17.969233,18.080822,20.000822,19.534771,18.116924,17.211079,17.178257,17.28,17.545847,18.359797,18.625643,18.290873,18.336823,19.016207,18.58954,17.942976,17.319386,16.305231,16.180513,16.282257,15.730873,14.582155,13.824001,0.26584616,0.2297436,0.26256412,0.3052308,0.34133336,0.38728207,0.3446154,0.29538465,0.27241027,0.27241027,0.256,0.2297436,0.23958977,0.26584616,0.29210258,0.28225642,0.29210258,0.31507695,0.34133336,0.37743592,0.4397949,0.43323082,0.37743592,0.47917953,0.6695385,0.58420515,0.6695385,0.761436,0.8336411,0.88615394,0.9189744,0.7778462,1.083077,1.5655385,2.231795,3.3608208,2.7470772,3.117949,3.3542566,3.245949,3.4789746,4.1747694,5.3825645,6.1440005,6.189949,5.9536414,5.83877,5.9503593,5.8420515,5.5171285,5.402257,5.428513,5.76,5.648411,4.955898,4.1550775,4.164923,4.4110775,4.4045134,4.197744,4.397949,5.10359,5.142975,5.353026,5.720616,5.3694363,5.586052,5.9503593,6.2884107,6.5378466,6.744616,7.125334,7.827693,8.992821,10.134975,10.14154,9.5146675,9.642668,9.682052,9.449026,9.403078,9.324308,8.966565,8.65477,8.549745,8.651488,8.687591,9.452309,9.737847,9.481847,9.787078,9.734565,9.478565,9.5606165,9.924924,9.90195,9.662359,8.684308,7.7718983,7.269744,7.066257,7.1647186,7.4010262,7.2336416,6.8332314,7.1089234,7.6209235,8.018052,8.218257,8.12636,7.6176414,7.00718,6.7216415,6.5772314,6.4295387,6.1538467,6.4065647,6.449231,6.5345645,6.6395903,6.445949,6.121026,6.173539,6.7577443,8.195283,10.965334,12.074668,11.559385,10.587898,10.282667,11.713642,14.86113,16.905848,17.26031,16.682669,17.289848,18.281027,18.14318,17.237335,16.774565,18.81272,20.33231,18.435284,16.049232,14.956308,15.80636,17.532719,18.530462,18.796309,18.281027,16.925539,15.602873,15.143386,14.920206,14.614976,14.217847,14.158771,13.771488,13.095386,12.301129,11.687386,12.179693,11.542975,10.532104,9.7673855,9.737847,9.508103,9.094564,8.4972315,7.906462,7.686565,6.091488,6.173539,6.3212314,5.927385,5.3727183,5.037949,4.4340515,4.135385,4.2469745,4.397949,4.0434875,4.1911798,4.338872,4.3684106,4.5423594,4.578462,4.5423594,4.604718,4.857436,5.3136415,5.156103,5.024821,4.850872,4.71959,4.886975,4.903385,5.175795,5.4153852,5.61559,6.052103,6.636308,6.2916927,5.7796926,5.622154,6.121026,5.2414365,4.788513,4.7491283,4.8016415,4.348718,4.2436924,4.8344617,5.8420515,6.4722056,5.402257,4.7294364,5.172513,5.9995904,6.485334,5.8945646,5.4153852,5.9470773,5.9470773,5.2348723,4.9952826,5.4186673,5.2545643,4.7360005,4.263385,4.417641,4.0008206,4.388103,5.3037953,6.1997952,6.242462,6.11118,5.687795,5.179077,4.785231,4.6933336,5.536821,6.3967185,6.7150774,6.2785645,5.211898,5.0674877,4.8607183,4.8049235,5.1167183,6.045539,6.626462,6.491898,6.3310776,6.186667,5.467898,4.955898,5.0084105,5.1298466,5.0904617,4.9132314,4.84759,4.9394875,4.962462,4.7327185,4.1222568,4.7392826,4.2174363,3.6102567,3.3247182,3.114667,3.1671798,3.4921029,4.201026,4.893539,4.6802053,4.493129,3.2131286,1.8018463,0.8205129,0.446359,0.25271797,0.36430773,0.7778462,1.2373334,1.2373334,1.5622566,1.1191796,0.8730257,1.024,0.9944616,2.484513,2.9407182,3.255795,3.564308,3.2656412,3.190154,4.4110775,5.1298466,5.3431797,6.8660517,3.7710772,2.6157951,2.6912823,3.31159,3.8071797,2.92759,1.7263591,0.86646163,0.6104616,0.8172308,0.38400003,0.3314872,0.4201026,0.48574364,0.43323082,0.35446155,0.17394873,0.07548718,0.09189744,0.098461546,0.09189744,0.101743594,0.17723078,0.318359,0.48902568,0.72861546,0.88615394,0.98461545,1.3981539,2.858667,4.020513,4.5128207,4.6539493,5.658257,9.626257,15.763694,16.538258,16.098463,16.54154,17.939693,15.629129,12.649027,12.898462,15.172924,13.170873,11.98277,11.572514,11.155693,10.538668,10.112,10.522257,10.266257,10.180923,10.499283,10.81436,11.539693,11.493745,11.385437,10.939077,8.910769,8.448001,8.392206,8.011488,7.4797955,7.8834877,7.496206,8.27077,9.209436,10.223591,12.12718,11.963078,10.522257,8.854975,7.200821,4.9985647,3.9975388,3.4002054,3.882667,5.405539,7.2205133,7.282872,7.712821,9.540924,12.018872,12.603078,5.0149746,2.0939488,1.3686155,2.0611284,5.097026,3.3608208,2.2416413,3.508513,5.8223596,4.7228723,3.0752823,1.2668719,1.913436,4.663795,6.1997952,5.2742567,5.037949,4.4734364,3.31159,2.048,3.0227695,2.425436,1.8904617,1.8904617,1.723077,1.0568206,0.86317956,0.955077,1.463795,2.8225644,5.504,7.056411,8.615385,9.531077,7.3780518,6.157129,3.2951798,2.6683078,4.7524104,6.6067696,7.4240007,6.121026,5.1364107,4.7458467,3.0785644,4.9493337,8.425026,8.854975,6.810257,8.080411,5.0149746,8.625232,12.553847,12.57354,6.5739493,3.9942567,3.876103,4.824616,5.6943593,5.602462,7.3649235,11.493745,12.757335,10.801231,10.125129,10.811078,10.781539,11.145847,12.028719,12.57354,8.864821,5.796103,5.0182567,6.7872825,9.947898,4.598154,3.2886157,4.384821,6.1472826,6.7183595,6.485334,7.1548724,7.565129,7.39118,7.1548724,5.428513,3.8432825,3.8104618,4.8311796,4.5095387,5.2709746,3.6758976,3.8301542,6.304821,8.136206,7.9163084,7.6701546,7.456821,7.315693,7.2894363,7.509334,6.875898,7.7390776,9.321027,7.7325134,8.845129,9.393231,8.887795,8.257642,9.852718,7.4174366,6.892308,7.0531287,6.7905645,5.110154,7.5552826,10.820924,13.380924,14.857847,16.019693,12.855796,20.719591,24.375797,19.846565,14.411489,14.8709755,13.459693,9.245539,5.9569235,11.992617,14.8020525,13.59754,11.802258,11.178667,11.828514,8.858257,7.6964107,8.379078,9.80677,9.737847,8.172308,7.4010262,7.640616,10.085744,16.91241,14.831591,13.430155,12.163283,10.817642,9.524513,5.149539,6.6002054,12.2847185,16.896002,11.434668,9.15036,12.274873,23.699694,33.58195,19.324718,9.409642,9.701744,10.5780525,9.153642,9.284924,6.633026,6.7872825,8.274052,9.475283,8.602257,10.082462,10.400822,10.131693,9.8363085,10.059488,9.744411,9.5606165,9.580308,10.095591,11.628308,11.211488,12.028719,12.320822,12.179693,13.564719,12.973949,13.718975,14.221129,13.144616,9.370257,19.682463,20.319181,19.157335,21.241438,28.757336,27.30995,30.099695,31.048208,30.181746,33.62462,35.08185,34.6158,34.27775,35.00308,36.581745,37.254566,36.28308,34.514053,32.610462,31.03836,30.303183,31.337029,32.57108,33.47036,34.533745,34.02503,33.079796,32.452927,32.518566,33.26359,33.529438,32.92226,30.848001,28.353643,28.117336,31.537233,32.932106,33.204514,32.994465,32.712208,31.320618,31.684925,32.01641,31.80308,31.822771,31.27795,30.82831,31.304207,32.39713,32.66626,33.155285,32.400414,30.765951,28.51118,25.787079,24.608822,24.753233,25.544207,25.849438,24.080412,22.889027,22.304823,21.700924,21.054361,20.949335,20.138668,19.876104,19.862976,20.246977,21.622156,21.454771,21.93395,22.596926,22.918566,22.324514,22.373745,22.672413,22.567387,22.183386,22.432823,21.064207,21.024822,21.888002,23.09908,23.96554,23.808002,24.87795,25.051899,24.323284,24.763079,27.27713,26.49272,24.776207,23.70954,24.113234,23.243488,23.975386,24.562874,23.903181,21.553232,20.397951,19.094976,18.12349,17.98236,19.190155,18.917746,18.198977,17.424412,16.994463,17.302977,17.348925,18.41559,18.930874,18.596104,18.379488,18.228514,17.319386,16.613745,16.17395,15.163078,15.343591,14.86113,14.247386,13.830565,13.75836,0.256,0.24943592,0.2855385,0.30851284,0.30851284,0.32820517,0.26256412,0.23302566,0.24287182,0.26584616,0.23958977,0.2297436,0.23630771,0.24943592,0.27241027,0.30851284,0.35446155,0.38400003,0.40369233,0.41682056,0.39712822,0.37415388,0.36102566,0.43323082,0.5546667,0.5481026,0.69251287,0.74830776,0.72861546,0.7056411,0.81066674,0.90912825,1.0929232,1.4867693,2.0906668,2.789744,3.373949,3.318154,3.2164104,3.2886157,3.3805132,4.44718,6.2030773,7.0432825,6.9021544,7.240206,6.51159,6.0258465,5.8092313,5.648411,5.0904617,5.028103,5.58277,5.8518977,5.3858466,4.1714873,3.757949,4.4307694,4.95918,4.9296412,4.7524104,5.2348723,5.2545643,5.7632823,6.557539,6.2916927,6.0291286,6.23918,6.436103,6.426257,6.3310776,6.629744,7.207385,8.293744,9.4916935,9.764103,9.810052,10.368001,10.643693,10.397539,9.938052,9.281642,8.891078,8.858257,9.02236,8.960001,8.812308,9.754257,10.233437,9.921641,9.682052,9.770667,9.895386,10.128411,10.43036,10.620719,10.345026,9.540924,8.500513,7.7292314,7.9228725,8.477539,8.536616,8.011488,7.466667,8.109949,8.231385,8.585847,8.667898,8.27077,7.4830775,6.685539,6.4722056,6.409847,6.232616,5.8125134,5.8978467,5.796103,6.0225644,6.6395903,7.2631803,7.4108725,7.6668725,8.041026,9.051898,11.736616,12.566976,11.490462,10.299078,9.852718,10.092308,12.947693,15.396104,17.299694,18.753643,20.112411,20.923079,19.56431,17.690258,16.705643,17.77559,20.374975,18.57313,16.420103,15.658668,15.701335,16.659693,18.028309,18.691284,17.99877,15.753847,12.704822,13.90277,15.711181,16.649847,17.385027,16.193642,15.130258,13.712411,12.09436,11.073642,11.303386,11.030975,10.072617,9.048616,9.3768215,9.43918,9.206155,8.953437,8.661334,7.9983597,6.5837955,6.3245134,6.193231,5.7698464,5.2709746,4.8836927,4.7983594,4.8672824,5.0051284,5.1659493,4.841026,4.4996924,4.2994876,4.2929235,4.450462,4.7983594,5.0510774,5.402257,5.789539,5.8978467,6.0783596,6.1440005,6.170257,6.2785645,6.6625648,5.799385,5.6287184,5.835488,6.3212314,7.1876926,7.2336416,6.764308,6.0028725,5.467898,5.9602056,5.3924108,5.0477953,5.10359,5.2414365,4.6572313,4.1780515,4.5390773,5.3136415,5.907693,5.579488,5.159385,5.684513,6.232616,6.311385,5.8518977,5.7632823,5.83877,5.8453336,5.651693,5.2381544,5.3037953,5.1987696,4.6802053,4.07959,4.3027697,4.640821,4.8771286,5.720616,6.8988724,7.13518,6.961231,6.0028725,5.2053337,5.0871797,5.7468724,6.5312824,7.1680007,7.2369237,6.629744,5.5729237,5.4908724,5.435077,5.7764106,6.5969234,7.6964107,7.6734366,7.4207187,7.020308,6.557539,6.124308,5.4974365,5.4153852,5.3924108,5.428513,6.0061545,6.432821,5.930667,5.408821,5.034667,4.2502565,4.640821,4.2929235,3.9548721,3.6824617,2.8356924,3.4198978,3.754667,4.1222568,4.578462,4.955898,5.0149746,3.7874875,2.1169233,0.77456415,0.45620516,0.36758977,0.3314872,1.0010257,1.9987694,1.9200002,1.5097437,1.1815386,1.1060513,1.4703591,2.4910772,4.9329233,5.5007186,5.3858466,4.5029745,1.4998976,5.1954875,6.626462,7.13518,7.433847,7.5946674,4.010667,2.8422565,2.793026,2.9407182,2.7273848,3.882667,2.5435898,1.0732309,0.56123084,0.7975385,0.6071795,0.40369233,0.34133336,0.36102566,0.19692309,0.21333335,0.13128206,0.098461546,0.14769232,0.17066668,0.16738462,0.18707694,0.30851284,0.51856416,0.7056411,0.76800007,0.7778462,0.77456415,1.3226668,3.4921029,4.4077954,5.723898,5.805949,6.3212314,12.265027,17.115898,15.520822,13.666463,14.506668,17.782156,14.624822,12.133744,12.740924,14.736411,12.25518,9.783795,10.55836,10.857026,9.645949,8.562873,9.353847,9.77395,10.125129,10.322052,9.888822,11.602052,11.881026,11.641437,11.050668,9.524513,8.822155,8.618668,8.103385,7.4469748,7.8080006,8.04759,8.858257,9.734565,10.811078,12.86236,12.507898,10.948924,9.147078,7.515898,5.920821,4.4964104,3.6857438,3.9089234,5.228308,7.3353853,6.6034875,7.0498466,8.513641,10.30236,11.204924,5.080616,2.678154,2.0217438,1.8281027,1.5327181,1.8773335,1.1716924,0.8205129,1.1881026,1.6049232,1.8379488,0.9911796,3.8596926,9.301334,10.249847,6.7314878,5.799385,5.976616,5.658257,3.1376412,4.0008206,3.006359,2.409026,2.5829747,2.0151796,1.3522053,1.3587693,1.9659488,3.0949745,4.6539493,8.690872,10.423796,9.875693,8.192,7.637334,4.2436924,2.6157951,2.2580514,3.0916924,5.4547696,7.030154,7.6734366,7.174565,5.3202057,1.8937438,3.2361028,6.157129,7.181129,6.4065647,7.515898,4.6276927,11.021129,17.762463,19.052309,12.248616,4.5817437,4.266667,7.574975,10.948924,10.971898,9.747693,9.035488,7.860513,7.066257,9.31118,10.505847,14.5263605,15.353437,12.274873,9.895386,12.645744,9.380103,6.5083084,6.8627696,9.711591,5.142975,3.2787695,4.020513,6.1407185,7.282872,6.12759,6.2490263,7.4108725,8.907488,9.563898,4.44718,2.6420515,3.3772311,5.2480006,6.2129235,6.1407185,4.827898,3.0654361,2.3138463,4.716308,6.3474874,5.175795,4.1714873,4.132103,3.6660516,3.370667,4.1222568,6.0192823,7.6668725,6.160411,6.616616,7.3058467,8.211693,8.851693,8.293744,7.6077952,6.701949,6.189949,6.377026,7.256616,4.2929235,3.8531284,5.034667,5.799385,2.9833848,3.8334363,6.2752824,6.9645133,5.98318,6.8299494,11.392001,14.916924,12.511181,7.207385,9.961026,17.08636,19.364103,17.06995,12.652308,10.7158985,8.65477,7.722667,11.434668,16.216616,11.405129,7.7456417,5.225026,3.5610259,4.5554876,12.081232,8.802463,5.6385646,4.9788723,6.892308,9.120821,5.7534366,6.157129,8.789334,9.770667,2.8849232,8.3364105,11.241027,19.295181,27.85477,19.974566,14.04718,10.994873,9.577026,9.337437,10.614155,7.256616,6.36718,7.512616,8.864821,7.177847,8.556309,8.356103,8.6580515,9.278359,7.785026,7.680001,7.860513,8.103385,8.661334,10.230155,10.089026,10.985026,11.218052,11.178667,13.344822,13.098668,12.819694,12.685129,11.926975,8.845129,14.480412,13.124924,12.425847,17.46708,30.772514,32.95508,35.150772,30.690464,23.414156,27.67426,31.251696,32.912415,33.38831,33.00759,31.684925,31.960617,32.518566,31.481438,29.06913,27.6119,26.791388,28.92472,31.130259,32.295387,33.06339,33.237335,31.382977,30.280207,30.775797,31.796515,30.007797,29.18072,28.71795,28.278156,27.769438,30.680618,31.471592,30.782362,29.607388,29.298874,30.546053,32.17067,32.47262,31.40595,30.569029,30.995695,31.012104,30.772514,30.148926,28.73108,29.239798,29.321848,28.800003,27.736618,26.456617,25.27508,24.612104,24.49395,24.070566,21.5959,20.821335,20.97231,21.353027,21.635284,21.865026,20.775387,19.62995,19.177027,20.023796,22.626463,22.144001,21.418669,21.054361,21.14954,21.287386,22.327797,23.003899,23.013746,22.426258,21.671387,20.489847,20.384823,21.435078,23.220514,24.805746,24.805746,25.061745,24.864822,24.392206,24.6679,25.46872,25.938053,26.210464,26.712618,28.182976,27.093336,26.59118,25.353848,23.430567,22.242464,21.861746,20.50954,19.219694,18.474669,18.208822,17.75918,17.893745,17.637745,17.184822,17.900309,17.61477,18.202257,18.786463,19.301744,20.470156,19.849848,18.011898,16.160822,14.78236,13.650052,13.840411,13.74195,13.755078,13.889642,13.771488,0.18379489,0.19692309,0.20676924,0.22646156,0.24287182,0.24287182,0.256,0.25928208,0.28225642,0.31507695,0.28882053,0.27897438,0.32164106,0.3708718,0.39384618,0.380718,0.41682056,0.43651286,0.42338464,0.38400003,0.33476925,0.4201026,0.46933338,0.47589746,0.46276927,0.48902568,0.9156924,0.93866676,0.9353847,1.0436924,1.1913847,1.3357949,1.5097437,1.8642052,2.4713848,3.3280003,3.6562054,2.986667,2.8488207,3.564308,4.273231,5.35959,6.4000006,7.138462,7.706257,8.621949,8.388924,7.955693,7.0892315,5.8486156,4.578462,4.3716927,5.077334,5.4514875,5.037949,4.197744,4.818052,4.9362054,5.280821,5.9470773,6.422975,6.1078978,6.2916927,6.6822567,7.0859494,7.4141545,6.2916927,6.6625648,7.174565,7.24677,7.066257,7.821129,7.515898,7.4863596,8.152616,9.019077,9.6525135,10.377847,10.725744,10.463181,9.596719,9.586872,9.609847,9.787078,9.83959,9.094564,9.094564,9.432616,9.517949,9.255385,9.048616,9.488411,10.026668,10.374565,10.594462,11.109744,10.66995,9.688616,8.864821,8.677744,9.399796,9.593436,8.976411,8.155898,7.7325134,8.27077,8.379078,8.598975,8.576,8.116513,7.200821,7.128616,6.99077,6.8332314,6.619898,6.23918,6.1308722,5.8190775,5.924103,6.49518,7.020308,7.5552826,7.837539,7.9228725,8.306872,9.91836,10.94236,10.459898,9.744411,9.324308,8.956718,11.605334,15.061335,18.392616,20.94277,22.324514,20.066463,17.634462,15.852309,15.346873,16.554668,18.898052,18.287592,17.417847,17.191385,16.679386,14.834873,16.233027,18.235079,19.085129,17.913437,15.763694,16.738462,17.506462,17.115898,16.984617,15.261539,15.445334,15.333745,14.102976,12.2847185,11.08677,10.240001,9.622975,9.147078,8.743385,8.999385,9.025641,8.818872,8.339693,7.522462,6.6428723,6.2490263,5.976616,5.648411,5.293949,4.6834874,4.6145644,4.9427695,5.21518,4.6539493,5.179077,4.9985647,4.594872,4.450462,5.034667,5.609026,5.8814363,6.0225644,6.180103,6.485334,6.889026,7.0334363,6.9349747,6.882462,7.430565,7.273026,7.0859494,6.9776416,7.0400004,7.3714876,6.8693337,6.498462,6.3868723,6.4000006,6.117744,5.717334,5.0477953,4.857436,5.218462,5.5236926,5.280821,5.1364107,4.850872,4.273231,3.3575387,4.381539,4.821334,5.3234878,5.937231,6.1341543,6.0717955,5.6352825,5.668103,6.1440005,6.180103,5.717334,5.21518,4.453744,3.9122055,4.7917953,4.8640003,4.6900516,4.768821,5.4875903,7.1122055,7.269744,6.5411286,5.7698464,5.720616,7.066257,6.882462,6.560821,6.114462,5.6943593,5.586052,5.658257,6.2818465,7.1089234,7.7948723,7.965539,7.90318,7.788308,7.000616,6.0750775,6.698667,6.491898,6.669129,6.875898,6.7610264,5.979898,6.2129235,5.940513,5.8880005,5.9470773,5.2020516,4.8607183,4.601436,4.594872,4.4964104,3.4330258,2.9801028,2.7208207,3.0227695,4.0533338,5.799385,4.529231,2.802872,1.5064616,0.8205129,0.19692309,0.44307697,0.35774362,1.0699488,2.284308,2.2744617,1.4933335,1.3784616,1.654154,2.8914874,6.5312824,7.6668725,5.1659493,3.879385,3.879385,0.47261542,6.4656415,8.073847,9.7903595,10.404103,3.006359,4.6178465,3.7185643,2.5238976,2.03159,2.044718,4.010667,2.5435898,0.86974365,0.44307697,0.9321026,1.2603078,0.702359,0.26256412,0.21989745,0.12143591,0.12143591,0.15097436,0.2100513,0.26912823,0.24287182,0.26912823,0.27569234,0.39712822,0.5940513,0.65641034,0.67938465,0.61374366,0.6301539,0.83035904,1.2209232,4.8705645,7.312411,7.5421543,7.2960005,11.030975,16.390566,16.439796,14.358975,12.852514,14.145642,12.022155,11.408411,12.914873,14.746258,12.694975,11.132719,11.585642,12.248616,12.018872,10.466462,9.4916935,9.18318,10.085744,11.303386,10.499283,11.401847,11.874462,11.72677,11.257437,11.244308,10.610872,9.803488,8.618668,7.64718,8.27077,8.648206,9.485129,10.082462,10.640411,12.251899,13.02318,11.30995,9.015796,7.066257,5.431795,4.2240005,3.1803079,3.6135387,5.61559,8.057437,8.54318,8.372514,8.3364105,8.641642,8.910769,5.3825645,4.2896414,3.6791797,2.5074873,0.64000005,1.0436924,0.9714873,0.82379496,0.7253334,0.51856416,2.9472823,1.6771283,2.3926156,5.8945646,8.103385,5.1954875,4.7360005,4.266667,3.1245131,2.4418464,4.6145644,3.0227695,2.8225644,4.9788723,6.2851286,2.9768207,2.425436,3.367385,4.7524104,5.7534366,6.889026,7.13518,6.688821,5.5991797,3.767795,3.5380516,3.9187696,3.5938463,2.6322052,2.487795,3.2820516,4.8082056,5.149539,4.716308,6.23918,4.640821,10.072617,14.332719,14.76595,14.267078,11.008,12.553847,18.372925,22.954668,15.839181,5.0477953,8.326565,14.749539,17.270155,12.740924,9.800206,6.701949,6.373744,9.970873,16.889437,14.55918,17.289848,18.110361,14.483693,8.329846,12.517745,11.277129,9.065026,7.965539,7.6603084,4.5456414,3.5314875,4.1911798,5.609026,6.377026,6.9021544,6.8594875,7.3714876,8.369231,8.576,5.106872,3.0424619,3.2000003,4.893539,5.920821,8.434873,11.270565,8.411898,1.9561027,2.0906668,2.7864618,5.093744,6.813539,6.764308,4.775385,5.0674877,8.592411,7.8014364,3.5478978,5.110154,6.3212314,6.675693,7.020308,6.9645133,4.9132314,5.7665644,6.9710774,6.3179493,4.522667,5.218462,5.586052,7.003898,6.678975,4.4865646,2.9604106,6.76759,5.973334,8.274052,12.921437,10.712616,7.39118,6.99077,7.6635904,8.421744,9.156924,21.986464,24.523489,19.794052,13.50236,14.037334,11.730052,9.324308,10.036513,12.99036,13.197129,7.5454364,3.0129232,1.4375386,2.097231,1.6935385,3.1113849,2.1825643,1.8970258,2.4648206,1.3423591,1.7460514,2.9538465,3.4921029,2.7634873,1.0535386,2.9702566,6.186667,10.427077,15.05477,19.058874,19.11795,20.726156,16.338053,8.625232,10.466462,8.136206,6.931693,6.8562055,7.568411,8.362667,9.107693,8.723693,8.516924,8.198565,5.904411,6.698667,7.2631803,7.4896417,7.6668725,8.484103,8.569437,9.242257,9.626257,10.026668,11.9171295,11.611898,12.461949,11.904001,10.932513,14.066873,19.695591,15.885129,10.525539,13.13477,34.852104,34.14318,29.06913,27.421541,29.344822,27.342772,28.393028,29.469542,30.923489,31.98031,30.74626,27.720207,27.474054,27.122873,25.96431,25.511387,28.49149,31.113848,31.619284,30.585438,30.913643,31.878567,32.531696,32.774567,32.50544,31.599592,28.721233,28.074669,28.032001,27.815386,27.510157,28.160002,29.144617,29.11508,27.762875,25.833027,28.983797,32.708927,33.00759,29.715694,26.505848,27.06708,26.98831,26.377848,25.619694,25.376822,25.816618,25.85272,25.54749,25.15036,25.10113,24.612104,23.345232,22.25231,21.362873,19.77436,19.872822,20.401232,21.664822,23.072823,23.14831,20.926361,19.656206,19.636515,20.52595,21.333336,21.30708,21.428514,21.129848,20.457027,20.066463,21.858463,21.704206,21.48431,21.658258,21.254566,21.07077,20.762259,21.769848,24.881233,30.227695,30.326157,28.353643,26.308926,25.4359,26.230156,29.256207,30.050465,29.988106,30.306463,32.08862,33.188107,29.423592,24.74995,21.471182,20.263386,21.205336,20.020514,18.376207,17.09949,16.160822,16.390566,16.30195,16.246155,16.633438,17.913437,17.266872,16.728617,16.925539,18.23836,20.81149,19.666052,17.152,14.772514,13.272616,12.649027,12.918155,13.167591,13.157744,13.138052,13.869949,0.15753847,0.20020515,0.24287182,0.27569234,0.29538465,0.3052308,0.27897438,0.24287182,0.23630771,0.26256412,0.27897438,0.2855385,0.34789747,0.38728207,0.4004103,0.4660513,0.512,0.48902568,0.44964105,0.42994875,0.45620516,0.571077,0.56123084,0.636718,0.78769237,0.7811283,1.1290257,1.024,1.0305642,1.270154,1.4473847,1.270154,1.1224617,1.4703591,2.2580514,2.8882053,3.4789746,3.6332312,3.9023592,4.5128207,5.346462,6.1308722,6.114462,6.436103,7.4174366,8.546462,8.579283,8.188719,6.997334,5.651693,5.8486156,5.4547696,5.3891287,5.5565133,5.6943593,5.3792825,5.0149746,4.955898,5.4186673,6.4689236,7.9983597,8.736821,8.841846,8.812308,8.960001,9.40636,7.6964107,6.7544622,6.9054365,7.5881033,7.3583593,7.9786673,8.41518,8.789334,9.019077,8.809027,8.418462,8.326565,8.697436,9.347282,9.731283,9.865847,10.023385,9.872411,9.3078985,8.434873,9.088,9.744411,10.039796,10.036513,10.220308,10.738873,11.575796,12.314258,12.721231,12.757335,11.818667,10.935796,10.55836,10.7158985,10.985026,10.929232,10.568206,9.915077,9.212719,8.930462,8.815591,9.02236,9.301334,9.258667,8.372514,7.450257,7.197539,6.8660517,6.4656415,6.741334,6.885744,6.498462,6.114462,6.0061545,6.189949,6.705231,7.4797955,8.034462,8.39877,9.101129,9.793642,10.683078,11.119591,11.001437,10.752001,11.428103,13.538463,16.370872,19.012924,20.38154,19.275488,17.073233,16.091898,16.745028,17.532719,18.645334,19.534771,19.879387,19.347694,17.591797,15.182771,16.059078,17.401438,17.828104,17.38831,15.993437,16.853334,17.296412,17.030565,18.166155,19.77436,19.24595,17.64759,15.684924,13.699283,12.025436,11.152411,10.525539,10.253129,11.109744,10.643693,9.760821,8.999385,8.320001,7.069539,7.4699492,7.3682055,6.7807183,5.910975,5.149539,5.0543594,5.3431797,5.622154,5.6418467,5.277539,5.412103,5.0084105,4.70318,4.7950773,5.2545643,5.730462,5.904411,6.0356927,6.193231,6.265436,6.550975,6.8660517,6.6592827,6.235898,6.73477,7.6701546,8.205129,7.9195905,7.2270775,7.3714876,7.181129,6.73477,6.7085133,6.99077,6.678975,6.9809237,6.304821,5.8518977,5.9963083,6.2818465,6.0849237,5.910975,5.661539,5.2644105,4.650667,4.2207184,4.2962055,4.8771286,5.6976414,6.242462,6.3179493,5.756718,5.21518,4.8311796,4.201026,4.7261543,4.6539493,4.3552823,4.2994876,5.07077,4.9394875,4.7228723,5.172513,6.422975,7.9885135,8.080411,6.820103,5.7403083,5.61559,6.491898,6.4065647,6.6067696,6.8955903,6.931693,6.2555904,6.1440005,6.8529234,7.466667,7.8736415,8.759795,8.63836,8.03118,7.243488,6.764308,7.259898,5.979898,5.8289237,6.232616,6.514872,5.920821,6.2194877,6.75118,6.7971287,6.308103,5.8880005,5.4383593,5.2545643,4.8377438,3.9712822,2.7142565,2.6617439,2.4352822,4.0041027,6.265436,5.041231,3.5478978,1.8740515,0.92225647,0.69907695,0.32164106,0.34133336,0.79097444,1.7591796,2.6223593,2.0545642,1.6049232,1.7952822,2.3926156,4.066462,8.39877,6.770872,5.579488,4.1846156,2.7864618,2.4385643,4.312616,4.8016415,5.477744,5.7665644,2.9702566,4.8738465,3.56759,2.5862565,2.789744,2.3630772,3.2131286,2.2514873,1.1027694,0.571077,0.6498462,0.88287187,0.48246157,0.15097436,0.101743594,0.072205134,0.09189744,0.14112821,0.190359,0.23302566,0.256,0.23302566,0.256,0.3446154,0.42994875,0.36430773,0.33805132,0.48574364,0.76800007,1.8281027,4.9920006,8.52677,9.304616,9.911796,10.906258,10.824206,15.159796,15.655386,13.988104,11.861334,11.008,10.125129,13.019898,11.995898,7.207385,6.688821,10.692924,14.053744,14.8939495,13.371078,11.664412,10.988309,10.118565,10.295795,11.053949,10.230155,10.57477,10.765129,10.870154,10.981745,11.185231,10.597744,10.226872,9.432616,8.470975,8.477539,8.953437,9.081436,9.593436,10.607591,11.641437,12.245335,10.9915905,9.035488,6.925129,4.565334,3.170462,2.740513,3.1245131,4.076308,5.2381544,6.0685134,7.9524107,9.6295395,10.299078,9.632821,7.059693,5.796103,4.699898,3.0523078,0.58092314,0.65969235,0.81394875,0.88615394,0.8369231,0.7253334,2.3729234,2.1398976,1.975795,2.4910772,2.9636924,4.785231,6.048821,4.8836927,2.4582565,2.9669745,5.684513,4.2469745,3.5610259,4.9788723,6.2752824,4.263385,3.436308,3.31159,3.2196925,2.28759,2.4057438,3.1540515,3.7776413,3.6726158,2.3893335,2.4320002,3.6857438,5.097026,5.5236926,3.757949,4.394667,5.169231,4.788513,4.266667,6.925129,6.0980515,9.465437,13.111795,16.393847,21.956924,22.613335,14.690463,11.575796,14.651078,13.275898,7.6996927,9.074872,12.025436,12.412719,7.3583593,8.303591,8.621949,12.248616,18.5239,22.212925,19.626669,21.402258,28.393028,33.552414,21.940514,12.202667,8.89436,8.448001,9.475283,12.773745,7.6110773,6.629744,5.986462,4.965744,5.986462,6.189949,6.294975,6.5247183,6.7150774,6.3179493,4.9099493,5.0149746,4.9394875,4.197744,3.515077,4.2929235,4.7950773,3.9811285,3.0391798,5.398975,4.46359,4.9854364,4.969026,4.194462,4.2272825,10.758565,11.611898,8.372514,4.4734364,5.1987696,6.4065647,6.1341543,6.695385,7.5520005,5.3169236,5.2709746,6.6395903,6.7807183,5.47118,4.8771286,3.436308,3.6069746,3.764513,3.751385,4.850872,6.872616,4.890257,15.9573345,30.834875,14.007796,11.625027,11.355898,11.818667,10.154668,2.0512822,4.775385,5.8912826,6.370462,6.75118,7.141744,4.5423594,4.1124105,4.2994876,4.4340515,4.7392826,3.2689233,3.4822567,4.1452312,4.4734364,4.1485133,4.2338467,5.3924108,6.2129235,5.674667,3.1376412,4.3027697,7.2237954,7.3025646,4.1813335,1.7591796,1.8018463,2.930872,5.6943593,10.312206,16.689232,18.917746,23.535591,24.58913,18.86195,5.901129,7.7981544,7.240206,6.36718,6.0324106,5.8092313,6.4590774,7.3550773,7.581539,6.744616,4.9788723,5.2644105,5.943795,6.2752824,6.47877,7.7259493,7.5881033,8.677744,9.347282,9.386667,10.049642,11.004719,11.940104,10.81436,11.142565,22.016,24.402054,20.224,15.182771,13.167591,16.262566,12.868924,20.86072,27.073643,28.832823,33.95939,31.894978,28.911592,28.274874,29.72554,29.489233,27.858053,26.154669,25.032207,24.579285,24.290462,28.100925,29.18072,28.563694,27.703796,28.471798,28.245335,29.08554,30.450874,31.481438,30.979284,28.681849,26.916105,25.924925,25.426054,24.595694,26.12185,27.362463,27.214771,25.62954,23.611078,27.024412,29.095387,28.944412,27.48718,27.431387,26.646976,25.951181,25.380104,24.71713,23.496206,23.584822,24.441439,24.979694,25.08472,25.600002,25.609848,24.484104,23.630772,23.102362,21.592617,22.09149,22.04554,21.91754,21.704206,20.93949,21.14954,20.594873,20.719591,21.635284,22.150566,21.979898,22.672413,22.71836,21.91754,21.372719,21.543386,20.814772,20.65395,21.13313,20.926361,21.612309,21.53354,21.320208,22.308104,26.54195,28.376617,28.232206,27.77272,28.104208,29.758362,33.575386,36.98544,39.33867,45.220104,64.436516,60.92472,42.348312,27.460926,22.71836,22.30154,20.762259,18.753643,17.125746,16.196924,15.75713,16.406975,16.636719,16.298668,15.898257,16.584206,16.180513,16.341335,16.531694,16.86318,18.090668,18.661745,17.801847,16.114874,14.14236,12.356924,11.969642,12.117334,12.698257,13.351386,13.4170265,0.18051283,0.21333335,0.23302566,0.27241027,0.318359,0.29210258,0.26256412,0.24287182,0.23958977,0.26912823,0.32820517,0.36430773,0.41025645,0.446359,0.47917953,0.54482055,0.5481026,0.5349744,0.61374366,0.7384616,0.73517954,0.7417436,0.80738467,0.92225647,1.0502565,1.148718,1.3095386,1.273436,1.2373334,1.2931283,1.4112822,1.2274873,1.3522053,1.7427694,2.4746668,3.7382567,4.1189747,4.2863593,4.585026,5.346462,6.87918,6.882462,6.3606157,6.413129,7.256616,8.228104,8.470975,7.8703594,7.0400004,6.616616,7.273026,6.8463597,6.3540516,6.3277955,6.5247183,5.933949,5.6287184,5.402257,5.792821,6.994052,8.841846,9.921641,10.010257,9.82318,9.80677,10.151385,8.5891285,7.6767187,7.515898,7.79159,7.788308,8.139488,8.946873,9.662359,9.7673855,8.749949,8.021334,7.7259493,8.234667,9.360411,10.341744,10.184206,9.872411,9.337437,8.736821,8.461129,9.961026,10.955488,11.319796,11.293539,11.457642,11.861334,12.796719,13.423591,13.443283,13.095386,12.583385,11.841642,11.539693,11.684103,11.631591,11.792411,11.575796,11.076924,10.5780525,10.512411,10.423796,10.676514,10.643693,10.154668,9.472001,8.549745,8.254359,7.88677,7.381334,7.27959,7.515898,6.9842057,6.3442054,5.933949,5.799385,6.0258465,6.701949,7.450257,7.9983597,8.172308,8.759795,9.878975,10.9226675,11.631591,12.068104,12.2387705,13.29559,15.038361,16.800821,17.480206,17.10277,16.567797,16.59077,17.237335,17.913437,18.776617,19.666052,19.99754,19.554462,18.471386,15.944206,15.442053,16.15754,17.286566,18.025026,17.703386,17.56554,17.30954,17.368616,18.930874,21.920822,22.50831,20.864002,17.929848,15.435489,14.073437,12.829539,12.3076935,12.42913,12.435693,11.67754,10.092308,8.769642,8.077128,7.643898,7.755488,7.6176414,7.1680007,6.38359,5.277539,5.4514875,6.088206,6.449231,6.2884107,5.861744,5.737026,5.504,5.287385,5.2512827,5.5762057,5.8223596,6.0192823,6.4032826,6.774154,6.485334,6.8233852,6.9349747,6.619898,6.1472826,6.2785645,7.397744,8.4512825,8.303591,7.1548724,6.564103,7.6176414,7.5585647,7.2960005,7.2894363,7.53559,7.6242056,7.0498466,6.47877,6.23918,6.3507695,5.3103595,5.5663595,5.927385,5.8912826,5.661539,4.8836927,4.493129,4.8377438,5.786257,6.7282057,6.567385,6.0324106,5.5269747,5.097026,4.420923,4.2962055,4.4406157,4.3618464,4.1222568,4.31918,4.7655387,4.923077,5.477744,6.5969234,7.936001,8.461129,7.962257,7.181129,6.678975,6.8430777,7.138462,7.39118,7.269744,6.810257,6.422975,6.3179493,7.1023593,7.8736415,8.470975,9.498257,8.907488,7.5979495,6.6822567,6.521436,6.7150774,5.786257,5.6320004,5.7829747,6.0192823,6.370462,7.194257,7.955693,7.565129,6.2818465,5.720616,5.4482055,4.785231,3.9876926,3.1934361,2.422154,2.4648206,2.8882053,4.965744,6.8430777,3.5511796,2.0742567,1.2668719,0.81394875,0.5284103,0.3511795,0.26912823,1.0699488,1.9954873,2.3860514,1.6705642,1.9922053,2.2416413,3.314872,5.3005133,7.4929237,6.045539,6.196513,5.7074876,4.516103,4.7327185,4.096,4.5128207,5.3760004,5.661539,3.948308,4.5128207,4.2174363,4.0303593,3.7448208,1.9561027,2.0020514,1.3522053,0.93866676,0.892718,0.56123084,0.50543594,0.27241027,0.098461546,0.052512825,0.032820515,0.036102567,0.08861539,0.14769232,0.190359,0.20348719,0.20348719,0.2231795,0.27569234,0.39384618,0.65641034,0.6498462,0.6695385,1.3193847,3.249231,7.171283,10.998155,11.264001,11.431385,12.491488,12.970668,14.572309,14.769232,13.51877,11.716924,11.201642,11.339488,13.292309,14.217847,14.011078,15.304206,14.276924,15.570052,15.42236,13.400617,12.393026,11.707078,10.427077,10.049642,10.358154,9.43918,10.473026,10.368001,10.246565,10.486155,10.722463,10.233437,10.016821,9.639385,9.114257,8.887795,8.832001,9.097847,9.846154,10.735591,10.932513,10.601027,8.937026,7.325539,5.9995904,4.0467696,2.540308,2.3827693,2.7273848,3.1573336,3.7087183,4.381539,6.918565,9.048616,9.737847,9.179898,8.87795,7.529026,5.405539,2.9604106,0.81066674,1.4473847,1.1979488,0.81066674,0.8336411,1.6114873,2.484513,2.8389745,2.8455386,2.6518977,2.3729234,5.5597954,6.5411286,4.926359,2.5600002,3.5183592,5.937231,3.9187696,3.3772311,5.8223596,8.369231,5.0116925,3.6102567,4.4406157,5.661539,3.3247182,2.537026,3.692308,3.820308,2.9571285,4.132103,7.568411,11.372309,13.659899,13.026463,8.533334,9.754257,8.812308,7.683283,8.3593855,12.852514,12.041847,11.490462,12.182976,15.891693,25.160208,23.289438,16.764719,11.812103,9.833026,7.433847,10.052924,12.747488,12.983796,11.017847,9.90195,13.35795,14.467283,16.321642,19.74154,23.2599,23.328823,23.384617,28.865643,37.776413,40.6679,28.882053,17.017437,10.299078,9.747693,12.166565,8.228104,6.9054365,6.3343596,5.835488,5.927385,6.1440005,6.36718,6.7183595,7.125334,7.3353853,6.554257,5.7731285,5.0576415,4.640821,4.9362054,6.173539,5.4153852,4.2371287,3.7710772,4.7327185,4.276513,6.173539,6.8463597,5.8190775,5.717334,7.9524107,8.172308,6.4032826,4.3552823,5.412103,6.2096415,5.533539,6.0685134,7.6143594,7.072821,4.9099493,4.9952826,5.333334,5.402257,6.1538467,4.5554876,3.5183592,2.8947694,2.8324106,3.767795,6.73477,4.4307694,12.980514,26.932514,19.242668,12.018872,10.456616,10.312206,8.027898,0.7220513,0.9485129,1.214359,2.2449234,3.692308,4.135385,3.5052311,3.5807183,3.5347695,3.2229745,3.1540515,3.5774362,4.46359,4.7950773,4.8672824,6.298257,4.4438977,4.5489235,4.585026,4.2502565,4.969026,4.7917953,5.218462,4.827898,3.5249233,2.5042052,2.1956925,2.4024618,3.9844105,6.409847,7.785026,11.237744,22.662565,26.194054,18.113642,6.8463597,6.1407185,6.3868723,6.6494365,6.2720003,4.8804107,5.113436,5.8945646,6.235898,5.927385,5.5138464,5.2644105,5.9995904,6.114462,5.7009234,6.557539,6.9710774,8.192,9.242257,9.619693,9.3078985,9.645949,9.90195,9.865847,12.06154,21.730463,26.089027,21.927387,16.452925,13.922462,15.61272,8.267488,20.870565,28.609644,25.974155,26.761848,27.703796,25.124104,24.6679,26.594463,25.777233,25.281643,23.873642,22.3639,21.270975,20.837746,24.884514,26.548515,26.41395,25.544207,25.491693,25.40636,26.630566,27.858053,28.49149,28.642464,26.12185,24.146053,22.692104,21.858463,21.858463,23.620924,24.595694,24.264208,23.030155,22.22277,24.421745,25.439182,25.442463,25.189745,26.026669,24.887796,24.372515,24.415182,24.201847,22.163694,21.973335,22.852924,24.336412,26.144823,28.18954,28.498053,26.5879,24.34954,22.885746,22.514874,23.217232,23.601233,23.161438,21.930668,20.476719,21.523693,21.300514,21.211899,22.01272,23.801437,23.922874,23.995079,23.502771,22.764309,22.92513,21.507284,20.63754,20.709745,21.43836,21.897848,22.14072,22.294975,21.48431,20.634258,22.478771,24.530054,25.984001,27.40513,29.023182,30.729849,34.497643,38.53785,42.912823,56.155903,95.26483,101.031395,73.406364,44.721233,29.748514,25.74113,21.530258,17.906874,16.06236,15.691488,14.979283,15.780104,15.701335,15.172924,14.76595,15.2155905,15.366566,15.488001,15.67836,15.980309,16.403694,16.95836,16.662975,16.02954,14.92677,12.593232,12.133744,12.212514,12.793437,13.4170265,13.233232,0.2231795,0.23302566,0.22646156,0.26256412,0.31507695,0.27569234,0.2986667,0.30194873,0.29538465,0.3052308,0.36758977,0.42994875,0.48246157,0.5152821,0.53825647,0.5874872,0.6432821,0.6170257,0.6498462,0.7515898,0.77128214,0.761436,0.9944616,1.1716924,1.2471796,1.4211283,1.3784616,1.4834872,1.6049232,1.6836925,1.7591796,1.5688206,1.7788719,2.038154,2.5632823,4.1156926,4.7950773,5.0510774,5.5269747,6.491898,7.817847,7.453539,6.820103,6.629744,7.066257,7.788308,7.9885135,7.785026,7.686565,7.90318,8.346257,7.765334,7.2270775,7.00718,6.882462,6.121026,5.72718,5.76,6.3179493,7.509334,9.452309,10.006975,9.91836,9.856001,10.036513,10.236719,9.160206,8.628513,8.3823595,8.329846,8.556309,8.402052,9.107693,9.905231,10.056206,8.87795,8.815591,8.730257,9.176616,10.164514,11.155693,10.794667,10.423796,9.862565,9.291488,9.242257,10.571488,11.204924,11.621744,11.979488,12.11077,12.422565,13.528616,14.214565,14.066873,13.466257,13.121642,12.616206,12.317539,12.248616,12.081232,12.343796,12.130463,11.779283,11.536411,11.546257,11.795693,12.035283,11.766154,11.076924,10.620719,9.944616,9.193027,8.605539,8.178872,7.634052,7.821129,7.4108725,6.931693,6.619898,6.413129,6.314667,6.5739493,7.194257,7.837539,7.817847,8.65477,9.908514,11.172104,12.317539,13.4859495,14.385232,15.123693,15.963899,16.617027,16.242872,16.190361,16.384,16.475899,16.662975,17.67713,18.22195,18.46154,18.599386,18.707693,18.71754,16.981335,15.852309,16.019693,17.552412,19.889233,19.5479,18.307283,17.88718,18.727386,19.984411,22.311386,23.906464,23.424002,20.969027,18.097233,16.20677,15.330462,14.693745,13.850258,12.668719,11.890873,10.722463,9.373539,8.326565,8.329846,8.073847,7.768616,7.5191803,7.0826674,5.83877,6.091488,6.6034875,6.73477,6.373744,5.937231,5.943795,5.8453336,5.6451287,5.4974365,5.691077,6.1440005,6.416411,6.7282057,7.0400004,7.059693,7.141744,7.056411,6.8397956,6.619898,6.6133337,7.5191803,8.549745,8.576,7.702975,7.24677,8.123077,7.936001,7.706257,7.8080006,7.9819493,8.306872,7.9130263,7.3550773,6.8988724,6.5083084,5.431795,5.8125134,6.3967185,6.482052,5.910975,5.277539,5.031385,5.2742567,5.927385,6.7216415,6.6494365,6.052103,5.684513,5.5630774,4.9362054,4.6539493,4.522667,4.201026,3.6857438,3.3050258,4.562052,4.9952826,5.435077,6.180103,6.9809237,7.9885135,8.615385,8.467693,7.762052,7.328821,7.765334,7.8670774,7.456821,6.875898,6.997334,6.803693,7.24677,8.044309,8.982975,9.938052,8.907488,7.8112826,7.24677,7.1548724,6.810257,6.3376417,6.363898,6.2523084,6.055385,6.5247183,7.5520005,8.011488,7.4043083,6.1341543,5.504,4.7228723,3.826872,3.131077,2.6256413,1.9889232,2.034872,3.8137438,6.0980515,6.741334,2.6551797,1.6410258,1.2668719,0.9156924,0.512,0.5152821,0.34789747,1.211077,1.8970258,1.8576412,1.1749744,2.044718,2.2186668,3.69559,6.47877,8.595693,6.4590774,6.117744,5.8814363,5.799385,7.6570263,6.370462,6.3212314,6.045539,5.0018463,3.5774362,4.076308,4.5554876,4.5554876,3.82359,2.3236926,2.3729234,1.3095386,0.75487185,0.892718,0.45292312,0.32164106,0.18051283,0.07548718,0.026256412,0.016410258,0.013128206,0.055794876,0.10502565,0.13128206,0.13784617,0.15753847,0.20348719,0.256,0.446359,1.0601027,1.1749744,1.3587693,2.681436,5.4186673,9.045334,12.947693,13.6697445,13.512206,13.35795,12.63918,13.269335,12.888617,11.523283,10.594462,12.898462,13.078976,14.171899,15.894976,17.552412,18.051283,15.812924,15.51754,14.956308,13.748514,13.331694,11.969642,10.70277,10.459898,10.683078,9.340718,10.440206,10.338462,10.059488,10.092308,10.417232,10.023385,9.90195,9.547488,9.074872,9.202872,8.835282,9.179898,9.833026,10.341744,10.200616,8.992821,7.269744,6.0619493,5.3858466,4.240411,2.678154,2.2646155,2.3762052,2.6880002,3.1638978,4.0500517,6.4000006,8.306872,8.979693,8.746667,10.59118,9.803488,6.994052,3.4789746,1.2832822,3.0818465,2.4516926,1.2635899,0.82379496,1.8674873,2.1103592,2.7142565,3.6693337,4.1846156,2.6551797,4.6834874,5.0051284,3.8564105,2.861949,5.037949,4.716308,3.7940516,4.3027697,6.121026,6.9776416,3.9351797,3.1737437,4.70318,6.4557953,4.2830772,4.086154,4.44718,4.673641,4.8082056,5.622154,13.164309,19.081848,20.821335,18.17272,13.269335,13.830565,10.7848215,9.334154,11.739899,17.302977,15.61272,12.550565,10.873437,12.757335,19.77436,17.913437,15.914668,12.425847,7.9425645,4.785231,13.029744,14.92677,12.711386,11.083488,17.207796,16.039387,14.87754,15.556924,18.323694,21.802668,24.979694,23.601233,25.600002,35.958157,56.710567,52.2437,33.83795,18.710976,12.786873,10.7158985,7.3747697,5.730462,5.664821,6.038975,4.6867695,5.658257,6.2785645,6.4689236,6.4557953,6.774154,6.3343596,7.1089234,6.5706673,5.1987696,6.482052,6.370462,5.720616,5.1167183,4.923077,5.2644105,4.457026,6.6133337,7.968821,7.755488,8.192,5.0477953,4.269949,4.4865646,5.100308,6.2785645,6.294975,5.586052,5.5630774,6.5772314,7.9163084,5.5663595,4.8082056,4.7261543,5.1298466,6.564103,5.037949,3.9844105,3.05559,2.3466668,2.3893335,5.914257,5.028103,7.8408213,13.781334,13.610668,7.145026,5.8223596,5.5072823,3.9844105,0.97805136,2.5074873,2.8422565,3.3608208,4.3684106,5.093744,5.366154,5.0018463,4.532513,4.1517954,3.7120004,4.5817437,4.713026,4.578462,4.8311796,6.3179493,4.4373336,4.332308,3.9417439,3.508513,5.5597954,5.0904617,4.4110775,4.1485133,4.2601027,4.013949,3.3411283,2.8192823,3.0818465,3.6726158,3.0358977,6.2555904,17.77559,21.612309,15.1466675,9.101129,7.6012316,6.6067696,6.2884107,5.9602056,4.086154,4.4767184,4.9952826,5.097026,5.0215387,5.796103,5.0510774,5.874872,6.189949,5.7534366,6.1538467,6.9152827,7.9819493,8.900924,9.209436,8.448001,8.070564,7.8506675,8.467693,11.296822,18.422155,24.74995,21.444925,15.944206,12.983796,14.5952835,7.8473854,18.707693,26.722464,24.894361,19.669334,23.975386,22.160412,21.730463,23.82113,23.19754,23.09908,22.587078,21.320208,19.790771,19.318155,21.707489,23.919592,24.585848,23.686565,22.554258,22.675694,23.840822,24.513643,24.454565,24.730259,22.688822,22.06195,21.441643,20.519386,20.096,20.588308,20.969027,21.379284,21.710772,21.632002,22.672413,22.675694,22.642874,23.105642,24.119797,23.75549,23.378054,22.79713,21.950361,20.913233,21.786259,22.022566,23.187695,25.455591,27.602053,27.621746,25.974155,24.165745,23.27631,23.955694,23.056412,23.739079,23.748924,22.416412,20.660515,22.403284,22.42954,22.245745,22.767591,24.306873,23.988514,23.32554,22.872618,22.918566,23.48636,21.612309,20.096,20.073027,21.425232,22.744617,22.111181,21.700924,20.634258,19.334566,19.524925,21.11672,22.695387,25.048616,27.812105,29.456413,32.134567,35.085133,39.66031,53.19549,89.00267,98.18585,77.46954,49.926567,30.408207,25.577028,22.317951,18.31713,15.90154,15.232001,14.293334,15.254975,14.834873,14.165335,13.791181,13.679591,14.490257,15.028514,15.340309,15.520822,15.721026,15.858873,15.435489,15.133539,14.844719,13.676309,12.882052,12.445539,12.576821,13.111795,13.5318985,0.26256412,0.24615386,0.24287182,0.26256412,0.29210258,0.28225642,0.35774362,0.36430773,0.36102566,0.3708718,0.4004103,0.48246157,0.5513847,0.58420515,0.5874872,0.61374366,0.7515898,0.65969235,0.5284103,0.48574364,0.5973334,0.702359,1.0568206,1.2931283,1.3587693,1.4933335,1.3784616,1.5721027,1.9068719,2.2121027,2.3269746,2.1267693,2.3040001,2.537026,2.92759,4.010667,5.3169236,5.943795,6.73477,7.6668725,7.821129,7.5487185,7.0892315,6.8594875,7.0137444,7.433847,7.515898,8.060719,8.5891285,8.854975,8.851693,8.260923,7.7718983,7.2894363,6.7872825,6.3212314,5.474462,6.1013336,7.0400004,8.077128,9.938052,9.842873,9.498257,9.6065645,10.095591,10.144821,9.537642,9.314463,9.255385,9.3078985,9.593436,8.832001,9.051898,9.639385,9.970873,9.416205,10.427077,10.778257,10.9456415,11.237744,11.805539,11.467488,11.588924,11.401847,10.817642,10.423796,10.706052,10.689642,11.172104,12.041847,12.291283,12.507898,13.705847,14.644514,14.7790785,14.257232,13.764924,13.482668,13.210258,12.908309,12.724514,12.822975,12.62277,12.507898,12.47836,12.156719,12.662155,12.642463,12.35036,12.035283,11.959796,11.428103,10.029949,9.045334,8.644924,7.893334,7.9491286,7.972103,7.968821,7.962257,7.975385,7.6701546,7.463385,7.7325134,8.310155,8.493949,9.6754875,11.07036,12.048411,12.747488,14.076719,16.17395,17.234053,17.713232,17.752617,17.171694,17.266872,17.220924,16.784412,16.515284,17.762463,17.7559,17.365335,17.365335,17.946259,18.710976,18.297438,17.792002,17.463797,18.12677,21.14954,20.427488,19.134361,19.15077,20.470156,21.205336,21.638565,23.177849,24.067284,23.22708,20.25354,17.499899,17.444103,16.613745,14.345847,12.813129,12.137027,12.084514,11.096616,9.38995,8.946873,8.539898,8.139488,8.064001,7.9425645,6.698667,6.8299494,6.8233852,6.5378466,6.0685134,5.7534366,6.009436,5.927385,5.7632823,5.687795,5.802667,6.47877,6.7314878,6.73477,6.882462,7.785026,7.4240007,7.3353853,7.3583593,7.430565,7.581539,8.139488,8.736821,8.930462,8.874667,9.321027,8.740103,8.057437,8.211693,8.786052,8.034462,8.851693,8.73354,8.346257,7.899898,7.128616,6.8233852,6.692103,6.8660517,6.9645133,6.088206,5.467898,5.72718,6.0619493,6.242462,6.62318,6.997334,6.265436,5.7632823,5.674667,5.0543594,5.3234878,4.781949,4.141949,3.626667,2.9768207,4.4274874,4.890257,5.3037953,5.924103,6.3245134,7.351795,8.408616,8.608821,8.050873,7.8145647,8.2215395,7.9786673,7.643898,7.584821,7.9917955,7.6307697,7.5191803,8.109949,9.212719,10.010257,8.953437,8.726975,8.73354,8.549745,7.9327188,7.4929237,7.506052,7.145026,6.442667,6.2916927,7.0531287,7.0925136,6.7314878,6.1374364,5.32677,3.4100516,2.8356924,2.7995899,2.5829747,1.5524104,1.7329233,4.279795,6.314667,6.0849237,2.9768207,2.4549747,1.6705642,0.9911796,0.6432821,0.7056411,0.4594872,1.0896411,1.4605129,1.2242053,0.7975385,1.5655385,1.6475899,3.4494362,7.138462,10.660104,7.318975,5.106872,4.2371287,5.2545643,9.032206,8.841846,8.064001,5.8978467,3.2098465,2.5435898,3.8038976,4.1911798,3.761231,3.1343591,3.4822567,3.5905645,2.156308,0.9878975,0.636718,0.37415388,0.318359,0.17723078,0.055794876,0.0032820515,0.013128206,0.02297436,0.052512825,0.068923086,0.072205134,0.07876924,0.101743594,0.19364104,0.28225642,0.5218462,1.3029745,1.6771283,2.4057438,4.663795,8.257642,11.628308,14.920206,16.357744,15.996719,13.929027,10.282667,11.451077,10.499283,8.822155,8.884514,14.227694,13.74195,14.404924,14.795488,14.096412,12.081232,14.572309,14.582155,14.224411,14.208001,13.843694,11.736616,11.011283,11.270565,11.460924,9.8592825,10.187488,10.371283,10.174359,9.898667,10.374565,10.075898,10.102155,9.501539,8.651488,9.248821,9.160206,9.078155,9.18318,9.403078,9.416205,7.906462,6.688821,5.924103,5.5007186,5.0510774,3.5971284,2.6551797,2.3696413,2.6518977,3.1803079,4.568616,6.5837955,8.214975,8.969847,8.871386,10.952206,10.834052,8.329846,4.535795,1.8084104,4.0303593,3.4198978,1.8838975,0.8467693,1.2504616,1.2406155,1.975795,3.8301542,5.395693,3.4888208,3.2886157,3.3608208,3.114667,3.3608208,6.311385,3.245949,4.0467696,5.431795,5.402257,3.259077,2.9538465,2.9538465,4.017231,5.172513,3.7316926,4.824616,3.8695388,5.21518,7.9097443,5.691077,14.342566,19.554462,19.495386,15.963899,14.381949,13.594257,9.366975,7.6964107,10.47959,15.501129,13.302155,10.282667,8.477539,8.648206,10.249847,10.837335,11.684103,10.902975,8.342975,5.5991797,13.722258,13.092104,9.974154,10.962052,23.000618,15.61272,11.533129,12.655591,16.81395,17.792002,22.682259,21.415386,21.159386,30.273643,58.305645,62.959595,46.628105,29.174156,18.290873,9.475283,6.1341543,4.716308,4.8114877,5.0215387,2.9538465,4.7655387,5.7764106,5.901129,5.5729237,5.7403083,5.0477953,8.598975,8.6580515,5.2578464,6.170257,3.751385,3.9023592,4.8640003,5.83877,6.9645133,5.3924108,6.4623594,7.433847,7.702975,8.802463,4.9788723,3.2065644,4.141949,6.488616,7.000616,6.2063594,5.7468724,5.1659493,5.074052,7.1515903,6.2588725,5.717334,5.1987696,4.962462,5.8518977,4.263385,4.0402055,3.5840003,2.5961027,2.0841026,4.1911798,5.179077,4.312616,2.2482052,1.024,0.73517954,1.1651284,1.3817437,1.2800001,1.5721027,4.1682053,5.0871797,5.5565133,6.245744,7.243488,6.7938466,5.9602056,5.152821,4.4996924,3.8498464,4.6802053,4.378257,4.4996924,5.142975,4.965744,4.5489235,5.5762057,5.7140517,4.775385,4.71959,5.5597954,6.0652313,6.1440005,5.8157954,5.221744,4.516103,3.5347695,2.6322052,2.4713848,4.007385,6.0947695,10.213744,12.793437,12.882052,12.140308,12.297847,8.018052,5.077334,4.644103,3.2820516,4.1550775,4.663795,4.4767184,4.2601027,5.671385,4.7261543,5.2315903,5.8978467,6.235898,6.5739493,7.328821,7.9130263,8.231385,8.067283,7.0990777,6.6527185,6.5050263,6.669129,8.533334,14.87754,20.394669,19.006361,15.944206,13.10195,9.045334,6.49518,11.749744,19.350975,23.502771,18.057848,23.77518,20.713028,18.960411,20.975592,21.56636,21.520412,21.398975,20.680206,19.718565,19.74154,19.75795,21.376001,22.28513,21.72718,20.480001,20.404514,20.821335,20.992002,20.808207,20.791796,19.643078,20.696617,21.5959,21.300514,20.073027,19.072002,18.49436,19.413334,21.00513,20.5719,21.582771,21.353027,21.215181,21.763283,22.836515,23.794874,23.18113,21.041233,18.894772,19.734976,22.04554,21.737028,21.80595,23.030155,23.94913,23.657028,23.332104,23.502771,24.237951,25.163488,22.216208,22.928411,23.40431,22.321232,20.923079,23.588104,23.781746,23.568413,23.620924,23.200823,21.96349,20.929642,21.26113,22.596926,23.043283,21.786259,19.590565,19.275488,21.047796,22.521437,21.336617,20.000822,18.838976,18.103796,17.952822,18.904617,19.324718,21.27754,24.480822,26.312206,27.11631,28.186258,31.015387,37.53026,50.113644,53.17908,49.250465,37.346466,23.716105,21.819078,22.134155,19.331284,16.66954,15.261539,14.070155,14.7561035,14.198155,13.689437,13.446565,12.603078,13.604104,14.887385,15.471591,15.376411,15.596309,15.461744,14.815181,14.224411,14.096412,14.680616,13.46954,12.504617,12.278154,12.924719,14.221129,0.27569234,0.23958977,0.27569234,0.28225642,0.256,0.3052308,0.29210258,0.27241027,0.3446154,0.48574364,0.5349744,0.6071795,0.6071795,0.6695385,0.761436,0.6859488,0.6498462,0.48574364,0.43651286,0.5481026,0.67282057,0.8533334,1.0666667,1.2537436,1.3587693,1.2964103,1.4572309,1.5491283,1.654154,1.8281027,2.1202054,2.1956925,3.1638978,4.2502565,4.97559,5.156103,6.0849237,6.885744,7.574975,7.8834877,7.24677,6.7610264,6.692103,7.0892315,7.5913854,7.4469748,7.896616,8.185436,8.582564,8.976411,8.864821,9.219283,8.228104,7.282872,6.954667,7.003898,6.1374364,7.0826674,8.146052,8.861539,10.010257,10.804514,10.505847,10.305642,10.450052,10.253129,9.764103,9.938052,10.246565,10.450052,10.55836,9.485129,9.068309,9.314463,10.016821,10.771693,11.772718,12.58995,12.544001,11.890873,11.841642,11.474052,11.933539,12.1698475,11.828514,11.23118,11.07036,11.664412,12.1698475,12.416001,12.87877,12.731078,13.37436,14.135796,14.660924,14.8939495,15.015386,14.697027,14.326155,14.007796,13.581129,13.581129,13.699283,14.096412,14.477129,14.099693,13.892924,13.108514,12.58995,12.763899,13.656616,13.046155,11.776001,10.538668,9.527796,8.454565,8.4053335,8.933744,9.31118,9.426052,9.780514,9.475283,9.051898,8.979693,9.458873,10.420513,11.398565,12.091078,11.877745,11.172104,11.428103,13.856822,15.271386,15.862155,16.489027,18.661745,19.137642,20.181335,20.450462,19.958155,20.079592,20.007385,19.505232,18.84554,18.635489,19.820309,20.004105,20.791796,19.925335,17.926565,18.097233,19.511797,20.755693,21.011694,20.729437,21.622156,20.657232,21.12,21.83549,21.451488,18.448412,17.129026,16.708925,16.183796,15.376411,14.936617,14.339283,14.36554,13.282462,11.204924,10.069334,8.812308,8.618668,8.881231,8.809027,7.430565,7.1614366,6.8562055,6.6428723,6.5083084,6.301539,6.117744,6.193231,6.3212314,6.436103,6.6067696,6.1308722,6.0291286,6.2687182,6.954667,8.346257,8.054154,8.172308,8.2215395,8.14277,8.300308,8.411898,8.786052,9.284924,9.80677,10.28595,9.626257,9.350565,9.813334,10.184206,8.438154,8.231385,8.572719,8.546462,8.129642,8.178872,7.77518,6.5870776,6.1407185,6.8562055,8.041026,6.6494365,6.5870776,6.892308,7.269744,8.086975,8.635077,7.9950776,6.816821,5.723898,5.3103595,5.139693,5.0215387,4.9920006,4.906667,4.457026,4.332308,4.8344617,5.8518977,7.141744,8.300308,8.372514,7.9425645,7.2369237,7.059693,8.805744,9.708308,8.661334,7.9819493,8.297027,8.530052,8.237949,8.172308,8.605539,9.363693,9.826463,9.472001,9.147078,8.809027,8.651488,9.078155,8.54318,7.748924,6.7774363,6.048821,6.3179493,6.7938466,7.1122055,7.1680007,6.5444107,4.532513,1.9922053,2.0808206,2.9735386,3.2623591,1.9692309,2.6157951,2.6945643,3.2262566,4.1747694,4.457026,3.4067695,1.8051283,0.8533334,0.7056411,0.47261542,0.27897438,0.44964105,0.5513847,0.57764107,0.9321026,0.77128214,0.8795898,3.1442053,6.4722056,6.7905645,6.242462,3.5872824,2.4155898,3.3805132,4.210872,6.373744,6.3179493,5.1987696,4.2174363,4.6080003,3.6332312,3.4527183,3.190154,2.9801028,3.9811285,2.1891284,2.5173335,2.1497438,0.79097444,0.65641034,0.26584616,0.08533334,0.01969231,0.0,0.0,0.013128206,0.032820515,0.04594872,0.04266667,0.029538464,0.09189744,0.17066668,0.26912823,0.54482055,1.3259488,2.1202054,3.3345644,6.4656415,11.250873,15.671796,17.329231,18.550156,17.158566,13.735386,11.611898,10.866873,9.481847,8.467693,9.173334,13.275898,12.701539,9.517949,10.161232,13.764924,12.1928215,15.169642,14.762668,13.551591,12.708103,11.963078,10.620719,10.896411,10.850462,10.056206,9.6295395,9.800206,10.197334,10.118565,9.764103,10.253129,10.118565,10.331899,9.875693,8.94359,8.956718,9.6295395,8.661334,8.185436,8.576,8.454565,7.39118,6.485334,6.0947695,6.1013336,5.904411,4.9887185,3.945026,3.3247182,3.2032824,3.2032824,4.388103,6.7183595,8.694155,9.590155,9.4457445,7.686565,6.7249236,5.98318,4.7261543,2.0906668,1.5786668,1.467077,1.2603078,0.8598975,0.58092314,1.020718,2.1070771,3.4166157,5.100308,7.9195905,6.47877,6.6592827,6.1078978,4.588308,3.9680004,4.601436,3.2689233,2.9144619,4.125539,5.1265645,7.213949,4.384821,4.2502565,6.6002054,3.4034874,3.4888208,3.1540515,5.3431797,8.267488,5.3858466,7.131898,6.1505647,3.9844105,3.370667,8.241231,8.507077,6.0685134,3.1606157,1.975795,4.6244106,4.965744,3.56759,4.269949,7.3714876,9.6295395,5.868308,6.045539,8.854975,10.348309,3.95159,5.405539,6.6395903,7.2237954,9.366975,17.900309,19.534771,17.168411,16.059078,15.606155,9.370257,13.312001,15.176207,14.601848,16.239592,29.741951,32.695797,31.721027,28.599796,21.64513,5.691077,5.677949,5.6943593,5.0051284,3.882667,3.6004105,4.650667,5.169231,6.75118,9.353847,11.306667,7.9983597,7.6110773,6.672411,4.6080003,3.754667,3.764513,3.767795,4.023795,4.450462,4.6080003,5.6320004,8.077128,7.906462,4.955898,2.930872,5.211898,5.5729237,5.799385,6.170257,5.4613338,4.4734364,4.2371287,4.457026,4.9526157,5.661539,4.135385,4.240411,4.4767184,4.6802053,6.012718,4.900103,4.5423594,4.1813335,3.5610259,2.9144619,1.585231,1.4244103,1.467077,1.5130258,2.1366155,1.7099489,2.353231,3.5413337,4.4996924,4.194462,3.367385,4.201026,4.5554876,4.2272825,4.95918,4.384821,4.3618464,4.348718,4.007385,3.190154,4.568616,5.0051284,5.3825645,5.805949,5.5991797,4.7327185,5.277539,5.8190775,5.3694363,3.3411283,5.0510774,5.2315903,4.4996924,3.5741541,3.2820516,5.074052,5.0477953,4.132103,3.2131286,3.1277952,4.824616,2.9801028,3.1638978,8.392206,19.134361,16.019693,8.625232,4.023795,3.7185643,3.6463592,3.9647183,4.2436924,4.391385,4.841026,6.560821,6.1341543,4.9821544,4.8672824,5.937231,6.744616,7.830975,7.525744,7.4765134,7.5388722,5.7665644,5.6320004,5.792821,5.169231,5.5269747,11.460924,13.059283,14.611693,19.446156,22.229336,8.973129,6.482052,5.172513,7.706257,13.505642,18.753643,25.078156,18.107079,13.725539,15.95077,16.951796,17.844515,16.564514,15.783386,16.482462,17.959387,18.533745,18.38277,18.517334,19.272207,20.309336,19.98113,19.10154,18.904617,19.48554,19.790771,17.851078,17.811693,18.901335,20.575182,22.550976,23.24677,21.060925,18.960411,17.851078,16.554668,19.265642,21.62872,22.360617,21.93395,22.567387,24.14277,23.05313,20.850874,19.03918,19.088411,19.990976,20.62113,21.146257,21.766565,22.705233,23.634052,23.745644,23.440413,23.122053,23.207386,22.098053,23.430567,23.23036,21.300514,21.241438,24.31672,24.287182,23.552002,22.895592,21.513847,20.562054,19.410053,20.14195,22.288412,22.81354,21.993027,21.028105,20.932924,21.385847,20.752413,20.007385,19.042463,17.857643,16.853334,16.83036,17.08636,16.712206,17.394873,19.43959,21.760002,20.598156,20.594873,20.886976,21.461334,23.135181,22.938257,23.328823,22.150566,19.856411,19.50195,20.184616,18.806156,17.716515,17.010874,14.555899,13.361232,12.777026,13.285745,14.14236,13.397334,13.128206,14.040616,14.998976,15.402668,15.182771,14.644514,14.49354,14.273643,13.863386,13.472821,12.924719,12.777026,13.210258,14.073437,14.8939495,0.3117949,0.33476925,0.318359,0.28225642,0.25271797,0.28225642,0.37743592,0.48246157,0.571077,0.60389745,0.5349744,0.6662565,0.67938465,0.84348726,1.0732309,0.9321026,0.6498462,0.67938465,0.8598975,1.017436,0.96492314,0.9714873,1.1979488,1.4342566,1.5360001,1.4080001,1.3522053,1.4506668,1.7001027,2.1267693,2.7798977,3.242667,3.6004105,4.2240005,5.146257,6.0717955,7.213949,7.4830775,8.090257,8.900924,8.43159,7.972103,7.4732313,7.5388722,8.15918,8.717129,8.982975,8.812308,8.392206,7.9195905,7.584821,8.093539,7.39118,6.806975,6.6494365,6.2096415,6.994052,8.395488,9.429334,10.177642,11.805539,11.815386,11.355898,11.23118,11.575796,11.841642,11.900719,11.664412,11.503591,11.441232,11.168821,10.358154,9.747693,9.570462,9.826463,10.272821,11.332924,11.71036,11.904001,11.995898,11.644719,11.464206,11.369026,11.405129,11.395283,10.912822,11.516719,11.874462,12.288001,12.829539,13.341539,13.791181,14.375385,15.041642,15.573335,15.599591,15.809642,15.537232,14.880821,14.299898,14.605129,14.536206,14.148924,13.824001,13.755078,13.952001,13.587693,12.983796,12.724514,13.088821,14.04718,13.653335,12.517745,11.408411,10.689642,10.308924,10.630565,10.696206,10.423796,10.003693,9.878975,9.593436,9.291488,9.212719,9.609847,10.752001,12.294565,12.859077,12.337232,11.490462,11.940104,13.344822,14.529642,15.104001,15.898257,18.980104,20.089437,20.07631,19.396925,18.569847,18.162872,18.38277,18.399181,18.576412,19.34113,21.188925,20.073027,19.423182,18.241642,17.122463,18.231796,20.096,20.791796,21.06749,20.73272,18.65518,20.384823,20.680206,21.044514,21.274258,19.472412,18.937437,17.552412,16.12472,14.890668,13.522053,13.216822,14.319591,13.745232,11.651283,11.424822,10.079181,9.481847,9.7214365,10.180923,9.554052,8.369231,7.50277,7.059693,6.872616,6.5083084,6.6002054,6.5378466,6.3376417,6.1472826,6.229334,5.8781543,5.904411,6.193231,6.8299494,8.113232,8.612103,8.592411,8.100103,7.748924,8.726975,8.868103,9.396514,9.869129,10.184206,10.601027,10.371283,10.213744,10.325335,10.253129,8.891078,7.5881033,8.119796,9.104411,9.701744,9.593436,9.258667,7.8145647,6.5444107,6.308103,7.5421543,6.73477,6.5312824,6.5050263,6.770872,7.9885135,7.6996927,7.0465646,6.931693,7.204103,6.6527185,5.973334,4.962462,4.4734364,4.650667,4.9329233,4.8377438,4.4964104,4.588308,5.408821,6.8594875,8.730257,9.005949,8.093539,7.0990777,7.827693,9.07159,8.28718,7.860513,8.247795,7.9917955,8.198565,8.369231,8.966565,10.013539,11.083488,10.134975,9.53436,9.242257,9.268514,9.665642,8.306872,7.322257,6.308103,5.549949,6.0225644,6.744616,7.1187696,6.7183595,5.540103,3.9942567,3.0752823,3.2984617,3.7087183,3.7152824,3.1048207,3.2918978,3.0654361,2.986667,3.170462,3.2951798,2.2646155,1.7558975,1.3161026,0.8041026,0.37415388,0.26912823,0.27897438,0.30851284,0.58092314,1.6377437,0.6892308,1.654154,4.70318,7.5979495,5.677949,6.518154,5.100308,4.5390773,4.8640003,3.0260515,6.4754877,6.5312824,6.0783596,5.543385,2.8882053,1.9495386,2.3368206,2.5140514,2.1989746,2.359795,2.156308,2.6945643,2.1891284,0.761436,0.4135385,0.19692309,0.13456412,0.101743594,0.055794876,0.036102567,0.08861539,0.059076928,0.02297436,0.01969231,0.055794876,0.18379489,0.24287182,0.26912823,0.8008206,2.8914874,4.788513,6.6067696,10.19077,14.854566,17.378464,17.78872,16.128002,14.634667,13.686155,11.795693,11.07036,10.33518,9.393231,9.015796,10.919386,10.19077,9.810052,11.418258,13.594257,11.861334,13.403898,12.914873,12.189539,11.871181,11.451077,11.113027,11.533129,11.431385,10.880001,11.313231,10.213744,10.633847,10.8996935,10.679795,10.975181,11.201642,10.758565,10.184206,9.750975,9.468719,9.5835905,8.845129,8.021334,7.4732313,7.1483083,6.5050263,6.2884107,5.8453336,5.3694363,5.904411,5.8092313,5.651693,5.3431797,4.8607183,4.2535386,4.9493337,6.2194877,7.709539,8.963283,9.432616,8.953437,7.9917955,7.75877,7.6964107,5.4580517,3.0424619,1.7526156,1.3029745,1.4244103,1.8871796,4.023795,3.5971284,3.767795,4.7360005,3.757949,4.571898,4.8114877,3.6660516,2.0841026,2.7602053,3.6069746,3.9253337,4.46359,4.8311796,3.4789746,3.9844105,7.4108725,7.8408213,5.2644105,5.549949,5.031385,5.9634876,6.6822567,6.419693,5.32677,5.6451287,4.3290257,3.8596926,5.0642056,7.1056414,4.013949,2.4746668,1.6804104,2.5928206,7.955693,5.671385,6.8463597,7.7423596,7.259898,6.931693,11.949949,10.154668,8.674462,9.563898,9.787078,6.2194877,10.217027,13.899488,14.381949,13.784616,21.474463,21.047796,19.472412,17.874052,11.529847,9.865847,8.749949,11.588924,17.273438,20.168207,17.61477,15.038361,16.193642,17.962667,10.368001,6.2720003,6.6592827,7.2237954,6.311385,4.906667,4.1025643,5.927385,7.860513,8.746667,8.805744,6.452513,5.2578464,6.2916927,7.4797955,3.6069746,4.565334,5.0477953,4.8114877,5.0543594,8.41518,4.7556925,3.889231,3.8531284,3.9614363,4.785231,6.2687182,5.9963083,6.3474874,7.5487185,7.6734366,7.171283,5.664821,4.2962055,3.7776413,4.378257,4.4340515,4.457026,4.33559,4.4045134,5.4613338,5.671385,4.95918,4.7261543,5.097026,4.9296412,3.8038976,3.511795,3.3903592,3.1934361,3.1113849,2.5862565,2.9669745,3.8137438,5.0149746,6.7610264,6.242462,6.058667,6.416411,6.8660517,6.2884107,5.618872,4.8082056,4.0303593,3.570872,3.8367183,4.650667,4.381539,4.2994876,4.9132314,5.9667697,5.412103,5.477744,5.579488,5.2578464,4.1583595,4.9493337,5.0543594,5.182359,5.4547696,5.4153852,5.139693,5.028103,4.194462,2.8258464,2.162872,3.5774362,2.7733335,3.8695388,9.465437,20.647387,13.02318,5.85518,2.8225644,3.6004105,3.8301542,3.6594875,4.125539,4.44718,4.6112823,5.366154,5.72718,5.2578464,5.1331286,5.8190775,7.072821,6.892308,6.8627696,7.066257,7.174565,6.439385,6.157129,5.901129,5.097026,4.5817437,6.5903597,21.986464,26.607592,24.592413,19.10154,12.327386,9.242257,7.1023593,6.633026,7.962257,10.624001,12.297847,12.603078,13.371078,14.785643,15.376411,16.94195,17.194668,16.433231,15.921232,17.88718,18.586258,18.248207,17.752617,17.650873,18.159592,18.369642,18.054565,17.34236,16.70236,16.95836,16.764719,16.807386,17.362053,18.65518,20.867283,21.93395,20.548925,18.336823,16.452925,15.579899,17.880617,18.556719,18.307283,18.208822,19.712002,20.155079,19.83672,18.691284,17.650873,18.635489,19.24595,19.61354,19.761232,19.820309,20.020514,21.766565,22.035694,22.3639,23.026873,23.013746,21.238155,23.013746,22.95795,20.778667,21.264412,23.929438,24.782772,23.876925,22.075079,21.028105,20.289642,20.22072,21.408823,22.99077,22.665848,21.799387,21.188925,20.772104,20.404514,19.849848,19.337847,18.609232,17.742771,16.948515,16.561232,16.282257,16.160822,16.610462,17.78872,19.610258,21.175797,23.338669,24.100105,22.934977,20.788515,20.516104,20.01395,18.75036,17.283283,17.289848,18.550156,18.688002,18.231796,17.19795,15.107284,14.368821,13.528616,13.801026,14.713437,14.106257,14.697027,15.031796,14.998976,14.815181,15.025232,15.179488,14.519796,13.909334,13.653335,13.4859495,12.95754,12.419283,12.22236,12.57354,13.538463,0.48574364,0.4201026,0.35446155,0.34789747,0.39056414,0.4201026,0.5218462,0.61374366,0.6892308,0.7318975,0.69907695,0.8960001,0.83035904,0.86317956,1.0272821,0.9911796,0.90584624,0.9682052,1.0010257,0.9714873,0.9911796,1.401436,1.5721027,1.7460514,1.9429746,1.9659488,1.9200002,2.0151796,2.2514873,2.6420515,3.2098465,4.0434875,4.1846156,4.4832826,5.290667,6.4295387,7.4371285,7.637334,8.1755905,9.133949,9.53436,8.136206,8.050873,8.241231,8.274052,8.310155,8.513641,8.39877,8.241231,8.103385,7.821129,7.5520005,7.0925136,6.987488,7.1187696,6.7249236,8.001641,9.6754875,10.765129,11.175385,11.713642,12.071385,12.242052,12.609642,13.15118,13.426873,13.00677,12.3306675,11.71036,11.290257,11.047385,10.112,9.5835905,9.468719,9.714872,10.220308,10.8996935,11.608616,12.084514,12.156719,11.753027,11.434668,11.385437,11.648001,12.068104,12.297847,12.688411,12.744206,12.649027,12.73436,13.495796,14.152206,14.775796,15.31077,15.635694,15.576616,15.8654375,15.579899,15.143386,14.880821,15.018668,14.7331295,14.119386,13.548308,13.193847,13.036308,12.911591,12.62277,12.888617,13.656616,14.099693,13.5089245,12.73436,12.228924,12.028719,11.769437,11.674257,11.648001,11.158976,10.31877,9.875693,9.645949,9.622975,9.645949,9.800206,10.420513,11.556104,12.1928215,12.694975,13.124924,13.223386,14.342566,15.29436,16.006565,17.007591,19.416616,20.06318,19.744822,18.648617,17.345642,16.777847,17.270155,17.641027,18.231796,19.035898,19.70872,18.70113,17.824821,17.073233,16.771284,17.588514,19.515078,20.420925,20.87713,20.581745,18.36308,19.961437,20.624413,20.598156,20.122257,19.426462,20.374975,19.06872,17.700104,16.728617,14.890668,13.22995,13.686155,13.53518,12.182976,11.178667,10.433641,10.033232,10.213744,10.650257,10.459898,9.015796,7.834257,7.381334,7.6077952,7.9425645,7.4207187,6.8004107,6.340924,6.193231,6.4000006,6.2588725,5.970052,6.1078978,6.8004107,7.7259493,8.772923,8.858257,8.257642,7.752206,8.605539,8.421744,8.969847,9.554052,9.954462,10.423796,10.20718,9.639385,9.284924,9.245539,9.176616,7.8736415,7.972103,8.887795,9.728001,9.317744,9.291488,8.277334,7.240206,6.803693,7.213949,7.4863596,7.837539,7.6635904,7.387898,8.441437,8.1755905,7.686565,7.387898,7.318975,7.13518,5.605744,4.906667,4.788513,4.8640003,4.6112823,5.1331286,4.7392826,4.8804107,5.7698464,6.380308,7.893334,8.792616,8.651488,7.7981544,7.2992826,8.293744,8.402052,8.503796,8.789334,8.756514,8.769642,8.470975,8.923898,10.125129,10.985026,10.180923,10.322052,10.486155,10.138257,9.107693,7.8736415,6.672411,5.651693,5.152821,5.720616,6.5247183,6.738052,6.416411,5.723898,4.9394875,4.384821,4.388103,4.3618464,4.0303593,3.4231799,3.2918978,2.993231,2.930872,3.131077,3.2525132,2.2777438,1.910154,1.4342566,0.7253334,0.23958977,0.27241027,0.39712822,0.6071795,0.8172308,0.86317956,1.4506668,3.1081028,6.38359,9.360411,7.643898,5.225026,4.378257,4.201026,4.4077954,5.3398976,6.5345645,5.835488,5.435077,5.3760004,3.5446157,2.9833848,3.4133337,3.4494362,2.7963078,2.2186668,2.8750772,2.8488207,1.8346668,0.47261542,0.34133336,0.18707694,0.15425642,0.12143591,0.07876924,0.16410258,0.08533334,0.03938462,0.013128206,0.006564103,0.032820515,0.108307704,0.2100513,0.6498462,1.8313848,4.2338467,6.764308,9.363693,12.258463,14.710155,15.025232,14.381949,13.423591,13.00677,12.950975,12.051693,11.579078,11.067078,10.223591,9.337437,9.288206,9.124104,10.509129,11.992617,12.455385,11.113027,12.57354,12.25518,11.72677,11.664412,11.844924,11.487181,11.441232,11.562668,11.700514,11.687386,10.256411,10.512411,10.952206,11.113027,11.585642,11.45436,11.250873,10.912822,10.509129,10.256411,9.91836,9.104411,8.067283,7.1154876,6.619898,5.927385,5.8092313,5.477744,5.0576415,5.5663595,5.8814363,6.1440005,6.2752824,6.0192823,4.9460516,5.425231,5.668103,6.193231,7.0400004,7.7718983,7.8769236,7.748924,7.899898,8.165744,7.683283,5.7435904,3.2918978,1.6705642,1.4276924,2.3236926,6.226052,4.9493337,3.4100516,3.2623591,2.8717952,3.4297438,3.2196925,2.806154,2.9604106,4.663795,4.775385,4.8738465,5.142975,5.333334,4.768821,4.2929235,5.044513,4.4701543,3.0818465,4.4767184,4.9329233,5.477744,6.36718,6.8332314,5.080616,9.07159,7.8506675,6.9743595,7.5520005,6.2162056,3.895795,2.8160002,3.1343591,5.5171285,11.142565,8.352821,9.655796,10.364718,8.861539,6.6034875,9.872411,8.78277,7.450257,7.9130263,10.128411,8.090257,11.575796,14.208001,13.292309,9.816616,13.522053,13.3251295,12.514462,12.727796,13.965129,15.205745,14.368821,14.933334,17.060104,17.575386,12.596514,10.157949,9.833026,10.640411,11.0605135,9.196308,9.488411,9.668923,8.917334,7.8703594,4.2863593,4.7589746,5.668103,5.481026,4.7261543,5.4514875,5.7107697,6.547693,7.145026,4.8344617,4.637539,7.4830775,7.722667,5.0543594,4.5456414,3.6069746,3.0752823,3.2032824,4.010667,5.284103,6.6625648,7.315693,7.955693,8.631796,8.726975,8.224821,7.0826674,5.405539,3.9876926,4.3060517,4.7589746,5.0642056,5.2381544,5.4449234,6.0028725,6.173539,5.353026,4.8738465,4.962462,4.7360005,3.9778464,3.698872,3.639795,3.620103,3.5413337,3.3345644,4.204308,5.1167183,5.681231,6.1472826,6.042257,6.1538467,6.47877,6.76759,6.5312824,5.717334,4.906667,4.2962055,4.0402055,4.2535386,4.2896414,4.4373336,4.8607183,5.3924108,5.536821,5.2578464,5.5991797,5.32677,4.5029745,4.457026,4.7458467,5.0838976,5.3891287,5.5762057,5.546667,4.95918,4.4964104,4.023795,3.4592824,2.802872,3.373949,3.0293336,3.2886157,5.5565133,11.113027,6.166975,3.8006158,3.4330258,3.9680004,3.8104618,3.3805132,3.820308,4.1452312,4.1846156,4.571898,4.955898,4.5029745,4.457026,5.21518,6.340924,6.3606157,6.518154,6.121026,5.4875903,5.9470773,5.6385646,5.228308,4.7556925,4.417641,4.5554876,13.407181,19.511797,21.27754,18.806156,13.873232,9.744411,7.958975,6.87918,6.2490263,7.207385,7.8539495,9.449026,11.211488,12.514462,12.914873,14.50995,14.989129,14.897232,14.91036,15.816206,16.836924,17.493334,17.178257,16.242872,16.01313,16.57436,16.83036,16.420103,15.645539,15.471591,15.737437,16.101746,16.357744,16.846771,18.451694,19.236105,18.146463,16.564514,15.317334,14.667488,15.172924,15.333745,15.360002,15.698052,17.046976,17.798565,18.625643,18.60595,18.133335,18.907898,19.62995,19.610258,19.042463,18.471386,18.789745,20.273232,20.12554,20.151796,20.686771,20.62113,20.276514,21.792822,21.622156,19.843283,20.171488,22.92513,25.232412,24.937027,22.107899,19.01949,19.088411,19.899078,21.142977,22.12431,21.776411,21.412104,21.093744,20.818052,20.5719,20.329027,19.662771,19.006361,18.17272,17.35877,17.109335,16.603899,16.311796,16.587488,17.539284,19.009642,21.658258,30.831593,39.86708,42.584618,33.266876,24.06072,19.104822,16.741745,15.954053,16.344616,17.572104,17.749334,16.659693,15.117129,14.959591,14.621539,14.112822,14.467283,15.29436,14.759386,15.8654375,16.055796,15.451899,14.63795,14.65436,15.012104,14.375385,13.833847,13.764924,13.846975,13.59754,12.524308,11.723488,11.661129,12.163283,0.6629744,0.41025645,0.38400003,0.42338464,0.45620516,0.50543594,0.5513847,0.571077,0.69579494,0.86646163,0.8402052,1.014154,0.9485129,0.86974365,0.8795898,0.9616411,1.0601027,1.1126155,1.0601027,1.0075898,1.2176411,1.6508719,1.8904617,2.1169233,2.3729234,2.5829747,2.7437952,2.7208207,2.8455386,3.2229745,3.7185643,4.4045134,4.4110775,4.647385,5.3103595,5.8945646,6.5411286,7.3386674,7.9130263,8.4053335,9.485129,8.704,8.953437,8.897642,8.214975,7.5946674,7.860513,8.100103,8.2904625,8.346257,8.139488,7.7718983,7.4141545,7.456821,7.8441033,8.086975,9.691898,11.208206,11.926975,11.871181,11.792411,11.776001,12.419283,13.259488,13.952001,14.283488,13.515489,12.704822,11.913847,11.195078,10.607591,9.67877,9.540924,9.645949,9.737847,9.865847,10.138257,11.021129,11.562668,11.523283,11.355898,11.1064625,11.332924,11.835078,12.448821,13.056001,13.259488,13.318565,13.184001,13.121642,13.682873,14.083283,14.63795,15.126975,15.40595,15.419078,15.717745,15.402668,14.772514,14.25395,14.372104,14.162052,13.453129,12.793437,12.438975,12.383181,12.645744,12.744206,13.115078,13.6237955,13.568001,12.698257,12.448821,12.78359,13.249642,12.983796,12.182976,12.107488,11.776001,10.994873,10.358154,9.819899,9.872411,10.003693,10.075898,10.312206,11.0375395,11.690667,12.547283,13.449847,13.814155,14.644514,15.82277,17.056822,18.208822,19.291899,17.942976,17.490053,16.981335,16.28554,16.075489,16.810667,17.345642,18.054565,18.714258,18.507488,18.005335,17.174976,16.695797,16.896002,17.739489,19.055592,20.178053,20.67036,20.250257,18.78318,19.941746,21.297232,20.742565,18.816002,18.67159,21.097027,20.329027,19.183592,18.612514,17.70995,14.34913,13.010053,12.501334,12.1238985,11.667693,10.981745,10.525539,10.571488,10.975181,11.18195,10.312206,8.6580515,7.893334,8.4053335,9.32759,8.195283,7.506052,7.2861543,7.3419495,7.240206,7.059693,6.6395903,6.5312824,6.8660517,7.3353853,8.228104,8.553026,8.214975,7.7259493,8.201847,8.185436,8.553026,9.143796,9.816616,10.456616,10.092308,8.868103,8.169026,8.441437,9.219283,8.628513,8.39877,8.595693,8.923898,8.713847,9.078155,8.375795,7.3419495,6.7150774,7.2270775,8.113232,8.838565,8.55959,7.781744,8.372514,8.585847,8.467693,7.9458466,7.276308,7.056411,5.4383593,5.097026,5.221744,5.221744,4.7261543,5.333334,5.1659493,5.61559,6.5969234,6.564103,7.5946674,8.576,9.133949,8.982975,7.958975,8.786052,9.468719,9.452309,9.091283,9.6295395,9.403078,8.848411,9.019077,9.852718,10.187488,9.895386,10.427077,10.676514,10.19077,9.186462,8.234667,6.311385,5.1167183,5.0838976,5.3727183,6.048821,6.301539,6.439385,6.432821,5.8978467,4.857436,4.6966157,4.535795,4.069744,3.5938463,2.9702566,2.7109745,2.9505644,3.2525132,2.5895386,2.1202054,1.7099489,1.1323078,0.5152821,0.31507695,0.4004103,0.71548724,0.955077,0.86317956,0.2100513,1.5064616,4.5128207,8.208411,10.180923,6.619898,4.6966157,5.5532312,8.077128,9.82318,7.00718,5.6418467,4.397949,4.059898,4.2863593,3.5938463,3.8400004,4.073026,3.9647183,3.2787695,1.8510771,2.412308,2.0939488,1.211077,0.32820517,0.24287182,0.15753847,0.14769232,0.10502565,0.055794876,0.16410258,0.052512825,0.016410258,0.026256412,0.09189744,0.23958977,0.27569234,0.6170257,1.595077,3.4297438,6.23918,9.104411,11.10318,12.763899,13.722258,12.73436,12.498053,12.291283,11.910565,11.313231,10.637129,10.315488,10.289231,10.033232,9.468719,8.969847,9.833026,10.896411,11.641437,11.730052,10.994873,11.979488,12.360206,12.130463,11.805539,12.422565,11.700514,11.529847,11.943385,12.3766165,11.67754,10.121847,10.184206,10.482873,10.709334,11.61518,11.369026,11.441232,11.592206,11.569232,11.093334,10.676514,9.603283,8.231385,7.000616,6.436103,5.5007186,5.044513,4.70318,4.598154,5.346462,5.943795,6.3606157,6.4722056,6.2227697,5.605744,5.792821,5.431795,5.395693,5.7107697,5.5630774,5.7468724,6.160411,6.3474874,6.485334,7.384616,6.889026,4.9427695,2.8127182,1.5556924,2.034872,5.5204105,4.9887185,3.8367183,3.511795,3.5314875,3.0293336,2.6420515,3.0884104,4.2338467,5.110154,4.8049235,4.818052,5.0609236,5.467898,5.98318,4.345436,2.5271797,2.4484105,4.309334,6.6133337,6.948103,5.4875903,5.7829747,7.512616,6.5017443,9.849437,9.015796,8.04759,7.6668725,5.2512827,5.139693,3.9154875,3.6726158,5.4514875,9.248821,7.200821,8.549745,9.153642,8.362667,9.03877,8.267488,6.180103,5.074052,5.85518,8.054154,7.4404106,9.521232,10.102155,8.576,7.9425645,7.6734366,6.567385,5.8256416,7.397744,13.978257,18.06113,16.955078,16.65313,17.306257,13.1872835,9.816616,10.095591,9.291488,7.1844106,8.064001,10.174359,11.565949,11.667693,10.282667,7.5913854,4.059898,3.7710772,3.5840003,2.858667,3.4625645,5.2348723,6.7183595,7.5552826,7.3780518,5.8223596,4.1025643,6.921847,7.515898,4.562052,2.1497438,3.1474874,3.4592824,4.007385,5.0477953,6.1768208,7.1483083,7.9786673,8.838565,9.340718,8.539898,7.5881033,7.4141545,6.5870776,5.287385,5.3005133,5.733744,5.648411,5.5597954,5.8125134,6.5903597,6.665847,6.2785645,5.8289237,5.425231,4.857436,4.2994876,3.948308,3.9154875,4.1550775,4.457026,4.2929235,5.3070774,6.055385,5.907693,5.024821,5.2611284,5.907693,6.2555904,6.1440005,5.9503593,5.533539,5.1364107,4.8049235,4.571898,4.457026,4.1517954,4.4865646,5.028103,5.362872,5.097026,4.7491283,5.172513,4.9427695,4.1813335,4.5423594,4.637539,5.32677,5.5302567,5.1626673,5.139693,5.146257,4.5489235,4.0336413,3.7874875,3.4921029,3.6004105,3.1507695,2.5928206,2.6026669,4.066462,2.6486156,3.3936412,4.2469745,4.273231,3.6824617,3.383795,3.6824617,3.9253337,4.0041027,4.352,4.535795,4.1747694,4.194462,4.778667,5.35959,5.920821,6.1768208,5.297231,4.059898,4.8607183,4.7425647,4.6178465,4.594872,4.519385,3.9778464,6.311385,13.387488,17.243898,15.488001,11.303386,8.576,8.477539,8.172308,7.384616,8.392206,8.572719,9.107693,10.069334,11.158976,11.700514,13.088821,13.302155,13.682873,14.355694,14.230975,14.880821,15.881847,16.28554,15.826053,14.913642,15.524104,15.862155,15.698052,15.133539,14.611693,14.828309,15.182771,15.415796,15.616001,16.22318,16.049232,15.448617,14.864411,14.418053,13.929027,13.1872835,13.371078,14.070155,14.946463,15.691488,16.31836,17.132309,17.572104,17.70995,18.244925,18.743795,18.822565,18.58954,18.330257,18.514053,19.8039,19.035898,18.034874,17.72636,18.14318,19.35754,20.404514,20.496412,19.968002,20.28636,22.44595,24.415182,24.192001,21.707489,18.82913,18.901335,19.360823,20.224,21.13313,21.343182,21.664822,21.540104,21.251284,20.978874,20.79836,19.859694,19.50195,18.819284,17.69354,16.81395,16.393847,16.347898,16.59077,17.204514,18.454975,21.257847,34.097233,49.555695,57.964314,47.382977,30.240824,20.407797,15.730873,14.513232,15.504412,16.794258,16.879591,15.524104,13.761642,13.896206,14.454155,14.601848,14.972719,15.484719,15.337027,16.784412,16.331488,15.153232,14.080001,13.59754,13.797745,13.817437,13.748514,13.525334,12.941129,13.033027,12.3306675,11.516719,11.024411,11.034257,0.6826667,0.34789747,0.4004103,0.44307697,0.39712822,0.49887183,0.50543594,0.46933338,0.62030774,0.8730257,0.82379496,0.9353847,0.9714873,0.9353847,0.8960001,0.9747693,1.1093334,1.1520001,1.1684103,1.273436,1.6114873,1.7558975,2.1530259,2.4976413,2.7208207,2.989949,3.4756925,3.3050258,3.2722054,3.6562054,4.2305646,4.2601027,4.240411,4.6572313,5.2512827,4.9920006,5.293949,6.688821,7.259898,7.0892315,8.251078,9.32759,9.42277,8.746667,7.8080006,7.427283,7.6734366,8.149334,8.385642,8.231385,7.8703594,7.975385,7.643898,7.6274877,8.260923,9.442462,11.398565,12.504617,12.63918,12.274873,12.47836,11.539693,12.097642,13.15118,14.050463,14.473847,13.99795,13.2562065,12.363488,11.369026,10.236719,9.819899,10.010257,10.069334,9.764103,9.373539,9.347282,10.006975,10.433641,10.453334,10.630565,10.788103,11.264001,11.785847,12.219078,12.586668,13.013334,13.387488,13.771488,14.112822,14.273643,14.171899,14.555899,15.094155,15.530668,15.675078,15.609437,15.012104,13.787898,12.635899,13.056001,13.367796,12.777026,12.032001,11.713642,12.22236,12.780309,13.344822,13.587693,13.387488,12.822975,11.648001,11.798975,12.747488,13.702565,13.636924,12.386462,12.120616,12.035283,11.723488,11.16554,10.246565,10.180923,10.348309,10.492719,10.732308,11.418258,12.015591,12.258463,12.504617,13.761642,14.303181,15.75713,17.165129,17.952822,17.946259,14.982565,14.546052,15.104001,15.681643,15.868719,16.83036,17.224207,17.782156,18.451694,18.422155,18.418873,17.64431,17.174976,17.595078,18.999796,18.947283,19.872822,20.230566,19.603693,18.714258,20.115694,22.104616,21.451488,18.799591,18.665028,21.113438,20.447182,19.360823,19.144207,19.698874,15.77354,12.836103,11.408411,11.526565,12.708103,11.785847,10.788103,10.453334,10.889847,11.552821,11.972924,10.272821,8.992821,9.058462,9.764103,8.667898,8.402052,8.635077,8.78277,8.027898,7.768616,7.5487185,7.282872,7.076103,7.2172313,7.4404106,7.8802056,7.890052,7.571693,7.79159,8.316719,8.5202055,8.996103,9.865847,10.752001,10.390975,8.792616,7.9950776,8.4053335,8.802463,8.989539,9.028924,8.78277,8.51036,8.87795,9.435898,8.726975,7.3091288,6.3179493,7.4765134,8.349539,8.960001,8.674462,7.834257,7.768616,8.362667,8.615385,8.3823595,7.7456417,7.026872,6.189949,5.61559,5.362872,5.35959,5.421949,5.6385646,5.651693,6.114462,6.8660517,6.941539,8.054154,8.73354,9.340718,9.6984625,9.110975,10.105436,10.948924,10.499283,9.399796,10.075898,9.91836,9.53436,9.366975,9.429334,9.31118,9.6,9.849437,9.865847,9.69518,9.6295395,8.720411,6.304821,5.0674877,5.333334,5.0871797,5.287385,5.8420515,6.4656415,6.705231,5.940513,4.667077,4.5587697,4.3651285,3.8498464,3.7874875,2.5895386,2.3893335,2.8258464,2.9768207,1.3653334,1.4309745,1.079795,0.5973334,0.31507695,0.5940513,0.574359,0.8763078,0.9288206,0.636718,0.38400003,1.017436,5.4416413,9.278359,9.186462,2.8488207,5.3070774,7.4436927,12.310975,15.67836,6.055385,3.748103,2.7208207,2.6190772,2.7733335,2.2219489,3.7743592,3.5905645,3.2820516,2.9013336,0.9419488,0.86646163,0.72861546,0.54482055,0.3249231,0.0951795,0.15425642,0.190359,0.12143591,0.006564103,0.036102567,0.016410258,0.03938462,0.18707694,0.4266667,0.6104616,0.7089231,1.404718,3.2361028,6.0324106,8.914052,11.211488,11.126155,11.506873,12.544001,11.798975,12.672001,11.979488,10.59118,9.028924,7.4797955,7.276308,7.9261546,8.700719,9.179898,9.284924,11.08677,10.896411,11.119591,11.963078,11.434668,11.562668,12.839386,12.977232,12.091078,12.704822,11.746463,11.894155,12.521027,12.865642,12.038565,10.246565,9.977437,9.990565,10.108719,11.23118,11.227899,11.441232,11.96636,12.304411,11.362462,11.23118,9.990565,8.339693,6.9054365,6.2720003,5.287385,4.634257,4.204308,4.2141542,5.1922054,6.091488,6.619898,6.449231,5.9470773,6.1768208,6.058667,5.546667,5.3234878,5.149539,3.8498464,4.0008206,4.4701543,4.450462,4.2568207,5.293949,6.301539,6.298257,4.919795,2.9505644,2.3236926,3.754667,4.493129,4.9362054,4.9821544,4.027077,3.0687182,2.937436,3.69559,4.4964104,3.5807183,3.43959,3.8071797,4.3651285,5.0084105,5.858462,3.2722054,1.8543591,3.239385,7.1876926,11.569232,10.04636,6.5837955,5.431795,7.1089234,8.418462,7.1122055,6.8562055,6.6560006,6.038975,5.041231,5.8847184,4.309334,2.6978464,2.4057438,3.767795,3.0818465,4.9952826,5.5236926,5.536821,10.771693,8.487385,4.650667,3.948308,6.308103,6.9021544,6.2030773,6.554257,6.4000006,6.4656415,9.754257,8.15918,5.7435904,4.135385,5.172513,10.893129,13.581129,11.618463,13.233232,16.07877,7.2303596,7.788308,11.063796,11.283693,7.722667,4.716308,8.306872,10.6469755,11.083488,9.186462,4.7294364,4.210872,4.5456414,3.5347695,2.2350771,4.955898,5.1298466,6.314667,7.5585647,7.7948723,5.835488,3.4100516,3.639795,3.9811285,3.7054362,3.9253337,4.020513,4.453744,5.421949,6.675693,7.5191803,7.890052,7.781744,8.277334,8.897642,7.6012316,6.1472826,6.5345645,6.8693337,6.564103,6.3310776,6.941539,6.173539,5.4482055,5.6451287,7.13518,7.207385,7.2336416,7.059693,6.5870776,5.7829747,5.1298466,4.601436,4.5423594,4.955898,5.4908724,5.1954875,5.796103,6.0258465,5.477744,4.601436,4.8771286,5.687795,6.0717955,5.7534366,5.152821,5.4580517,5.5236926,5.225026,4.71959,4.4242053,4.2896414,4.2896414,4.381539,4.59159,5.0215387,4.391385,4.450462,4.6145644,4.650667,4.6802053,4.7589746,5.536821,5.674667,5.0838976,4.896821,5.356308,4.8640003,4.0434875,3.4888208,3.7743592,3.7907696,3.2065644,2.5632823,2.4320002,3.4100516,3.5610259,4.2305646,4.5456414,4.2240005,3.5610259,3.56759,3.7218463,3.889231,4.0500517,4.315898,4.4701543,4.535795,4.644103,4.8016415,4.857436,5.6976414,5.8880005,4.965744,3.6890259,4.0369234,4.0533338,4.3749747,4.6834874,4.706462,4.2338467,5.9602056,12.987078,15.094155,10.86359,7.6964107,7.4732313,9.271795,10.108719,9.800206,10.971898,10.213744,9.875693,10.157949,11.011283,12.166565,13.272616,13.177437,13.472821,14.102976,13.338258,13.479385,14.165335,15.186052,15.809642,14.795488,15.0777445,14.9398985,14.811898,14.677335,14.080001,14.001232,14.309745,14.834873,15.16636,14.63795,13.50236,13.492514,13.715693,13.732103,13.581129,12.76718,12.941129,14.024206,15.363283,15.747283,15.694771,15.468308,15.55036,16.042667,16.705643,16.748308,17.362053,18.116924,18.579693,18.33354,19.472412,18.57313,17.027283,16.059078,16.748308,18.166155,18.714258,19.56431,20.880411,21.80595,23.026873,23.30913,22.95795,22.229336,21.300514,19.984411,19.19672,19.426462,20.457027,21.382566,22.288412,22.180105,21.654976,21.090464,20.667078,19.423182,19.314873,18.921026,17.719797,16.09518,15.747283,16.187078,16.384,16.426668,17.529438,19.524925,29.128208,43.185234,53.89457,48.804108,33.437542,22.764309,16.111591,13.124924,13.755078,15.465027,15.940925,15.356719,14.194873,13.262771,14.749539,15.632411,16.019693,16.114874,16.249437,17.391592,15.842463,14.158771,13.2562065,12.42913,12.35036,13.545027,14.267078,13.732103,12.114052,12.058257,12.09436,11.661129,10.86359,10.469745,0.36758977,0.39056414,0.38728207,0.33805132,0.32820517,0.5481026,0.6235898,0.60389745,0.5316923,0.48246157,0.58092314,0.8008206,0.8467693,1.0601027,1.3522053,1.204513,1.401436,1.3751796,1.3653334,1.463795,1.6475899,2.2711797,2.6551797,2.868513,2.9801028,3.0523078,3.8564105,3.7842054,3.570872,3.6791797,4.3027697,3.6693337,4.066462,4.8016415,5.297231,5.1265645,5.4186673,5.8880005,6.058667,6.1046157,6.8365135,7.860513,7.4043083,6.560821,6.439385,8.149334,7.9163084,7.8408213,8.034462,8.103385,7.125334,6.4295387,6.2916927,6.7085133,7.7456417,9.55077,11.273847,12.297847,12.560411,12.406155,12.58995,12.393026,12.455385,13.430155,14.805334,14.87754,15.182771,14.152206,12.527591,11.017847,10.28595,11.139283,10.811078,10.023385,9.472001,9.826463,9.435898,9.93477,10.390975,10.532104,10.725744,11.372309,11.930258,12.186257,12.1468725,12.025436,12.842668,13.512206,14.227694,14.992412,15.638975,15.323898,15.645539,16.249437,16.771284,16.846771,15.491283,13.860104,12.547283,11.956513,12.297847,13.46954,13.489232,12.701539,11.831796,11.979488,12.527591,13.679591,14.628103,14.592001,12.849232,11.113027,11.047385,11.680821,12.402873,12.941129,12.071385,11.460924,11.204924,11.250873,11.398565,10.994873,11.030975,11.080206,11.099898,11.428103,12.22236,12.905026,12.983796,13.016617,14.601848,15.602873,16.118155,15.681643,14.749539,14.726565,14.79877,15.090873,15.652103,16.101746,15.625848,16.820515,16.571077,16.613745,17.385027,18.021746,18.678156,18.422155,18.372925,19.062155,20.417643,18.340103,18.609232,18.901335,18.38277,17.700104,19.495386,21.490873,22.400002,22.166977,21.973335,20.788515,18.569847,17.526155,17.831387,17.624617,15.914668,13.722258,11.943385,11.155693,11.595488,11.864616,10.220308,8.976411,9.101129,10.223591,12.225642,12.442257,11.195078,9.432616,8.713847,8.713847,8.493949,8.352821,8.12636,7.1876926,7.5421543,7.5552826,7.4765134,7.499488,7.765334,7.6570263,7.6570263,7.6012316,7.522462,7.643898,8.024616,8.546462,9.035488,9.616411,10.725744,10.886565,9.964309,9.317744,8.960001,7.568411,7.6767187,8.87795,9.842873,10.220308,10.633847,10.794667,10.148104,8.956718,7.8047185,7.5979495,8.454565,8.720411,8.795898,8.612103,7.6603084,7.8441033,8.044309,8.507077,8.835282,7.9786673,7.893334,6.380308,5.106872,4.896821,5.7534366,6.3507695,6.3277955,6.117744,6.160411,6.882462,7.9917955,8.746667,8.674462,8.198565,8.635077,9.941334,11.303386,11.69395,11.040821,10.223591,10.502565,10.20718,9.665642,9.163487,8.956718,9.665642,9.67877,10.049642,10.240001,8.103385,6.9809237,6.2687182,5.907693,5.661539,5.110154,4.2568207,5.106872,5.661539,5.284103,4.6834874,5.1954875,5.280821,4.5522056,3.5446157,3.6758976,2.3236926,2.1497438,2.2088206,1.9987694,1.4506668,0.8041026,0.44964105,0.28882053,0.36430773,0.8402052,0.5349744,0.27569234,0.17066668,0.39712822,1.1913847,1.8609232,5.7829747,7.785026,6.2030773,2.8849232,5.47118,3.5478978,2.477949,3.2984617,2.6847181,1.6475899,1.6344616,1.6311796,1.2570257,0.79425645,4.210872,3.114667,1.8642052,1.6640002,0.56451285,0.3708718,0.24615386,0.15425642,0.08205129,0.04594872,0.3511795,0.446359,0.27569234,0.0,0.0,0.0,0.17394873,0.7187693,1.2340513,0.7318975,1.0371283,1.8904617,5.674667,10.732308,11.369026,10.843898,8.549745,7.9786673,9.55077,10.650257,10.5780525,9.120821,7.9130263,6.8693337,4.197744,4.5390773,5.2447186,6.9120007,8.684308,8.27077,10.102155,11.099898,12.199386,12.888617,11.21477,11.897437,13.3251295,13.453129,12.3995905,12.435693,11.641437,11.818667,12.514462,13.223386,13.380924,11.306667,10.220308,10.249847,10.939077,11.23118,11.119591,11.871181,11.98277,11.1064625,10.056206,10.276103,9.432616,8.152616,6.882462,5.904411,5.5762057,5.832206,5.6418467,4.923077,4.532513,5.7632823,6.633026,6.875898,6.5903597,6.226052,6.2752824,5.72718,4.7622566,3.82359,3.6168208,4.240411,4.9985647,4.9854364,4.342154,4.2568207,6.4065647,7.683283,7.9524107,7.2172313,5.6287184,6.741334,6.1768208,5.0182567,3.8334363,2.6847181,2.9669745,3.0654361,3.436308,3.895795,3.6168208,3.446154,3.2196925,3.2000003,3.6627696,4.8836927,3.1376412,1.7591796,1.4342566,3.9417439,12.130463,8.418462,6.1538467,4.9526157,4.916513,6.636308,6.698667,7.125334,7.2237954,7.0793853,7.568411,5.431795,4.2469745,2.8816411,1.7066668,2.609231,3.5610259,5.3727183,5.277539,3.7382567,4.4701543,4.5817437,4.535795,8.982975,14.641232,10.282667,11.808822,8.858257,10.801231,16.928822,16.479181,11.437949,8.218257,6.235898,5.3858466,6.058667,3.3345644,3.6890259,5.6418467,7.8145647,8.92718,11.378873,12.47836,9.43918,4.9985647,7.4141545,6.0717955,4.850872,4.3060517,4.6080003,5.5236926,7.4765134,8.119796,5.9667697,3.0030773,4.699898,3.515077,2.8160002,2.9571285,3.8564105,5.0051284,3.3312824,2.3729234,1.9167181,2.6322052,6.0717955,6.547693,7.0334363,7.6734366,8.152616,7.6898465,8.470975,7.8703594,6.6133337,5.8190775,7.003898,5.733744,5.287385,5.5269747,5.904411,5.477744,6.9054365,6.961231,6.813539,7.2205133,8.513641,7.64718,6.672411,6.2851286,6.370462,5.9667697,4.9887185,4.388103,4.493129,4.9788723,4.8672824,5.149539,5.4843082,5.21518,4.565334,4.637539,4.345436,4.841026,5.07077,4.893539,5.0674877,5.431795,5.6418467,5.2348723,4.4242053,4.1189747,4.132103,4.0336413,4.1025643,4.4964104,5.2644105,4.716308,4.4045134,4.8311796,5.536821,5.097026,5.1954875,5.1922054,5.549949,5.8486156,4.775385,4.276513,3.7185643,3.255795,3.249231,4.2863593,3.639795,3.9351797,3.5774362,2.737231,3.370667,3.895795,4.578462,4.4996924,3.7809234,3.5872824,3.4756925,3.5872824,3.7809234,3.8498464,3.508513,4.0467696,4.667077,5.0510774,5.211898,5.4941545,6.2752824,6.0750775,5.221744,4.391385,4.6244106,4.073026,4.276513,4.709744,5.110154,5.477744,3.8662567,7.722667,12.291283,14.214565,11.503591,9.3078985,10.827488,12.12718,11.336206,8.651488,7.456821,7.8802056,9.032206,10.640411,13.046155,13.692719,13.341539,13.147899,12.911591,11.093334,12.534155,14.093129,14.598565,14.221129,14.464001,14.027489,13.203693,13.482668,14.496821,14.007796,13.128206,14.503386,15.691488,15.445334,13.686155,12.980514,12.757335,12.859077,13.239796,13.945437,13.545027,13.203693,13.827283,15.258258,16.295385,16.662975,16.141129,15.461744,15.264822,16.082052,16.338053,17.263592,17.47036,16.94195,17.014154,16.856617,17.345642,17.906874,17.906874,16.662975,15.940925,15.809642,17.499899,20.548925,22.78072,24.598976,25.071592,26.404104,27.66113,24.77949,20.936207,19.689028,19.39036,19.528206,20.736002,21.88472,21.540104,21.031385,20.752413,20.14195,18.468103,17.595078,17.306257,17.352207,17.424412,16.508718,16.472616,16.259283,15.980309,16.905848,16.33477,16.886156,19.446156,22.472206,22.019283,25.731283,24.021336,19.075283,13.4859495,10.240001,12.534155,13.75836,14.690463,15.547078,15.960617,16.948515,18.405745,19.328001,19.265642,18.326975,17.385027,15.31077,13.771488,13.200411,12.770463,12.675283,15.195899,16.896002,16.656412,15.655386,14.106257,13.08554,12.458668,11.88759,10.850462,0.46276927,0.63343596,0.54482055,0.49887183,0.5907693,0.6826667,0.74830776,0.8369231,0.7581539,0.5874872,0.6662565,1.0305642,1.1782565,1.2077949,1.1946667,1.1946667,1.3292309,1.3423591,1.3357949,1.4539489,1.8806155,2.1103592,2.6551797,3.7120004,4.6112823,3.7973337,3.7021542,3.4724104,3.4494362,3.6332312,3.6791797,3.3575387,3.9811285,4.4373336,4.4701543,4.699898,5.080616,4.926359,5.169231,5.789539,5.8092313,7.2172313,8.041026,8.067283,7.6701546,7.8080006,7.6242056,8.027898,8.2904625,7.9524107,6.820103,6.5050263,7.2927184,8.237949,9.07159,10.174359,11.552821,12.458668,12.645744,12.209231,11.562668,11.319796,12.035283,13.259488,14.477129,15.097437,15.471591,14.9628725,13.909334,12.747488,12.005745,12.373334,11.050668,9.842873,9.465437,9.547488,9.741129,10.364718,10.817642,10.9226675,10.9226675,11.579078,11.881026,12.087796,12.422565,13.062565,13.751796,14.112822,14.6871805,15.333745,15.248411,15.225437,15.409232,15.281232,14.998976,15.40595,14.381949,13.384206,12.698257,12.35036,12.114052,12.251899,12.649027,13.193847,13.59754,13.3940525,13.308719,13.564719,14.050463,14.198155,12.970668,12.320822,12.100924,12.025436,11.900719,11.608616,10.148104,9.613129,9.852718,10.640411,11.703795,11.739899,11.447796,11.136001,10.985026,11.050668,11.569232,11.798975,12.251899,13.190565,14.601848,15.182771,15.632411,15.688207,15.744001,16.810667,16.436514,16.46277,17.043694,17.67713,17.211079,17.792002,17.434258,17.959387,19.433027,20.145233,20.178053,19.662771,18.983387,18.816002,20.112411,20.65395,21.093744,20.936207,20.306053,19.945026,22.347488,23.02031,22.298258,20.716309,19.006361,18.691284,18.842258,18.648617,17.864206,16.817232,16.055796,15.95077,15.484719,14.244103,12.438975,11.536411,10.453334,9.508103,9.07159,9.590155,11.562668,12.475078,12.12718,10.880001,9.6525135,9.340718,9.481847,9.452309,9.170052,9.078155,8.54318,7.972103,7.8736415,8.293744,8.815591,8.687591,8.4053335,7.958975,7.634052,8.011488,8.12636,8.395488,8.39877,8.162462,8.152616,9.258667,10.689642,11.674257,11.670976,10.374565,8.697436,9.252103,10.282667,10.771693,10.463181,8.434873,7.578257,7.4929237,7.571693,7.0137444,7.243488,7.9327188,8.900924,9.563898,8.953437,8.786052,8.444718,8.487385,8.684308,8.004924,7.702975,6.672411,5.9930263,5.8781543,5.677949,6.5805135,6.6034875,6.741334,7.3419495,8.090257,7.8441033,8.615385,9.275078,9.255385,8.562873,9.488411,10.564924,11.119591,10.781539,9.465437,10.410667,10.368001,10.177642,9.924924,8.94359,8.5202055,8.477539,9.26195,9.872411,7.834257,6.3606157,5.1856413,4.1878977,3.4756925,3.4166157,4.6802053,6.1538467,6.8660517,6.5739493,5.7698464,5.110154,4.0500517,3.121231,2.5796926,2.4188719,2.0512822,2.1300514,2.1792822,1.975795,1.5721027,0.78769237,0.6268718,0.62030774,0.57764107,0.5940513,0.80738467,0.60389745,0.39384618,0.9353847,3.3509746,6.2096415,5.5597954,6.245744,8.4972315,7.899898,7.6274877,4.4734364,2.8258464,3.1113849,1.8182565,1.1126155,1.1684103,1.4473847,1.6771283,1.8674873,1.9364104,1.4900514,1.1093334,0.8763078,0.380718,0.20676924,0.11158975,0.08205129,0.0951795,0.108307704,0.31507695,0.2100513,0.06235898,0.0,0.0,0.009846155,0.3249231,0.7844103,1.1946667,1.3193847,2.1792822,4.565334,7.9163084,10.115283,7.499488,7.6668725,7.817847,8.441437,9.199591,8.930462,8.211693,7.50277,6.6560006,5.618872,4.4406157,5.4547696,6.6461544,9.137232,11.437949,9.429334,8.946873,11.336206,13.069129,12.714667,10.935796,10.981745,11.611898,11.936821,11.71036,11.336206,11.168821,11.720206,12.924719,13.991385,13.4170265,11.654565,10.9686165,10.824206,10.925949,11.218052,9.43918,10.394258,10.981745,10.325335,9.77395,9.895386,9.586872,8.891078,7.6964107,5.733744,5.149539,5.10359,5.2447186,5.661539,6.8627696,6.9842057,7.4108725,8.01477,8.2215395,7.00718,5.924103,4.71959,3.3903592,2.2678976,2.028308,2.553436,3.2525132,3.7940516,3.9154875,3.43959,5.3431797,7.0892315,7.8145647,7.785026,8.36595,7.7259493,6.3967185,4.8738465,3.5610259,2.7470772,2.3433847,2.1103592,2.2022567,2.477949,2.481231,2.2121027,3.1770258,3.9417439,4.322462,5.408821,4.2272825,3.0490258,2.0676925,2.5928206,7.0531287,7.1515903,7.8441033,7.9885135,7.197539,5.832206,5.8847184,4.857436,6.5083084,9.26195,6.226052,6.5411286,10.217027,11.208206,8.930462,8.260923,6.311385,4.397949,4.1156926,5.612308,7.5946674,4.141949,9.750975,15.842463,16.44636,8.2215395,7.9130263,5.0084105,5.684513,10.112,12.465232,9.179898,12.120616,14.221129,13.522053,13.138052,15.494565,14.759386,11.628308,8.329846,8.608821,10.673231,8.766359,7.584821,7.8441033,6.2555904,7.686565,6.2030773,4.781949,4.824616,6.170257,8.809027,9.527796,6.9120007,2.9735386,3.1376412,2.5961027,3.0326157,3.3214362,3.0194874,2.3794873,2.5435898,2.3663592,2.15959,3.0424619,6.9645133,7.213949,7.512616,7.9130263,8.2904625,8.326565,8.139488,8.086975,6.8463597,5.0149746,5.1232824,5.35959,6.0652313,7.1122055,7.8408213,7.0531287,6.5378466,6.7282057,7.574975,9.002667,10.932513,9.019077,7.1680007,6.5378466,6.7905645,6.0750775,4.972308,4.420923,4.562052,5.169231,5.6254363,5.9536414,5.76,4.906667,3.9384618,4.089436,3.6693337,3.9122055,4.276513,4.4832826,4.529231,4.2994876,4.3618464,4.2305646,3.8301542,3.4855387,3.5380516,3.5511796,3.5511796,3.5446157,3.5446157,3.3247182,3.4133337,3.7284105,4.0500517,4.010667,4.585026,5.024821,5.1954875,4.841026,3.5807183,3.0391798,3.4855387,4.128821,4.4340515,4.1058464,3.8301542,3.5741541,3.636513,3.826872,3.446154,3.69559,3.7874875,3.7349746,3.5807183,3.4133337,3.186872,3.1015387,3.3936412,3.8006158,3.5446157,3.8400004,4.2305646,4.3552823,4.4274874,5.2381544,6.114462,6.9087186,6.6560006,5.4383593,4.391385,4.397949,4.276513,4.634257,5.474462,6.2227697,5.031385,7.4141545,11.474052,13.991385,10.43036,7.9786673,9.31118,19.702156,30.119387,17.207796,9.810052,8.500513,8.966565,9.83959,12.691693,13.075693,13.046155,12.416001,11.37559,10.496001,12.3076935,13.620514,14.401642,14.887385,15.599591,14.358975,13.827283,13.794462,14.263796,15.435489,13.912617,13.702565,13.712411,13.659899,14.089848,13.4400015,13.5778475,13.666463,13.499078,13.495796,13.062565,13.633642,14.050463,14.080001,14.404924,14.674052,15.028514,14.729847,13.820719,13.105232,14.41477,15.954053,17.096207,17.618053,17.723078,17.562258,16.889437,16.571077,16.472616,15.442053,14.769232,16.305231,18.927591,21.054361,20.634258,21.162668,21.819078,22.711796,22.882463,20.325745,19.603693,19.961437,19.587284,18.628925,19.160616,19.429745,19.620104,19.538054,19.163898,18.6519,17.828104,17.385027,16.932104,16.531694,16.692514,16.052513,15.622565,15.642258,16.098463,16.722052,16.91241,16.708925,16.850052,17.286566,17.19795,20.772104,20.059898,17.69354,14.959591,11.802258,13.02318,13.801026,14.588719,15.396104,15.803078,16.233027,17.536001,18.881643,19.239386,17.362053,17.621334,15.540514,13.689437,13.315283,14.332719,15.251694,15.977027,15.898257,15.126975,14.496821,14.506668,13.827283,12.750771,11.713642,11.300103,0.6170257,0.60389745,0.512,0.512,0.62030774,0.7187693,0.764718,0.8763078,0.84348726,0.69579494,0.69579494,0.9878975,1.1027694,1.1585642,1.2635899,1.5195899,1.5753847,1.4933335,1.4867693,1.6443079,1.9298463,2.3860514,2.9111798,3.9318976,4.95918,4.588308,3.9680004,3.7776413,3.767795,3.9253337,4.457026,4.493129,4.4734364,4.3749747,4.348718,4.7294364,4.585026,4.568616,4.8672824,5.3037953,5.3431797,6.806975,7.9327188,8.372514,8.162462,7.7390776,7.532308,8.146052,8.4053335,7.9917955,7.456821,7.6570263,8.27077,9.268514,10.502565,11.720206,12.721231,13.02318,12.855796,12.337232,11.45436,10.722463,11.08677,12.343796,13.860104,14.565744,15.931078,16.036104,15.136822,13.850258,13.1872835,13.407181,11.825232,10.5780525,10.381129,10.518975,10.289231,10.614155,10.788103,10.817642,11.418258,11.904001,12.268309,12.521027,12.681848,12.770463,13.971693,14.536206,15.074463,15.648822,15.737437,15.573335,15.340309,14.92677,14.55918,14.808617,14.227694,13.817437,13.564719,13.275898,12.583385,12.3076935,12.658873,13.367796,13.879796,13.37436,12.973949,12.675283,12.744206,12.928001,12.461949,12.563693,12.425847,12.304411,12.100924,11.35918,9.974154,9.737847,10.059488,10.735591,11.972924,12.461949,11.910565,11.122872,10.604308,10.551796,10.962052,11.414975,12.343796,13.682873,14.867694,15.694771,14.949745,14.49354,15.130258,16.610462,16.567797,16.049232,15.858873,15.996719,15.648822,16.544823,16.935387,17.910154,19.456001,20.427488,21.303797,20.844309,19.492104,18.290873,18.898052,19.744822,20.821335,22.196514,23.013746,21.48759,21.38913,21.014977,20.09272,18.806156,17.778873,18.773335,19.236105,19.239386,18.428719,16.022976,14.290052,14.454155,15.638975,16.426668,14.864411,13.659899,11.930258,10.43036,9.69518,10.023385,12.025436,12.964104,12.855796,12.015591,11.040821,10.341744,10.41395,10.482873,10.269539,10.010257,9.334154,8.628513,8.448001,8.825437,9.271795,8.953437,8.592411,8.356103,8.329846,8.513641,9.032206,9.842873,10.276103,9.783795,7.936001,7.860513,9.6295395,11.296822,11.733335,10.6469755,8.904206,9.337437,10.06277,9.915077,8.444718,7.200821,6.5378466,6.948103,7.6110773,6.4000006,6.2687182,7.4732313,8.766359,9.366975,8.976411,9.416205,9.009232,8.677744,8.677744,8.605539,8.149334,7.1876926,6.5805135,6.2588725,5.2315903,6.163693,6.229334,6.4590774,7.1680007,7.962257,7.3386674,7.785026,8.835282,9.563898,8.582564,8.848411,9.396514,9.800206,9.816616,9.3768215,10.417232,10.30236,10.33518,10.394258,8.960001,7.6307697,7.7948723,8.155898,7.9195905,6.813539,6.8693337,5.910975,4.263385,2.9013336,3.4297438,4.4110775,4.8836927,5.1265645,5.1856413,4.844308,4.007385,2.9440002,2.2153847,1.910154,1.657436,2.0709746,2.477949,2.231795,1.4802053,1.1716924,0.81394875,0.6301539,0.6498462,0.81066674,0.94523084,1.142154,0.72861546,1.4506668,3.6791797,6.426257,8.2215395,5.146257,4.2469745,7.0793853,9.714872,7.259898,6.0028725,6.4000006,6.678975,2.8553848,1.3193847,0.9878975,1.1158975,1.3718976,1.8445129,1.3817437,1.7723079,1.6738462,0.8960001,0.4004103,0.19364104,0.11158975,0.09189744,0.12143591,0.23958977,0.17394873,0.15097436,0.18379489,0.19692309,0.0,0.25271797,0.74830776,1.3423591,1.9232821,2.409026,3.2196925,4.818052,5.8781543,6.183385,6.6494365,7.174565,7.4929237,7.680001,7.5979495,6.9152827,7.0400004,6.954667,6.432821,6.0324106,7.1089234,6.38359,7.0465646,8.500513,9.419488,7.762052,9.255385,11.329642,12.360206,12.209231,12.209231,10.738873,10.8537445,11.290257,11.260718,10.476309,11.050668,11.424822,12.406155,13.5318985,13.088821,12.458668,11.493745,10.889847,10.683078,10.243283,9.176616,9.672206,10.059488,9.90195,10.023385,9.55077,9.429334,8.973129,7.8473854,6.0849237,6.157129,5.5893335,5.356308,5.9667697,7.456821,8.139488,7.650462,7.79159,8.457847,7.6603084,5.7501545,3.698872,2.1956925,1.5195899,1.5327181,2.156308,2.7109745,3.2164104,3.5610259,3.4921029,4.381539,5.3202057,6.0160003,6.7807183,8.52677,7.7981544,6.3606157,4.886975,3.8465643,3.501949,3.0162053,2.2121027,1.8215386,1.9462565,2.041436,1.6311796,2.4385643,3.498667,4.4832826,5.6943593,5.156103,3.7973337,3.9680004,5.4383593,5.398975,5.106872,6.5739493,7.906462,8.195283,7.515898,7.273026,7.145026,7.830975,9.120821,9.882257,8.933744,10.407386,10.886565,9.688616,8.858257,6.4722056,4.854154,5.612308,7.768616,7.765334,3.2623591,9.465437,15.796514,15.163078,3.9351797,5.9995904,6.8233852,7.1056414,7.171283,7.000616,6.961231,12.274873,15.31077,14.464001,14.148924,17.401438,17.447386,14.598565,10.752001,9.380103,10.417232,8.155898,7.79159,9.760821,9.764103,8.549745,8.113232,7.4174366,6.117744,4.5489235,7.6274877,7.250052,5.287385,3.3509746,2.809436,3.170462,2.9801028,3.7054362,4.57518,2.556718,1.8412309,2.034872,3.0916924,4.460308,5.07077,6.226052,6.705231,7.0334363,7.5421543,8.3823595,7.312411,7.256616,6.7872825,5.76,5.3234878,5.7435904,6.701949,7.4732313,7.79159,7.857231,6.3507695,5.5007186,5.7435904,7.1089234,9.209436,7.529026,6.4623594,6.2227697,6.226052,5.0871797,4.4274874,4.332308,4.601436,5.1922054,6.2162056,6.3179493,5.8814363,4.778667,3.5282054,3.2754874,2.7634873,2.7109745,3.0752823,3.6102567,3.8728209,3.9187696,3.9942567,3.9154875,3.5872824,3.006359,2.9210258,2.9801028,2.9472823,2.8521028,2.993231,3.006359,2.865231,2.8160002,3.0391798,3.6660516,4.2436924,4.923077,5.10359,4.571898,3.4921029,3.2656412,3.5511796,3.9811285,4.2535386,4.1222568,3.692308,3.3936412,3.5249233,3.7842054,3.2820516,3.2131286,3.114667,3.1507695,3.2787695,3.2525132,3.114667,2.9111798,2.92759,3.0982566,3.0326157,3.2131286,3.436308,3.7973337,4.4734364,5.7140517,5.789539,6.3540516,6.4590774,5.7468724,4.453744,4.95918,5.0838976,5.284103,5.5762057,5.540103,4.519385,6.4656415,8.644924,9.55077,8.891078,6.688821,10.348309,26.020105,39.712822,17.289848,9.747693,9.997129,10.292514,9.202872,11.634872,12.20595,13.026463,12.803283,11.61518,10.893129,11.641437,12.760616,13.751796,14.201437,13.778052,12.448821,12.27159,12.918155,13.896206,14.575591,13.827283,13.243078,12.750771,12.550565,13.111795,12.521027,13.078976,13.692719,13.810873,13.446565,13.019898,13.226667,13.528616,13.774771,14.214565,13.791181,13.413745,13.400617,13.571283,13.24636,13.410462,14.880821,16.187078,16.78113,17.027283,17.220924,16.718771,16.315079,16.075489,15.346873,15.2155905,16.856617,19.121233,20.407797,18.678156,18.848822,20.145233,20.696617,19.70872,17.480206,20.148514,21.195488,20.25354,18.36636,17.962667,17.929848,17.99877,18.054565,18.097233,18.225233,17.70995,17.184822,16.272411,15.284514,15.218873,14.119386,13.8765135,14.5263605,15.629129,16.275694,16.088617,15.589745,15.228719,15.097437,14.920206,16.452925,16.265848,15.563488,14.693745,13.154463,13.495796,14.194873,15.176207,15.996719,15.835898,15.688207,17.660719,18.953848,18.340103,16.167385,16.518566,14.923489,13.423591,13.387488,15.520822,16.17395,15.894976,16.154257,16.521847,14.674052,15.126975,14.78236,13.338258,11.500309,10.965334,0.77456415,0.5874872,0.5218462,0.574359,0.7089231,0.8763078,0.79425645,0.90912825,0.9321026,0.8402052,0.8467693,1.020718,1.204513,1.4145643,1.6771283,2.044718,1.782154,1.5688206,1.5556924,1.7690258,2.1103592,2.4024618,3.006359,3.7973337,4.4898467,4.6605134,4.1846156,3.8137438,3.620103,3.7349746,4.3552823,4.9296412,4.6966157,4.565334,4.775385,4.8836927,4.378257,4.3552823,4.699898,5.2381544,5.7403083,6.6395903,7.387898,7.719385,7.716103,7.8014364,8.3593855,8.92718,8.874667,8.310155,8.064001,8.329846,8.769642,9.475283,10.450052,11.611898,12.301129,12.327386,12.064821,11.605334,10.774975,10.312206,10.502565,11.54954,13.098668,14.230975,15.737437,15.872002,15.140103,14.194873,13.833847,13.4170265,12.06154,11.237744,11.208206,11.063796,10.397539,10.896411,11.283693,11.346052,11.926975,12.150155,12.340514,12.402873,12.360206,12.356924,14.158771,15.130258,15.835898,16.42995,16.646564,16.338053,15.885129,15.27795,14.706873,14.555899,14.41477,14.342566,14.076719,13.653335,13.4170265,13.131488,13.236514,13.620514,13.889642,13.354668,12.586668,11.920411,11.71036,11.88759,11.959796,12.327386,12.386462,12.566976,12.747488,12.242052,11.372309,11.008,10.8767185,11.008,11.746463,12.514462,12.281437,11.61518,10.988309,10.765129,11.008,11.720206,12.970668,14.575591,16.108309,16.278976,14.6642065,13.791181,14.447591,15.701335,16.36431,16.059078,15.494565,14.956308,14.299898,14.795488,15.192616,16.167385,17.604925,18.57313,19.994259,19.91877,18.993233,17.992207,17.811693,18.090668,19.449438,21.664822,23.35508,21.999592,20.78195,20.004105,19.19672,18.432001,18.33354,18.937437,18.947283,19.055592,18.724104,16.210052,14.168616,13.426873,14.227694,15.540514,15.048206,13.6697445,11.933539,10.827488,10.742155,11.477334,12.668719,13.344822,13.069129,12.100924,11.395283,10.857026,10.656821,10.676514,10.765129,10.71918,10.164514,9.609847,9.344001,9.45559,9.833026,9.544206,9.465437,9.645949,9.77395,9.16677,9.747693,10.709334,11.421539,11.250873,9.5606165,8.280616,9.189744,10.499283,10.889847,9.531077,7.7325134,7.8539495,8.320001,8.100103,6.698667,6.7150774,6.4754877,6.9710774,7.6012316,6.186667,6.0061545,7.213949,8.5891285,9.3078985,8.969847,9.481847,9.386667,8.976411,8.55959,8.464411,8.04759,7.250052,6.7905645,6.5345645,5.504,6.012718,6.124308,6.38359,7.000616,7.8506675,7.509334,7.4010262,8.123077,9.078155,8.464411,8.379078,8.277334,8.260923,8.356103,8.523488,9.508103,9.737847,9.990565,10.118565,9.032206,7.571693,7.515898,7.1647186,6.229334,5.8256416,6.498462,5.8125134,4.4274874,3.242667,3.4067695,3.495385,3.436308,4.568616,6.1308722,5.277539,4.342154,3.0326157,2.0151796,1.5360001,1.4145643,2.2449234,2.7076926,2.3236926,1.4506668,1.2931283,1.4145643,0.88287187,0.636718,0.94523084,1.3981539,1.6902566,1.7296412,2.5173335,4.138667,5.7796926,6.4754877,4.2929235,2.9702566,3.9548721,6.419693,4.785231,6.091488,8.034462,8.438154,5.2480006,1.6213335,0.8369231,0.9517949,1.0732309,1.3686155,1.4244103,2.1924105,2.048,0.9485129,0.44307697,0.190359,0.1148718,0.08861539,0.0951795,0.2100513,0.0951795,0.23302566,0.38728207,0.39712822,0.15753847,1.0272821,1.9331284,2.733949,3.367385,3.8432825,3.1967182,3.698872,4.1025643,4.6080003,6.8496413,7.138462,7.4141545,7.686565,7.4765134,5.8486156,6.2555904,6.485334,6.2720003,6.2096415,7.765334,8.257642,8.579283,8.231385,7.384616,6.8693337,10.902975,12.045129,11.867898,11.749744,12.875488,10.709334,10.86359,11.113027,10.656821,10.098872,10.496001,10.5780525,11.378873,12.550565,12.393026,12.465232,11.497026,10.555078,9.911796,9.035488,9.124104,9.278359,9.504821,9.872411,10.505847,9.393231,9.048616,8.4053335,7.2927184,6.452513,7.1581545,6.304821,5.8945646,6.51159,7.3321033,8.54318,7.860513,7.4043083,7.6767187,7.581539,5.159385,2.9046156,1.591795,1.339077,1.6114873,2.1497438,2.4582565,2.8521028,3.3312824,3.5938463,3.9844105,4.2141542,4.7524104,5.989744,8.257642,7.640616,6.4065647,5.1364107,4.2896414,4.194462,3.7087183,2.6190772,1.9561027,1.9790771,2.1891284,1.7296412,1.8937438,2.7273848,4.1452312,5.914257,5.717334,5.179077,6.1341543,7.509334,5.3005133,5.9470773,6.2884107,6.7544622,7.1647186,6.7117953,7.4469748,8.024616,8.65477,9.4916935,10.620719,9.288206,9.95118,9.242257,7.0432825,6.485334,7.394462,8.27077,9.114257,9.281642,7.463385,3.2131286,9.396514,13.3940525,10.341744,3.121231,7.2172313,10.8307705,10.722463,8.018052,8.178872,8.5202055,12.432411,14.083283,12.708103,12.586668,13.095386,13.272616,12.25518,10.348309,9.032206,9.964309,9.317744,9.32759,10.394258,11.07036,8.805744,9.153642,9.701744,8.493949,4.017231,6.0783596,5.2480006,4.263385,3.9417439,3.190154,3.5413337,2.7995899,3.4691284,4.84759,3.0162053,1.4244103,2.156308,4.1682053,5.536821,3.4855387,5.0543594,5.937231,6.47877,6.997334,7.8080006,7.3025646,6.997334,6.6034875,6.1046157,5.756718,6.419693,7.138462,7.3649235,7.259898,7.706257,6.482052,4.854154,4.2174363,5.031385,6.810257,5.543385,5.080616,5.031385,4.926359,4.201026,3.8564105,4.315898,4.821334,5.3366156,6.5706673,6.925129,6.2490263,4.97559,3.6758976,3.0654361,2.484513,2.1891284,2.3926156,2.92759,3.239385,3.6594875,3.757949,3.7185643,3.5347695,2.986667,2.6322052,2.5632823,2.4746668,2.428718,2.8356924,2.5698464,2.2383592,2.1202054,2.412308,3.239385,3.7874875,4.4996924,4.775385,4.4800005,3.9351797,3.9581542,3.9089234,3.8596926,3.889231,4.086154,3.3772311,3.2000003,3.259077,3.239385,2.806154,2.6847181,2.6551797,2.8258464,3.0884104,3.117949,2.9538465,2.6683078,2.4451284,2.3794873,2.4648206,2.7109745,2.930872,3.623385,4.775385,5.8847184,5.47118,5.543385,5.5729237,5.3136415,4.8049235,5.5105643,5.612308,5.546667,5.356308,4.6900516,3.8071797,5.35959,6.166975,5.940513,7.27959,6.0652313,9.787078,24.684309,37.569645,15.835898,9.616411,10.781539,11.178667,9.409642,10.840616,11.145847,12.212514,12.310975,11.211488,10.167795,10.394258,11.680821,12.786873,13.02318,12.258463,11.040821,11.477334,12.530872,13.407181,13.548308,12.852514,12.773745,12.737642,12.553847,12.409437,11.713642,12.511181,13.259488,13.3251295,12.970668,12.560411,12.675283,13.174155,13.830565,14.342566,14.063591,12.895181,12.461949,12.987078,13.285745,12.790154,14.17518,15.369847,15.803078,16.423386,16.403694,16.233027,15.908104,15.55036,15.409232,15.924514,17.060104,18.258053,18.579693,16.705643,16.754873,18.244925,18.6519,17.47036,16.200207,19.02277,20.447182,20.089437,18.635489,17.814976,18.110361,17.926565,17.870771,18.130053,18.474669,17.670565,16.951796,16.022976,15.012104,14.486976,13.22995,13.115078,13.958565,15.100719,15.432206,14.818462,14.093129,13.787898,13.929027,14.070155,14.815181,14.815181,14.41477,13.948719,13.781334,13.692719,14.070155,14.956308,15.724309,15.113848,14.900514,17.11918,18.136618,16.807386,14.470565,14.683899,13.899488,13.197129,13.5778475,15.96718,16.584206,16.246155,16.836924,17.578669,15.031796,15.117129,14.690463,13.13477,11.076924,10.417232,0.7778462,0.6235898,0.58092314,0.67938465,0.8566154,0.97805136,0.8566154,1.0502565,1.1257436,1.0338463,1.1126155,1.1881026,1.5130258,1.8445129,2.1070771,2.3696413,1.7460514,1.6443079,1.7624617,2.0250258,2.553436,2.2186668,2.917744,3.5183592,3.751385,4.1846156,4.197744,3.626667,3.3509746,3.5183592,3.5249233,4.5817437,4.706462,4.8344617,5.10359,4.8311796,4.565334,4.4077954,4.821334,5.7140517,6.422975,6.672411,6.9645133,6.9349747,6.8594875,7.650462,9.206155,9.577026,9.386667,8.996103,8.513641,8.490667,8.858257,9.094564,9.255385,10.003693,10.620719,10.771693,10.597744,10.171078,9.508103,10.006975,10.499283,11.303386,12.547283,14.158771,14.8250265,14.516514,14.053744,13.869949,14.04718,12.763899,11.999181,11.815386,11.825232,11.221334,10.6469755,11.634872,12.373334,12.297847,12.11077,12.2157955,12.051693,11.936821,12.137027,12.875488,14.680616,15.826053,16.682669,17.289848,17.365335,16.948515,16.597334,15.9573345,15.117129,14.605129,14.989129,14.998976,14.385232,13.659899,14.106257,14.004514,13.761642,13.620514,13.558155,13.269335,12.566976,11.940104,11.631591,11.611898,11.588924,12.015591,12.406155,13.013334,13.643488,13.659899,13.321847,12.383181,11.536411,11.145847,11.247591,12.058257,12.406155,12.3995905,12.1698475,11.851488,11.995898,12.678565,13.840411,15.481437,17.686975,16.695797,15.24513,14.670771,15.113848,15.537232,16.804104,17.401438,17.007591,15.839181,14.631386,14.198155,13.515489,13.827283,15.012104,15.602873,16.57436,16.987898,17.293129,17.414566,16.764719,16.725334,17.870771,19.492104,20.841026,21.139694,21.257847,20.880411,20.230566,19.662771,19.649643,18.504206,18.01518,18.110361,18.185848,17.06995,15.852309,14.011078,12.816411,12.626052,12.885334,11.329642,10.381129,10.512411,11.638155,13.131488,13.243078,13.748514,13.223386,11.779283,11.0375395,10.929232,10.729027,10.81436,11.18195,11.451077,11.155693,10.866873,10.476309,10.184206,10.486155,10.633847,10.850462,11.34277,11.556104,10.157949,10.098872,10.338462,10.673231,10.893129,10.794667,9.521232,9.613129,10.210463,10.217027,8.310155,6.1505647,5.661539,5.9503593,6.3310776,6.3212314,6.5280004,6.626462,6.987488,7.2205133,6.1768208,6.2884107,7.0334363,8.323282,9.498257,9.350565,9.347282,9.544206,9.209436,8.316719,7.5454364,7.177847,6.6461544,6.5411286,6.741334,6.4065647,6.38359,6.5312824,6.7183595,7.0925136,8.096821,8.3593855,7.6635904,7.522462,8.060719,8.021334,7.9425645,7.315693,6.941539,7.0334363,7.240206,8.1755905,9.065026,9.386667,9.127385,8.763078,7.571693,6.9710774,6.265436,5.4547696,5.2315903,5.044513,4.637539,4.2338467,3.7284105,2.6715899,2.6026669,4.466872,7.890052,10.522257,8.064001,6.567385,4.3027697,2.349949,1.3357949,1.401436,2.176,2.4320002,2.3105643,2.097231,2.2416413,2.5764105,1.4998976,0.90912825,1.3456411,1.9823592,2.162872,3.3214362,3.318154,2.4648206,3.511795,2.9538465,2.9997952,2.349949,1.1191796,0.8336411,1.8674873,5.4514875,7.3058467,6.8627696,7.256616,1.657436,0.62030774,0.88287187,0.90584624,0.8795898,1.654154,2.2547693,1.8215386,0.7056411,0.4955898,0.2297436,0.101743594,0.04594872,0.032820515,0.068923086,0.20020515,0.40369233,0.5021539,0.49230772,0.5481026,2.3663592,4.06318,4.5554876,4.086154,4.2502565,2.3105643,3.0949745,4.535795,5.61559,6.3573337,6.186667,6.9152827,8.057437,8.303591,5.5204105,5.2315903,5.32677,5.3431797,5.3103595,5.72718,9.741129,10.249847,8.434873,6.445949,7.427283,12.882052,13.065847,11.841642,11.45436,12.527591,10.466462,10.843898,10.883283,10.082462,10.240001,9.609847,9.645949,10.469745,11.503591,11.493745,11.753027,11.211488,10.115283,8.881231,8.113232,8.769642,8.891078,9.219283,9.944616,10.7158985,9.275078,8.530052,7.4732313,6.294975,6.3901544,7.2205133,6.547693,6.491898,7.276308,7.253334,8.149334,8.004924,7.2927184,6.6395903,6.8266673,4.2371287,2.412308,1.5163078,1.4145643,1.6869745,1.9265642,2.100513,2.605949,3.2886157,3.4494362,3.945026,4.059898,4.532513,5.7698464,7.857231,6.9776416,6.042257,5.172513,4.588308,4.601436,4.069744,3.0916924,2.359795,2.156308,2.3696413,2.2088206,1.9200002,2.2580514,3.5511796,5.7009234,5.943795,6.7905645,7.2664623,6.928411,5.861744,8.257642,7.8047185,6.9152827,6.3179493,5.0543594,8.277334,7.207385,8.096821,10.712616,8.356103,7.9294367,10.433641,9.426052,5.1331286,4.417641,9.878975,12.379898,11.300103,8.205129,6.8627696,4.397949,9.796924,10.052924,4.594872,5.3070774,9.153642,12.980514,12.186257,9.032206,12.642463,12.868924,14.14236,14.122667,12.425847,10.630565,8.608821,7.893334,7.4075904,7.2237954,8.562873,8.717129,10.003693,10.712616,10.04636,8.109949,7.712821,8.228104,10.262975,11.434668,6.38359,5.093744,4.647385,4.663795,4.663795,4.082872,3.2984617,2.5698464,2.5928206,3.062154,2.6584618,1.3751796,2.5862565,4.33559,5.080616,3.6627696,4.5489235,5.8190775,6.8594875,7.315693,7.0957956,8.083693,7.6603084,6.6822567,5.914257,6.0192823,7.056411,7.4174366,7.387898,7.210667,7.0957956,6.813539,5.297231,4.135385,4.125539,5.2644105,4.6112823,3.9909747,3.6660516,3.748103,4.204308,3.876103,4.670359,5.3891287,5.8223596,6.7544622,7.6143594,6.744616,5.4514875,4.388103,3.5347695,3.0293336,2.6354873,2.556718,2.7437952,2.8816411,3.5380516,3.754667,3.8465643,3.8465643,3.495385,2.809436,2.3893335,2.1530259,2.1891284,2.737231,2.0151796,1.6902566,1.7624617,2.1398976,2.6354873,3.255795,3.876103,4.2535386,4.345436,4.2896414,4.2371287,4.1813335,4.0041027,3.8038976,3.879385,3.1277952,3.0030773,2.9210258,2.6387694,2.2613335,2.2547693,2.3335385,2.5796926,2.878359,2.917744,2.5993848,2.300718,2.0644104,1.9790771,2.162872,2.5238976,2.8849232,3.7448208,4.8640003,5.284103,5.2447186,5.0674877,4.7261543,4.519385,5.110154,5.664821,5.477744,5.1331286,4.854154,4.4996924,3.8400004,4.6211286,5.0838976,5.146257,6.3967185,6.8463597,7.817847,16.479181,26.450054,17.80513,9.744411,10.06277,11.155693,10.499283,10.660104,9.724719,10.43036,10.676514,9.816616,8.651488,8.848411,10.535385,11.805539,12.120616,12.320822,10.896411,11.697231,12.626052,12.895181,13.026463,11.661129,12.27159,13.115078,13.292309,12.737642,11.684103,12.35036,12.829539,12.566976,12.35036,11.881026,12.570257,13.7386675,14.690463,14.726565,15.392821,13.988104,12.727796,12.514462,12.937847,12.750771,13.696001,14.385232,14.690463,15.740719,15.2155905,14.995693,14.841437,14.818462,15.281232,16.377438,17.112617,17.211079,16.521847,15.038361,14.930053,15.82277,16.105026,15.645539,15.77354,16.324924,17.972515,19.213129,19.383797,18.642054,19.190155,18.799591,18.438566,18.438566,18.507488,17.391592,16.784412,16.295385,15.66195,14.739694,14.011078,13.755078,14.201437,14.874257,14.598565,13.860104,12.921437,12.517745,12.86236,13.650052,15.14995,15.29436,14.424617,13.380924,13.492514,13.590976,13.453129,13.856822,14.486976,13.932309,14.171899,15.616001,16.141129,15.015386,12.898462,13.193847,13.512206,13.715693,14.086565,15.333745,16.725334,17.332514,17.450668,16.787693,14.464001,14.424617,13.63036,12.114052,10.482873,9.941334,0.3511795,0.508718,0.4955898,0.6104616,0.761436,0.44307697,0.8566154,1.3456411,1.4736412,1.2832822,1.2964103,1.2832822,1.4834872,1.6836925,1.7985642,1.847795,1.4080001,2.1103592,2.8127182,3.0785644,3.190154,2.6387694,2.9965131,3.2525132,3.367385,4.2568207,4.1846156,4.1747694,4.5587697,5.0149746,4.562052,5.405539,5.4580517,4.893539,4.20759,4.2568207,4.8804107,5.4186673,6.0061545,6.3868723,5.937231,6.8397956,7.4863596,7.4141545,6.8562055,6.7610264,7.5520005,7.778462,8.805744,10.161232,9.55077,9.626257,9.140513,8.89436,9.186462,9.796924,10.834052,10.817642,10.233437,9.521232,9.094564,9.924924,10.607591,11.585642,12.76718,13.548308,13.892924,13.590976,13.197129,13.193847,14.024206,13.02318,13.164309,13.285745,13.016617,12.770463,12.882052,13.476104,13.200411,12.097642,11.595488,12.071385,12.045129,12.619488,13.948719,15.241847,15.622565,16.118155,16.594053,16.948515,17.11918,16.315079,16.150976,16.12472,15.911386,15.350155,16.633438,16.676104,15.872002,14.726565,13.88636,13.971693,13.29559,12.3076935,11.523283,11.536411,12.708103,13.128206,12.87877,12.087796,10.939077,11.96636,12.973949,13.974976,14.647796,14.342566,13.978257,12.612924,11.45436,11.067078,11.382154,12.068104,12.11077,12.475078,13.184001,13.305437,13.866668,14.25395,14.657642,15.540514,17.637745,17.322668,17.050259,17.611488,18.405745,17.440823,18.697847,19.67918,19.111385,17.316103,16.20349,16.338053,14.421334,13.384206,13.797745,13.869949,13.735386,14.306462,14.903796,15.067899,14.54277,15.225437,16.20349,17.001026,17.624617,18.54031,20.115694,20.883694,21.028105,20.627693,19.636515,18.208822,17.302977,16.692514,16.459488,16.984617,16.07877,14.280207,12.698257,11.920411,11.992617,10.761847,9.819899,10.026668,11.460924,13.413745,14.217847,15.00554,14.55918,13.065847,12.100924,11.513436,12.327386,13.190565,13.206975,11.963078,12.304411,12.225642,11.542975,10.643693,10.499283,11.487181,11.155693,11.621744,12.685129,11.85477,10.71918,9.586872,8.940309,8.595693,7.706257,7.975385,8.966565,9.974154,10.128411,8.408616,6.6494365,5.7632823,5.622154,6.160411,7.3714876,6.11118,5.9995904,6.189949,6.12759,5.5532312,6.311385,6.8299494,7.702975,8.887795,9.705027,9.984001,9.764103,9.110975,8.155898,7.0793853,6.2752824,5.6320004,5.7665644,6.4557953,6.636308,6.8693337,7.0367184,6.76759,6.6067696,8.011488,8.891078,7.827693,7.017026,7.0793853,7.0793853,6.885744,6.2588725,6.2096415,6.8955903,7.6307697,8.411898,9.347282,9.156924,7.968821,7.3091288,5.504,4.9329233,4.9493337,5.07077,4.97559,4.1452312,4.5128207,4.525949,3.501949,1.6311796,3.0490258,11.139283,16.38072,15.570052,11.808822,9.124104,5.651693,2.7109745,1.083077,1.024,1.1815386,1.3587693,1.9626669,2.9013336,3.5872824,3.7316926,2.294154,1.8904617,2.861949,3.2656412,1.8248206,3.8367183,4.141949,3.4756925,8.467693,3.0358977,1.5130258,1.0732309,0.56451285,0.5021539,1.4309745,7.5487185,8.52677,4.4734364,5.9503593,1.3357949,0.38400003,0.45292312,0.40369233,0.6104616,2.3926156,2.7470772,1.6902566,0.2986667,0.702359,0.4955898,0.17723078,0.0,0.032820515,0.16738462,0.571077,0.58092314,0.4397949,0.48902568,1.1585642,4.0402055,7.030154,5.651693,1.2603078,1.0535386,1.8937438,5.7403083,6.5345645,4.0008206,3.6463592,3.817026,4.8311796,6.0028725,6.2884107,4.2863593,3.5314875,2.9210258,2.9636924,3.5807183,4.1058464,7.2172313,7.9491286,6.0685134,4.069744,7.171283,13.298873,12.596514,10.9915905,11.158976,12.527591,9.596719,9.416205,9.938052,10.28595,10.725744,9.383386,9.91836,10.509129,10.564924,10.712616,11.713642,11.395283,10.059488,8.454565,7.781744,8.283898,8.306872,8.704,9.504821,9.93477,8.736821,7.9425645,6.73477,5.4383593,5.5236926,5.914257,5.901129,6.488616,7.522462,7.706257,7.5454364,7.499488,7.131898,6.498462,6.117744,3.761231,2.1300514,1.4276924,1.3587693,1.1126155,1.1881026,1.782154,2.7208207,3.498667,3.2656412,3.4133337,3.5774362,4.1517954,5.0642056,5.7829747,4.5489235,3.9220517,3.9942567,4.5522056,5.0674877,4.699898,3.9023592,2.8717952,1.9396925,1.5885129,2.4549747,2.3696413,2.4713848,3.1737437,4.1517954,6.1046157,6.665847,5.7731285,4.923077,7.1548724,5.5565133,8.828718,11.099898,10.827488,10.801231,16.905848,10.082462,6.9349747,10.614155,10.834052,8.854975,9.898667,10.417232,9.153642,7.141744,12.182976,11.136001,6.166975,1.5786668,3.8006158,6.363898,5.4482055,4.056616,3.5872824,3.8301542,5.832206,8.677744,7.1187696,3.0720003,5.5991797,14.293334,16.774565,18.021746,17.490053,9.140513,11.98277,11.119591,7.9819493,6.3179493,12.176412,6.1078978,7.056411,9.705027,9.69518,3.6168208,3.639795,4.562052,8.871386,13.915898,11.900719,4.381539,3.748103,4.969026,5.5729237,5.6451287,3.3378465,2.294154,1.6771283,1.339077,1.8149745,1.657436,2.231795,2.0545642,2.0250258,5.431795,4.9329233,6.242462,7.9524107,8.717129,7.27959,8.267488,8.339693,7.650462,6.8594875,7.141744,7.4469748,7.6701546,7.9819493,8.083693,7.2172313,6.9842057,6.2851286,4.900103,3.6036925,4.164923,5.4482055,4.6145644,3.8400004,4.1550775,5.4613338,5.2315903,5.786257,6.419693,6.803693,6.9743595,7.3747697,6.7249236,6.0061545,5.32677,3.9351797,3.9614363,3.6726158,3.2820516,3.0260515,3.1737437,4.210872,4.9920006,5.284103,5.031385,4.348718,3.3608208,2.4155898,1.8543591,1.9331284,2.8225644,2.5304618,2.0644104,1.9593848,2.2580514,2.5009232,3.1113849,3.6758976,4.135385,4.3027697,3.876103,3.314872,3.623385,3.8662567,3.7316926,3.5249233,3.2820516,3.0260515,2.6354873,2.2383592,2.2121027,1.9790771,1.8871796,1.972513,2.1956925,2.4418464,2.1234872,2.034872,1.9626669,1.9429746,2.2744617,2.5173335,2.9801028,3.7251284,4.3552823,4.013949,5.0871797,4.972308,4.420923,4.1222568,4.6834874,4.854154,4.962462,4.565334,4.197744,5.356308,5.024821,4.8049235,5.1232824,6.0783596,7.4469748,9.888822,8.979693,9.386667,14.450873,26.167797,8.418462,7.8473854,11.1064625,11.867898,10.817642,7.5585647,8.402052,9.366975,9.153642,9.140513,7.722667,9.449026,11.260718,12.173129,13.259488,10.781539,10.528821,11.510155,12.5374365,12.20595,11.644719,12.035283,12.836103,13.590976,13.945437,12.2387705,12.324103,13.019898,13.436719,12.983796,12.251899,13.423591,15.816206,17.765745,16.633438,17.558975,16.12472,14.805334,14.572309,14.87754,14.194873,13.00677,12.11077,12.0549755,13.154463,13.312001,12.721231,13.298873,14.890668,15.24513,16.866463,17.831387,17.555695,16.17395,14.5263605,14.368821,14.089848,13.804309,13.856822,14.8480015,15.799796,17.24718,19.18031,20.62113,19.606976,18.875078,18.14318,17.385027,16.820515,16.905848,16.649847,16.889437,16.626873,15.740719,14.982565,15.192616,14.739694,14.746258,15.14995,14.710155,13.794462,12.905026,12.202667,12.002462,12.770463,14.017642,14.677335,14.217847,13.026463,12.406155,13.430155,13.24636,13.24636,13.712411,13.8075905,14.516514,14.217847,13.771488,13.4629755,12.983796,13.584412,15.425642,16.170668,15.136822,13.305437,15.91795,18.458258,17.834667,14.388514,11.88759,13.791181,12.993642,11.30995,9.954462,9.55077,0.5218462,0.62030774,0.67282057,0.7384616,0.85005134,0.9911796,1.0666667,1.1454359,1.1552821,1.142154,1.2603078,1.6771283,1.9396925,1.9265642,1.9593848,2.7995899,2.3696413,2.0873847,2.4024618,2.934154,2.4582565,2.4648206,2.9243078,3.1638978,3.1474874,3.4527183,3.5938463,3.5511796,4.0041027,4.824616,5.074052,5.8190775,6.114462,5.9569235,5.481026,4.9526157,4.8836927,5.2053337,5.674667,6.1472826,6.5837955,6.547693,6.9743595,7.322257,7.499488,7.8703594,8.018052,8.274052,8.766359,9.143796,8.562873,8.608821,8.979693,8.914052,8.717129,9.747693,10.883283,10.210463,9.216001,8.582564,8.214975,9.366975,10.614155,11.483898,11.999181,12.681848,12.4685135,12.62277,12.763899,12.905026,13.4629755,14.257232,14.454155,14.086565,13.620514,13.942155,13.39077,13.019898,12.704822,12.504617,12.658873,12.832822,13.2562065,14.034052,15.07118,16.072206,15.983591,15.593027,15.688207,16.216616,16.288822,16.256,15.970463,15.635694,15.353437,15.094155,14.76595,14.194873,13.37436,12.521027,12.07795,11.762873,11.487181,11.434668,11.877745,13.157744,13.492514,13.042872,12.406155,11.884309,11.477334,10.978462,11.145847,12.028719,13.042872,12.950975,12.750771,12.087796,11.034257,10.154668,10.492719,11.487181,12.442257,13.190565,13.7386675,14.27036,14.989129,14.720001,14.477129,14.79877,15.747283,17.227488,17.345642,18.179283,19.685745,19.698874,19.754667,20.033642,18.704412,16.613745,17.289848,16.38072,14.854566,14.309745,14.775796,14.713437,14.78236,15.222155,15.694771,15.658668,14.381949,15.632411,17.417847,18.553438,18.73395,18.527182,18.822565,18.730669,18.681437,18.41231,16.964924,15.616001,14.411489,13.817437,14.057027,15.126975,14.057027,13.636924,13.082257,12.189539,11.332924,10.834052,10.026668,9.964309,11.313231,14.339283,15.048206,14.867694,14.14236,13.541744,14.040616,13.5318985,12.872206,12.324103,11.805539,10.912822,11.52,11.848206,11.497026,10.66995,10.180923,10.916103,10.604308,10.417232,10.666668,10.794667,11.759591,12.173129,11.940104,10.965334,9.147078,8.329846,8.408616,8.3364105,7.965539,8.041026,7.466667,6.925129,6.3967185,6.0783596,6.370462,5.464616,5.8190775,6.5411286,6.820103,5.943795,6.048821,6.5050263,7.0104623,7.5454364,8.372514,8.802463,9.347282,9.133949,8.12636,7.141744,6.5805135,6.1472826,5.9569235,6.045539,6.3573337,6.5706673,6.7314878,6.8594875,7.0465646,7.4732313,8.723693,8.297027,7.702975,7.427283,6.9087186,6.1078978,6.012718,6.0849237,6.2523084,6.8955903,7.6012316,8.730257,9.015796,8.326565,7.686565,7.1023593,6.8299494,6.695385,6.298257,4.9985647,3.757949,3.7120004,4.1124105,5.7829747,11.093334,12.3536415,15.100719,14.851283,11.352616,8.598975,4.7327185,2.540308,1.5097437,1.0305642,0.37415388,0.61374366,0.72861546,1.0108719,1.3554872,1.2668719,1.1191796,1.1552821,1.9331284,3.1638978,3.7054362,4.95918,7.565129,8.812308,7.256616,2.7208207,4.1222568,6.1308722,4.5029745,0.4266667,0.5513847,3.5413337,10.473026,11.250873,5.618872,3.1803079,0.77128214,0.71548724,0.7384616,0.24287182,0.29210258,1.0699488,0.99774367,0.82379496,0.8730257,1.0305642,0.62030774,0.21989745,0.01969231,0.07876924,0.3511795,0.8992821,1.142154,1.1191796,1.2964103,2.5632823,4.644103,3.7349746,2.048,0.9714873,1.0765129,2.4188719,3.2229745,3.7087183,3.9187696,3.7316926,4.644103,4.5489235,4.5522056,4.6112823,3.5052311,4.194462,3.2951798,2.4188719,2.2908719,2.737231,4.844308,6.432821,5.668103,4.6178465,9.222565,12.626052,13.036308,12.501334,11.923694,11.073642,10.223591,10.482873,10.633847,10.509129,10.95877,10.387693,10.397539,10.289231,10.427077,12.212514,12.278154,11.300103,9.557334,8.064001,8.562873,8.848411,8.461129,8.192,8.421744,9.104411,8.553026,6.9743595,5.61559,4.9920006,4.900103,5.106872,5.464616,6.052103,6.695385,6.9842057,7.450257,7.250052,6.4032826,5.5072823,5.7632823,3.6135387,2.2383592,1.585231,1.467077,1.5524104,1.7427694,2.1333334,2.7076926,3.3476925,3.8400004,4.4832826,4.076308,4.1485133,4.8607183,5.0149746,4.1517954,4.092718,4.5456414,4.9788723,4.6145644,4.1714873,3.9680004,3.3608208,2.4418464,2.038154,2.3958976,2.8455386,3.626667,4.342154,3.9417439,5.858462,6.2687182,5.668103,5.330052,7.3386674,10.358154,11.270565,9.370257,6.6494365,7.77518,9.682052,7.5421543,6.422975,7.138462,6.245744,9.842873,8.625232,9.140513,11.175385,7.762052,7.200821,5.792821,4.9821544,5.428513,6.997334,7.207385,5.080616,4.2601027,4.8836927,3.5741541,3.9745643,4.338872,4.017231,3.751385,5.674667,7.2172313,9.340718,11.168821,12.934566,16.000002,13.90277,9.908514,7.3025646,7.6143594,10.601027,5.648411,6.629744,9.334154,10.70277,8.851693,9.570462,6.1407185,4.5128207,5.8289237,6.419693,4.457026,4.493129,5.211898,5.080616,2.349949,3.3936412,5.428513,6.088206,4.699898,2.2678976,4.20759,2.6256413,1.394872,2.2711797,4.893539,5.4875903,6.518154,7.430565,7.857231,7.6077952,6.994052,6.9743595,6.7938466,6.0750775,4.8344617,5.2676926,6.114462,6.701949,6.925129,7.2303596,7.213949,7.072821,6.2687182,5.097026,4.70318,5.7107697,5.543385,4.9460516,4.663795,5.4153852,5.8157954,6.4722056,6.6395903,6.5936418,7.643898,7.5585647,6.8463597,6.2227697,5.756718,4.8640003,4.5095387,4.2863593,3.9154875,3.5446157,3.761231,4.201026,4.0434875,3.7743592,3.7448208,4.1550775,3.515077,3.0129232,2.5304618,2.156308,2.1891284,2.2580514,1.8937438,1.7460514,1.8970258,1.8674873,1.9396925,2.481231,3.1737437,3.7284105,3.876103,3.2164104,3.2525132,3.4855387,3.7415388,4.1583595,3.5840003,2.8947694,2.284308,1.8576412,1.6377437,1.3095386,1.2635899,1.6771283,2.2153847,2.0512822,1.654154,1.7591796,1.9790771,2.162872,2.3958976,2.4746668,2.8455386,3.4100516,3.9056413,3.9154875,4.3651285,4.276513,4.276513,4.562052,4.8804107,3.8990772,4.57518,4.781949,4.273231,4.673641,5.211898,5.3398976,5.907693,6.5903597,5.8945646,6.0619493,5.2709746,5.3694363,7.4469748,11.851488,5.9569235,7.0367184,9.878975,11.277129,10.013539,8.5891285,9.019077,9.127385,8.582564,8.884514,7.643898,8.201847,9.6,10.948924,11.441232,10.282667,9.055181,9.642668,11.477334,11.54954,11.280411,11.500309,12.301129,13.00677,12.189539,11.867898,11.749744,12.386462,13.213539,12.547283,12.409437,12.937847,14.034052,15.796514,18.546873,18.392616,17.345642,16.01641,14.92677,14.500104,14.372104,13.879796,13.275898,12.708103,12.225642,12.78359,13.111795,13.705847,14.63795,15.547078,15.855591,16.54154,16.777847,16.193642,14.867694,14.319591,14.434463,14.171899,13.761642,14.713437,15.117129,16.580925,18.051283,18.70113,17.923283,17.23077,17.46708,17.457232,17.017437,16.955078,16.436514,16.278976,16.331488,16.259283,15.520822,15.153232,14.70359,14.611693,14.7790785,14.562463,13.958565,12.813129,11.949949,11.844924,12.626052,13.108514,13.525334,13.384206,12.924719,13.111795,13.63036,13.430155,13.331694,13.5318985,13.6008215,14.096412,14.188309,13.869949,13.334975,12.983796,13.896206,15.254975,16.06236,15.484719,12.842668,13.755078,15.629129,15.415796,12.95754,10.981745,12.389745,11.894155,10.522257,9.29477,9.235693,0.6104616,0.69579494,0.67938465,0.7417436,0.8992821,1.0010257,1.1716924,1.1257436,1.1552821,1.276718,1.2340513,2.028308,2.3401027,2.3663592,2.3827693,2.7634873,2.3794873,2.2186668,2.4615386,2.8127182,2.5206156,3.2229745,3.501949,3.626667,3.5872824,3.0851285,3.515077,4.135385,4.6539493,5.0510774,5.5893335,5.8453336,5.83877,5.7731285,5.5138464,4.578462,4.6276927,5.142975,5.924103,6.47877,6.038975,6.445949,6.9677954,7.194257,7.2237954,7.680001,8.093539,8.523488,9.209436,9.803488,9.370257,9.252103,9.613129,9.632821,9.3768215,9.780514,10.515693,10.617436,10.203898,9.622975,9.452309,10.069334,10.935796,11.625027,11.953232,11.98277,11.700514,12.009027,12.347078,12.681848,13.522053,14.086565,14.191591,13.659899,13.003489,13.430155,12.937847,12.363488,12.173129,12.4685135,12.970668,13.83713,14.670771,15.14995,15.392821,15.960617,15.737437,15.392821,15.42236,15.734155,15.642258,15.940925,15.43877,14.759386,14.306462,14.260514,14.122667,13.764924,13.157744,12.504617,12.258463,12.356924,12.471796,12.760616,13.35795,14.378668,14.368821,13.380924,12.511181,12.265027,12.5374365,12.009027,11.667693,11.625027,11.785847,11.844924,12.022155,12.265027,12.058257,11.651283,12.071385,13.5778475,14.611693,14.943181,14.70359,14.401642,14.345847,14.421334,14.555899,14.91036,15.914668,17.191385,17.240616,17.54913,18.848822,21.097027,20.260103,19.672617,18.44513,16.840206,16.272411,15.465027,14.86113,14.641232,14.851283,15.399385,16.085335,16.62031,16.551386,15.734155,14.332719,15.924514,18.628925,20.158361,19.672617,17.792002,17.056822,16.62031,16.426668,16.36431,16.249437,16.114874,14.355694,13.285745,13.653335,14.674052,15.333745,15.970463,15.304206,13.676309,13.036308,12.836103,12.140308,11.552821,11.667693,13.042872,13.814155,13.74195,13.718975,14.582155,17.125746,17.414566,14.92677,12.800001,12.140308,12.015591,12.76718,12.724514,12.245335,11.641437,11.1983595,11.96636,12.340514,12.07795,11.382154,10.9226675,11.290257,11.588924,11.972924,12.209231,11.667693,10.125129,9.426052,9.18318,9.068309,8.809027,7.9228725,7.1187696,6.2588725,5.5302567,5.421949,5.0674877,5.5236926,6.1013336,6.3376417,5.979898,5.7501545,6.3540516,7.000616,7.450257,7.9950776,8.201847,8.470975,8.323282,7.712821,7.020308,6.380308,6.2490263,6.157129,5.973334,5.920821,6.1505647,6.091488,6.485334,7.3452315,7.9524107,8.605539,9.078155,8.746667,7.6274877,6.373744,5.7731285,5.9667697,6.1997952,6.2720003,6.547693,6.806975,7.896616,8.434873,8.178872,8.021334,7.2270775,6.8627696,6.6461544,6.0980515,4.519385,3.4921029,5.1856413,8.470975,12.484924,16.643284,15.081027,13.315283,10.072617,6.091488,4.1091285,2.4943593,2.1300514,1.8543591,1.339077,1.083077,0.6662565,0.45620516,0.44964105,0.5284103,0.4660513,0.41682056,0.55794877,1.7624617,3.5413337,4.069744,6.8627696,7.958975,7.9195905,6.547693,2.8914874,2.674872,3.387077,2.8324106,2.041436,5.287385,8.306872,9.728001,7.680001,3.6168208,2.3236926,0.5907693,0.4660513,0.50543594,0.26256412,0.3052308,0.6170257,0.5152821,0.69251287,1.0994873,0.93866676,0.79097444,0.42994875,0.24287182,0.38728207,0.77128214,1.6935385,1.8379488,1.8084104,1.8051283,1.6344616,2.3860514,1.9331284,1.3259488,1.2242053,1.8970258,3.7809234,3.3280003,3.0949745,3.629949,3.4691284,3.9614363,3.6627696,3.367385,3.0752823,2.028308,3.9220517,3.3345644,2.6518977,2.4943593,1.7362052,3.2262566,5.1200004,5.504,5.6943593,10.256411,11.208206,11.881026,11.884309,10.9915905,9.156924,9.8592825,10.676514,11.093334,11.096616,11.155693,11.208206,11.227899,10.752001,10.486155,12.288001,12.629334,12.160001,11.057232,9.718155,8.730257,8.749949,8.277334,7.9491286,7.968821,8.090257,7.50277,6.0816417,5.1298466,4.926359,4.7261543,4.7983594,5.287385,5.8092313,6.3376417,7.2172313,8.79918,8.251078,6.8266673,5.618872,5.5565133,4.086154,2.6584618,1.8773335,1.910154,2.477949,1.9364104,1.9954873,2.231795,2.546872,3.1671798,4.345436,4.6211286,5.0215387,5.4941545,4.8771286,3.9023592,4.263385,4.650667,4.5456414,4.2174363,4.135385,4.194462,3.9417439,3.383795,2.9768207,2.986667,3.186872,3.9942567,4.84759,4.210872,5.799385,5.7796926,5.0543594,4.706462,5.9930263,7.4371285,9.110975,9.472001,8.792616,9.170052,10.443488,8.621949,8.474257,9.570462,6.294975,7.8670774,8.966565,9.862565,10.368001,9.82318,5.9470773,5.4482055,6.439385,7.4075904,7.2303596,8.556309,7.834257,5.6451287,3.4625645,3.6463592,3.9384618,5.3234878,7.0137444,8.402052,9.051898,10.029949,9.613129,8.648206,9.527796,16.196924,15.241847,10.262975,6.117744,5.077334,6.810257,4.450462,5.182359,7.0104623,8.300308,7.755488,8.484103,9.347282,8.004924,5.2578464,5.024821,6.186667,7.6635904,6.5411286,3.3772311,2.2022567,3.5840003,6.2490263,6.3245134,4.089436,3.9745643,3.6857438,1.8313848,2.0939488,4.46359,5.2381544,5.7731285,6.3573337,6.75118,7.072821,7.8080006,8.165744,7.9228725,7.2303596,6.117744,4.4865646,4.2830772,4.8804107,5.87159,6.8660517,7.4797955,7.2172313,6.7183595,6.636308,6.5411286,4.9099493,5.0871797,5.4449234,5.540103,5.346462,5.2447186,5.8880005,6.7314878,6.918565,6.629744,7.0793853,7.0859494,6.7150774,6.4590774,6.3343596,5.901129,5.612308,5.408821,5.0477953,4.571898,4.325744,4.1517954,3.7842054,3.442872,3.4198978,4.066462,4.010667,3.6791797,3.370667,2.9735386,1.9561027,1.8937438,1.5491283,1.467077,1.6869745,1.7263591,1.9659488,2.2580514,2.6912823,3.186872,3.4625645,3.1376412,3.1803079,3.2229745,3.2853336,3.751385,3.1343591,2.6453335,2.2711797,1.9462565,1.5688206,1.3095386,1.4867693,2.3630772,3.1474874,1.9987694,1.4375386,1.6147693,2.0676925,2.3991797,2.2613335,2.3138463,2.5271797,2.9013336,3.2754874,3.314872,3.8695388,4.135385,4.5128207,5.0609236,5.477744,4.604718,5.074052,5.208616,4.8016415,5.1331286,5.927385,6.3343596,6.820103,6.885744,5.0674877,4.965744,4.854154,4.493129,4.342154,5.543385,5.549949,7.8408213,9.977437,10.541949,9.143796,8.809027,8.891078,8.986258,8.726975,7.7948723,7.499488,7.785026,8.224821,8.79918,9.888822,10.230155,9.298052,9.747693,11.477334,11.638155,11.188514,11.076924,11.45436,12.038565,12.143591,12.028719,11.815386,12.143591,12.632616,11.867898,12.225642,12.832822,13.774771,15.090873,16.794258,17.355488,17.027283,16.026258,14.828309,14.165335,14.14236,13.66318,13.213539,12.931283,12.58995,12.740924,13.4859495,14.122667,14.506668,15.067899,15.37313,16.393847,16.981335,16.426668,14.477129,13.551591,13.574565,13.656616,13.50236,13.4170265,14.437745,15.468308,16.134565,16.288822,16.000002,15.442053,15.931078,16.30195,16.091898,15.540514,15.0777445,15.491283,16.101746,16.331488,15.701335,15.238565,14.772514,14.247386,13.801026,13.7386675,13.545027,12.662155,11.867898,11.730052,12.6063595,13.39077,13.633642,13.262771,12.786873,13.308719,13.676309,13.515489,13.338258,13.3940525,13.659899,13.909334,14.037334,13.666463,13.095386,13.305437,13.692719,14.237539,15.07118,15.51754,14.080001,13.499078,13.61395,13.453129,12.389745,10.144821,10.496001,10.561642,10.345026,9.947898,9.577026,0.5546667,0.7056411,0.76800007,0.86646163,1.0010257,1.0436924,1.211077,1.204513,1.3357949,1.5327181,1.3620514,2.0217438,2.300718,2.546872,2.7864618,2.7437952,2.3269746,2.2449234,2.5238976,2.9505644,3.0818465,3.8695388,4.197744,4.2141542,3.9318976,3.2262566,3.4264617,4.2371287,4.7392826,4.890257,5.5204105,5.6287184,5.6418467,5.5729237,5.221744,4.1452312,4.4307694,4.955898,6.0947695,7.312411,7.125334,7.2336416,7.27959,7.0859494,6.928411,7.5520005,8.303591,8.868103,9.380103,9.632821,9.074872,9.340718,9.6,10.056206,10.545232,10.561642,10.276103,10.538668,10.886565,11.0375395,10.909539,10.906258,11.083488,11.280411,11.382154,11.329642,11.424822,11.684103,12.09436,12.685129,13.5089245,13.449847,13.568001,13.131488,12.3306675,12.2847185,12.265027,11.88759,11.864616,12.347078,12.914873,14.060308,14.828309,15.110565,15.179488,15.67836,15.770258,15.596309,15.212309,14.923489,15.27795,15.530668,14.880821,14.211283,13.929027,13.961847,14.237539,14.135796,13.705847,13.1872835,13.010053,13.213539,13.29559,13.380924,13.564719,13.922462,14.080001,13.4859495,12.865642,12.547283,12.475078,12.11077,11.828514,11.460924,11.142565,11.313231,11.608616,12.166565,12.740924,13.289026,13.965129,15.291079,16.085335,16.032822,15.222155,14.132514,13.748514,14.122667,14.460719,14.720001,15.586463,16.04595,16.518566,16.853334,17.667284,20.322464,19.899078,19.879387,19.528206,18.471386,16.705643,15.642258,15.304206,15.238565,15.366566,15.990155,16.833643,17.109335,16.577642,15.428925,14.273643,15.218873,17.375181,18.75036,18.389336,16.387283,15.320617,14.949745,14.985847,15.38954,16.341335,16.472616,14.582155,13.574565,14.214565,15.130258,16.607182,17.828104,17.6279,16.341335,15.819489,15.189335,14.329437,13.351386,12.501334,12.133744,12.511181,12.544001,13.5318985,15.885129,19.114668,19.272207,16.09518,13.522053,13.095386,13.991385,15.43877,14.345847,12.980514,12.36677,12.291283,12.458668,12.849232,13.200411,13.210258,12.540719,11.395283,10.955488,11.050668,11.336206,11.277129,10.154668,9.662359,9.711591,9.91836,9.590155,7.88677,6.5805135,5.658257,5.077334,4.7392826,4.7261543,5.106872,5.5204105,5.8256416,6.0816417,5.76,6.262154,7.0367184,7.6996927,8.044309,8.027898,7.75877,7.381334,7.0104623,6.764308,6.0192823,6.193231,6.3442054,6.124308,5.799385,5.901129,5.7468724,6.196513,7.250052,8.03118,8.172308,8.851693,8.572719,7.2303596,6.0685134,5.5302567,5.7665644,6.173539,6.442667,6.554257,6.62318,7.2992826,7.683283,7.5454364,7.318975,6.6625648,5.973334,5.346462,4.7228723,3.8728209,3.0194874,5.467898,9.852718,14.36554,16.718771,12.678565,9.074872,5.7829747,3.18359,2.1792822,2.487795,2.6584618,2.1497438,1.2668719,1.1618463,0.56123084,0.27241027,0.23958977,0.33805132,0.4004103,0.4594872,0.40369233,1.394872,3.1934361,4.1682053,6.0717955,6.042257,6.491898,6.944821,4.027077,1.6443079,1.4966155,2.4582565,3.9220517,5.7764106,7.79159,6.2490263,3.620103,1.7985642,2.1202054,0.5316923,0.2231795,0.32820517,0.39384618,0.36758977,0.44964105,0.4397949,0.6826667,1.020718,0.8172308,0.86974365,0.5546667,0.42338464,0.8008206,1.7723079,2.2022567,2.0841026,1.8445129,1.522872,0.7778462,0.8795898,1.3784616,1.8248206,2.3860514,3.8334363,4.8836927,4.194462,3.698872,3.8104618,3.4133337,3.1442053,2.6584618,2.5140514,2.3991797,1.1027694,3.2918978,2.9735386,2.9472823,3.3411283,1.6147693,2.7766156,4.273231,5.579488,7.3616414,11.457642,10.066052,9.750975,9.905231,9.728001,8.241231,9.747693,10.712616,11.218052,11.346052,11.142565,11.516719,11.313231,10.614155,10.299078,12.048411,12.225642,12.245335,11.864616,10.948924,9.468719,9.03877,8.4053335,7.9983597,7.7357955,7.0531287,6.426257,5.2709746,4.6178465,4.667077,4.788513,4.6769233,5.156103,5.7009234,6.2851286,7.3747697,9.265231,8.592411,7.125334,5.98318,5.654975,4.420923,2.934154,2.1464617,2.2022567,2.4352822,1.6344616,1.6804104,1.9298463,2.2186668,2.868513,4.204308,4.8049235,5.1922054,5.349744,4.71959,4.1156926,4.6112823,4.647385,4.027077,3.9056413,4.266667,4.453744,4.466872,4.3290257,4.0992823,3.8071797,3.7284105,4.2994876,5.037949,4.5423594,5.349744,5.218462,4.969026,5.1167183,5.87159,5.208616,6.5706673,7.975385,8.582564,8.700719,11.316514,8.786052,8.753231,11.437949,9.632821,8.470975,9.55077,10.28595,9.895386,9.38995,6.23918,5.7796926,6.8496413,7.515898,5.0871797,6.7282057,6.918565,4.7950773,2.9571285,7.4797955,6.7216415,7.574975,8.615385,9.750975,12.232206,16.961643,14.28677,9.793642,8.470975,14.742975,17.857643,16.370872,11.208206,5.540103,4.772103,4.578462,5.2545643,5.865026,6.1308722,6.442667,6.11118,8.556309,9.07159,6.7150774,4.273231,5.668103,7.0137444,5.674667,2.7470772,3.058872,3.318154,4.9788723,5.0182567,3.5183592,3.6627696,2.2121027,2.300718,3.9286156,5.9602056,6.12759,6.117744,6.0717955,6.0324106,6.3606157,7.722667,9.193027,8.960001,7.9983597,6.820103,5.4580517,4.457026,4.397949,5.3005133,6.6395903,7.3386674,6.997334,6.012718,6.377026,7.3485136,5.435077,5.3169236,5.7042055,6.183385,6.3212314,5.648411,5.87159,6.619898,6.8397956,6.442667,6.3179493,6.409847,6.4623594,6.5083084,6.485334,6.2490263,5.9602056,5.8190775,5.61559,5.2414365,4.699898,4.309334,4.1550775,3.8104618,3.4002054,3.6036925,4.141949,3.9909747,3.7710772,3.4231799,2.2186668,1.7952822,1.4834872,1.3522053,1.3915899,1.5327181,1.9954873,2.1202054,2.3401027,2.7569232,3.1277952,3.0916924,3.0490258,2.8980515,2.7667694,3.0227695,2.5862565,2.2678976,1.9922053,1.719795,1.4572309,1.332513,1.5589745,2.4976413,3.3476925,2.1530259,1.5031796,1.6377437,2.0545642,2.2613335,1.7985642,1.9364104,2.1825643,2.553436,2.9210258,3.0162053,3.56759,4.082872,4.4307694,4.640821,4.886975,4.5587697,4.9132314,5.1200004,5.106872,5.586052,6.377026,7.1089234,7.177847,6.4065647,5.0215387,5.4843082,5.835488,5.3070774,4.4110775,4.926359,6.547693,8.694155,9.734565,9.301334,8.264206,8.477539,8.3823595,8.516924,8.562873,7.3353853,7.0990777,7.059693,7.076103,7.453539,8.946873,10.036513,9.409642,9.524513,10.893129,12.068104,11.605334,11.208206,10.988309,11.076924,11.618463,11.592206,11.23118,11.411694,11.884309,11.270565,11.802258,12.583385,13.889642,15.133539,14.854566,15.340309,15.671796,15.53395,14.933334,14.208001,14.158771,13.636924,13.049437,12.668719,12.642463,12.675283,13.659899,14.375385,14.467283,14.450873,15.435489,16.466053,16.748308,15.911386,14.007796,13.111795,13.115078,13.200411,13.065847,12.950975,13.925745,14.358975,14.473847,14.378668,14.04718,13.958565,14.464001,14.887385,14.8709755,14.368821,14.785643,15.212309,15.510976,15.530668,15.097437,14.65436,14.244103,13.604104,12.993642,13.157744,12.76718,12.297847,11.910565,11.861334,12.507898,13.46954,13.764924,13.403898,12.895181,13.236514,13.505642,13.22995,13.010053,13.177437,13.774771,13.869949,14.201437,13.991385,13.397334,13.51877,13.74195,13.833847,14.280207,14.92677,15.002257,14.083283,13.062565,12.672001,12.514462,11.067078,10.650257,10.624001,10.794667,10.840616,10.30236,0.47589746,0.73517954,1.0436924,1.1881026,1.1716924,1.2274873,1.2274873,1.2964103,1.5261539,1.7558975,1.5885129,1.7755898,2.048,2.4713848,2.8980515,2.9702566,2.5140514,2.3171284,2.605949,3.2131286,3.570872,3.9286156,4.5029745,4.4832826,3.9122055,3.698872,3.31159,3.639795,4.1058464,4.5489235,5.2020516,5.6418467,5.8978467,5.6976414,5.028103,4.125539,4.562052,4.7491283,5.924103,7.955693,9.340718,8.444718,7.958975,7.565129,7.325539,7.6668725,8.592411,9.330873,9.3078985,8.585847,7.857231,8.618668,9.005949,9.941334,11.195078,11.392001,10.473026,10.20718,10.840616,11.766154,11.536411,11.355898,11.090053,10.791386,10.696206,11.1983595,11.510155,11.651283,12.09436,12.747488,12.95754,12.954257,13.302155,13.003489,12.045129,11.382154,11.848206,11.815386,11.946668,12.373334,12.71795,13.334975,13.804309,14.260514,14.788924,15.455181,15.839181,15.668514,14.729847,13.843694,14.857847,14.982565,14.401642,14.043899,14.112822,14.102976,14.25395,14.152206,13.889642,13.587693,13.413745,13.272616,13.056001,12.793437,12.57354,12.534155,13.00677,13.1872835,13.016617,12.455385,11.464206,10.965334,11.024411,11.149129,11.224616,11.510155,11.592206,11.835078,12.63918,13.824001,14.63795,15.087591,15.619284,15.566771,14.838155,13.883078,13.781334,14.017642,14.070155,13.978257,14.352411,14.539488,15.977027,17.09949,17.604925,18.44513,18.881643,20.109129,20.788515,20.345438,18.960411,16.91241,16.026258,16.039387,16.479181,16.66954,17.092924,16.600616,15.816206,15.05477,14.319591,14.01436,14.313026,14.943181,15.379693,14.854566,14.096412,13.810873,14.162052,15.100719,16.377438,15.766975,14.214565,13.718975,14.680616,15.8884115,16.78113,17.877335,18.720821,18.901335,18.041437,16.410257,15.064616,14.290052,13.840411,12.934566,12.484924,12.068104,13.426873,16.328207,18.569847,17.808413,15.980309,14.746258,14.854566,16.144411,17.844515,15.891693,13.666463,12.757335,12.980514,11.953232,11.661129,12.586668,13.994668,13.912617,12.297847,11.54954,10.873437,9.944616,8.900924,8.349539,8.704,9.193027,9.488411,9.682052,7.456821,5.805949,5.0642056,4.955898,4.598154,4.5587697,4.8311796,5.2676926,5.7534366,6.2096415,6.114462,6.3868723,6.997334,7.712821,8.090257,7.9228725,7.2861543,6.685539,6.409847,6.5444107,5.8847184,6.1046157,6.373744,6.3212314,6.0192823,5.7632823,5.72718,6.1374364,6.8529234,7.394462,7.7325134,7.972103,7.5487185,6.6560006,6.2588725,5.6385646,5.6320004,5.9667697,6.422975,6.8299494,6.957949,6.9809237,6.918565,6.7117953,6.245744,5.970052,4.906667,3.8104618,3.1540515,3.1507695,2.4352822,3.8629746,6.5870776,9.567181,11.575796,7.253334,4.844308,3.5249233,2.8422565,2.7208207,3.2262566,2.7437952,1.7723079,0.8467693,0.5316923,0.35446155,0.21661541,0.26584616,0.46276927,0.6104616,0.6235898,0.4955898,0.9682052,2.176,3.6332312,3.4166157,3.498667,6.3245134,9.301334,4.8114877,3.508513,3.8137438,5.362872,6.0717955,2.1431797,2.8914874,2.4516926,1.6410258,1.1716924,1.6475899,0.45292312,0.25928208,0.42338464,0.5316923,0.38400003,0.34789747,0.4594872,0.6301539,0.77128214,0.78769237,0.8041026,0.5415385,0.54482055,1.2077949,2.7569232,2.2613335,1.7558975,1.2274873,0.8205129,0.82379496,1.2800001,1.8510771,2.9144619,4.450462,6.0324106,5.3366156,5.0510774,4.8049235,4.3716927,3.6529233,2.809436,2.1530259,2.353231,2.6978464,1.083077,2.4615386,2.4188719,2.986667,3.7940516,2.0906668,2.930872,3.9187696,5.9634876,9.137232,12.678565,10.020103,8.3593855,8.277334,8.969847,8.228104,9.737847,10.584617,11.0375395,11.23118,11.172104,11.45436,10.811078,10.052924,10.095591,11.959796,11.1983595,10.8767185,10.748719,10.71918,10.866873,10.006975,8.956718,8.195283,7.5487185,6.193231,5.72718,4.673641,4.059898,4.2338467,4.8738465,4.568616,4.827898,5.5696416,6.4754877,6.9743595,8.132924,7.765334,6.8397956,6.055385,5.8190775,4.453744,3.0851285,2.3729234,2.166154,1.4933335,1.2373334,1.5064616,1.9692309,2.546872,3.4264617,4.588308,4.7458467,4.57518,4.4865646,4.6145644,4.70318,4.9099493,4.493129,3.69559,3.7152824,4.3651285,4.6966157,4.906667,5.0084105,4.821334,4.529231,4.4045134,4.6539493,5.028103,4.821334,4.630975,4.6539493,5.2545643,6.226052,6.7971287,6.11118,5.8912826,5.8256416,5.976616,6.7971287,9.862565,6.9021544,6.160411,9.32759,11.546257,10.433641,9.590155,9.724719,9.990565,7.9917955,7.3550773,5.970052,6.0980515,6.7117953,3.5216413,3.2689233,2.681436,2.2219489,4.076308,12.1468725,9.370257,8.064001,6.8529234,6.8988724,11.897437,23.591387,19.272207,11.74318,8.628513,12.3536415,17.736206,24.631796,21.937233,11.247591,6.875898,7.145026,7.762052,7.020308,5.7698464,7.4371285,5.179077,4.57518,5.7632823,6.744616,3.3772311,3.6726158,3.2525132,3.0227695,3.495385,4.8016415,4.397949,3.5544617,3.508513,3.6594875,1.5721027,1.3489232,3.9187696,5.8486156,6.2851286,6.9382567,6.550975,5.973334,5.5204105,5.72718,7.3583593,9.380103,9.248821,8.385642,7.499488,6.5772314,5.2053337,4.601436,5.0018463,6.0192823,6.6461544,6.803693,5.8157954,6.1341543,7.312411,6.0324106,6.3540516,6.363898,6.6822567,7.059693,6.38359,5.933949,6.422975,6.5411286,6.091488,5.989744,6.0028725,6.2884107,6.5050263,6.442667,6.0356927,5.5236926,5.4580517,5.549949,5.5302567,5.179077,4.8377438,4.781949,4.312616,3.4560003,2.9472823,3.7973337,3.8334363,3.5774362,3.259077,2.806154,2.0250258,1.7788719,1.522872,1.1913847,1.2012309,1.591795,1.7165129,1.9954873,2.5107694,3.0162053,3.058872,2.8455386,2.609231,2.4746668,2.4681027,2.1891284,1.8346668,1.4375386,1.1388719,1.1848207,1.1388719,1.2209232,1.8084104,2.5238976,2.2514873,1.7493335,1.7985642,1.9429746,1.847795,1.2931283,1.5589745,1.9364104,2.3958976,2.8455386,3.1507695,3.4198978,3.9351797,3.9975388,3.6102567,3.4691284,3.5807183,4.06318,4.5522056,4.9296412,5.330052,6.3507695,7.27959,6.7610264,5.290667,5.218462,6.193231,6.6494365,6.3868723,6.012718,6.9382567,7.8506675,8.78277,8.700719,7.8112826,7.565129,7.755488,7.643898,7.5618467,7.5454364,7.315693,6.4689236,6.0160003,6.173539,7.000616,8.395488,9.6984625,9.232411,8.792616,9.544206,12.048411,11.792411,11.47077,11.008,10.532104,10.354873,10.57477,10.115283,10.289231,11.030975,10.896411,11.300103,12.137027,13.63036,14.943181,14.165335,13.505642,14.14236,14.959591,15.156514,14.250668,14.293334,14.211283,13.479385,12.383181,12.025436,12.317539,13.321847,14.083283,14.267078,14.12595,15.392821,15.95077,15.67836,14.815181,13.955283,13.302155,13.226667,12.947693,12.632616,13.426873,13.499078,13.482668,13.46954,13.279181,12.442257,13.078976,13.99795,14.506668,14.486976,14.391796,15.875283,15.317334,14.378668,13.827283,13.512206,13.059283,12.931283,12.701539,12.435693,12.694975,11.9860525,11.71036,11.733335,11.940104,12.258463,12.777026,13.029744,13.013334,12.918155,13.121642,13.22995,12.816411,12.642463,13.016617,13.801026,13.840411,14.506668,14.65436,14.063591,13.426873,13.869949,13.971693,13.830565,13.850258,14.726565,14.6182575,13.466257,12.649027,12.635899,12.99036,12.435693,11.88759,11.621744,11.565949,11.323078,0.67282057,0.9878975,1.4900514,1.6246156,1.3620514,1.1913847,1.2865642,1.2931283,1.5064616,1.8084104,1.6640002,1.8576412,2.412308,2.5993848,2.481231,2.8849232,2.6518977,2.986667,3.1967182,3.117949,3.1442053,3.5216413,3.9548721,3.9680004,3.7349746,4.089436,3.6758976,3.6332312,4.240411,5.2414365,5.874872,6.705231,6.3540516,5.579488,4.8705645,4.457026,5.225026,5.031385,5.540103,7.1187696,8.864821,8.438154,9.291488,9.718155,8.923898,7.020308,8.326565,9.613129,9.796924,9.078155,8.956718,8.79918,9.38995,9.816616,9.90195,10.20718,11.172104,11.569232,11.533129,11.280411,11.109744,11.487181,11.490462,11.569232,11.956513,12.665437,11.871181,11.992617,12.3536415,12.383181,11.628308,12.885334,13.656616,13.167591,11.871181,11.444513,11.907283,12.199386,12.484924,12.678565,12.435693,12.35036,13.216822,14.119386,14.660924,14.953027,14.588719,14.477129,13.909334,13.1872835,13.627078,14.053744,13.88636,13.63036,13.492514,13.380924,12.918155,12.76718,12.960821,13.243078,13.046155,12.937847,12.908309,12.914873,12.937847,12.983796,13.203693,12.793437,12.416001,12.150155,11.490462,10.893129,10.752001,11.201642,11.9860525,12.452104,12.317539,12.337232,12.619488,13.026463,13.200411,12.954257,13.259488,13.449847,13.505642,14.053744,13.784616,13.745232,13.545027,13.364513,13.961847,15.340309,17.434258,19.167181,19.800617,18.921026,17.93313,17.969233,18.707693,19.669334,20.217438,17.250463,15.852309,16.059078,17.168411,17.729643,17.80513,16.331488,15.261539,15.087591,14.831591,14.185027,13.226667,13.029744,13.673027,14.221129,13.843694,13.016617,12.832822,13.791181,15.793232,15.376411,14.04718,13.308719,13.984821,16.20349,16.961643,16.896002,17.67713,18.822565,17.700104,15.113848,13.147899,13.689437,15.753847,15.471591,14.447591,13.000206,12.836103,13.991385,14.8480015,14.309745,16.170668,18.107079,18.87836,18.340103,17.217642,16.233027,15.012104,13.820719,13.564719,11.759591,11.378873,11.250873,11.044104,11.277129,12.373334,12.806565,12.822975,12.235488,10.390975,7.778462,8.077128,8.969847,9.242257,8.805744,6.948103,5.549949,4.965744,5.0871797,5.356308,5.0018463,5.2348723,5.6352825,5.904411,5.8453336,6.5411286,7.125334,7.27959,7.2369237,7.7981544,7.3583593,6.5805135,6.304821,6.5805135,6.6527185,6.3967185,5.976616,5.979898,6.311385,6.163693,5.3234878,5.4875903,6.0619493,6.6002054,6.820103,8.260923,8.493949,7.962257,7.210667,6.882462,6.954667,6.3606157,5.858462,6.0258465,7.2336416,7.0367184,6.5870776,6.196513,6.235898,7.125334,5.4908724,4.2207184,3.5183592,3.1015387,2.1989746,2.2350771,2.481231,3.062154,3.6168208,3.31159,1.5786668,2.2613335,2.665026,2.0644104,1.7099489,1.6475899,1.404718,1.086359,0.8730257,1.0075898,0.95835906,0.6268718,0.32164106,0.34133336,0.97805136,0.8041026,0.54482055,0.7318975,1.3751796,1.9364104,2.0118976,2.678154,5.970052,9.718155,7.584821,10.243283,8.832001,9.101129,9.977437,3.570872,3.3641028,2.231795,1.083077,0.4135385,0.3052308,0.34133336,0.54482055,0.63343596,0.5546667,0.45620516,0.46933338,0.8205129,0.85005134,0.58092314,0.702359,0.64000005,0.5349744,0.827077,1.522872,2.1825643,2.3040001,1.1815386,0.61374366,0.9353847,1.0075898,2.2646155,3.1737437,5.0051284,7.020308,6.485334,5.4482055,6.2030773,5.976616,4.457026,3.8006158,2.7995899,2.9243078,3.515077,3.511795,1.4506668,1.1552821,2.162872,2.8488207,2.6518977,2.0906668,2.1398976,3.892513,6.7905645,10.003693,12.419283,11.687386,10.505847,9.665642,9.009232,7.4469748,8.264206,9.567181,10.70277,11.428103,11.9171295,11.611898,11.122872,10.70277,10.752001,11.825232,10.361437,8.4283085,7.9458466,9.416205,11.9171295,11.172104,9.494975,8.254359,7.460103,5.7534366,5.3727183,4.519385,4.06318,4.263385,4.775385,4.420923,4.0303593,5.159385,6.9349747,6.058667,6.2884107,6.6395903,6.340924,5.5630774,5.4153852,4.634257,3.5872824,2.674872,1.9692309,1.2373334,1.6640002,1.7887181,2.0512822,2.7798977,4.197744,5.356308,5.0609236,4.585026,4.637539,5.3694363,5.1889234,4.5095387,3.761231,3.3476925,3.6758976,4.348718,4.955898,5.3694363,5.297231,4.273231,4.906667,4.781949,4.562052,4.663795,5.2480006,4.493129,4.1846156,4.5456414,5.293949,5.661539,6.5772314,7.3353853,8.349539,9.590155,10.604308,9.091283,5.2709746,2.8291285,2.878359,3.95159,5.7698464,8.891078,9.114257,7.955693,12.619488,10.020103,8.700719,7.6209235,6.9021544,7.8441033,4.97559,2.6190772,2.3696413,4.578462,8.362667,4.9821544,4.7655387,5.280821,5.3169236,4.9132314,26.873438,19.685745,9.462154,6.5312824,5.431795,4.9920006,23.67672,30.244104,19.826874,13.932309,12.294565,11.969642,9.593436,6.692103,9.659078,5.398975,4.644103,4.460308,3.9384618,4.197744,5.612308,4.0533338,2.7044106,3.945026,9.353847,11.063796,5.6385646,1.8116925,1.8281027,1.4506668,2.097231,3.9876926,5.979898,7.13518,6.744616,6.806975,6.4000006,5.5696416,5.172513,6.882462,9.908514,9.31118,7.906462,6.954667,6.1505647,5.3924108,4.9296412,5.1987696,5.8420515,5.7074876,7.1220517,7.072821,6.8233852,6.5936418,5.5696416,6.4000006,6.1407185,6.0619493,6.38359,6.2851286,5.9930263,6.6527185,6.7249236,6.1505647,6.3310776,6.3442054,6.485334,6.931693,7.2336416,6.3179493,5.5597954,5.435077,5.76,6.2523084,6.5444107,5.8256416,4.9788723,4.31918,3.7907696,2.9604106,3.4494362,3.3772311,3.1048207,2.9669745,3.2951798,2.356513,2.1398976,2.0053334,1.654154,1.1290257,1.0666667,1.2373334,1.7723079,2.5009232,2.930872,3.0030773,2.8849232,2.7503593,2.6157951,2.3335385,1.8215386,1.5097437,1.1815386,0.90256417,1.0371283,0.9156924,0.9485129,1.2603078,1.7165129,1.9232821,1.9462565,1.9790771,1.9265642,1.7329233,1.404718,1.6968206,1.8707694,2.1333334,2.5764105,3.1737437,3.4067695,3.7940516,3.8432825,3.5807183,3.5544617,3.7251284,4.023795,4.312616,4.414359,4.135385,6.2096415,6.764308,5.802667,4.3651285,4.5456414,5.366154,6.055385,6.3540516,6.6100516,7.781744,7.893334,8.073847,7.640616,6.941539,7.3714876,6.7117953,6.619898,6.2162056,5.605744,5.874872,5.8518977,5.7698464,5.6320004,5.8814363,7.430565,9.800206,10.31877,9.475283,8.717129,10.436924,10.033232,10.584617,11.017847,10.817642,10.026668,10.148104,9.984001,9.856001,10.029949,10.725744,10.935796,11.920411,12.652308,13.078976,14.129231,13.275898,13.656616,14.444309,14.667488,13.213539,13.617231,14.907078,14.785643,13.049437,11.595488,11.644719,12.025436,12.645744,13.430155,14.296617,13.942155,14.17518,14.375385,14.418053,14.6642065,13.686155,12.645744,12.245335,12.560411,13.062565,12.829539,12.852514,12.872206,12.599796,11.733335,12.967385,15.455181,16.754873,16.38072,15.80636,16.784412,14.867694,12.744206,11.572514,10.985026,10.571488,11.162257,11.621744,11.523283,11.168821,11.670976,11.017847,10.686359,11.158976,11.9171295,11.575796,10.896411,10.939077,11.913847,13.184001,13.13477,13.049437,13.078976,13.285745,13.640206,13.640206,14.145642,14.424617,14.086565,13.062565,12.977232,13.019898,12.928001,12.885334,13.51877,14.385232,13.154463,11.802258,11.513436,12.711386,12.465232,12.35036,12.3076935,12.383181,12.724514,1.2077949,1.1355898,1.2668719,1.2406155,1.1585642,1.591795,1.7493335,1.6016412,1.5655385,1.7394873,1.8937438,1.6508719,2.3138463,2.7011285,2.5993848,2.737231,2.9440002,3.2722054,3.318154,3.18359,3.4592824,3.2131286,3.2853336,3.5216413,3.9417439,4.7360005,3.6463592,3.6430771,4.06318,4.466872,4.640821,4.965744,5.6287184,5.904411,5.756718,5.858462,6.442667,6.445949,6.547693,7.0925136,8.096821,8.536616,9.051898,9.275078,9.488411,10.630565,10.072617,9.970873,10.151385,10.28595,9.908514,8.598975,8.835282,9.199591,9.416205,10.354873,11.71036,11.831796,11.651283,11.644719,11.815386,11.805539,11.657847,11.923694,12.616206,13.226667,12.629334,11.904001,11.54954,11.913847,13.226667,14.592001,13.909334,12.816411,12.186257,12.140308,11.569232,11.306667,11.336206,11.670976,12.373334,12.727796,13.633642,14.204719,14.27036,14.368821,14.263796,14.089848,13.682873,13.331694,13.761642,15.018668,14.969437,14.050463,13.056001,13.161027,13.226667,12.744206,12.422565,12.517745,12.839386,13.315283,13.515489,13.633642,13.63036,13.22995,12.678565,12.396309,11.956513,11.418258,11.293539,10.902975,11.260718,11.756309,11.956513,11.621744,11.88759,12.347078,12.612924,12.3306675,11.172104,10.998155,11.23118,11.680821,12.3306675,13.35795,13.410462,13.810873,14.592001,15.501129,16.000002,15.855591,17.824821,19.24595,19.27877,18.898052,17.253744,16.49559,16.54154,17.473642,19.5479,18.67159,16.68595,15.780104,16.49559,17.729643,17.207796,16.361027,15.619284,15.113848,14.660924,14.8250265,13.4400015,12.422565,12.635899,13.866668,12.931283,11.789129,11.418258,12.097642,13.423591,13.380924,12.507898,11.897437,12.163283,13.459693,14.821745,15.579899,16.141129,16.265848,15.074463,14.03077,13.302155,13.781334,15.317334,16.705643,15.553642,13.846975,13.883078,15.432206,15.750566,16.01313,20.70318,23.758772,22.79713,19.14749,18.569847,17.736206,17.877335,18.23836,16.068924,13.312001,12.340514,11.762873,11.23118,11.434668,12.317539,13.312001,13.869949,13.6467705,12.47836,9.26195,8.602257,9.668923,11.119591,11.099898,8.500513,6.560821,5.920821,6.0816417,5.3924108,5.037949,5.431795,5.7468724,5.72718,5.684513,7.0925136,7.88677,8.214975,8.228104,8.067283,7.6668725,7.637334,7.6110773,7.450257,7.240206,7.5585647,6.747898,6.058667,5.924103,5.933949,5.284103,5.1856413,5.5302567,6.0783596,6.4557953,7.893334,8.267488,7.565129,6.370462,5.85518,6.045539,6.2851286,6.3474874,6.482052,7.4141545,6.62318,6.6395903,6.6100516,6.3376417,6.2720003,5.0642056,3.9187696,2.7667694,1.9068719,1.9889232,2.9144619,3.1934361,3.0030773,2.789744,3.2754874,3.1245131,3.3509746,3.1245131,2.3466668,1.6607181,0.96492314,1.1848207,1.4276924,1.2570257,0.67610264,1.0010257,0.5316923,0.4266667,0.86974365,1.0732309,1.1093334,0.9911796,1.3587693,2.0676925,2.2186668,5.756718,3.7120004,3.5216413,5.9470773,5.080616,4.6769233,5.405539,5.277539,3.6791797,1.3620514,1.7690258,1.719795,1.3653334,1.0272821,1.2209232,0.7975385,0.45292312,0.28225642,0.26584616,0.2855385,0.41682056,0.57764107,0.8763078,1.1257436,0.8467693,0.62030774,0.64000005,0.7844103,1.3456411,3.0490258,2.1169233,1.0436924,0.9156924,1.7066668,2.2777438,1.6968206,2.097231,4.4898467,6.8594875,4.1550775,2.9013336,4.5062566,5.35959,4.578462,4.007385,3.4560003,4.7622566,5.861744,5.3070774,2.2678976,2.3368206,3.249231,3.6463592,2.9013336,1.1388719,1.6278975,3.4297438,6.193231,9.216001,11.457642,11.300103,9.93477,8.763078,8.385642,8.582564,9.127385,10.404103,11.16554,11.424822,12.491488,11.178667,11.093334,10.9456415,10.381129,9.984001,10.43036,10.026668,9.7673855,10.328616,12.051693,10.738873,8.848411,8.3364105,8.700719,6.9743595,5.609026,4.7491283,4.854154,5.398975,4.886975,4.7261543,5.0084105,5.395693,5.5565133,5.1659493,5.037949,5.8847184,6.232616,5.723898,5.100308,4.562052,4.2272825,3.629949,2.6945643,1.7493335,1.6968206,2.097231,2.7766156,3.6004105,4.4898467,5.044513,5.1298466,5.3924108,5.986462,6.5903597,6.3606157,5.1659493,4.086154,3.7251284,4.1911798,4.568616,5.0871797,5.3858466,5.4186673,5.4580517,5.280821,5.208616,5.0642056,4.824616,4.637539,4.818052,4.519385,4.525949,4.9296412,5.100308,5.467898,5.914257,6.889026,8.119796,8.615385,9.015796,9.202872,8.454565,7.0826674,6.416411,7.250052,5.9634876,4.1025643,3.1474874,4.4898467,5.7665644,6.442667,6.245744,5.208616,3.6693337,6.4065647,6.803693,7.5454364,8.982975,9.153642,4.6112823,5.346462,10.282667,14.122667,7.3419495,10.387693,8.011488,6.23918,6.705231,6.6395903,5.9963083,11.71036,14.729847,13.29559,12.954257,6.7872825,7.752206,7.6603084,5.106872,5.4843082,3.4198978,4.916513,4.6244106,2.4516926,3.5478978,8.5891285,8.080411,6.7905645,7.6603084,11.818667,7.6307697,3.8465643,1.7755898,1.6475899,2.5961027,4.4045134,5.4974365,6.304821,6.75118,6.242462,7.204103,7.9885135,7.958975,7.4732313,7.8834877,8.792616,9.238976,8.884514,7.830975,6.626462,6.1407185,5.717334,5.6943593,6.114462,6.7314878,6.7807183,7.3583593,6.8594875,5.9503593,7.571693,6.370462,5.5302567,5.5138464,6.0750775,6.262154,4.857436,5.654975,6.2588725,6.0750775,6.294975,5.7501545,5.9634876,6.6461544,7.2336416,6.9021544,6.7905645,6.5345645,6.0356927,5.5236926,5.533539,5.2315903,4.906667,4.84759,4.6244106,3.0818465,2.7798977,2.7766156,2.9440002,3.1409233,3.1967182,2.5600002,2.228513,2.2383592,2.3236926,1.9331284,2.546872,2.356513,2.409026,2.8225644,2.7700515,2.7963078,2.9505644,2.789744,2.353231,2.1398976,2.0742567,1.723077,1.2274873,0.78769237,0.65969235,0.7515898,0.92553854,1.3161026,1.785436,1.9364104,2.0184617,1.8970258,1.7099489,1.6213335,1.8182565,2.1989746,2.2416413,2.2613335,2.4549747,2.917744,3.2164104,3.6594875,3.6824617,3.2853336,3.0194874,3.190154,3.6562054,3.9778464,3.9187696,3.4625645,4.3290257,4.5817437,4.1058464,3.370667,3.436308,3.9909747,5.149539,6.4295387,7.4240007,7.7948723,7.397744,7.269744,6.8562055,6.3179493,6.5411286,6.2720003,6.4590774,6.3310776,5.8420515,5.691077,5.0904617,5.7107697,6.180103,6.308103,7.076103,8.713847,9.321027,9.005949,8.553026,9.42277,9.6754875,10.469745,10.742155,10.292514,9.793642,9.271795,9.724719,9.980719,9.829744,10.006975,10.331899,11.552821,12.363488,12.626052,13.37436,12.859077,13.384206,14.578873,15.432206,14.299898,14.431181,14.647796,14.322873,13.308719,11.963078,12.596514,12.586668,12.86236,13.63036,14.372104,14.39836,14.198155,13.965129,13.906053,14.237539,13.971693,13.249642,12.757335,12.675283,12.658873,13.10195,13.059283,12.4685135,11.378873,9.964309,11.703795,13.551591,15.126975,15.747283,14.391796,14.10954,13.50236,13.131488,12.872206,11.913847,11.313231,10.627283,10.345026,10.463181,10.509129,11.090053,11.195078,10.817642,10.338462,10.548513,9.662359,9.078155,9.330873,10.532104,12.3766165,12.632616,12.570257,12.898462,13.522053,13.545027,14.217847,14.053744,13.794462,13.676309,13.453129,13.131488,12.924719,12.691693,12.363488,11.933539,12.632616,12.386462,12.107488,12.2157955,12.649027,12.327386,12.389745,12.586668,12.678565,12.445539,1.332513,1.1848207,1.2668719,1.4112822,1.5163078,1.585231,1.7165129,1.6836925,1.654154,1.7263591,1.9068719,1.8018463,2.0545642,2.3401027,2.481231,2.4451284,2.5796926,2.7208207,2.8914874,3.114667,3.4133337,2.993231,3.373949,4.0369234,4.562052,4.6145644,4.332308,4.013949,4.007385,4.378257,4.9296412,4.7425647,5.100308,5.3366156,5.356308,5.6254363,6.695385,7.056411,7.0990777,7.1548724,7.509334,8.602257,8.815591,8.4512825,8.411898,10.200616,9.780514,9.659078,9.911796,10.200616,9.800206,8.500513,8.6580515,9.386667,9.990565,9.961026,11.480617,11.684103,11.483898,11.313231,11.152411,11.296822,11.244308,11.529847,12.100924,12.304411,12.196103,11.45436,11.162257,11.792411,13.203693,14.385232,13.561437,12.744206,12.619488,12.544001,11.963078,11.585642,11.300103,11.191795,11.546257,12.22236,12.901745,13.282462,13.305437,13.15118,13.1872835,13.269335,13.200411,13.157744,13.702565,14.998976,15.366566,14.519796,13.10195,12.704822,12.379898,12.251899,12.360206,12.668719,13.069129,13.180719,13.039591,12.914873,12.740924,12.117334,11.191795,11.401847,11.579078,11.30995,10.935796,10.630565,10.971898,11.451077,11.815386,12.091078,12.304411,12.668719,12.809847,12.35036,10.912822,11.332924,11.392001,11.503591,11.828514,12.294565,12.826258,13.912617,15.350155,16.718771,17.371899,16.456207,17.227488,18.031591,18.149744,17.792002,17.207796,16.420103,16.426668,17.61477,19.780924,19.990976,18.62236,16.666258,15.205745,15.42236,16.554668,16.528412,15.8884115,14.857847,13.344822,13.11836,12.780309,12.475078,12.570257,13.650052,12.885334,11.162257,10.368001,10.978462,12.071385,12.100924,11.490462,10.9456415,10.912822,11.59877,13.092104,14.565744,15.717745,16.108309,15.169642,14.907078,14.742975,14.8020525,15.556924,17.85436,16.899282,14.838155,14.368821,15.448617,15.317334,15.845745,18.596104,20.548925,20.850874,20.81149,20.145233,18.530462,18.70113,19.908924,17.920002,15.133539,13.705847,12.681848,11.815386,11.546257,11.35918,11.953232,12.507898,12.458668,11.480617,9.613129,8.749949,9.357129,10.975181,12.242052,8.835282,6.5411286,5.651693,5.6418467,5.146257,5.0477953,5.5630774,5.943795,5.9963083,6.0750775,7.194257,8.264206,8.710565,8.464411,7.9327188,7.9228725,7.9458466,7.830975,7.6143594,7.532308,8.067283,7.3321033,6.452513,5.9602056,5.7731285,5.408821,5.146257,5.221744,5.730462,6.629744,7.958975,8.841846,8.152616,6.304821,5.2611284,5.5893335,5.930667,6.514872,7.13518,7.131898,6.1046157,6.058667,6.2129235,6.1407185,5.7829747,4.713026,3.7973337,2.6289232,1.7788719,2.789744,3.239385,3.3542566,3.2525132,3.1343591,3.2820516,3.2656412,3.2525132,3.318154,3.1737437,2.1792822,1.142154,1.2898463,1.3357949,0.96492314,0.82379496,1.020718,0.86974365,0.8960001,1.1618463,1.2832822,1.6738462,1.3522053,1.7624617,2.6486156,2.0611284,3.6693337,2.9078977,4.0434875,6.491898,4.8311796,4.71959,5.333334,3.945026,1.270154,1.4506668,1.0962052,1.2307693,1.3095386,1.1979488,1.2012309,1.0896411,0.57764107,0.32820517,0.42338464,0.36430773,0.5218462,0.6629744,0.8730257,1.0535386,0.892718,0.5874872,0.69251287,0.9878975,1.5721027,2.8717952,2.1891284,1.2471796,1.595077,2.9801028,3.3542566,1.7099489,2.4418464,4.4242053,5.618872,3.1113849,2.3991797,3.692308,4.919795,5.031385,4.013949,3.0982566,3.9384618,4.3618464,3.8334363,3.4527183,3.8137438,3.889231,3.3542566,2.2547693,1.020718,2.297436,4.076308,6.3540516,8.595693,9.731283,9.235693,8.388924,7.939283,8.044309,8.260923,8.979693,10.6469755,11.644719,11.641437,11.592206,10.597744,10.440206,10.492719,10.387693,10.006975,11.0375395,10.889847,10.696206,10.902975,11.270565,10.541949,9.156924,8.490667,8.674462,8.5891285,6.186667,5.3202057,5.32677,5.481026,5.0051284,5.6287184,6.1997952,6.042257,5.297231,4.9362054,4.391385,4.6933336,5.034667,4.9985647,4.5522056,4.0336413,4.312616,4.0369234,2.9571285,1.913436,2.0709746,2.8455386,3.56759,4.0369234,4.516103,4.9493337,5.4514875,5.874872,6.2096415,6.5870776,6.3212314,5.425231,4.6605134,4.4701543,4.9788723,5.349744,5.435077,5.395693,5.3825645,5.533539,4.84759,4.667077,4.827898,4.9362054,4.3684106,5.1265645,5.0116925,4.8672824,4.9887185,5.1232824,4.8804107,4.8377438,5.228308,5.940513,6.5247183,7.9327188,9.350565,9.711591,9.084719,8.681026,8.556309,7.325539,6.235898,5.1856413,2.7044106,2.9801028,5.5072823,7.1515903,6.51159,3.9351797,8.021334,7.433847,7.0498466,8.28718,9.114257,6.918565,7.315693,12.412719,16.249437,4.827898,7.0826674,9.38995,9.777231,7.9163084,5.139693,8.904206,11.638155,10.962052,10.295795,18.881643,7.253334,8.146052,9.803488,7.529026,3.6726158,4.6834874,7.2237954,6.373744,3.2689233,5.106872,6.1407185,6.5903597,6.626462,6.7938466,7.9885135,5.5729237,3.2098465,2.4484105,3.5314875,5.3825645,5.9602056,6.5837955,6.928411,6.8693337,6.49518,7.906462,8.900924,9.091283,8.710565,8.635077,8.51036,8.946873,8.996103,8.425026,7.7325134,7.5585647,6.688821,5.8420515,5.805949,7.456821,7.171283,7.4371285,6.813539,5.7074876,6.3868723,5.989744,5.7501545,5.7501545,6.0356927,6.62318,4.9952826,5.2348723,6.0619493,6.6067696,6.416411,5.920821,5.904411,6.380308,6.9349747,6.738052,7.145026,6.764308,6.0324106,5.2512827,4.585026,4.240411,4.2568207,4.5587697,4.6900516,3.826872,2.9604106,2.4746668,2.5435898,3.0358977,3.5216413,2.7700515,2.7241027,2.806154,2.8258464,2.9768207,3.4756925,2.8816411,2.4746668,2.605949,2.6847181,2.7109745,2.6157951,2.4352822,2.2514873,2.172718,1.9889232,1.6705642,1.211077,0.7318975,0.49230772,0.57764107,0.8205129,1.1815386,1.5425643,1.7001027,2.0250258,2.1366155,2.0611284,1.9659488,2.1792822,2.3040001,2.2383592,2.3335385,2.6289232,2.8356924,2.9636924,3.0293336,2.9111798,2.6190772,2.297436,2.6453335,3.1606157,3.5380516,3.620103,3.4067695,3.6463592,3.7842054,3.6430771,3.3575387,3.3772311,3.9614363,4.778667,5.5729237,6.2884107,7.072821,6.806975,6.5280004,6.442667,6.550975,6.672411,6.6395903,6.4656415,6.11118,5.786257,5.937231,5.648411,5.5007186,5.805949,6.564103,7.4830775,8.011488,8.283898,8.050873,7.8014364,8.776206,9.865847,10.31877,10.112,9.540924,9.186462,8.474257,8.710565,9.478565,10.226872,10.28595,10.213744,11.155693,11.861334,12.130463,12.809847,12.521027,12.045129,12.379898,13.6008215,14.874257,13.63036,13.883078,14.191591,13.8075905,12.649027,13.190565,13.059283,12.911591,13.069129,13.51877,13.978257,13.705847,13.249642,13.157744,13.965129,14.267078,14.060308,13.696001,13.371078,13.144616,12.721231,12.2617445,11.756309,11.283693,11.024411,11.155693,11.175385,11.9171295,12.993642,12.78359,12.514462,12.63918,12.826258,12.731078,11.98277,11.707078,11.093334,10.880001,11.050668,10.840616,10.604308,10.630565,10.548513,10.164514,9.485129,8.467693,8.3823595,8.871386,9.8363085,11.444513,12.009027,11.999181,12.143591,12.524308,12.593232,13.019898,13.010053,12.793437,12.599796,12.635899,12.235488,11.877745,11.818667,11.926975,11.700514,11.920411,11.618463,11.579078,12.018872,12.580104,12.209231,12.219078,12.176412,12.045129,12.199386,1.394872,1.2406155,1.3489232,1.5392822,1.657436,1.5721027,1.6508719,1.6771283,1.5983591,1.5130258,1.6377437,1.9003079,1.8346668,2.1103592,2.6715899,2.7076926,2.861949,2.9604106,3.1507695,3.4231799,3.636513,3.3608208,3.8531284,4.46359,4.6867695,4.1452312,4.5095387,4.2896414,4.194462,4.516103,5.1298466,5.100308,5.280821,5.2480006,4.9920006,4.903385,5.907693,6.7938466,7.3485136,7.568411,7.6570263,8.4053335,8.598975,8.530052,8.595693,9.265231,9.278359,9.32759,9.642668,10.082462,10.134975,9.291488,8.805744,9.29477,10.213744,9.849437,10.758565,11.093334,11.155693,11.0145645,10.515693,10.774975,10.679795,10.886565,11.372309,11.431385,11.667693,11.37559,11.319796,11.772718,12.521027,13.584412,13.659899,13.354668,12.977232,12.524308,12.182976,11.766154,11.257437,10.8307705,10.866873,11.572514,11.972924,12.235488,12.356924,12.186257,12.179693,12.438975,12.58995,12.786873,13.725539,14.746258,15.120412,14.490257,13.197129,12.294565,12.0549755,12.458668,12.993642,13.361232,13.472821,13.003489,12.557129,12.212514,11.907283,11.460924,11.096616,11.730052,12.137027,11.881026,11.293539,11.1294365,11.451077,11.904001,12.301129,12.62277,12.921437,13.216822,13.456411,13.302155,12.133744,12.337232,12.235488,12.048411,11.88759,11.72677,12.248616,13.627078,15.140103,16.426668,17.522873,17.299694,17.234053,17.165129,17.168411,17.572104,17.427694,17.066668,17.024002,17.575386,18.730669,19.626669,18.930874,17.24718,15.353437,14.178463,15.9573345,16.23631,15.629129,14.470565,12.78359,11.969642,12.12718,12.511181,12.809847,13.11836,12.78359,11.10318,10.262975,10.804514,11.634872,11.552821,11.027693,10.584617,10.594462,11.257437,12.389745,13.656616,15.126975,16.341335,16.31836,16.311796,16.07877,15.66195,15.629129,17.092924,16.754873,14.880821,14.057027,14.592001,14.523078,15.025232,15.530668,16.167385,17.335796,19.689028,19.820309,18.271181,18.340103,19.74154,18.592821,17.161848,15.885129,14.562463,13.410462,13.08554,11.099898,10.564924,10.8767185,11.395283,11.457642,10.394258,9.4916935,9.399796,10.368001,12.245335,9.393231,7.072821,5.658257,5.139693,5.10359,5.172513,5.5696416,5.989744,6.2818465,6.4295387,7.3386674,8.362667,8.805744,8.493949,7.762052,8.123077,8.264206,8.3364105,8.4283085,8.549745,8.940309,8.129642,7.0826674,6.3277955,5.9634876,5.681231,5.2447186,5.0510774,5.402257,6.5247183,7.8080006,8.769642,8.28718,6.5772314,5.1987696,5.467898,5.6976414,6.636308,7.7948723,7.4732313,6.688821,6.1440005,5.8157954,5.5893335,5.2447186,4.1911798,3.3411283,2.4385643,1.9364104,2.9735386,2.9801028,2.9997952,3.0818465,3.1376412,2.937436,2.7503593,2.7602053,3.0227695,3.186872,2.484513,1.9823592,1.8149745,1.5097437,1.0962052,1.1093334,1.0929232,1.1848207,1.2438976,1.2964103,1.5688206,2.034872,4.138667,4.5456414,2.9965131,2.3105643,1.8642052,1.847795,3.9122055,6.5706673,5.221744,4.896821,4.1813335,2.5271797,0.8992821,1.7624617,0.92225647,0.8566154,1.0568206,1.1585642,0.90912825,0.92553854,0.63343596,0.47589746,0.5513847,0.6071795,0.75487185,0.8795898,0.86646163,0.7778462,0.86974365,0.7122052,0.8566154,1.1454359,1.595077,2.4188719,2.0775387,1.8510771,2.7569232,4.204308,4.013949,2.3433847,2.674872,3.764513,4.8672824,5.737026,4.532513,4.1747694,4.4373336,4.571898,3.3050258,2.9604106,3.4133337,2.9505644,2.15959,3.9089234,4.4734364,4.0402055,3.0752823,2.0808206,1.6114873,3.9975388,5.533539,7.0925136,8.546462,8.779488,7.785026,7.4075904,7.5979495,7.9097443,7.4863596,8.5661545,10.532104,12.015591,12.419283,11.936821,11.201642,10.633847,10.525539,10.729027,10.660104,11.418258,11.451077,11.418258,11.457642,11.1983595,10.81436,9.498257,8.546462,8.539898,9.330873,7.2861543,6.4590774,6.058667,5.664821,5.218462,6.1013336,6.8332314,6.5017443,5.3760004,4.9362054,4.31918,4.46359,4.778667,4.7458467,3.9253337,3.9417439,4.2994876,4.1517954,3.4198978,2.7864618,2.8225644,3.383795,3.8728209,4.128821,4.4307694,5.4580517,6.265436,6.550975,6.436103,6.4754877,6.2063594,5.684513,5.287385,5.277539,5.8125134,6.058667,5.730462,5.4449234,5.3727183,5.2512827,4.6834874,4.57518,4.84759,5.0674877,4.44718,5.10359,5.110154,4.9099493,4.8377438,5.1364107,4.493129,4.194462,4.1517954,4.315898,4.663795,6.5969234,7.8506675,8.907488,9.810052,10.14154,9.826463,9.622975,9.143796,7.9786673,5.6943593,2.8750772,4.6834874,6.5805135,6.5312824,5.0084105,8.835282,8.1755905,6.987488,6.8988724,7.2172313,6.2720003,7.53559,10.630565,11.953232,4.663795,8.868103,12.327386,11.904001,7.9524107,4.309334,11.149129,15.097437,14.729847,14.759386,26.016823,11.972924,12.087796,14.267078,11.720206,2.9571285,5.1626673,7.3419495,6.413129,4.0402055,6.62318,4.890257,4.6539493,4.70318,4.4734364,4.06318,5.605744,4.8016415,3.9909747,4.6112823,7.200821,5.874872,6.1341543,6.7117953,7.0104623,7.1056414,8.480822,9.206155,9.275078,9.045334,9.229129,9.340718,9.232411,8.713847,8.03118,7.8441033,8.139488,7.276308,6.117744,5.7632823,7.5454364,7.4863596,7.4240007,6.8233852,5.8125134,5.2020516,6.0160003,6.363898,6.3540516,6.3245134,6.8365135,5.297231,4.844308,5.425231,6.3212314,6.1538467,6.045539,5.7501545,5.8814363,6.439385,6.8233852,7.4797955,6.747898,5.8256416,5.07077,3.9844105,3.6496413,3.8301542,4.2601027,4.6276927,4.578462,3.5314875,2.5895386,2.3401027,2.8356924,3.6004105,3.1081028,3.121231,3.242667,3.3542566,3.6069746,3.764513,3.1770258,2.6945643,2.6026669,2.612513,2.5107694,2.231795,2.0676925,2.0578463,1.9954873,1.7165129,1.467077,1.1388719,0.7417436,0.42338464,0.5415385,0.8008206,1.086359,1.5425643,2.5435898,2.7700515,2.5009232,2.2449234,2.1858463,2.2022567,2.172718,2.176,2.4352822,2.7864618,2.681436,2.740513,2.4549747,2.2186668,2.1169233,1.9003079,2.1202054,2.4713848,2.7766156,3.0194874,3.3509746,3.4789746,3.5840003,3.4625645,3.2196925,3.2623591,3.8498464,4.2535386,4.594872,5.179077,6.482052,6.183385,5.9503593,6.0980515,6.498462,6.5805135,6.7150774,6.3212314,5.9470773,5.901129,6.2818465,6.2096415,5.5565133,5.612308,6.6560006,7.972103,7.6701546,7.5191803,7.27959,7.2237954,8.123077,9.481847,10.010257,9.649232,8.704,7.8670774,7.7292314,7.824411,8.5891285,9.747693,10.295795,10.5780525,11.395283,11.940104,12.084514,12.379898,11.9171295,11.0145645,10.768411,11.628308,13.384206,11.923694,12.99036,13.869949,13.59754,12.967385,13.5318985,13.197129,12.731078,12.550565,12.721231,13.252924,13.367796,13.124924,13.00677,13.892924,14.634667,14.483693,13.83713,13.180719,13.065847,12.245335,11.713642,11.792411,12.396309,13.013334,11.736616,10.70277,10.683078,11.460924,11.83836,11.907283,12.248616,12.324103,12.022155,11.657847,11.405129,10.981745,11.001437,11.336206,11.132719,10.387693,10.075898,10.167795,10.226872,9.399796,8.717129,8.55959,8.704,9.26195,10.699488,11.2672825,11.296822,11.392001,11.716924,11.98277,12.012309,11.782565,11.516719,11.457642,11.877745,11.447796,11.0605135,11.050668,11.32636,11.37559,11.431385,11.208206,11.286975,11.785847,12.3536415,12.071385,11.926975,11.641437,11.447796,12.104206,1.5491283,1.332513,1.3915899,1.4309745,1.4408206,1.6771283,1.7624617,1.6836925,1.5163078,1.3751796,1.4145643,1.8773335,1.7887181,2.2055387,3.1015387,3.3641028,3.6135387,4.0402055,4.1780515,4.0402055,4.1189747,4.135385,4.394667,4.565334,4.4274874,3.889231,4.0336413,4.2601027,4.3651285,4.394667,4.6539493,5.356308,5.832206,5.805949,5.3366156,4.7983594,5.2545643,6.413129,7.515898,8.14277,8.218257,7.955693,8.172308,8.923898,9.590155,8.891078,8.937026,8.966565,9.31118,9.993847,10.758565,10.325335,8.864821,8.553026,9.481847,9.672206,9.787078,10.226872,10.617436,10.692924,10.282667,10.312206,10.14154,10.345026,10.94236,11.395283,11.716924,11.930258,11.972924,11.963078,12.189539,13.272616,14.41477,14.404924,13.285745,12.360206,11.98277,11.487181,10.952206,10.594462,10.758565,11.122872,11.382154,11.651283,11.861334,11.759591,11.539693,11.74318,11.963078,12.360206,13.676309,14.358975,14.326155,13.774771,12.954257,12.156719,12.632616,13.298873,13.879796,14.135796,13.860104,13.08554,12.655591,12.25518,11.871181,11.795693,12.422565,13.233232,13.426873,12.918155,12.35036,12.320822,12.704822,13.029744,13.02318,12.6063595,13.138052,13.482668,13.935591,14.250668,13.653335,12.780309,12.517745,12.337232,12.012309,11.654565,11.858052,12.921437,13.935591,14.851283,16.469334,17.93641,18.054565,17.588514,17.427694,18.599386,17.913437,17.716515,17.266872,16.607182,16.587488,18.235079,18.146463,17.641027,16.91241,15.025232,16.068924,16.305231,15.596309,14.280207,13.1872835,12.140308,12.09436,12.658873,13.147899,12.576821,12.294565,11.313231,10.86359,11.221334,11.67754,11.58236,11.044104,10.781539,11.136001,12.058257,12.658873,13.200411,14.49354,16.357744,17.634462,17.729643,17.076513,16.190361,15.409232,14.8939495,15.199181,14.10954,13.512206,13.879796,14.28677,14.54277,14.313026,14.326155,15.028514,16.577642,17.7559,17.299694,17.811693,19.252514,18.924309,19.104822,18.28431,16.94195,15.842463,16.04595,12.662155,10.545232,10.089026,11.067078,12.616206,11.2672825,10.44677,9.93477,9.96759,11.218052,10.108719,8.165744,6.3540516,5.3202057,5.4153852,5.35959,5.5171285,5.8912826,6.314667,6.432821,7.4929237,8.326565,8.713847,8.52677,7.719385,8.188719,8.598975,9.088,9.626257,10.033232,9.980719,8.740103,7.515898,6.8332314,6.5280004,6.117744,5.428513,4.916513,4.972308,5.933949,7.177847,7.722667,7.5421543,6.747898,5.5893335,5.61559,5.943795,7.0367184,8.375795,8.474257,8.15918,6.774154,5.5171285,4.8607183,4.5489235,3.4855387,2.6486156,2.172718,2.1398976,2.5665643,2.4024618,2.353231,2.4418464,2.5337439,2.3138463,2.294154,2.4516926,2.5304618,2.5009232,2.5632823,2.937436,2.4648206,2.0053334,1.7920002,1.4309745,1.3653334,1.3915899,1.3981539,1.4605129,1.8510771,2.487795,8.116513,8.448001,3.8334363,5.2611284,3.1606157,1.4769232,2.0742567,4.1846156,4.381539,3.0720003,1.5261539,0.9616411,1.401436,1.6672822,0.96492314,0.65969235,0.74830776,0.9616411,0.76800007,0.56123084,0.69579494,0.8008206,0.81394875,0.9878975,1.0535386,1.0469744,0.8795898,0.69907695,0.88943595,0.9124103,1.0765129,1.2307693,1.4473847,2.0512822,1.9987694,2.5993848,3.948308,5.1331286,4.2305646,3.3903592,2.7011285,3.6004105,6.5050263,10.817642,7.003898,5.5171285,4.6769233,3.6004105,2.1989746,3.045744,3.5774362,2.7667694,1.7394873,3.7973337,4.1714873,3.767795,3.0949745,2.550154,2.4516926,5.435077,6.7117953,7.653744,8.546462,8.618668,7.778462,7.4699492,7.634052,7.768616,6.9349747,8.211693,10.213744,12.163283,13.423591,13.505642,12.576821,11.667693,11.067078,10.866873,10.981745,11.257437,11.634872,11.844924,11.920411,12.20595,11.32636,9.796924,8.963283,9.032206,9.068309,8.726975,7.8769236,7.13518,6.5739493,5.7074876,5.87159,6.6625648,6.5870776,5.5696416,4.95918,4.6769233,5.169231,5.5072823,5.080616,3.623385,4.414359,4.309334,3.9975388,3.8596926,3.9548721,3.56759,3.6594875,3.9154875,4.1911798,4.5390773,6.170257,7.131898,7.4240007,7.2303596,6.921847,6.7840004,6.416411,6.0717955,5.9963083,6.4065647,6.3507695,5.933949,5.671385,5.5532312,5.034667,4.8311796,4.97559,5.2315903,5.280821,4.7392826,4.9526157,5.0018463,4.7655387,4.5390773,5.0149746,4.266667,3.8728209,3.6791797,3.5741541,3.4855387,5.5893335,6.4754877,7.827693,9.613129,10.079181,10.328616,10.722463,10.049642,8.891078,9.636104,5.1889234,4.013949,4.20759,4.673641,5.10359,8.008205,9.094564,8.536616,6.8332314,4.824616,3.4198978,5.7829747,7.174565,6.6428723,7.026872,10.066052,11.201642,9.43918,6.1440005,5.034667,10.486155,16.636719,20.502975,23.16472,29.794464,16.705643,15.763694,17.959387,15.75713,3.1081028,4.0336413,5.034667,4.594872,3.754667,6.12759,5.973334,4.325744,3.239385,3.131077,2.7700515,6.2555904,6.6494365,5.586052,4.95918,6.9120007,4.7655387,4.9132314,5.973334,7.0367184,7.6570263,8.756514,8.953437,8.78277,8.78277,9.501539,10.272821,9.672206,8.39877,7.2664623,7.2205133,7.765334,7.3550773,6.547693,6.1341543,7.138462,7.24677,7.177847,6.7314878,5.943795,5.077334,6.3245134,6.6494365,6.6560006,6.698667,6.885744,5.4580517,4.562052,4.6145644,5.3366156,5.7435904,6.0947695,5.671385,5.5105643,6.0225644,6.9842057,7.453539,6.3310776,5.2676926,4.644103,3.5905645,3.3476925,3.623385,4.076308,4.522667,4.9132314,4.1682053,3.18359,2.6847181,2.8849232,3.4691284,3.5052311,3.2951798,3.367385,3.6890259,3.6693337,3.5905645,3.4067695,3.2131286,2.9735386,2.5435898,2.2580514,2.048,1.8576412,1.6804104,1.5786668,1.4276924,1.2504616,1.0568206,0.827077,0.49887183,0.7417436,0.9321026,1.142154,2.0808206,5.0871797,5.290667,3.3772311,2.1070771,2.1267693,1.9823592,2.0086155,2.1530259,2.4615386,2.7241027,2.4582565,2.5140514,2.0808206,1.785436,1.782154,1.7394873,1.6607181,1.7394873,1.847795,2.1464617,3.0752823,3.4756925,3.5807183,3.245949,2.7700515,2.8816411,3.370667,3.56759,3.9154875,4.6867695,5.973334,5.4383593,5.431795,5.618872,5.7764106,5.802667,5.9634876,5.8420515,5.910975,6.232616,6.4754877,6.4557953,6.0619493,6.0028725,6.6461544,8.011488,7.6077952,7.3714876,7.256616,7.3091288,7.6701546,8.746667,9.586872,9.396514,8.116513,6.4295387,7.0859494,7.381334,7.8080006,8.5891285,9.705027,10.673231,11.608616,12.176412,12.25518,11.926975,11.080206,10.696206,10.614155,10.696206,10.807796,10.581334,12.3766165,13.220103,12.586668,12.416001,13.522053,12.918155,12.251899,12.133744,12.156719,12.445539,13.072412,13.275898,13.184001,13.810873,14.70359,14.14236,12.967385,12.038565,12.258463,12.120616,11.936821,12.484924,13.53518,13.830565,12.560411,12.045129,12.002462,12.038565,11.625027,11.825232,12.028719,11.766154,11.250873,11.362462,10.837335,10.322052,10.374565,10.8767185,11.044104,10.781539,10.381129,10.213744,10.203898,9.826463,9.741129,9.127385,8.704,8.999385,10.328616,10.617436,10.617436,10.860309,11.434668,11.992617,11.926975,10.94236,10.308924,10.571488,11.536411,11.355898,10.935796,10.57477,10.456616,10.6469755,10.71918,10.988309,11.332924,11.657847,11.884309,11.877745,11.67754,11.418258,11.408411,12.1238985,1.7690258,1.4145643,1.2996924,1.2865642,1.3850257,1.7394873,2.0086155,1.7624617,1.8051283,2.1366155,1.9528207,2.0151796,1.9922053,2.3958976,3.1081028,3.387077,3.1803079,4.4373336,4.926359,4.315898,4.1813335,4.460308,4.706462,4.890257,4.900103,4.5456414,3.8137438,3.9614363,3.8695388,3.5052311,3.9220517,5.093744,5.5597954,5.976616,6.409847,6.3474874,7.177847,7.512616,7.8670774,8.218257,8.011488,7.4732313,7.072821,7.1647186,7.584821,7.643898,7.680001,7.939283,8.280616,8.805744,9.842873,9.537642,8.086975,7.5191803,8.011488,7.890052,8.766359,9.45559,9.626257,9.488411,9.780514,9.255385,9.547488,10.095591,10.84718,12.2387705,12.580104,12.885334,12.901745,12.822975,13.275898,14.299898,15.2155905,15.02195,13.801026,12.724514,11.762873,11.273847,10.998155,10.893129,11.122872,10.794667,11.234463,11.851488,12.11077,11.54954,11.0375395,11.067078,11.431385,12.051693,12.954257,13.29559,13.13477,12.553847,12.035283,12.452104,13.206975,13.459693,13.906053,14.434463,14.129231,13.581129,13.423591,13.052719,12.491488,12.406155,12.855796,13.682873,14.155488,13.948719,13.167591,12.973949,13.190565,13.036308,12.448821,12.068104,12.386462,12.530872,12.763899,13.115078,13.397334,11.808822,11.277129,11.264001,11.349334,11.21477,11.789129,12.1238985,12.393026,13.039591,14.785643,17.335796,18.5239,19.554462,20.371695,19.636515,19.026052,17.631182,16.354464,15.730873,15.914668,18.747078,20.086155,19.538054,17.795284,16.646564,18.064411,18.993233,17.713232,14.785643,13.075693,12.235488,13.029744,13.830565,13.833847,13.075693,11.674257,11.221334,11.136001,11.175385,11.444513,11.858052,11.369026,11.32636,12.009027,12.619488,13.180719,14.10954,15.346873,16.938667,19.026052,19.551182,18.668308,17.142155,15.504412,14.037334,14.099693,13.896206,14.102976,14.8020525,15.471591,15.179488,14.887385,14.76595,15.186052,16.722052,16.420103,16.643284,18.281027,20.5719,21.13313,20.424206,19.295181,18.36308,18.120207,18.950565,16.679386,12.826258,10.240001,9.980719,11.323078,10.003693,9.885539,9.872411,9.5835905,9.337437,9.412924,8.277334,7.066257,6.304821,5.8912826,5.3760004,5.5893335,5.874872,5.979898,6.042257,7.0925136,8.333129,8.835282,8.438154,7.765334,7.975385,8.208411,8.618668,9.32759,10.436924,9.777231,7.9458466,6.957949,7.1614366,7.24677,6.7610264,5.720616,4.716308,4.345436,5.2480006,6.1997952,6.5050263,6.5017443,6.38359,6.163693,6.042257,6.9743595,8.109949,8.900924,9.110975,8.851693,6.436103,4.716308,4.3684106,3.892513,2.8160002,2.4385643,2.4320002,2.674872,3.249231,2.284308,1.8149745,1.9495386,2.300718,1.9823592,2.5698464,2.6880002,2.6387694,2.7109745,3.1737437,3.0884104,2.5435898,2.2514873,2.2482052,1.9068719,2.0644104,1.7755898,1.7099489,1.9495386,1.9987694,4.0992823,8.323282,8.369231,6.7249236,14.647796,7.0793853,2.0939488,0.06235898,0.12143591,0.18379489,0.46276927,0.96492314,1.7099489,2.3138463,1.9823592,1.0666667,0.702359,0.50543594,0.47589746,0.97805136,0.8172308,1.1979488,1.7493335,2.0250258,1.5261539,1.3062565,0.9944616,0.9714873,1.1815386,1.1454359,0.8763078,1.0568206,1.4703591,1.8182565,1.7099489,2.8192823,2.9046156,4.1550775,5.8157954,4.1813335,4.3749747,3.8564105,7.13518,12.806565,13.564719,4.6539493,6.4623594,7.384616,4.1517954,1.847795,2.1136413,2.2547693,2.1464617,2.428718,4.516103,3.748103,3.242667,2.8717952,2.6453335,2.7306669,4.1714873,5.730462,6.7216415,7.1548724,7.752206,8.582564,8.011488,7.4371285,7.276308,6.957949,7.837539,9.760821,12.005745,13.636924,13.505642,12.576821,12.07795,10.998155,9.770667,10.28595,10.686359,10.880001,11.122872,11.805539,13.426873,11.365745,10.820924,10.834052,10.459898,8.789334,9.947898,8.763078,8.14277,8.293744,6.744616,5.4153852,5.9503593,6.5247183,6.2162056,5.0215387,5.21518,5.3825645,5.280821,4.8672824,4.31918,4.8049235,4.1124105,3.370667,3.1606157,3.5413337,3.501949,4.1911798,4.6769233,4.8311796,5.293949,5.8945646,6.931693,7.9983597,8.592411,8.116513,8.457847,8.152616,7.4141545,6.636308,6.3934364,6.173539,6.2194877,6.298257,6.048821,4.97559,4.2896414,4.5489235,5.21518,5.618872,4.95918,5.398975,5.618872,5.3202057,4.8311796,5.110154,4.453744,3.5840003,3.058872,3.0949745,3.570872,5.3037953,6.6527185,7.7259493,8.274052,7.6767187,8.480822,9.718155,9.7903595,8.779488,8.438154,8.195283,4.8016415,3.1343591,4.027077,4.273231,4.8344617,6.633026,7.939283,7.7292314,5.691077,5.4974365,4.788513,7.5487185,10.870154,4.97559,7.427283,6.265436,4.1714873,3.387077,5.7074876,4.97559,13.725539,21.40554,24.546463,26.77826,14.657642,12.580104,16.449642,18.025026,4.9296412,3.6824617,4.086154,3.9089234,2.733949,1.9528207,5.041231,4.604718,4.1846156,4.4800005,3.3575387,3.882667,3.748103,5.4449234,7.571693,4.8377438,4.7524104,5.58277,6.491898,7.145026,7.706257,8.805744,8.182155,7.8408213,8.388924,9.048616,8.999385,8.6580515,8.2904625,8.064001,8.024616,7.719385,7.259898,6.7183595,6.3934364,6.820103,6.294975,6.301539,6.1013336,5.5171285,4.9427695,5.907693,5.58277,5.7107697,6.629744,7.2631803,5.9930263,5.0904617,4.8640003,5.32677,6.196513,6.8299494,6.557539,6.245744,6.1440005,5.874872,5.533539,4.594872,3.9811285,3.6890259,2.8225644,2.3335385,2.8258464,3.442872,3.9253337,4.6080003,4.6933336,4.266667,3.8334363,3.6758976,3.8596926,3.7021542,3.515077,3.308308,3.2164104,3.508513,3.3641028,3.5380516,3.6102567,3.31159,2.5173335,2.3105643,2.1956925,1.7493335,1.1749744,1.2964103,1.273436,1.1552821,1.0535386,0.98461545,0.8992821,1.2406155,1.1716924,1.3259488,3.2196925,9.26195,10.873437,5.737026,2.0644104,2.0676925,1.9823592,2.0578463,2.028308,2.1136413,2.3105643,2.3958976,2.103795,1.654154,1.276718,1.0929232,1.1290257,1.3259488,1.3193847,1.276718,1.5622566,2.7470772,3.626667,3.7907696,3.3214362,2.7208207,2.930872,3.370667,3.3772311,3.5380516,4.020513,4.59159,4.312616,4.663795,4.890257,4.7622566,4.59159,4.420923,4.965744,5.7698464,6.3901544,6.377026,7.062975,6.9677954,6.675693,6.6428723,7.2172313,7.6931286,8.224821,8.43159,8.303591,8.195283,9.232411,9.242257,8.950154,8.28718,6.3934364,6.636308,7.1483083,7.8802056,8.641642,9.094564,9.009232,9.810052,10.9456415,11.69395,11.168821,10.400822,10.518975,10.725744,10.712616,10.650257,11.457642,12.461949,12.504617,11.54954,10.679795,12.842668,12.320822,11.398565,11.109744,11.23118,11.437949,11.930258,12.173129,12.33395,13.275898,13.679591,12.898462,11.851488,11.293539,11.85477,12.685129,12.721231,12.586668,12.281437,11.168821,11.414975,12.635899,13.4859495,13.161027,11.428103,11.45436,11.385437,10.935796,10.555078,11.460924,11.227899,10.758565,10.581334,10.765129,10.909539,12.278154,12.491488,11.457642,9.862565,9.156924,9.458873,9.353847,9.494975,9.987283,10.390975,10.453334,10.338462,10.407386,10.906258,11.992617,12.248616,10.840616,9.803488,9.984001,11.047385,11.949949,11.224616,10.010257,9.3768215,10.328616,9.708308,10.266257,10.870154,11.076924,11.139283,11.592206,11.703795,11.808822,11.989334,12.100924,1.5753847,1.3193847,1.1913847,1.0962052,1.1881026,1.8740515,1.8412309,1.7526156,1.9790771,2.300718,1.9528207,2.169436,1.9167181,2.5206156,3.8596926,4.3749747,4.089436,4.516103,4.525949,4.263385,5.146257,5.464616,5.146257,4.460308,3.9318976,4.338872,4.204308,5.0609236,4.785231,3.5774362,3.9811285,5.1626673,6.3277955,6.944821,6.872616,6.370462,6.616616,7.4436927,8.434873,9.104411,8.87795,7.2861543,6.87918,6.9710774,7.145026,7.253334,7.515898,6.8988724,6.692103,7.4896417,9.170052,8.484103,8.323282,8.6580515,9.304616,9.915077,9.796924,9.40636,9.554052,10.394258,11.428103,10.289231,10.066052,10.151385,10.200616,10.125129,11.736616,12.960821,13.328411,13.075693,13.115078,13.371078,14.106257,14.001232,13.157744,13.128206,12.028719,11.59877,10.9456415,10.134975,10.220308,10.722463,11.008,11.250873,11.464206,11.539693,11.493745,11.0375395,10.712616,10.758565,11.122872,11.250873,11.414975,11.608616,11.956513,12.731078,13.430155,13.74195,14.057027,14.313026,14.007796,13.925745,13.272616,12.58995,12.104206,11.746463,11.85477,12.530872,13.065847,13.223386,13.252924,12.970668,12.704822,12.36677,12.002462,11.789129,11.628308,11.674257,11.733335,11.848206,12.288001,10.71918,10.482873,10.660104,10.870154,11.250873,11.201642,10.712616,10.683078,11.602052,13.551591,17.138874,19.626669,21.06749,21.62872,21.579489,19.718565,17.69354,15.832617,14.828309,15.744001,21.280823,22.800411,20.844309,17.913437,18.454975,17.749334,19.242668,19.43631,17.266872,14.102976,12.967385,12.219078,12.425847,13.098668,12.675283,10.9686165,10.476309,10.571488,10.929232,11.529847,11.730052,11.808822,12.081232,12.5374365,12.813129,12.642463,13.659899,14.916924,16.262566,18.320412,18.894772,18.297438,17.09949,15.77354,14.710155,14.644514,14.795488,14.309745,13.607386,14.385232,15.117129,14.437745,14.667488,16.292105,17.956104,17.066668,16.90913,18.297438,20.168207,19.606976,17.473642,17.007591,16.25272,16.101746,20.28308,20.266668,16.836924,13.003489,10.7158985,10.857026,10.272821,9.869129,9.800206,9.80677,9.193027,8.562873,7.968821,7.6110773,7.3025646,6.4754877,5.612308,5.8289237,6.052103,5.933949,5.858462,5.874872,6.961231,8.011488,8.39877,7.962257,7.1844106,7.1056414,7.4896417,8.100103,8.704,8.2215395,6.8955903,6.304821,6.7314878,7.138462,6.4065647,5.474462,4.644103,4.309334,4.969026,5.228308,5.7665644,6.301539,6.636308,6.6395903,6.7905645,7.4240007,8.208411,8.697436,8.329846,8.129642,6.701949,5.622154,5.179077,4.378257,3.3345644,2.9768207,2.8553848,2.7175386,2.5304618,2.228513,2.2186668,2.1333334,2.03159,2.3991797,2.740513,2.300718,2.4746668,3.0523078,2.1989746,2.1891284,1.7394873,2.100513,3.6102567,5.691077,3.3214362,1.8215386,1.2438976,1.4211283,1.9364104,13.548308,9.156924,5.930667,8.008205,6.5083084,4.31918,2.2514873,1.6016412,1.7952822,0.40369233,0.83035904,0.8763078,1.2012309,1.6672822,1.3489232,0.73517954,0.7450257,0.9353847,1.1913847,1.719795,3.367385,2.9210258,2.166154,1.8806155,1.8182565,1.276718,1.3522053,1.5688206,1.463795,0.6071795,1.1782565,1.3259488,1.7427694,2.2022567,1.5753847,1.7394873,2.1136413,3.879385,5.8781543,4.630975,5.228308,5.3136415,6.009436,7.069539,6.889026,3.7973337,4.9952826,5.937231,4.9526157,3.249231,2.2383592,5.0051284,5.293949,3.4756925,6.518154,5.3005133,3.5478978,3.3903592,3.9942567,1.5589745,3.6069746,5.681231,6.7774363,6.73477,6.23918,7.6143594,7.5454364,7.568411,7.896616,7.433847,7.7259493,10.089026,12.130463,12.773745,12.258463,11.808822,11.204924,10.44677,9.8592825,10.089026,11.126155,11.762873,12.081232,12.25518,12.560411,11.825232,10.962052,10.463181,10.121847,9.045334,10.594462,9.816616,9.350565,9.412924,7.7948723,6.961231,6.245744,6.157129,6.308103,5.421949,5.297231,5.21518,5.356308,5.5204105,5.1364107,4.7655387,4.0992823,4.0434875,4.384821,3.7973337,4.453744,4.667077,4.8311796,5.0051284,4.9526157,5.865026,7.4108725,8.621949,8.940309,8.241231,8.612103,8.172308,7.466667,6.941539,6.941539,6.7117953,6.6461544,6.449231,5.920821,4.962462,5.146257,5.2644105,5.106872,4.841026,5.0215387,5.333334,4.890257,4.138667,3.6463592,4.1222568,4.4406157,3.9844105,3.2886157,2.917744,3.4592824,3.945026,5.5007186,6.770872,7.0498466,6.294975,7.8145647,8.2904625,8.592411,8.792616,8.155898,8.060719,7.499488,5.671385,3.7054362,4.663795,5.0084105,7.1056414,8.070564,7.529026,7.6209235,8.546462,8.004924,9.110975,10.036513,3.9745643,6.436103,6.11118,5.0084105,4.2994876,4.3027697,9.330873,9.990565,14.001232,19.124514,13.144616,7.056411,10.331899,14.690463,13.945437,4.0008206,5.664821,4.634257,4.2830772,4.6276927,2.3302567,3.1934361,3.6135387,3.8367183,3.9417439,3.8465643,3.82359,4.716308,5.7435904,6.2129235,5.5204105,5.72718,6.3179493,6.8266673,7.1187696,7.387898,8.448001,7.9195905,7.3616414,7.77518,9.596719,8.641642,7.4436927,6.944821,7.4371285,8.562873,7.857231,7.2172313,7.131898,7.2664623,6.4557953,6.3901544,6.5378466,6.6067696,6.4032826,5.858462,5.651693,5.0543594,4.841026,5.113436,5.297231,4.9854364,4.7327185,4.709744,5.2381544,6.76759,6.564103,5.796103,5.169231,4.916513,4.8114877,4.900103,4.092718,3.6036925,3.5478978,2.9440002,3.4921029,3.5314875,3.639795,4.059898,4.706462,4.352,4.210872,4.0303593,3.754667,3.5052311,3.4166157,3.7973337,4.086154,4.141949,4.2305646,3.761231,3.2623591,3.0752823,3.1934361,3.249231,3.0523078,2.7864618,2.3138463,1.7493335,1.4309745,1.3292309,1.2898463,1.2931283,1.2832822,1.1684103,0.9944616,0.98461545,2.1530259,4.46359,6.8332314,5.152821,3.0260515,1.9823592,2.156308,2.2777438,2.409026,2.2186668,2.169436,2.284308,2.176,1.5327181,1.3686155,1.2406155,1.020718,0.90912825,1.1520001,1.3718976,1.5261539,1.7296412,2.2580514,3.058872,3.5774362,3.4822567,3.0096412,2.9538465,3.3345644,3.564308,3.9778464,4.4865646,4.5817437,4.5456414,4.824616,5.0609236,5.3005133,6.009436,5.5926156,5.5991797,5.796103,5.805949,5.110154,6.0750775,6.1997952,6.2030773,6.377026,6.5706673,7.719385,8.411898,8.937026,9.232411,8.891078,8.726975,8.152616,8.123077,8.539898,8.247795,7.5552826,7.5520005,8.293744,9.3078985,9.593436,8.982975,9.015796,8.969847,8.841846,9.350565,10.679795,10.725744,10.604308,10.860309,11.444513,11.136001,10.971898,11.008,11.096616,10.86359,10.604308,11.283693,11.82195,11.897437,11.949949,11.004719,11.588924,12.314258,12.458668,11.98277,11.759591,11.674257,11.772718,12.058257,12.504617,12.63918,12.337232,11.871181,11.808822,13.013334,13.216822,13.157744,12.901745,12.150155,10.220308,10.272821,10.735591,11.040821,11.155693,11.58236,11.211488,10.210463,9.458873,9.544206,10.774975,11.34277,11.707078,11.657847,11.18195,10.473026,9.947898,10.233437,10.341744,9.990565,9.622975,9.96759,10.354873,10.564924,10.752001,11.467488,12.133744,11.565949,10.916103,10.79795,11.303386,11.113027,10.706052,10.249847,10.023385,10.440206,9.193027,9.212719,9.895386,10.781539,11.565949,12.163283,12.612924,13.046155,13.190565,12.379898,1.6738462,1.7099489,1.5983591,1.4211283,1.3751796,1.7690258,1.7394873,1.7985642,2.044718,2.422154,2.7044106,2.2350771,2.3466668,3.0194874,3.9548721,4.588308,5.0642056,4.955898,4.8147697,4.9493337,5.431795,5.3792825,5.5302567,5.2020516,4.57518,4.6802053,5.0215387,5.802667,5.602462,4.571898,4.417641,4.644103,5.330052,5.9963083,6.452513,6.816821,7.318975,8.182155,8.989539,9.317744,8.720411,7.463385,6.820103,6.813539,7.1548724,7.24677,7.4108725,7.1023593,6.8397956,7.181129,8.700719,7.9195905,8.136206,8.602257,9.061745,9.744411,9.31118,8.828718,9.124104,10.085744,10.66995,9.947898,10.118565,10.292514,10.105436,9.724719,10.525539,11.411694,12.294565,13.078976,13.653335,13.745232,13.515489,12.816411,11.913847,11.506873,10.804514,11.011283,11.063796,10.561642,9.77395,10.269539,10.341744,10.597744,11.149129,11.59877,11.739899,11.2672825,10.975181,10.9456415,10.555078,11.011283,11.050668,11.1064625,11.516719,12.5374365,13.082257,13.590976,13.974976,14.158771,14.096412,13.919181,13.049437,12.393026,12.245335,12.2847185,12.288001,12.540719,12.57354,12.3306675,12.166565,11.700514,11.421539,11.0145645,10.55836,10.509129,10.089026,10.236719,10.289231,10.262975,10.86359,10.003693,9.622975,9.622975,9.974154,10.729027,10.985026,10.817642,10.94236,11.736616,13.252924,16.439796,17.47036,18.002052,18.694565,19.236105,18.087385,17.749334,17.125746,16.216616,16.114874,19.236105,20.552206,20.696617,20.676924,21.897848,20.54236,19.748104,18.91118,17.604925,15.586463,13.909334,12.534155,12.340514,12.996924,12.977232,11.546257,11.490462,11.874462,12.232206,12.557129,11.392001,11.533129,11.923694,12.06154,11.992617,12.944411,14.004514,15.120412,16.617027,19.19672,19.67918,19.30831,18.409027,17.34236,16.479181,15.891693,16.269129,16.787693,16.433231,13.994668,13.774771,13.24636,13.636924,14.916924,15.793232,15.904821,15.921232,16.361027,17.152,17.604925,16.534975,16.600616,16.508718,16.561232,18.65518,21.526976,20.256823,16.436514,12.386462,11.145847,11.444513,10.200616,9.452309,9.521232,9.019077,8.425026,8.152616,8.086975,7.8473854,6.7971287,6.0192823,5.8945646,5.943795,5.8880005,5.6385646,5.5991797,6.3376417,7.5454364,8.562873,8.369231,7.9885135,7.433847,7.3747697,7.837539,8.188719,7.702975,6.554257,6.042257,6.4295387,6.954667,6.226052,5.4514875,4.637539,4.194462,4.916513,5.2644105,5.7468724,6.3245134,6.7282057,6.4656415,6.7150774,7.2664623,7.8539495,8.136206,7.6767187,7.1187696,6.245744,5.412103,4.71959,4.023795,3.9023592,3.6758976,3.4921029,3.3312824,3.0194874,2.6420515,2.537026,2.2580514,1.910154,2.1464617,1.9856411,2.1497438,3.0030773,4.027077,3.8038976,4.3060517,4.1583595,4.378257,4.781949,4.010667,2.2153847,1.3357949,0.95835906,2.6453335,9.915077,10.039796,7.3780518,8.03118,11.605334,11.188514,3.7284105,1.8510771,1.6705642,1.1946667,0.33805132,0.8533334,1.1060513,1.1290257,1.0502565,1.1093334,0.9878975,1.1782565,1.4572309,1.8313848,2.5665643,3.620103,3.4133337,2.8882053,2.3236926,1.3718976,1.7788719,1.8510771,1.6935385,1.4211283,1.1520001,1.3620514,1.719795,1.6902566,1.5556924,2.4484105,2.9538465,3.4198978,4.2568207,4.9329233,3.9680004,6.2884107,6.088206,6.5936418,7.2631803,3.7710772,4.31918,5.684513,6.0816417,5.044513,3.4264617,2.930872,5.4186673,7.3353853,7.8145647,8.667898,5.431795,3.4330258,2.7569232,2.5665643,1.083077,3.698872,5.2676926,6.3573337,6.8430777,5.914257,6.872616,6.741334,7.450257,8.759795,8.267488,8.326565,10.456616,12.383181,13.072412,12.724514,11.283693,10.256411,10.056206,10.453334,10.59118,10.893129,11.316514,11.67754,11.913847,12.087796,12.1238985,11.565949,11.0375395,10.594462,9.741129,11.280411,10.778257,10.154668,9.856001,8.835282,7.788308,6.6395903,6.1078978,6.0783596,5.5893335,5.579488,5.3366156,5.4580517,5.7435904,5.211898,5.0215387,3.8695388,3.6660516,4.345436,3.8596926,4.565334,4.785231,5.2480006,5.8912826,5.8912826,6.2063594,7.351795,8.274052,8.470975,7.9786673,7.7981544,7.529026,7.069539,6.547693,6.301539,6.3343596,6.7840004,6.633026,5.83877,5.333334,5.7074876,5.6352825,5.2709746,5.0149746,5.4941545,5.041231,4.4767184,4.164923,4.161641,4.197744,4.266667,3.8662567,3.2787695,2.9571285,3.5249233,3.4231799,4.5489235,5.1987696,5.0609236,5.182359,6.314667,6.8627696,7.5454364,8.205129,7.8112826,7.9852314,8.077128,6.9710774,5.1200004,4.5489235,6.170257,7.351795,7.4896417,7.204103,8.339693,9.432616,8.024616,7.955693,8.989539,6.816821,8.310155,8.224821,6.931693,5.074052,3.5774362,9.540924,9.468719,12.402873,17.670565,14.887385,7.138462,9.895386,13.331694,11.670976,3.18359,5.3792825,5.8223596,5.277539,4.5489235,4.5029745,4.7524104,4.453744,4.2535386,4.273231,4.1222568,3.370667,4.076308,4.7327185,4.7622566,4.529231,6.0324106,6.6592827,6.485334,6.0225644,6.2096415,7.640616,7.857231,7.7981544,8.021334,8.681026,8.018052,7.4010262,6.8463597,6.921847,8.723693,8.182155,7.2270775,6.803693,6.7840004,5.9602056,6.193231,6.052103,6.088206,6.3868723,6.5378466,5.612308,5.2676926,5.0084105,4.6244106,4.1846156,4.132103,3.9318976,3.9581542,4.529231,5.904411,5.0149746,4.7556925,4.650667,4.5390773,4.601436,5.0904617,4.1189747,3.383795,3.383795,3.4330258,4.325744,3.9187696,3.8465643,4.325744,4.161641,4.073026,4.013949,3.8498464,3.6004105,3.446154,3.3345644,3.6562054,3.9220517,3.9647183,3.9417439,3.892513,3.0949745,2.6912823,2.9604106,3.3247182,3.3050258,3.245949,3.0030773,2.5271797,1.8576412,1.657436,1.2471796,1.0601027,1.148718,1.1815386,0.98461545,1.1881026,2.0611284,3.259077,3.817026,2.5829747,1.9528207,1.8904617,2.1300514,2.1858463,2.8882053,2.6880002,2.3138463,2.0775387,1.8740515,1.5360001,1.3686155,1.214359,1.014154,0.80738467,0.8467693,1.0272821,1.404718,1.8149745,1.8806155,2.6322052,3.5347695,3.895795,3.623385,3.2065644,3.308308,3.4133337,3.6102567,3.9187696,4.266667,4.466872,4.7392826,5.1200004,5.477744,5.5105643,5.4449234,5.7829747,5.8945646,5.7501545,5.907693,6.6395903,6.1768208,6.170257,6.7085133,6.3442054,7.515898,8.283898,8.763078,9.097847,9.458873,8.487385,8.054154,8.096821,8.241231,7.778462,8.139488,8.65477,9.186462,9.5835905,9.6754875,9.252103,9.084719,8.65477,8.165744,8.546462,9.156924,9.728001,10.28595,10.8767185,11.569232,11.057232,10.689642,10.423796,10.151385,9.682052,9.137232,10.256411,11.16554,11.237744,11.113027,10.066052,10.299078,11.132719,11.733335,11.145847,10.94236,11.168821,11.831796,12.714667,13.377642,13.305437,13.092104,12.603078,12.530872,14.41477,15.783386,14.55918,12.642463,11.099898,10.148104,9.842873,10.423796,10.870154,10.8996935,10.971898,11.300103,11.139283,10.843898,10.834052,11.611898,11.890873,11.920411,11.720206,11.306667,10.692924,10.656821,11.057232,11.250873,10.857026,9.731283,9.905231,10.233437,10.305642,10.43036,11.638155,12.182976,11.746463,11.369026,11.441232,11.697231,11.644719,11.063796,10.390975,9.96759,10.036513,9.540924,9.563898,9.895386,10.381129,10.912822,11.644719,12.173129,12.921437,13.423591,12.340514,1.7329233,1.9035898,1.8806155,1.8346668,1.785436,1.5885129,1.7526156,1.8116925,2.03159,2.4549747,2.868513,2.156308,2.7470772,3.4789746,3.9154875,4.3716927,5.2480006,5.21518,5.139693,5.3727183,5.7501545,5.356308,5.605744,5.677949,5.32677,4.857436,5.356308,5.8453336,5.835488,5.218462,4.273231,4.46359,4.7425647,5.2480006,6.045539,7.1483083,7.958975,8.598975,8.868103,8.661334,7.955693,7.213949,6.6395903,6.701949,7.24677,7.509334,7.059693,7.0957956,7.0367184,7.02359,7.9130263,7.8112826,8.008205,8.36595,8.786052,9.199591,9.012513,8.979693,9.189744,9.508103,9.570462,9.747693,10.151385,10.308924,10.059488,9.5606165,9.741129,10.177642,11.0605135,12.166565,12.885334,12.560411,11.959796,11.385437,10.86359,10.164514,9.793642,9.990565,10.289231,10.266257,9.517949,9.521232,9.396514,9.846154,10.735591,11.073642,11.45436,11.2672825,11.119591,10.994873,10.256411,11.067078,11.428103,11.739899,12.179693,12.708103,12.914873,13.302155,13.607386,13.682873,13.499078,13.078976,12.363488,11.910565,11.874462,12.025436,11.943385,12.104206,12.018872,11.634872,11.32636,10.686359,10.305642,9.93477,9.6754875,9.980719,9.593436,9.573745,9.458873,9.301334,9.662359,9.501539,9.242257,9.156924,9.45559,10.308924,10.9226675,11.011283,11.303386,12.074668,13.11836,14.976001,15.05477,15.264822,16.229744,17.289848,17.194668,17.99549,18.313848,17.769028,16.968206,18.067694,18.668308,19.570873,20.982155,22.514874,21.028105,18.930874,17.499899,16.922258,16.305231,15.00554,13.689437,13.4629755,14.116103,14.112822,12.891898,12.481642,12.409437,12.458668,12.685129,11.516719,11.897437,12.47836,12.553847,12.035283,13.341539,14.267078,15.176207,16.692514,19.695591,20.027079,19.705437,19.06872,18.405745,17.962667,16.607182,17.024002,18.546873,19.006361,14.720001,12.95754,12.652308,13.108514,13.718975,13.98154,15.356719,15.698052,15.126975,14.5263605,15.537232,16.026258,17.194668,17.801847,17.64431,17.575386,21.297232,22.964514,21.123283,16.512001,12.084514,12.6063595,10.955488,9.609847,9.238976,8.736821,8.641642,8.598975,8.379078,7.8112826,6.7840004,6.4656415,6.117744,5.970052,5.976616,5.8157954,5.664821,6.229334,7.4043083,8.539898,8.441437,8.293744,7.5421543,7.2336416,7.6668725,8.395488,7.6077952,6.6461544,6.088206,6.1472826,6.6625648,6.193231,5.5991797,4.818052,4.263385,4.818052,5.349744,5.8486156,6.36718,6.7216415,6.47877,6.941539,7.387898,7.752206,7.8506675,7.387898,6.445949,5.7829747,5.028103,4.2436924,3.9286156,4.381539,4.069744,3.7152824,3.511795,3.114667,2.5829747,2.4516926,2.172718,1.7755898,1.8412309,1.7394873,2.5009232,3.1606157,3.5347695,4.2240005,6.298257,5.8256416,4.9788723,4.1485133,1.9396925,1.2504616,1.142154,2.9243078,6.9087186,12.412719,5.0510774,7.5585647,12.993642,16.44636,15.061335,3.9384618,2.0151796,1.7788719,0.5546667,0.5284103,0.7253334,1.1158975,1.1355898,0.8730257,1.0666667,1.6672822,2.03159,2.678154,3.5249233,3.9023592,4.0369234,3.8006158,3.2853336,2.4385643,1.083077,2.034872,1.7132308,1.467077,1.6246156,1.5097437,1.785436,1.7723079,1.7362052,2.0053334,2.9833848,4.325744,5.074052,4.906667,4.4242053,5.139693,6.875898,7.276308,7.8834877,7.8736415,4.082872,3.7021542,4.571898,4.916513,4.46359,4.4274874,3.9023592,4.923077,7.634052,10.555078,10.571488,6.189949,3.2886157,1.785436,1.2307693,0.8336411,4.135385,5.156103,5.907693,6.7150774,6.2129235,6.5050263,6.23918,7.0859494,8.661334,8.536616,8.648206,10.233437,11.910565,12.921437,13.111795,11.529847,10.358154,10.266257,10.880001,10.765129,10.450052,10.57477,10.9686165,11.431385,11.72677,12.028719,11.848206,11.431385,11.053949,11.011283,12.084514,12.104206,11.437949,10.387693,9.18318,8.162462,7.256616,6.747898,6.482052,5.8453336,5.6943593,5.408821,5.402257,5.5630774,5.2480006,4.893539,3.8596926,3.3641028,3.748103,4.4832826,5.2709746,5.674667,6.419693,7.351795,7.4240007,6.76759,7.351795,7.8473854,7.748924,7.3714876,6.810257,6.6428723,6.6034875,6.4656415,6.038975,5.989744,6.692103,6.6494365,5.874872,5.8847184,5.7698464,5.5893335,5.284103,5.0543594,5.353026,4.716308,4.204308,4.2371287,4.5489235,4.1714873,3.8432825,3.4067695,2.9735386,2.8127182,3.370667,3.6660516,4.417641,4.6145644,4.4077954,5.10359,5.21518,5.8518977,6.806975,7.4929237,6.928411,7.3583593,8.306872,8.267488,6.7971287,4.5390773,5.6254363,6.0685134,6.3507695,6.803693,7.634052,9.032206,9.07159,7.936001,6.7577443,7.5979495,9.120821,8.4972315,7.6996927,7.197539,5.970052,8.530052,10.459898,14.969437,20.26995,19.590565,8.595693,7.9917955,9.856001,9.101129,3.43959,4.7655387,6.882462,6.518154,4.4340515,5.4514875,5.4908724,4.598154,3.9876926,3.9876926,4.0500517,3.4592824,4.1780515,5.031385,5.2578464,4.535795,5.297231,5.605744,5.3103595,4.8836927,5.4153852,6.5903597,7.3321033,7.955693,8.339693,7.9327188,7.5552826,7.3058467,6.7807183,6.6067696,8.418462,7.837539,7.0432825,6.626462,6.498462,5.8814363,5.687795,5.3891287,5.543385,6.1013336,6.4032826,5.4875903,5.431795,5.280821,4.634257,3.6594875,3.3444104,3.249231,3.4625645,3.9680004,4.6605134,4.0336413,4.204308,4.2929235,4.1682053,4.4307694,5.031385,4.3552823,3.639795,3.5183592,4.0303593,4.9296412,4.578462,4.457026,4.650667,3.8498464,4.128821,4.089436,3.7710772,3.367385,3.255795,3.0687182,3.2754874,3.383795,3.3378465,3.515077,3.8400004,3.0720003,2.556718,2.6322052,2.6453335,2.9571285,3.259077,3.2754874,2.8980515,2.169436,1.7263591,1.1290257,0.84348726,0.892718,0.88287187,1.083077,1.3522053,1.5491283,1.6278975,1.6443079,1.4441026,1.5753847,1.8084104,1.9528207,1.8248206,3.0424619,3.0030773,2.4320002,1.8773335,1.7165129,1.6082052,1.6311796,1.585231,1.3456411,0.86317956,0.9353847,0.93866676,1.276718,1.8182565,1.8740515,2.3138463,3.18359,3.692308,3.6758976,3.5905645,3.5183592,3.3509746,3.308308,3.495385,3.889231,4.312616,4.772103,5.1889234,5.402257,5.1331286,5.47118,6.1013336,6.1538467,5.930667,6.9152827,7.1680007,6.7117953,6.7085133,7.056411,6.4000006,7.0925136,7.6307697,8.096821,8.681026,9.672206,7.939283,7.752206,8.008205,8.008205,7.4436927,8.533334,9.350565,9.609847,9.465437,9.527796,9.462154,9.350565,8.910769,8.303591,8.12636,7.824411,8.598975,9.616411,10.397539,10.807796,10.650257,10.502565,10.210463,9.737847,9.176616,8.779488,9.586872,10.06277,9.8363085,9.691898,9.222565,9.117539,9.705027,10.541949,10.417232,10.266257,10.525539,11.339488,12.4685135,13.292309,13.098668,13.482668,13.938873,14.296617,14.70359,15.333745,13.948719,11.946668,10.55836,10.837335,10.049642,10.374565,10.729027,10.686359,10.489437,11.313231,11.848206,11.936821,11.792411,12.032001,12.488206,12.281437,11.703795,11.126155,11.017847,10.86359,11.004719,11.395283,11.516719,10.397539,10.075898,10.164514,10.131693,10.194052,11.339488,12.038565,11.690667,11.273847,11.218052,11.392001,12.022155,11.67754,10.893129,10.059488,9.419488,9.478565,9.6754875,9.911796,10.102155,10.203898,10.95877,11.602052,12.409437,13.052719,12.586668,1.5458462,1.719795,1.8248206,2.028308,2.1366155,1.6180514,1.9298463,1.8149745,1.8970258,2.2350771,2.3171284,2.1464617,3.0687182,3.7940516,3.9220517,3.9351797,4.650667,5.1167183,5.2053337,5.2742567,6.173539,5.835488,5.5926156,5.5597954,5.4613338,4.6539493,5.146257,5.579488,5.786257,5.4383593,4.0303593,4.8016415,5.110154,5.402257,6.0225644,7.210667,7.9163084,8.211693,8.01477,7.499488,7.0892315,6.3245134,6.232616,6.6461544,7.3025646,7.830975,6.9021544,6.8365135,6.7840004,6.567385,6.665847,7.4797955,7.5946674,7.975385,8.677744,8.87795,9.07159,9.4457445,9.360411,8.920616,8.982975,9.760821,10.023385,10.026668,9.816616,9.235693,9.435898,9.691898,10.105436,10.581334,10.820924,9.938052,9.833026,10.059488,10.184206,9.764103,9.429334,8.946873,8.763078,8.917334,9.025641,8.681026,8.605539,9.284924,10.299078,10.30236,10.781539,10.94236,10.971898,10.827488,10.256411,11.063796,11.956513,12.842668,13.364513,12.914873,12.839386,12.905026,12.960821,12.819694,12.258463,11.930258,11.54954,11.201642,10.932513,10.748719,10.532104,10.893129,11.162257,11.113027,10.965334,10.338462,9.744411,9.442462,9.5835905,10.217027,10.112,9.6984625,9.31118,9.104411,9.065026,9.18318,9.281642,9.291488,9.412924,10.108719,10.617436,10.47959,10.860309,11.926975,12.836103,13.51877,13.948719,14.739694,15.96718,17.168411,17.536001,18.002052,18.215385,18.051283,17.604925,18.609232,18.579693,18.277744,18.477951,19.961437,18.688002,17.273438,16.400412,16.190361,16.200207,15.75713,14.710155,14.523078,15.238565,15.442053,14.260514,12.882052,11.769437,11.234463,11.447796,11.687386,12.855796,13.892924,14.152206,13.397334,13.794462,14.352411,15.041642,16.226463,18.661745,18.868515,18.596104,18.38277,18.428719,18.58954,16.820515,16.768002,17.98236,18.648617,15.576616,13.082257,12.842668,13.193847,13.397334,13.633642,15.494565,16.154257,15.192616,13.676309,14.148924,15.589745,17.824821,18.770052,18.225233,17.877335,20.33231,24.054155,25.465437,22.514874,14.670771,13.725539,12.173129,10.768411,9.731283,8.736821,9.173334,9.186462,8.54318,7.450257,6.554257,6.747898,6.5411286,6.2752824,6.193231,6.416411,5.8945646,6.4689236,7.5421543,8.438154,8.39877,7.7357955,7.1089234,6.948103,7.522462,8.92718,7.890052,7.131898,6.4689236,6.0291286,6.226052,6.173539,5.7435904,5.0674877,4.516103,4.713026,5.225026,5.8847184,6.3540516,6.567385,6.7314878,7.453539,7.817847,8.041026,8.04759,7.4863596,6.308103,5.4843082,4.7491283,4.1780515,4.1813335,4.4701543,3.9548721,3.4527183,3.1277952,2.4746668,2.1103592,2.1136413,1.9561027,1.6640002,1.8215386,2.2350771,2.9046156,2.6945643,2.281026,4.135385,7.4929237,5.943795,3.764513,2.6026669,1.4867693,1.214359,1.2603078,4.9854364,9.744411,6.8955903,4.073026,10.095591,16.633438,18.100513,11.667693,3.826872,3.045744,2.4976413,0.65641034,1.3259488,0.7515898,0.8763078,1.0699488,1.1355898,1.3062565,2.5928206,3.121231,4.07959,5.356308,5.533539,5.182359,4.2994876,3.2065644,2.1267693,1.148718,1.6935385,1.1027694,1.2307693,1.9790771,1.3029745,2.2153847,1.4703591,1.8838975,3.4888208,3.508513,5.405539,5.976616,5.152821,4.562052,7.532308,6.8463597,7.939283,8.018052,6.6625648,5.802667,3.9876926,2.678154,2.6486156,3.9318976,5.792821,4.926359,4.535795,6.482052,9.961026,11.503591,7.827693,3.5413337,1.3226668,1.2077949,0.58092314,4.1452312,5.2644105,5.792821,6.452513,6.8332314,6.5706673,6.4065647,6.8955903,7.79159,8.057437,8.421744,9.468719,10.781539,11.9860525,12.744206,12.058257,11.280411,10.981745,10.962052,10.272821,9.908514,9.829744,10.197334,10.7848215,10.985026,11.34277,11.428103,11.254155,11.319796,12.599796,13.039591,13.410462,12.668719,10.824206,8.946873,8.3593855,7.972103,7.7325134,7.3485136,6.2720003,5.5762057,5.280821,5.1298466,5.0510774,5.142975,4.4012313,4.164923,3.570872,3.2196925,5.142975,6.2129235,6.987488,7.824411,8.556309,8.484103,7.315693,7.4732313,7.5487185,7.0892315,6.629744,6.2194877,6.058667,6.3573337,6.738052,6.242462,5.901129,6.4295387,6.449231,5.927385,6.196513,5.4153852,5.2053337,4.9526157,4.578462,4.5423594,4.4373336,4.0336413,3.9745643,4.1550775,3.7185643,3.3542566,2.937436,2.6518977,2.6453335,3.0424619,4.135385,4.781949,4.9821544,5.0510774,5.609026,4.778667,5.293949,6.301539,6.8365135,5.8190775,6.36718,8.43159,9.271795,7.88677,5.0149746,4.1025643,4.010667,5.225026,6.8266673,6.4590774,7.4010262,9.980719,8.78277,4.7950773,5.402257,8.598975,7.2960005,8.241231,11.877745,12.337232,10.174359,11.273847,16.295385,21.700924,19.748104,9.872411,6.2851286,6.3343596,7.017026,4.972308,4.8836927,7.6077952,7.5454364,4.706462,4.71959,4.6900516,3.95159,3.2065644,2.9669745,3.5478978,3.8728209,4.972308,6.3606157,7.0826674,5.7468724,4.092718,3.8038976,4.0467696,4.4964104,5.32677,5.723898,6.5280004,7.509334,8.129642,7.5487185,7.1647186,6.816821,6.432821,6.422975,7.6701546,6.8660517,6.5378466,6.5805135,6.6428723,6.1341543,5.225026,5.0543594,5.5138464,6.0980515,5.917539,5.169231,5.1954875,5.2512827,4.8049235,3.501949,2.8356924,2.9965131,3.4921029,3.9122055,3.9187696,4.1025643,4.161641,3.948308,3.7316926,4.2240005,4.6605134,4.598154,4.276513,4.07959,4.519385,5.3366156,5.4580517,5.297231,4.9329233,4.1025643,4.378257,4.2994876,3.8498464,3.2886157,3.1638978,2.8849232,3.0030773,2.9440002,2.7798977,3.2000003,3.4888208,2.9768207,2.553436,2.3827693,1.9003079,2.4648206,2.858667,2.8717952,2.550154,2.172718,1.5064616,1.0601027,0.8467693,0.74830776,0.54482055,1.1782565,1.3357949,1.1126155,0.79097444,0.8467693,0.94523084,1.4933335,1.8707694,1.8642052,1.6640002,2.802872,2.8553848,2.3433847,1.7887181,1.6968206,1.6640002,2.048,2.1924105,1.8182565,1.0338463,1.4145643,1.2242053,1.2504616,1.6705642,2.048,2.162872,2.5895386,2.8849232,3.114667,3.8596926,3.7907696,3.383795,3.242667,3.446154,3.5610259,4.1682053,4.8344617,5.142975,5.113436,5.179077,5.5630774,6.183385,6.2555904,6.1078978,7.174565,6.941539,7.13518,7.3485136,7.256616,6.619898,6.7249236,6.8332314,7.2927184,8.165744,9.232411,7.3747697,7.145026,7.5520005,7.9163084,7.8506675,8.612103,9.051898,9.088,8.976411,9.314463,9.357129,9.442462,9.163487,8.457847,7.634052,7.3091288,7.8769236,8.835282,9.6754875,9.872411,9.947898,9.898667,9.974154,10.06277,9.682052,9.235693,9.317744,9.074872,8.503796,8.461129,8.818872,8.749949,8.992821,9.5146675,9.494975,9.225847,9.452309,10.266257,11.434668,12.416001,12.120616,13.128206,14.916924,15.980309,13.830565,12.347078,11.848206,11.293539,10.8537445,11.913847,10.843898,10.65354,10.676514,10.5780525,10.328616,11.178667,11.867898,12.051693,11.88759,12.045129,12.626052,12.235488,11.329642,10.70277,11.467488,10.637129,10.390975,10.886565,11.54954,11.076924,10.338462,10.292514,10.256411,10.144821,10.482873,11.759591,11.753027,11.18195,10.656821,10.709334,11.85477,12.081232,11.500309,10.381129,9.153642,9.120821,9.344001,9.691898,9.964309,9.892103,10.679795,11.421539,12.009027,12.488206,13.072412,1.024,1.4867693,1.6672822,1.8018463,2.0086155,2.28759,2.3368206,1.9298463,1.5130258,1.4736412,2.1202054,2.681436,3.7284105,4.161641,3.7874875,3.31159,4.164923,4.854154,5.0510774,5.1232824,6.1505647,6.550975,6.2030773,5.618872,5.0215387,4.348718,5.2020516,6.121026,6.5739493,6.363898,5.6320004,5.093744,5.353026,5.7632823,6.235898,7.24677,7.259898,7.197539,6.997334,6.747898,6.698667,5.172513,5.651693,6.672411,7.453539,7.90318,8.149334,7.716103,6.8004107,5.7731285,5.1889234,5.5893335,5.737026,6.4590774,7.6209235,8.132924,8.119796,8.136206,7.9786673,7.8834877,8.530052,8.615385,8.982975,9.288206,9.40636,9.429334,8.917334,8.871386,9.140513,9.465437,9.4916935,8.979693,9.38995,9.6295395,9.42277,9.337437,8.874667,8.228104,7.830975,7.755488,7.706257,8.083693,8.674462,9.540924,10.400822,10.620719,10.328616,10.57477,11.277129,11.930258,11.611898,11.782565,12.071385,12.396309,12.438975,11.657847,11.913847,12.189539,12.120616,11.723488,11.369026,12.015591,11.680821,10.9686165,10.322052,10.039796,9.6984625,9.888822,10.203898,10.354873,10.148104,9.938052,9.531077,9.219283,9.193027,9.521232,9.777231,9.301334,8.946873,9.025641,9.3078985,9.173334,9.084719,9.084719,9.252103,9.705027,9.472001,9.028924,9.645949,11.273847,12.544001,13.860104,14.319591,15.29436,16.718771,17.060104,17.033848,16.699078,16.38072,16.324924,16.679386,17.056822,17.83795,17.96595,17.58195,18.021746,17.897026,17.335796,16.659693,16.213335,16.374155,15.225437,13.948719,13.075693,13.318565,15.563488,14.683899,13.338258,11.802258,10.44677,9.750975,10.420513,12.980514,14.815181,15.16636,15.107284,14.946463,14.9628725,15.432206,16.01313,15.730873,15.940925,16.15754,16.968206,18.136618,18.599386,17.818258,16.20349,14.880821,14.283488,14.158771,13.170873,12.813129,12.668719,12.691693,13.22995,14.04718,15.067899,15.097437,14.368821,14.5263605,16.12472,17.430975,18.005335,17.913437,17.729643,19.305027,21.80595,25.6919,27.730053,20.978874,15.671796,13.840411,13.11836,12.009027,9.872411,10.299078,9.885539,8.786052,7.4108725,6.409847,6.5903597,6.892308,6.7216415,6.380308,7.066257,6.550975,6.9349747,7.8834877,8.874667,9.216001,7.6668725,7.1220517,7.325539,8.119796,9.475283,9.084719,8.198565,7.2894363,6.49518,5.61559,5.943795,5.5893335,5.031385,4.699898,4.9427695,5.35959,6.1046157,6.3245134,6.11118,6.5017443,7.072821,7.702975,8.300308,8.523488,7.765334,6.4590774,4.9526157,4.1911798,4.1550775,3.876103,3.7185643,3.4034874,3.1967182,2.92759,1.9987694,2.2678976,2.15959,1.910154,1.7985642,2.1530259,2.5042052,2.162872,2.1530259,3.7809234,8.651488,9.6754875,6.921847,4.5587697,3.5380516,1.5721027,1.1815386,0.892718,0.7384616,0.92553854,1.8149745,6.6002054,11.195078,12.288001,8.772923,1.7558975,2.487795,4.4110775,3.4691284,0.8369231,2.8980515,1.3489232,0.8795898,0.9944616,1.4408206,2.1956925,3.5511796,4.0467696,4.0041027,4.3618464,6.669129,5.7042055,4.2174363,2.989949,2.1234872,1.0371283,0.84348726,1.1060513,1.5425643,1.7165129,1.024,1.8149745,1.2537436,1.723077,3.754667,6.012718,7.4404106,5.681231,4.027077,4.322462,6.957949,6.6034875,5.07077,4.3060517,4.6900516,5.0215387,11.782565,6.0291286,2.6190772,4.8640003,4.5456414,5.8420515,4.8836927,5.113436,7.4765134,10.407386,8.818872,4.6145644,2.2383592,2.0578463,0.33476925,2.484513,4.7524104,6.294975,7.0531287,7.7357955,7.017026,7.328821,7.716103,7.716103,7.384616,8.093539,8.900924,10.000411,11.23118,12.084514,11.339488,11.457642,11.565949,11.027693,9.429334,9.025641,8.651488,8.805744,9.275078,9.140513,9.908514,10.331899,10.8307705,11.85477,13.869949,14.112822,13.459693,11.897437,10.023385,9.032206,8.677744,8.408616,7.9983597,7.394462,6.698667,5.464616,4.9920006,4.706462,4.348718,3.9811285,4.2863593,4.5390773,4.0434875,3.31159,4.0434875,5.2512827,6.9087186,7.9228725,7.9950776,7.6307697,7.5454364,7.256616,6.9152827,6.554257,6.1046157,6.3967185,6.442667,6.521436,6.436103,5.5072823,5.5696416,6.052103,6.117744,5.730462,5.6451287,5.024821,4.713026,4.322462,3.9056413,3.9680004,4.1878977,4.066462,3.8006158,3.5216413,3.3280003,3.2656412,2.9472823,2.930872,3.1638978,3.006359,3.8367183,4.3716927,4.640821,4.778667,5.034667,4.3027697,4.8344617,5.7009234,6.1505647,5.5991797,5.989744,7.1581545,8.192,8.162462,6.1505647,5.7468724,3.9712822,5.1232824,8.218257,6.9743595,3.764513,4.2141542,6.088206,6.9776416,4.3027697,10.138257,9.472001,12.658873,20.040207,21.956924,19.295181,10.236719,7.2205133,11.434668,12.803283,14.168616,11.398565,9.419488,9.097847,7.2172313,5.8978467,8.352821,7.8145647,4.269949,4.4406157,5.110154,4.84759,3.69559,2.4385643,2.609231,3.242667,4.007385,5.540103,6.9677954,5.904411,3.9384618,3.5478978,4.3552823,5.435077,5.32677,5.7042055,6.4656415,6.997334,6.961231,6.301539,6.2523084,6.4689236,6.377026,6.1308722,6.6067696,6.2030773,5.720616,5.737026,6.121026,6.012718,5.5236926,5.5007186,6.1078978,6.8463597,6.5772314,4.7458467,4.644103,5.0609236,4.969026,3.5413337,3.1376412,3.245949,3.748103,4.309334,4.394667,4.345436,3.9220517,3.69559,3.9417439,4.637539,4.919795,4.7524104,4.788513,5.0084105,4.716308,5.533539,5.865026,5.622154,5.041231,4.699898,4.273231,3.945026,3.7185643,3.6890259,4.0434875,3.7251284,3.3641028,2.9801028,2.674872,2.6387694,2.5173335,2.3401027,2.3466668,2.5107694,2.546872,2.8291285,2.4320002,1.8281027,1.4900514,1.8937438,1.4408206,1.1815386,1.0043077,0.8598975,0.761436,1.2012309,1.3128207,1.270154,1.1749744,1.0535386,1.211077,1.8543591,2.300718,2.3958976,2.5173335,2.5042052,2.0644104,1.8051283,1.8051283,1.5885129,2.0512822,2.422154,2.3138463,1.7558975,1.204513,1.7427694,1.4736412,1.1618463,1.2307693,1.7558975,2.3269746,2.3335385,2.3466668,2.7241027,3.6168208,3.5544617,3.1015387,2.8816411,3.0490258,3.2820516,3.9778464,4.4077954,4.6145644,4.5817437,4.2272825,3.9942567,4.6966157,5.504,6.088206,6.636308,6.1013336,6.3245134,7.02359,7.5585647,6.9120007,6.948103,6.8660517,6.8660517,7.1187696,7.765334,7.962257,7.2336416,7.000616,7.496206,7.752206,7.9950776,7.6996927,7.637334,8.155898,9.156924,8.789334,9.291488,9.347282,8.425026,6.7905645,6.889026,7.581539,8.562873,9.580308,10.420513,9.580308,8.946873,9.478565,10.525539,9.842873,9.609847,9.202872,8.667898,8.169026,8.011488,8.914052,9.55077,9.846154,9.517949,8.103385,7.785026,8.228104,9.242257,10.6469755,12.2847185,12.173129,12.786873,14.427898,15.478155,12.389745,11.559385,12.176412,12.383181,12.097642,13.000206,12.242052,11.477334,10.548513,9.793642,10.026668,10.939077,11.946668,12.619488,12.888617,13.046155,12.727796,11.503591,9.984001,9.258667,10.896411,10.834052,10.633847,10.794667,11.175385,11.017847,10.59118,10.70277,10.617436,10.226872,10.056206,11.802258,12.337232,12.081232,11.503591,11.122872,11.867898,11.943385,11.237744,10.240001,10.056206,9.993847,9.787078,9.69518,9.7673855,9.842873,11.001437,11.457642,11.723488,12.196103,13.121642,0.9353847,1.204513,1.467077,1.9003079,2.3729234,2.4484105,2.6912823,2.5796926,2.0775387,1.6869745,2.4516926,3.1015387,3.4658465,4.076308,4.4307694,3.0194874,5.221744,5.7042055,5.4153852,5.080616,5.1987696,5.464616,5.668103,5.3005133,4.568616,4.384821,5.034667,6.1013336,6.196513,5.504,5.7764106,6.0028725,5.5958977,5.549949,6.2063594,7.259898,7.4863596,7.466667,7.4699492,7.351795,6.5411286,5.3070774,5.435077,5.730462,5.9930263,7.000616,8.320001,7.955693,7.026872,6.1440005,5.431795,5.687795,5.865026,6.9021544,8.4512825,8.864821,7.8769236,7.515898,7.3780518,7.4043083,7.893334,7.8047185,8.188719,8.963283,9.852718,10.394258,10.026668,9.29477,8.694155,8.533334,8.930462,8.612103,8.326565,8.086975,7.8539495,7.5454364,7.430565,7.3714876,7.13518,6.9743595,7.6209235,8.4283085,9.196308,9.567181,9.494975,9.265231,9.724719,10.423796,11.1983595,11.798975,11.881026,12.393026,12.937847,13.11836,12.754052,11.864616,11.828514,11.687386,11.457642,11.296822,11.490462,11.414975,10.975181,10.289231,9.642668,9.478565,9.6754875,9.924924,10.003693,9.803488,9.340718,9.252103,8.89436,8.530052,8.3364105,8.421744,8.297027,8.195283,8.2904625,8.644924,9.199591,8.986258,8.94359,8.956718,8.874667,8.4972315,8.585847,7.8802056,7.5946674,8.192,9.393231,11.073642,12.675283,13.90277,14.7331295,15.435489,16.065641,16.311796,16.262566,16.210052,16.640001,15.983591,15.540514,16.31836,17.877335,18.326975,20.069746,19.10154,17.368616,15.904821,14.834873,14.25395,13.640206,13.558155,13.883078,13.794462,14.145642,13.840411,12.793437,11.277129,9.895386,10.089026,12.09436,13.971693,14.621539,13.787898,13.269335,14.585437,15.497848,15.163078,14.119386,14.680616,15.474873,16.534975,17.578669,18.01518,16.73518,15.507693,14.723283,14.214565,13.282462,12.6063595,12.22236,11.897437,11.716924,12.117334,12.018872,12.550565,14.007796,15.734155,16.137848,16.964924,17.457232,17.956104,18.674873,19.682463,19.784206,19.928617,21.586054,24.064001,24.520206,19.15077,15.058052,12.691693,11.72677,11.044104,11.579078,11.365745,10.102155,8.36595,7.6307697,6.9054365,6.9054365,6.7872825,6.5345645,6.954667,6.892308,6.928411,7.5421543,8.516924,8.937026,7.532308,7.4863596,7.955693,8.500513,9.07159,8.87795,8.057437,7.3025646,6.675693,5.5893335,5.910975,5.654975,5.077334,4.634257,4.955898,5.7042055,6.619898,6.9645133,6.8693337,7.318975,7.0432825,7.3714876,8.03118,8.369231,7.3386674,6.432821,4.8738465,4.138667,4.1517954,3.2656412,3.6529233,3.2131286,2.5698464,2.176,2.3040001,2.0742567,1.5195899,1.2373334,1.6902566,3.2262566,2.231795,2.0086155,2.176,3.4231799,7.50277,6.957949,4.9821544,3.1015387,1.9954873,1.4736412,1.2898463,0.8369231,0.6170257,4.2272825,18.379488,6.810257,5.0477953,8.15918,9.714872,1.8149745,1.4441026,1.7066668,2.1103592,2.231795,1.7263591,1.8970258,1.7394873,1.6968206,2.0053334,2.674872,3.1113849,5.287385,6.2588725,5.9634876,7.2172313,5.421949,3.3345644,2.3762052,2.4057438,1.719795,1.2635899,1.0929232,1.204513,1.6902566,2.7306669,1.3357949,1.1815386,3.383795,6.12759,4.6572313,5.5007186,5.080616,4.5423594,4.630975,5.723898,6.5050263,4.886975,2.8225644,1.5589745,1.6147693,2.7241027,2.7864618,3.1048207,3.764513,3.6332312,5.910975,6.416411,6.0192823,5.835488,7.2205133,7.1187696,5.32677,4.6572313,4.391385,0.2855385,1.3620514,4.240411,6.2129235,6.7544622,7.515898,7.450257,7.24677,7.197539,7.325539,7.397744,7.6077952,8.329846,9.596719,11.080206,12.071385,11.730052,11.579078,11.395283,10.952206,10.026668,9.330873,8.612103,8.247795,8.201847,8.027898,8.418462,9.291488,10.138257,11.122872,13.088821,12.76718,12.097642,11.057232,10.098872,10.154668,9.449026,8.710565,7.906462,7.174565,6.820103,6.232616,5.5236926,5.0149746,4.8836927,5.1922054,3.7087183,3.5577438,3.623385,3.6332312,4.141949,4.6769233,5.5269747,6.419693,6.928411,6.49518,5.8223596,5.5007186,5.412103,5.543385,5.979898,6.363898,6.803693,6.8594875,6.426257,5.7534366,5.228308,5.3202057,5.5269747,5.5630774,5.3891287,4.630975,4.086154,3.8334363,3.8695388,4.125539,4.0533338,3.9844105,3.751385,3.4231799,3.3280003,3.245949,2.8882053,2.930872,3.3509746,3.3969233,3.7382567,4.161641,4.857436,5.5302567,5.3760004,4.4800005,4.397949,4.388103,4.276513,4.4406157,5.7698464,6.262154,7.145026,8.241231,8.004924,7.6307697,5.658257,4.916513,5.756718,6.045539,6.5083084,5.8912826,5.8157954,5.910975,3.8038976,6.747898,6.7938466,12.0549755,19.810463,16.512001,18.274464,9.360411,7.312411,13.308719,12.156719,17.447386,16.538258,14.250668,12.097642,8.254359,4.397949,8.618668,11.034257,8.149334,2.8521028,4.3060517,4.1058464,3.2918978,2.4320002,1.6443079,2.5632823,3.2131286,3.6036925,3.6004105,2.937436,3.5314875,5.362872,5.940513,5.1987696,5.5072823,6.0619493,6.0783596,6.242462,6.554257,6.314667,4.525949,5.3037953,6.088206,6.0980515,6.3507695,6.485334,6.0160003,5.408821,5.041231,5.2053337,4.7360005,4.604718,4.788513,5.0149746,4.7458467,3.9187696,3.9089234,4.086154,4.023795,3.501949,3.511795,3.4888208,4.096,5.146257,5.602462,5.113436,4.397949,3.892513,3.9351797,4.7491283,4.532513,4.634257,4.709744,4.7458467,5.0674877,5.0674877,4.841026,4.8705645,5.159385,5.2381544,4.906667,4.3552823,4.1682053,4.378257,4.457026,4.647385,4.3552823,3.5971284,2.6715899,2.1267693,1.847795,1.7001027,1.8313848,2.1431797,2.2678976,2.5107694,2.2777438,1.8937438,1.7099489,2.1234872,1.2537436,1.0338463,1.014154,0.93866676,0.761436,1.086359,1.2406155,1.2931283,1.2800001,1.1881026,1.5425643,1.8149745,2.1891284,2.6322052,2.9210258,3.0949745,2.5206156,2.231795,2.2153847,1.4408206,1.7296412,2.5829747,2.9243078,2.3630772,1.2176411,1.394872,1.7755898,2.2055387,2.422154,2.0611284,2.097231,2.409026,2.6978464,2.989949,3.6168208,3.515077,3.314872,3.1343591,3.0687182,3.18359,3.8498464,4.2568207,4.522667,4.571898,4.128821,3.5249233,4.568616,5.612308,6.2030773,7.066257,6.5772314,6.232616,6.432821,7.0367184,7.3747697,7.5388722,7.686565,7.529026,7.0367184,6.422975,6.7938466,6.7774363,6.7117953,6.5247183,5.737026,6.636308,7.177847,7.64718,8.280616,9.252103,8.4972315,8.375795,8.434873,8.260923,7.4863596,7.3386674,7.650462,8.274052,9.048616,9.77395,9.636104,9.478565,9.586872,9.731283,9.18318,9.147078,9.235693,8.786052,7.837539,7.131898,8.651488,9.419488,9.209436,8.27077,7.3321033,7.9524107,8.812308,9.645949,10.564924,12.064821,12.921437,12.42913,12.137027,12.163283,11.195078,11.369026,12.156719,12.704822,12.790154,12.806565,11.608616,10.712616,9.964309,9.567181,10.06277,10.732308,11.628308,12.278154,12.62277,12.996924,12.905026,11.657847,10.541949,9.856001,8.89436,9.350565,9.7214365,10.397539,11.355898,12.163283,12.07795,11.933539,11.30995,10.522257,10.604308,12.07795,13.279181,13.466257,12.566976,11.172104,11.096616,11.16554,10.8767185,10.315488,10.14154,9.688616,9.580308,9.636104,9.6754875,9.524513,10.128411,10.758565,11.323078,11.881026,12.635899,1.0075898,1.276718,1.4769232,1.7657437,2.1464617,2.4516926,2.281026,2.3893335,2.1858463,1.9593848,2.861949,4.2601027,4.2830772,4.056616,3.7842054,2.7536411,4.962462,5.730462,5.622154,5.2709746,5.3792825,5.349744,5.4974365,5.139693,4.338872,3.9187696,4.699898,5.832206,6.2916927,6.0750775,6.196513,6.5903597,5.76,5.32677,5.874872,6.951385,7.282872,7.0367184,6.8955903,6.9382567,6.6461544,5.8223596,5.5565133,5.3136415,5.225026,6.0783596,7.2992826,7.3682055,6.99077,6.4065647,5.3924108,5.2315903,5.467898,6.6002054,8.264206,9.242257,9.340718,9.179898,8.973129,8.690872,8.073847,7.6635904,7.762052,8.237949,8.900924,9.4916935,9.396514,8.651488,8.41518,8.779488,8.763078,8.251078,7.7948723,7.6176414,7.6077952,7.3058467,7.3386674,7.27959,7.1089234,7.1647186,8.155898,8.786052,9.271795,9.199591,8.786052,8.897642,9.970873,10.66995,11.293539,11.930258,12.452104,13.371078,13.61395,13.722258,13.718975,13.13477,11.707078,11.37559,11.444513,11.539693,11.621744,11.109744,10.463181,9.90195,9.468719,9.019077,8.533334,8.772923,8.976411,8.861539,8.598975,8.379078,8.090257,7.762052,7.5421543,7.7357955,7.8473854,7.824411,7.9195905,8.14277,8.274052,8.113232,8.201847,8.027898,7.5946674,7.387898,7.1647186,6.875898,6.8955903,7.4174366,8.43159,10.049642,12.025436,13.443283,14.106257,14.5263605,15.445334,15.668514,15.419078,15.304206,16.311796,15.996719,14.513232,14.25395,15.126975,14.529642,19.009642,20.374975,19.183592,16.564514,14.247386,13.692719,13.37436,13.400617,13.682873,13.919181,13.83713,13.988104,13.571283,12.458668,11.178667,11.346052,12.058257,12.905026,13.279181,12.386462,11.572514,13.193847,14.54277,14.427898,13.1872835,12.905026,13.571283,14.762668,15.849027,16.02954,14.608412,13.426873,13.167591,13.46954,12.941129,12.504617,12.563693,12.544001,12.379898,12.517745,12.2387705,11.296822,12.5374365,15.271386,15.258258,16.170668,16.902565,17.723078,18.888206,20.611284,19.912207,19.183592,19.249231,20.312616,21.96349,19.24595,17.690258,15.721026,13.233232,11.621744,11.2672825,11.1294365,10.515693,9.488411,8.868103,7.653744,7.3091288,7.145026,6.8496413,6.514872,6.4557953,6.445949,6.9382567,7.6767187,7.722667,7.5487185,7.6570263,7.899898,8.320001,9.147078,8.385642,7.8080006,7.269744,6.5969234,5.586052,5.579488,5.6287184,5.356308,4.9788723,5.3070774,6.0849237,7.020308,7.5520005,7.77518,8.4283085,7.6767187,7.578257,7.857231,8.018052,7.351795,6.436103,5.293949,4.7294364,4.5095387,3.370667,3.2361028,2.8455386,2.28759,1.847795,2.0053334,1.5786668,1.2898463,1.5524104,2.1956925,2.4582565,1.8838975,1.4867693,1.4802053,2.176,3.9778464,3.8432825,3.045744,2.1924105,1.5885129,1.2471796,0.90912825,3.2623591,5.0051284,8.956718,24.06072,7.578257,3.0260515,3.6332312,4.161641,0.9156924,1.8051283,1.2865642,2.2088206,4.1452312,3.3936412,6.0652313,4.4701543,2.878359,2.9407182,3.698872,3.5774362,5.2578464,6.3179493,6.432821,7.3550773,5.5269747,3.4855387,2.2219489,1.8018463,1.3620514,1.0502565,0.86646163,1.0043077,1.3554872,1.529436,0.67938465,1.4178462,3.6791797,5.602462,3.5478978,4.955898,3.761231,4.2371287,6.5870776,6.9349747,8.064001,4.9985647,2.8356924,2.5829747,1.1651284,1.1323078,2.156308,2.7700515,2.8291285,3.511795,4.6834874,5.664821,5.8420515,5.546667,6.058667,5.549949,4.322462,4.5817437,4.969026,0.57764107,1.0601027,3.3444104,5.32677,6.2687182,6.7938466,7.138462,6.675693,6.678975,7.4207187,8.178872,7.972103,8.260923,9.245539,10.5780525,11.382154,11.959796,11.405129,10.505847,9.865847,9.895386,8.999385,8.356103,8.067283,7.962257,7.604513,7.9195905,9.127385,10.289231,11.195078,12.373334,11.864616,11.277129,10.610872,10.085744,10.154668,9.504821,9.147078,8.392206,7.450257,7.4108725,7.194257,6.5969234,5.924103,5.3366156,4.8607183,3.9942567,3.7809234,3.748103,3.7251284,3.8531284,4.2207184,4.4077954,4.699898,4.9788723,4.7458467,4.132103,4.7458467,5.5269747,5.924103,5.8945646,6.0061545,6.36718,6.380308,5.917539,5.3366156,4.7917953,4.6933336,4.7622566,4.821334,4.7950773,4.7491283,4.4274874,4.2962055,4.420923,4.4865646,4.201026,3.757949,3.3542566,3.0523078,2.7963078,2.937436,3.2295387,3.501949,3.6463592,3.6036925,3.639795,4.0336413,4.716308,5.221744,4.667077,3.8367183,3.7152824,3.7973337,3.8662567,3.9942567,4.8836927,5.865026,6.5805135,7.062975,7.7456417,8.55959,7.269744,5.4383593,4.3290257,4.890257,7.177847,5.6418467,4.818052,5.3760004,4.135385,6.8332314,6.931693,8.769642,12.002462,11.592206,10.197334,10.476309,16.79754,23.972105,17.24718,16.308514,16.393847,14.805334,11.027693,6.7282057,3.1015387,4.97559,8.182155,9.242257,5.35959,4.9132314,4.1550775,3.748103,3.6135387,2.9243078,2.2482052,2.7766156,3.1770258,2.8192823,1.7657437,3.5347695,6.042257,6.1078978,3.889231,2.8914874,4.44718,5.8125134,6.226052,5.973334,6.380308,5.3169236,4.8672824,5.3037953,6.180103,6.3310776,6.432821,5.586052,4.7983594,4.529231,4.70318,4.1156926,3.7087183,3.6004105,3.698872,3.692308,3.1048207,3.370667,3.5905645,3.5282054,3.623385,3.3509746,3.442872,3.8432825,4.4800005,5.2644105,4.7622566,4.6966157,4.4242053,4.1091285,4.7294364,5.024821,4.923077,4.785231,4.893539,5.4416413,4.5095387,4.4865646,4.598154,4.519385,4.3651285,4.900103,4.670359,4.59159,4.824616,4.7622566,4.854154,4.9362054,4.4865646,3.4756925,2.3663592,1.6672822,1.4769232,1.5655385,1.7788719,2.0512822,2.3335385,2.4057438,2.2678976,2.041436,1.9429746,1.2373334,1.148718,1.148718,1.017436,0.8467693,1.0075898,1.0929232,1.1782565,1.3128207,1.5491283,1.595077,1.5556924,1.7362052,2.156308,2.5435898,2.934154,2.4582565,2.2547693,2.3729234,1.7887181,1.8346668,4.6178465,5.7665644,4.092718,1.6049232,1.4572309,1.7755898,2.100513,2.2547693,2.3663592,1.9659488,2.097231,2.2482052,2.3729234,2.8750772,3.1376412,3.1770258,3.1081028,3.1245131,3.4888208,3.620103,3.82359,3.9778464,3.9680004,3.7021542,3.4822567,4.2338467,4.896821,5.0642056,4.955898,4.972308,5.2742567,6.11118,7.207385,7.75877,7.4240007,7.213949,7.0957956,6.8627696,6.124308,5.5663595,5.2020516,5.464616,6.0160003,5.72718,6.7971287,7.8014364,8.237949,8.283898,8.802463,8.539898,8.04759,7.8703594,7.9885135,7.8145647,8.004924,8.333129,8.41518,8.549745,9.714872,9.728001,9.783795,9.764103,9.544206,9.019077,8.78277,9.301334,9.005949,7.939283,7.762052,9.5606165,10.322052,9.691898,8.372514,8.139488,8.201847,8.838565,9.810052,10.79795,11.37559,12.3306675,12.160001,11.756309,11.516719,11.372309,11.608616,11.795693,12.143591,12.1698475,10.732308,9.449026,8.940309,8.828718,9.107693,10.154668,10.259693,10.712616,11.300103,11.953232,12.737642,13.266052,12.186257,10.925949,10.138257,9.691898,9.412924,9.6065645,10.423796,11.405129,11.480617,11.437949,11.61518,11.506873,11.349334,12.1238985,12.619488,13.15118,12.872206,11.792411,10.781539,10.57477,10.620719,10.604308,10.512411,10.6469755,10.433641,10.256411,10.180923,10.154668,9.984001,10.059488,10.601027,11.270565,11.877745,12.373334,1.1651284,1.3423591,1.6278975,1.8576412,2.0184617,2.2383592,1.9889232,2.156308,2.166154,2.2121027,3.2525132,4.6933336,4.7556925,4.2141542,3.5610259,2.989949,4.97559,5.7501545,5.658257,5.2315903,5.1856413,5.353026,5.3792825,5.0051284,4.309334,3.7185643,4.394667,5.405539,6.2851286,6.705231,6.4590774,6.560821,5.8518977,5.3694363,5.536821,6.157129,6.5936418,6.491898,6.485334,6.695385,6.7249236,6.048821,5.7698464,5.2578464,4.713026,5.156103,6.2162056,6.7085133,6.957949,6.8693337,5.910975,5.211898,5.481026,6.363898,7.515898,8.576,9.563898,9.990565,10.164514,9.849437,8.251078,7.5421543,7.2336416,7.5552826,8.267488,8.65477,8.310155,8.116513,8.484103,9.005949,8.461129,7.571693,7.181129,7.204103,7.3386674,7.062975,6.9054365,6.8562055,6.961231,7.351795,8.260923,8.700719,8.992821,8.904206,8.726975,9.284924,10.217027,10.889847,11.510155,12.173129,12.852514,13.587693,13.620514,13.692719,13.879796,13.581129,11.782565,11.61518,11.723488,11.493745,11.067078,10.620719,10.144821,9.783795,9.43918,8.772923,8.2215395,8.39877,8.402052,8.034462,7.8080006,7.77518,7.5552826,7.13518,6.7117953,6.685539,7.138462,7.427283,7.568411,7.574975,7.466667,7.6110773,7.7292314,7.3452315,6.738052,6.941539,6.948103,6.921847,6.9645133,7.2270775,7.899898,9.731283,11.900719,13.37436,13.869949,13.879796,14.690463,15.402668,15.445334,15.241847,16.219898,16.003283,14.043899,13.010053,13.124924,12.173129,16.088617,19.213129,19.410053,16.86318,14.076719,12.885334,12.603078,12.918155,13.581129,14.395078,14.211283,15.051488,15.261539,14.273643,12.612924,12.3995905,11.976206,11.730052,11.707078,11.592206,10.95877,12.258463,13.617231,13.955283,12.983796,11.779283,12.025436,13.065847,13.978257,13.604104,12.393026,11.58236,11.605334,12.209231,12.465232,11.976206,12.317539,12.616206,12.691693,13.049437,13.15118,12.173129,12.5374365,13.994668,13.610668,14.943181,16.452925,17.542566,18.297438,19.482258,18.865232,18.54031,18.09395,17.923283,19.236105,18.130053,18.809437,18.602669,16.512001,13.220103,11.300103,10.673231,10.35159,9.911796,9.501539,8.418462,7.522462,7.1909747,7.1515903,6.491898,5.940513,5.7435904,5.976616,6.452513,6.701949,7.066257,7.4404106,7.634052,7.716103,8.004924,7.4929237,7.4404106,7.250052,6.6527185,5.7009234,5.3103595,5.47118,5.5236926,5.3891287,5.5893335,6.3310776,7.145026,7.64718,7.9524107,8.661334,8.234667,7.706257,7.5388722,7.5913854,7.1187696,5.9930263,5.152821,4.637539,4.1813335,3.1967182,2.9505644,2.609231,2.1234872,1.6410258,1.4998976,1.1093334,1.3883078,2.1169233,2.5435898,1.3718976,1.4276924,1.6705642,2.7208207,3.8531284,2.986667,2.2186668,1.7788719,1.6738462,3.5478978,10.676514,2.7667694,3.6004105,6.8955903,11.286975,20.342155,7.197539,4.315898,3.8564105,2.3269746,0.5973334,2.930872,2.0151796,2.7667694,5.1954875,4.388103,7.6110773,5.9569235,4.2272825,4.201026,4.650667,4.0992823,5.2053337,5.9470773,6.114462,7.2992826,5.5663595,3.6036925,2.0775387,1.2438976,0.9288206,0.8041026,0.8566154,1.020718,1.0371283,0.41682056,0.9517949,2.6420515,4.457026,5.1659493,3.370667,4.3716927,2.5009232,3.5347695,7.3025646,7.680001,7.9261546,4.1583595,2.428718,3.2918978,1.8018463,2.3138463,2.2908719,2.0545642,2.1989746,3.6168208,4.1682053,4.4996924,4.713026,5.0510774,5.910975,4.962462,3.7710772,3.6529233,3.6758976,0.6268718,0.92225647,2.3893335,4.2338467,5.7829747,6.488616,6.931693,6.3868723,6.6002054,7.8736415,9.074872,8.425026,8.500513,9.18318,10.105436,10.656821,11.529847,10.758565,9.639385,9.002667,9.179898,8.346257,8.008205,7.8670774,7.752206,7.6176414,7.9524107,9.058462,10.269539,11.306667,12.297847,11.487181,11.286975,10.860309,10.121847,9.757539,9.557334,9.531077,9.035488,8.211693,7.965539,7.765334,7.4929237,6.954667,6.0356927,4.6966157,4.391385,4.1452312,3.95159,3.82359,3.817026,4.0041027,3.9318976,3.889231,4.020513,4.3060517,4.2436924,5.1298466,5.8781543,6.0258465,5.720616,5.8880005,6.009436,5.8847184,5.4416413,4.7392826,4.276513,4.023795,4.056616,4.269949,4.3618464,4.6572313,4.516103,4.3290257,4.197744,3.948308,3.879385,3.4100516,2.9013336,2.5829747,2.550154,2.868513,3.4231799,3.6791797,3.570872,3.5183592,3.5052311,3.9548721,4.529231,4.772103,4.092718,3.2820516,3.062154,3.2951798,3.69559,3.8071797,4.414359,5.5893335,6.196513,6.3573337,7.4141545,8.503796,7.9195905,6.4656415,4.969026,4.2601027,7.1581545,5.425231,4.2830772,5.1626673,5.7042055,6.5903597,7.1909747,7.1154876,7.381334,10.407386,6.688821,14.007796,22.744617,25.682053,17.99877,25.445745,21.658258,15.638975,11.556104,8.723693,4.4077954,3.2918978,4.7556925,6.6592827,5.3169236,5.3037953,5.097026,4.788513,4.706462,5.395693,3.501949,3.0687182,3.0851285,2.809436,1.7723079,3.751385,4.962462,4.955898,4.31918,4.6769233,5.4153852,6.3245134,6.0849237,4.890257,4.4340515,5.4153852,4.565334,4.3585644,5.293949,5.868308,6.1505647,5.3070774,4.4077954,3.9909747,4.092718,3.7251284,3.2164104,3.1081028,3.3280003,3.2032824,2.6880002,3.4034874,3.8859491,3.748103,3.6726158,3.3411283,3.3411283,3.3509746,3.570872,4.7261543,4.420923,4.7261543,4.667077,4.2338467,4.4077954,4.7458467,4.5423594,4.309334,4.4373336,5.1922054,4.096,4.3027697,4.4307694,4.06318,3.7284105,5.0904617,4.9493337,4.6112823,4.5489235,4.384821,4.240411,4.6145644,4.6244106,3.9680004,2.9210258,2.0217438,1.6607181,1.5885129,1.6311796,1.6902566,2.0873847,2.4713848,2.5632823,2.3236926,1.9626669,1.3456411,1.1716924,1.1651284,1.1716924,1.1520001,1.0535386,0.95835906,1.0469744,1.3259488,1.6311796,1.5425643,1.3489232,1.4834872,1.9265642,2.2219489,2.2777438,1.9856411,2.0742567,2.5009232,2.4484105,2.225231,5.425231,7.059693,5.549949,2.7109745,2.28759,2.5238976,2.4976413,2.162872,2.3466668,1.9232821,2.0151796,2.1202054,2.162872,2.5140514,2.8553848,2.8750772,2.8882053,3.0785644,3.4756925,3.1671798,3.1638978,3.31159,3.4297438,3.3247182,3.4100516,3.7415388,4.073026,4.20759,3.9680004,3.9975388,4.785231,6.0619493,7.2631803,7.5388722,7.138462,6.7183595,6.619898,6.688821,6.2523084,5.21518,4.420923,4.588308,5.398975,5.477744,6.3507695,7.6274877,8.165744,7.936001,8.008205,8.362667,8.093539,7.8637953,7.9228725,8.096821,8.385642,8.825437,8.809027,8.704,9.852718,10.043077,10.236719,10.167795,9.718155,8.907488,8.779488,9.324308,9.124104,8.300308,8.513641,9.780514,10.220308,9.728001,8.897642,9.035488,8.36595,8.65477,9.6754875,10.850462,11.254155,11.841642,12.301129,12.320822,12.012309,11.913847,11.680821,11.421539,11.585642,11.661129,10.157949,9.163487,8.726975,8.809027,9.271795,9.878975,9.291488,9.636104,10.453334,11.457642,12.553847,13.115078,12.219078,10.998155,10.266257,10.522257,10.233437,10.164514,10.729027,11.572514,11.559385,11.575796,11.634872,11.618463,11.844924,13.069129,12.800001,12.616206,11.926975,10.857026,10.233437,10.102155,10.253129,10.443488,10.59118,10.781539,10.807796,10.735591,10.610872,10.456616,10.266257,10.184206,10.555078,11.247591,11.956513,12.173129,1.3554872,1.394872,1.8806155,2.172718,2.100513,1.972513,2.041436,2.1530259,2.176,2.3794873,3.4100516,4.2962055,4.7917953,4.650667,4.073026,3.6857438,5.3924108,5.865026,5.5958977,5.024821,4.535795,5.2414365,5.297231,5.0510774,4.70318,4.2994876,4.5062566,5.139693,6.038975,6.7150774,6.3474874,6.0717955,5.8486156,5.661539,5.5007186,5.362872,5.8420515,6.0783596,6.304821,6.488616,6.3474874,5.858462,6.0160003,5.681231,4.900103,4.9296412,5.8157954,6.311385,6.7150774,6.957949,6.6002054,5.901129,5.976616,6.2884107,6.619898,7.062975,8.01477,8.992821,9.728001,9.682052,8.04759,7.5487185,6.8397956,7.0892315,8.077128,8.182155,7.450257,7.962257,8.5661545,8.576,7.755488,6.7216415,6.5444107,6.695385,6.75118,6.3934364,5.973334,6.048821,6.4590774,7.062975,7.752206,8.267488,8.65477,8.950154,9.3078985,9.980719,10.381129,11.044104,11.680821,12.199386,12.698257,13.036308,13.282462,13.361232,13.266052,13.069129,12.1238985,12.212514,11.926975,10.962052,10.105436,9.924924,9.842873,9.659078,9.235693,8.500513,8.530052,8.621949,8.2215395,7.466667,7.197539,7.4929237,7.3025646,6.8332314,6.2588725,5.7074876,6.186667,6.8594875,7.145026,7.020308,7.0367184,7.5388722,7.6176414,7.197539,6.698667,7.066257,7.716103,7.584821,7.200821,7.0334363,7.499488,9.321027,11.58236,13.249642,13.906053,13.7386675,14.201437,15.602873,16.390566,16.38072,16.771284,15.940925,14.076719,13.078976,13.098668,12.530872,13.384206,16.28554,17.529438,16.144411,13.906053,12.07795,11.67754,12.383181,13.61395,14.50995,15.07118,16.613745,17.174976,16.059078,13.840411,12.71795,11.651283,10.889847,10.738873,11.562668,11.277129,11.848206,12.793437,13.453129,12.996924,11.503591,11.575796,12.3306675,12.78359,11.848206,10.817642,10.706052,10.870154,11.168821,11.956513,11.628308,11.851488,12.058257,12.248616,12.977232,13.768207,14.086565,13.794462,13.115078,12.629334,14.296617,16.15754,17.132309,17.174976,17.257027,17.214361,17.910154,17.903591,17.56882,19.088411,17.562258,18.034874,19.081848,18.865232,15.126975,12.120616,10.755282,10.213744,9.90195,9.478565,9.035488,7.6603084,7.0104623,7.24677,7.0400004,5.9503593,5.4383593,5.277539,5.504,6.409847,6.564103,7.1483083,7.387898,7.0137444,6.2555904,6.6592827,7.056411,7.194257,6.921847,6.183385,5.481026,5.402257,5.5663595,5.723898,5.7534366,6.3540516,7.0432825,7.3649235,7.50277,8.27077,8.5891285,7.7390776,7.181129,7.1187696,6.47877,5.1200004,4.2502565,3.6693337,3.2131286,2.733949,2.8422565,2.3958976,1.8051283,1.3226668,1.0371283,0.9517949,1.5327181,2.3401027,2.5271797,0.86317956,1.3522053,2.7831798,5.1889234,6.882462,4.4406157,2.1202054,1.2964103,1.4276924,5.7534366,21.31036,5.100308,1.5885129,4.6539493,9.314463,11.71036,5.2578464,6.180103,7.1220517,5.146257,1.7460514,3.6069746,2.806154,3.7382567,5.904411,3.9384618,5.7009234,5.536821,5.2447186,5.3103595,4.8738465,4.391385,5.3136415,5.677949,5.5696416,7.145026,5.297231,3.2886157,1.8248206,1.0994873,0.8041026,0.8336411,1.079795,1.1290257,0.8402052,0.3446154,1.7723079,4.1091285,5.58277,5.3891287,3.6758976,3.1409233,2.0086155,3.373949,6.669129,7.6734366,5.868308,2.5173335,1.276718,2.281026,2.156308,3.2951798,2.353231,1.5195899,1.8642052,3.3214362,4.6211286,3.8432825,3.1967182,3.7809234,5.5893335,4.716308,3.9745643,2.9538465,1.654154,0.48246157,0.7515898,1.6771283,3.2754874,5.172513,6.5772314,6.685539,6.3179493,6.918565,8.536616,9.852718,8.615385,8.661334,9.206155,9.741129,10.043077,10.459898,10.013539,9.429334,8.92718,8.241231,7.785026,7.8539495,7.785026,7.5618467,7.8080006,8.303591,8.950154,9.8363085,11.0375395,12.596514,11.605334,11.82195,11.405129,10.148104,9.508103,9.810052,9.819899,9.645949,9.248821,8.448001,7.896616,7.9852314,7.830975,6.9743595,5.3924108,4.824616,4.414359,4.1813335,4.128821,4.2207184,4.1091285,4.073026,4.1189747,4.388103,5.139693,5.5991797,5.8880005,5.85518,5.6320004,5.6320004,5.9995904,5.8125134,5.5072823,5.113436,4.2469745,3.817026,3.43959,3.5544617,4.0467696,4.2338467,4.2929235,4.1156926,3.764513,3.3247182,2.8882053,3.1737437,2.9702566,2.5009232,2.2186668,2.7634873,2.9702566,3.2361028,3.2623591,3.1245131,3.249231,3.314872,3.82359,4.33559,4.493129,4.020513,3.2886157,2.7995899,2.858667,3.3312824,3.6627696,4.601436,5.467898,6.0947695,6.6494365,7.64718,7.88677,7.686565,7.515898,6.8955903,4.4012313,7.0137444,6.3343596,5.3891287,5.7534366,7.571693,5.504,6.7117953,7.6964107,8.375795,12.087796,9.298052,16.170668,19.462566,16.344616,14.41477,39.565132,29.659899,16.876308,13.817437,13.505642,6.6527185,4.1091285,3.18359,2.550154,2.2350771,4.6112823,6.2030773,6.308103,6.3442054,9.869129,8.12636,4.7917953,2.861949,2.7241027,2.172718,3.446154,2.7766156,4.0369234,7.6143594,10.381129,8.293744,7.6931286,6.9743595,5.353026,2.878359,4.2994876,3.9975388,3.498667,3.7349746,5.0477953,5.799385,5.2578464,4.2207184,3.3936412,3.4002054,3.6594875,3.3312824,3.4297438,3.8662567,3.4592824,2.937436,3.8301542,4.453744,4.2305646,3.692308,3.629949,3.3280003,2.9735386,3.0424619,4.315898,4.2863593,4.522667,4.4996924,4.1452312,3.8498464,3.4494362,3.4592824,3.501949,3.6857438,4.6112823,3.948308,4.089436,4.2469745,4.0992823,3.8038976,5.3037953,5.037949,4.240411,3.626667,3.3936412,3.131077,3.6562054,4.066462,3.945026,3.3903592,2.6945643,2.0676925,1.8116925,1.8018463,1.4834872,1.9856411,2.4484105,2.5337439,2.294154,2.1431797,1.4736412,1.0732309,1.0469744,1.2800001,1.4244103,1.1520001,0.8960001,0.9911796,1.3357949,1.3915899,1.4539489,1.3357949,1.591795,2.103795,2.0873847,1.5458462,1.4211283,1.7887181,2.4385643,2.861949,2.5435898,4.31918,5.7107697,5.504,3.7218463,3.4034874,3.8006158,3.508513,2.484513,2.0611284,1.8806155,2.103795,2.3466668,2.4976413,2.7208207,2.7602053,2.6551797,2.6945643,2.8980515,3.0227695,2.6617439,2.5796926,2.8258464,3.170462,3.1081028,3.2032824,3.3509746,3.639795,4.082872,4.6244106,4.4274874,5.182359,6.232616,6.957949,6.774154,6.820103,6.5936418,6.49518,6.498462,6.166975,5.5729237,4.8607183,4.5587697,4.630975,4.466872,5.0051284,6.1997952,7.1056414,7.4010262,7.3780518,8.086975,8.362667,8.28718,8.152616,8.461129,8.52677,8.920616,9.120821,9.219283,9.90195,10.410667,10.765129,10.725744,10.138257,8.940309,9.18318,9.242257,8.835282,8.264206,8.425026,8.838565,8.825437,8.769642,8.907488,9.330873,8.484103,8.536616,9.373539,10.660104,11.808822,11.723488,12.4685135,12.757335,12.356924,12.114052,11.707078,11.605334,11.766154,11.946668,11.67754,10.807796,10.023385,9.7214365,9.67877,9.061745,8.155898,8.87795,10.157949,11.414975,12.576821,12.599796,11.759591,10.886565,10.394258,10.272821,11.224616,11.237744,11.303386,11.828514,12.63918,12.842668,12.3766165,11.848206,11.85477,12.980514,12.534155,12.09436,11.372309,10.433641,9.731283,9.567181,9.895386,10.266257,10.44677,10.381129,10.456616,10.686359,10.765129,10.57477,10.180923,10.217027,10.459898,11.073642,11.776001,11.835078,1.5261539,1.782154,2.2022567,2.2383592,1.9593848,2.044718,2.0086155,2.0906668,2.1956925,2.409026,3.006359,4.312616,5.6451287,5.4875903,4.2469745,4.273231,4.893539,5.4613338,5.586052,5.2414365,4.7917953,5.402257,5.5269747,5.7107697,5.9963083,5.933949,5.5926156,5.5630774,5.83877,6.12759,5.858462,5.7501545,5.684513,5.874872,6.0947695,5.691077,5.9470773,5.7107697,5.2447186,4.8705645,4.9427695,5.674667,6.4557953,6.99077,7.1122055,6.7610264,6.4656415,6.11118,5.586052,5.2348723,5.8453336,6.8332314,6.173539,5.7403083,5.9503593,5.7665644,6.5739493,7.433847,7.8112826,7.680001,7.522462,8.546462,7.522462,6.747898,6.8397956,6.7282057,6.889026,7.568411,7.837539,7.4010262,6.6067696,6.3277955,6.62318,6.810257,6.5903597,6.0258465,5.930667,5.858462,5.927385,6.3245134,7.325539,8.155898,8.763078,9.416205,10.066052,10.345026,11.126155,11.467488,11.536411,11.526565,11.674257,12.832822,13.745232,13.88636,13.420309,13.213539,12.63918,12.442257,11.703795,10.518975,9.993847,9.4457445,9.189744,8.999385,8.585847,7.584821,7.1089234,7.1154876,7.062975,6.951385,7.3550773,7.1844106,6.948103,6.997334,7.0990777,6.439385,6.304821,6.619898,6.741334,6.5739493,6.560821,6.9645133,7.174565,7.1122055,6.9349747,7.020308,7.276308,7.0925136,7.00718,7.3747697,8.375795,8.267488,10.089026,12.763899,14.946463,15.044924,15.251694,15.809642,16.761436,17.798565,18.248207,16.784412,15.192616,14.208001,13.689437,12.603078,13.702565,14.8939495,15.16636,14.418053,13.443283,12.406155,11.844924,12.032001,12.973949,14.388514,15.573335,16.554668,16.800821,16.20677,15.120412,13.033027,11.579078,11.139283,11.513436,11.9171295,11.122872,10.660104,11.155693,12.156719,12.130463,11.300103,12.117334,12.911591,12.859077,11.992617,10.417232,10.637129,11.237744,11.67754,12.297847,13.590976,13.420309,12.750771,12.232206,12.20595,13.673027,13.98154,14.037334,14.03077,13.459693,15.058052,15.428925,15.724309,16.331488,16.89272,16.915693,18.149744,18.852104,19.160616,21.103592,18.894772,17.552412,16.246155,14.920206,14.296617,12.685129,11.385437,10.965334,10.84718,9.3078985,9.577026,8.52677,7.3550773,6.918565,7.7357955,6.9677954,6.5378466,6.1768208,6.055385,6.774154,7.653744,7.5979495,7.13518,6.7314878,6.806975,6.9152827,6.889026,6.948103,7.1581545,7.4141545,6.488616,5.907693,5.8289237,6.0685134,6.117744,6.1440005,6.9809237,7.3714876,7.4896417,8.940309,9.222565,8.257642,7.2336416,6.5411286,5.7829747,4.31918,3.2656412,2.7602053,2.733949,2.930872,2.4910772,1.657436,1.0043077,0.7450257,0.7318975,1.3292309,1.2340513,1.7690258,2.5009232,1.204513,2.6715899,4.197744,4.8082056,4.2929235,3.2196925,1.719795,1.1946667,1.3850257,2.7437952,6.4557953,1.6705642,1.2340513,2.0217438,3.0785644,5.6320004,2.665026,3.9548721,4.8771286,4.2962055,4.578462,2.0644104,2.6256413,6.0061545,8.713847,4.013949,4.916513,4.9952826,5.2578464,5.3727183,3.6758976,4.7261543,4.6867695,4.7917953,5.5696416,6.8496413,4.70318,2.8389745,1.6672822,1.148718,0.79425645,1.1355898,1.1651284,0.9944616,0.67282057,0.19692309,1.2832822,3.6529233,4.9460516,4.4077954,2.868513,1.463795,2.9078977,5.21518,7.3583593,9.26195,4.818052,1.6311796,0.6170257,1.2176411,1.3883078,2.8291285,2.5107694,1.8642052,1.6475899,1.9528207,4.5522056,3.6758976,2.3204105,2.1989746,3.7218463,2.674872,3.3805132,2.989949,1.3128207,0.82379496,0.81066674,1.4966155,2.5632823,4.0008206,6.088206,5.2578464,5.58277,7.1089234,9.232411,10.696206,8.595693,8.172308,8.648206,9.248821,9.199591,9.275078,10.098872,10.397539,9.5606165,7.643898,7.8408213,8.3364105,8.484103,8.188719,7.9195905,9.028924,9.3078985,9.521232,10.30236,12.1468725,12.06154,11.992617,11.145847,9.888822,9.764103,9.947898,10.112,10.272821,10.167795,9.278359,8.080411,8.329846,8.457847,7.8080006,6.636308,5.904411,5.172513,4.8016415,4.7950773,4.8049235,4.598154,4.4274874,4.5128207,4.857436,5.2480006,5.297231,5.3825645,5.6320004,5.973334,6.117744,5.7632823,5.080616,4.7327185,4.637539,3.9680004,3.6758976,3.3444104,3.314872,3.6594875,4.197744,4.2568207,3.9614363,3.6496413,3.4231799,3.1442053,3.0227695,2.477949,2.0742567,2.1792822,2.9604106,2.5698464,2.737231,2.8291285,2.7864618,3.1277952,3.05559,3.4494362,3.889231,4.1058464,3.9811285,3.895795,3.4100516,3.05559,3.1113849,3.6004105,4.8344617,5.9569235,6.7610264,7.256616,7.6603084,7.5881033,7.6242056,7.8441033,7.50277,5.034667,6.4754877,8.602257,9.291488,8.339693,7.460103,6.3507695,6.4656415,7.4075904,9.07159,11.674257,9.488411,8.960001,8.4972315,9.544206,16.587488,33.348927,24.372515,14.198155,12.383181,13.51877,4.096,2.6453335,2.809436,2.0742567,1.7690258,2.7109745,5.930667,8.375795,11.053949,19.012924,18.546873,8.956718,2.7175386,2.674872,2.0151796,1.3554872,1.4375386,6.380308,13.200411,11.808822,7.171283,9.4457445,12.074668,11.789129,8.5891285,4.1222568,2.9407182,2.861949,3.1934361,4.7294364,5.609026,4.713026,3.698872,3.2525132,3.0818465,4.0336413,4.0336413,4.2305646,4.8147697,5.034667,3.9844105,3.9253337,3.9417439,3.8137438,3.9975388,3.826872,3.4560003,3.045744,2.8750772,3.3280003,3.620103,4.2502565,4.3060517,3.7382567,3.370667,2.297436,2.6617439,3.4855387,4.2568207,4.9296412,4.0500517,3.948308,4.1682053,4.279795,3.876103,4.352,4.5522056,3.8629746,2.6978464,2.5009232,2.2580514,3.1113849,3.9548721,4.1222568,3.4034874,3.1967182,2.3368206,2.0086155,2.300718,2.228513,2.6912823,2.6157951,2.103795,1.5819489,1.8018463,1.4834872,1.148718,0.9944616,1.020718,1.024,1.0699488,0.955077,1.0666667,1.3423591,1.2832822,1.3062565,1.522872,1.8707694,2.0644104,1.5885129,1.3193847,1.3062565,1.4145643,1.6410258,2.1070771,2.2153847,3.0227695,3.3017437,2.8947694,2.6847181,3.4789746,4.125539,3.6857438,2.4516926,1.9364104,1.6804104,1.6344616,1.8937438,2.356513,2.7470772,2.5862565,2.8225644,2.8717952,2.6584618,2.609231,2.546872,2.6157951,2.7995899,2.9735386,2.8980515,3.0818465,3.5413337,3.889231,4.06318,4.31918,5.100308,5.943795,6.5312824,6.629744,6.1046157,6.226052,6.3573337,6.422975,6.180103,5.2020516,5.362872,5.464616,5.0084105,4.1878977,3.9056413,4.2962055,4.568616,5.661539,7.243488,7.719385,8.52677,8.78277,8.674462,8.536616,8.864821,8.999385,9.005949,8.864821,8.87795,9.659078,10.292514,10.8537445,11.116308,10.834052,9.734565,9.819899,8.999385,7.719385,6.705231,6.9743595,7.6701546,7.5881033,7.256616,7.4404106,9.124104,8.795898,8.667898,9.252103,10.587898,12.22236,11.063796,11.579078,11.864616,11.503591,11.54954,12.504617,13.170873,13.2562065,12.983796,13.108514,11.093334,10.177642,9.517949,8.707283,7.765334,7.7292314,8.956718,10.496001,11.805539,12.770463,12.698257,11.664412,10.985026,10.686359,9.4916935,12.005745,12.652308,12.274873,11.871181,12.603078,13.029744,12.744206,12.199386,11.9171295,12.465232,12.294565,11.785847,11.040821,10.197334,9.416205,8.937026,9.258667,9.783795,10.089026,9.91836,10.102155,10.505847,11.047385,11.2672825,10.315488,10.203898,10.433641,10.696206,10.896411,11.139283,1.5261539,1.6738462,1.9593848,2.1333334,1.9987694,1.4112822,1.7920002,2.3401027,2.5600002,2.5042052,2.7634873,3.6004105,4.588308,4.9362054,4.637539,4.457026,5.106872,5.024821,5.0510774,5.3070774,5.156103,5.211898,5.5926156,5.8256416,5.7665644,5.618872,5.618872,5.4843082,5.5171285,5.7074876,5.7140517,5.408821,5.3103595,5.346462,5.3792825,5.1922054,5.280821,5.536821,5.664821,5.5532312,5.284103,5.0018463,5.7107697,6.6428723,7.2336416,7.1122055,7.017026,6.055385,5.4186673,5.6320004,6.564103,6.7117953,6.6428723,6.774154,7.072821,7.02359,6.6100516,5.677949,5.792821,6.928411,7.4732313,8.050873,7.197539,6.5903597,6.6133337,6.373744,6.7085133,6.7544622,6.554257,6.3212314,6.436103,5.861744,5.930667,6.170257,6.245744,5.9667697,5.586052,5.3858466,5.32677,5.671385,6.994052,8.477539,9.508103,10.249847,10.778257,11.076924,11.16554,10.952206,10.771693,10.873437,11.441232,11.946668,12.6063595,12.84595,12.550565,12.07795,12.471796,12.905026,12.452104,11.1983595,10.213744,8.999385,8.740103,8.841846,8.822155,8.280616,7.276308,7.1680007,7.2336416,7.177847,7.1220517,6.76759,6.5444107,6.5050263,6.567385,6.5247183,6.0291286,6.2818465,6.6034875,6.747898,6.9021544,6.9645133,7.0531287,6.9776416,6.701949,6.3474874,6.3507695,6.485334,6.885744,7.6242056,8.681026,9.101129,9.865847,11.211488,13.180719,15.632411,16.259283,16.193642,16.170668,16.321642,16.187078,14.155488,13.292309,13.696001,14.621539,14.470565,14.79877,15.232001,15.07118,14.473847,14.444309,13.426873,13.285745,13.676309,14.36554,15.241847,15.140103,16.400412,17.152,16.89272,16.502155,13.5548725,11.034257,10.545232,11.976206,13.492514,12.327386,11.257437,10.752001,10.686359,10.361437,10.781539,12.166565,12.964104,12.73436,12.140308,11.424822,11.162257,10.86359,10.788103,11.956513,13.689437,14.106257,13.453129,12.63918,13.220103,12.888617,12.750771,12.970668,13.515489,14.155488,16.328207,16.662975,16.30195,16.216616,17.207796,17.778873,17.552412,17.536001,18.835693,22.639591,20.969027,19.288616,16.882874,14.385232,13.771488,12.895181,11.851488,12.12718,12.819694,10.637129,10.036513,9.416205,8.815591,8.264206,7.7718983,7.3058467,7.1483083,7.056411,7.2664623,8.484103,9.097847,8.736821,8.185436,7.762052,7.318975,7.253334,7.0498466,7.1581545,7.4863596,7.39118,6.8627696,6.2523084,5.9667697,6.0980515,6.413129,6.875898,7.532308,7.8047185,7.7357955,7.9786673,8.385642,7.768616,6.928411,6.121026,5.0642056,4.2830772,3.114667,2.5206156,2.5731285,2.4648206,1.9593848,1.1815386,0.7515898,0.90912825,1.4998976,1.2800001,1.1520001,1.1913847,1.2373334,0.8992821,1.0962052,1.8313848,2.3105643,2.3138463,2.2055387,1.585231,1.332513,1.5064616,3.5840003,10.456616,4.4438977,8.070564,11.073642,10.308924,9.744411,8.1066675,5.5762057,3.69559,2.868513,2.3696413,1.7887181,3.4691284,5.366154,5.989744,4.4045134,6.9677954,5.9602056,4.9887185,5.32677,5.924103,5.7632823,5.0084105,5.041231,5.98318,6.7282057,4.6867695,3.436308,2.3958976,1.4900514,1.148718,1.4211283,1.0962052,0.82379496,0.67282057,0.13784617,1.2537436,2.7142565,3.754667,3.6168208,1.5491283,1.142154,3.4658465,4.650667,5.5696416,11.83836,7.325539,2.6256413,0.6071795,1.0765129,0.7778462,1.6049232,1.8510771,1.467077,0.9682052,1.4408206,5.3103595,6.1768208,4.893539,3.2361028,3.892513,2.3860514,2.1136413,2.1924105,1.8838975,0.60389745,0.54482055,1.404718,2.5764105,3.8367183,5.3694363,5.044513,6.2129235,7.778462,9.091283,9.938052,8.602257,8.192,8.454565,8.845129,8.54318,8.996103,9.833026,9.9282055,8.910769,7.1680007,7.325539,8.024616,8.425026,8.247795,7.7718983,8.766359,9.4916935,9.908514,10.33518,11.424822,12.005745,11.497026,10.706052,10.272821,10.66995,10.345026,10.266257,9.885539,9.255385,9.009232,8.438154,8.720411,8.753231,8.162462,7.282872,6.2194877,5.1200004,4.6145644,4.6834874,4.634257,4.4865646,4.4110775,4.6244106,4.8836927,4.5029745,4.5029745,5.2676926,5.9963083,6.363898,6.5083084,5.737026,5.0576415,4.713026,4.4832826,3.6758976,3.498667,3.2853336,3.5183592,4.017231,3.9384618,4.2436924,4.1846156,3.9876926,3.7284105,3.3509746,3.062154,2.9013336,2.8160002,2.8389745,3.0818465,2.7602053,2.733949,2.7011285,2.6945643,3.05559,2.9144619,2.989949,3.4297438,3.9023592,3.6036925,3.7054362,3.6004105,3.4592824,3.4592824,3.7710772,4.466872,5.4941545,6.2588725,6.616616,6.8529234,6.567385,7.0925136,7.6734366,7.79159,7.171283,4.4406157,3.2361028,4.0467696,6.088206,7.2894363,7.565129,6.806975,5.412103,4.6572313,6.6822567,5.717334,7.1548724,9.386667,12.160001,16.587488,23.318975,14.25395,7.827693,9.980719,14.14236,4.023795,2.878359,3.7809234,3.3444104,1.719795,2.2514873,3.6102567,3.9778464,4.3618464,8.598975,14.483693,7.453539,2.294154,2.9604106,2.5632823,1.6016412,2.1497438,5.3234878,9.4457445,10.075898,9.265231,11.464206,14.953027,16.160822,9.6525135,4.578462,2.5731285,2.353231,2.986667,3.8990772,4.604718,3.9122055,3.3509746,3.3476925,3.2164104,4.5095387,4.414359,4.086154,4.0369234,4.1189747,3.3050258,3.4494362,3.7251284,3.9647183,4.644103,4.201026,4.381539,4.647385,4.6802053,4.4012313,4.164923,4.1452312,4.0402055,3.7907696,3.5905645,2.1267693,2.1792822,2.8324106,3.3575387,3.2196925,3.767795,4.0434875,4.135385,4.1025643,3.9745643,3.6496413,3.7743592,3.495385,2.7700515,2.3794873,2.6354873,3.186872,3.5577438,3.5183592,3.1113849,2.609231,2.0808206,2.0151796,2.2908719,2.1792822,2.0676925,1.9856411,1.6344616,1.1454359,1.0929232,1.1848207,1.3029745,1.2307693,1.0108719,0.9616411,1.1355898,1.1027694,1.086359,1.2077949,1.4900514,1.6607181,1.8116925,1.8904617,1.8018463,1.404718,1.3193847,1.4933335,1.4900514,1.3751796,1.7033848,2.1366155,2.6190772,2.6157951,2.4057438,3.0752823,4.007385,4.276513,3.6824617,2.7175386,2.5961027,1.9987694,1.9396925,2.1956925,2.5304618,2.6847181,2.537026,2.6420515,2.6847181,2.6387694,2.7569232,2.7044106,2.8192823,2.8849232,2.878359,2.9604106,2.9571285,3.4264617,3.9614363,4.263385,4.1485133,5.3103595,5.933949,6.38359,6.6527185,6.370462,6.5247183,6.2162056,6.4689236,6.961231,6.0324106,5.097026,4.7983594,5.0215387,5.284103,4.699898,4.768821,4.4242053,4.9887185,6.5280004,7.8539495,8.484103,8.720411,8.556309,8.172308,7.9261546,8.530052,8.884514,8.700719,8.146052,7.8637953,8.51036,9.43918,10.06277,10.052924,9.344001,8.766359,8.123077,7.27959,6.6067696,6.9743595,7.4929237,7.243488,6.948103,7.1056414,7.9885135,8.644924,8.530052,8.868103,9.741129,10.098872,9.5835905,11.270565,12.06154,11.234463,10.453334,12.107488,12.996924,13.174155,12.852514,12.386462,10.7158985,10.164514,10.036513,9.662359,8.388924,7.8047185,8.786052,10.515693,12.189539,13.026463,13.072412,11.83836,10.614155,10.059488,10.210463,11.428103,11.815386,11.759591,11.588924,11.579078,11.867898,11.401847,11.122872,11.329642,11.674257,11.122872,10.971898,11.090053,11.178667,10.758565,9.6754875,9.055181,9.163487,9.665642,9.6,9.199591,8.999385,9.416205,10.213744,10.509129,10.233437,10.200616,10.249847,10.266257,10.187488,1.6640002,1.7263591,1.8412309,2.0217438,2.0578463,1.5064616,1.7690258,2.3072822,2.7109745,2.937436,3.3050258,3.761231,4.644103,5.1922054,5.10359,4.529231,5.1298466,4.8114877,4.70318,5.0642056,5.3136415,5.1922054,5.280821,5.654975,5.979898,5.5302567,5.7042055,5.8880005,5.87159,5.681231,5.5926156,5.6352825,5.924103,5.9602056,5.5269747,4.6900516,4.95918,5.5729237,5.917539,5.8486156,5.7009234,5.037949,5.927385,6.8529234,7.125334,6.882462,6.8988724,6.7216415,6.38359,6.1374364,6.4590774,6.669129,6.560821,6.7216415,7.456821,8.776206,6.6067696,5.2709746,5.113436,5.8486156,6.554257,6.8365135,6.8266673,6.7117953,6.5444107,6.2785645,6.5312824,6.6592827,6.692103,6.744616,6.997334,6.518154,6.3540516,6.518154,6.7544622,6.5083084,6.042257,6.0980515,6.564103,7.4043083,8.661334,9.7214365,10.469745,10.837335,10.850462,10.620719,10.9456415,10.738873,10.909539,11.588924,12.153437,12.143591,11.949949,11.956513,12.202667,12.3995905,12.36677,11.949949,11.503591,11.116308,10.59118,9.475283,9.094564,8.736821,8.103385,7.318975,6.9743595,6.957949,6.944821,6.76759,6.416411,6.0717955,5.9963083,6.0750775,6.189949,6.226052,6.232616,6.1472826,6.1472826,6.265436,6.3934364,6.5312824,6.6494365,6.636308,6.439385,6.0685134,6.1472826,6.166975,6.3606157,6.954667,8.155898,9.222565,9.504821,9.829744,10.8307705,12.947693,13.873232,14.716719,14.8020525,14.185027,13.656616,13.459693,12.84595,13.387488,14.903796,15.442053,14.887385,15.169642,14.966155,14.227694,14.171899,13.59754,13.581129,14.441027,15.783386,16.49231,14.811898,14.795488,15.694771,16.754873,17.23077,14.404924,11.867898,11.277129,12.635899,14.306462,13.282462,12.3536415,12.051693,12.265027,12.196103,12.688411,13.167591,13.190565,12.694975,12.002462,11.956513,12.452104,12.626052,12.317539,12.071385,13.892924,14.736411,14.549335,13.8765135,13.840411,12.274873,11.569232,12.038565,13.29559,14.273643,15.75713,16.505438,16.423386,16.190361,17.26031,19.016207,18.625643,17.808413,18.057848,20.644104,21.435078,20.404514,18.17272,15.77354,14.657642,14.086565,13.161027,13.426873,14.421334,13.643488,10.971898,9.96759,9.3768215,8.677744,8.067283,7.4765134,7.509334,7.653744,8.064001,9.55077,9.639385,9.426052,9.133949,8.854975,8.546462,8.333129,7.9163084,7.709539,7.64718,7.194257,7.204103,6.669129,6.2129235,6.1308722,6.38359,7.2960005,7.817847,8.093539,8.132924,7.8473854,7.1122055,6.554257,6.3310776,6.12759,5.1298466,4.4406157,2.9144619,2.100513,2.1924105,2.038154,1.3751796,0.86317956,0.8992821,1.2832822,1.2077949,1.014154,0.90256417,1.020718,1.3620514,1.7493335,1.8018463,2.0545642,3.8564105,5.792821,3.6660516,1.8412309,3.0785644,3.2886157,3.3214362,8.950154,5.901129,5.7501545,6.1538467,6.232616,6.5805135,6.87918,4.585026,2.5764105,1.9954873,2.2449234,3.5413337,4.772103,5.225026,5.5565133,7.8047185,9.435898,7.3550773,6.193231,6.9645133,7.0531287,6.47877,5.477744,5.3398976,6.117744,6.626462,4.9099493,4.2929235,3.4560003,2.2580514,1.7394873,1.3587693,0.86317956,0.5284103,0.34789747,0.049230773,0.90912825,1.6311796,2.2482052,2.3696413,1.1749744,1.5786668,4.670359,6.1997952,7.194257,13.955283,5.1856413,1.4441026,0.51856416,0.6235898,0.37743592,1.8051283,4.3585644,4.1058464,1.5360001,1.5589745,4.3552823,4.8114877,3.948308,3.4198978,5.4843082,2.1825643,1.4178462,1.5688206,1.4473847,0.29210258,0.61374366,1.1520001,2.7733335,4.8377438,5.1987696,6.3573337,6.9710774,7.318975,7.8736415,9.301334,8.631796,8.546462,8.5661545,8.467693,8.283898,8.835282,9.478565,9.573745,8.937026,7.8637953,7.4404106,7.5191803,7.6964107,7.6077952,6.9677954,7.5585647,8.576,9.330873,9.665642,9.944616,11.392001,11.109744,10.473026,10.31877,10.932513,10.699488,10.368001,9.964309,9.531077,9.124104,8.3364105,8.060719,8.008205,7.8539495,7.243488,6.0980515,5.333334,4.8771286,4.634257,4.5029745,4.4340515,4.4307694,4.453744,4.394667,4.069744,4.6802053,5.349744,5.730462,5.8518977,6.121026,5.5958977,4.900103,4.266667,3.7316926,3.1540515,2.989949,2.930872,3.1638978,3.623385,3.9778464,4.4734364,4.352,4.066462,3.7940516,3.4494362,3.170462,3.2065644,3.2262566,3.1507695,3.1573336,2.5107694,2.4418464,2.3630772,2.228513,2.5140514,2.3860514,2.6026669,3.1245131,3.623385,3.508513,3.3345644,3.2328207,3.1770258,3.2623591,3.7152824,4.7458467,5.5007186,6.23918,6.7150774,6.186667,5.609026,6.1472826,7.1056414,7.9195905,8.162462,5.0051284,3.8564105,3.9647183,4.4734364,4.391385,4.896821,4.7950773,4.273231,4.082872,5.5138464,4.5095387,6.954667,9.662359,10.889847,10.325335,18.907898,13.088821,6.5739493,6.055385,11.195078,4.007385,4.532513,7.273026,7.968821,3.5872824,1.8084104,4.309334,5.218462,3.9122055,5.0084105,8.664616,4.6539493,2.4713848,3.8301542,2.665026,1.7427694,2.1300514,3.3903592,4.972308,6.2030773,6.5969234,7.4108725,9.685334,11.349334,7.1909747,4.3027697,2.6354873,2.3236926,2.917744,3.3805132,3.9318976,3.757949,3.4855387,3.4067695,3.4527183,3.7973337,3.626667,3.3050258,3.0490258,2.9210258,2.7634873,3.2689233,3.7743592,4.1714873,4.896821,5.221744,5.398975,5.2578464,4.9526157,4.972308,4.562052,4.453744,4.3618464,4.20759,4.1222568,3.0818465,2.789744,2.8127182,2.8882053,2.9472823,3.7185643,4.0434875,4.007385,3.9023592,4.197744,3.367385,3.2525132,3.0982566,2.7044106,2.4320002,2.678154,2.9997952,3.117949,2.9407182,2.5600002,2.353231,1.8510771,1.6902566,1.8281027,1.5524104,1.5392822,1.5392822,1.3456411,1.0338463,0.9714873,0.99774367,1.0666667,1.014154,0.8763078,0.88287187,1.1257436,1.2438976,1.2274873,1.2570257,1.6968206,2.0151796,1.8806155,1.8806155,1.9495386,1.3686155,1.2274873,1.2504616,1.2209232,1.2209232,1.6377437,2.2547693,2.6289232,2.6912823,2.6190772,2.8455386,3.6332312,4.2207184,4.0008206,3.2722054,3.255795,2.4713848,2.225231,2.300718,2.546872,2.8717952,2.865231,2.6715899,2.5731285,2.681436,2.9210258,3.2656412,3.3542566,3.2525132,3.114667,3.186872,3.121231,3.4264617,3.5741541,3.4494362,3.3345644,4.388103,5.175795,5.6976414,5.9667697,6.0192823,6.409847,6.445949,6.7249236,7.059693,6.498462,5.179077,4.7360005,4.841026,5.093744,5.024821,4.71959,4.9920006,5.5302567,6.311385,7.5881033,7.8145647,7.8441033,7.64718,7.509334,8.021334,8.211693,8.500513,8.195283,7.200821,6.0061545,6.550975,7.9524107,8.854975,8.763078,8.067283,8.083693,8.280616,8.050873,7.427283,7.066257,7.026872,6.5345645,6.294975,6.629744,7.466667,8.218257,8.283898,8.395488,8.572719,8.139488,8.277334,10.026668,10.427077,9.045334,7.9983597,10.459898,11.290257,11.35918,11.339488,11.703795,10.476309,10.066052,10.072617,10.026668,9.396514,8.388924,9.101129,10.752001,12.511181,13.4859495,13.11836,11.723488,10.20718,9.334154,9.714872,10.098872,10.312206,10.240001,9.95118,9.711591,10.9915905,10.70277,10.41395,10.765129,11.483898,11.401847,11.424822,11.392001,11.063796,10.14154,9.567181,9.07159,9.012513,9.321027,9.501539,9.012513,8.674462,8.858257,9.42277,9.718155,9.632821,9.577026,9.370257,9.091283,9.078155,1.7920002,1.9528207,2.0151796,2.166154,2.3269746,2.1431797,2.2416413,2.3860514,2.678154,3.1474874,3.751385,4.096,4.8049235,5.3858466,5.405539,4.4865646,4.8771286,4.709744,4.706462,5.0543594,5.3924108,5.5204105,5.5302567,5.9503593,6.432821,5.756718,5.425231,6.2162056,6.738052,6.4295387,5.5565133,5.6976414,5.868308,5.691077,5.110154,4.378257,4.565334,5.3924108,5.9995904,6.163693,6.298257,5.6320004,6.245744,6.9743595,7.2664623,7.1614366,6.9349747,7.0400004,6.764308,6.1997952,6.242462,6.363898,6.170257,6.4065647,7.259898,8.356103,6.052103,4.9427695,4.7524104,5.1987696,5.970052,5.7534366,6.048821,6.2818465,6.2720003,6.229334,6.121026,6.3376417,6.7807183,7.240206,7.381334,7.240206,6.9842057,6.9710774,7.128616,6.941539,6.813539,6.99077,7.634052,8.759795,10.223591,11.011283,11.648001,11.795693,11.277129,10.039796,10.7158985,10.893129,11.273847,11.992617,12.629334,12.58995,11.989334,11.782565,12.12718,12.412719,12.22236,11.040821,10.289231,10.308924,10.358154,9.412924,8.992821,8.310155,7.322257,6.7249236,6.7872825,6.678975,6.550975,6.409847,6.1046157,5.7435904,5.684513,5.730462,5.7435904,5.664821,5.930667,5.865026,5.8125134,5.858462,5.83877,5.9930263,6.1046157,6.0849237,5.9569235,5.83877,5.9503593,5.5696416,5.333334,5.6976414,6.9382567,8.303591,8.625232,8.713847,9.120821,10.148104,11.254155,12.301129,12.800001,12.694975,12.343796,12.836103,13.161027,13.745232,14.624822,15.42236,14.76595,15.491283,15.760411,14.956308,13.679591,13.699283,13.692719,14.464001,15.786668,16.387283,14.352411,13.748514,14.477129,15.8654375,16.66954,14.775796,13.344822,13.141335,13.906053,14.336001,13.774771,13.817437,14.503386,15.38954,15.553642,15.586463,15.067899,14.536206,13.948719,12.698257,12.960821,14.057027,14.907078,14.821745,13.495796,14.267078,14.880821,15.090873,14.795488,14.070155,12.57354,11.828514,12.097642,13.121642,14.12595,15.025232,16.114874,16.748308,17.027283,17.80513,19.094976,18.773335,17.690258,17.24718,19.373951,21.169233,20.151796,18.468103,17.089642,15.816206,15.284514,14.884104,15.360002,16.384,16.548103,12.268309,10.742155,10.056206,9.26195,8.375795,7.6143594,7.8539495,8.234667,8.681026,9.911796,9.6,9.508103,9.580308,9.737847,9.875693,10.240001,9.6065645,8.641642,7.7948723,7.273026,7.269744,6.941539,6.73477,6.8463597,7.2270775,7.821129,8.132924,8.39877,8.651488,8.717129,6.99077,6.0816417,6.0324106,6.235898,5.428513,4.381539,2.6847181,1.8116925,1.8576412,1.5458462,0.95835906,0.8402052,1.467077,2.176,1.3489232,1.4145643,1.1388719,1.0765129,1.4145643,1.9561027,2.0053334,2.1497438,4.2174363,6.4754877,3.6332312,3.1277952,4.056616,4.716308,5.6418467,9.622975,7.387898,4.9854364,4.7622566,7.066257,10.217027,7.4929237,4.3290257,2.3433847,2.3466668,4.3651285,5.2414365,5.4843082,5.4875903,6.3442054,9.826463,9.288206,8.280616,8.267488,8.723693,7.138462,6.5345645,5.543385,5.4580517,6.3868723,7.259898,5.789539,5.211898,4.394667,3.131077,2.15959,1.1552821,0.7450257,0.4594872,0.14769232,0.0,1.1093334,2.3794873,2.6322052,1.7723079,0.80738467,1.4473847,5.5204105,9.206155,11.080206,12.087796,3.0260515,0.73517954,0.56123084,0.30194873,0.20020515,1.9495386,5.9930263,5.9503593,2.100513,1.3883078,3.4330258,3.4330258,3.308308,4.1878977,6.3934364,2.7798977,2.169436,1.9167181,1.017436,0.098461546,0.81394875,1.1782565,2.5928206,4.4996924,4.384821,6.518154,7.145026,7.0859494,7.259898,8.690872,8.553026,8.854975,8.694155,8.12636,8.155898,8.4283085,8.838565,9.137232,9.084719,8.4512825,7.7423596,7.141744,6.7872825,6.6133337,6.3376417,6.675693,7.6668725,8.684308,9.206155,8.828718,10.345026,10.633847,10.381129,10.249847,10.889847,11.067078,10.564924,10.230155,10.108719,9.472001,8.385642,7.8112826,7.5946674,7.3780518,6.6100516,5.8092313,5.2348723,4.7589746,4.378257,4.2141542,4.204308,4.1517954,4.1025643,4.092718,4.1517954,4.854154,5.280821,5.533539,5.618872,5.4580517,5.028103,4.4767184,3.8662567,3.2951798,2.934154,2.8192823,2.8521028,2.9669745,3.2295387,3.8367183,4.397949,4.4274874,4.3027697,4.1550775,3.8629746,3.498667,3.4921029,3.4067695,3.1573336,3.0194874,2.231795,2.166154,2.1497438,2.0118976,2.0676925,1.9429746,2.1956925,2.5895386,2.9538465,3.2032824,2.937436,2.8225644,2.8488207,3.0687182,3.623385,4.5456414,5.041231,5.5991797,6.0324106,5.4547696,5.093744,5.504,6.4000006,7.53559,8.707283,6.872616,5.9963083,5.1626673,4.204308,3.7152824,3.190154,3.249231,3.7316926,4.6539493,6.229334,4.893539,5.8781543,8.306872,9.662359,5.7829747,13.574565,12.760616,7.394462,2.9243078,6.2063594,3.5282054,4.95918,9.081436,12.100924,7.8637953,3.6758976,5.6287184,8.618668,9.691898,8.054154,6.117744,2.861949,3.761231,7.968821,8.333129,7.463385,5.6320004,3.7415388,2.7536411,3.692308,3.4691284,3.8137438,5.2381544,6.62318,5.225026,4.240411,3.0949745,2.540308,2.7076926,3.0884104,3.3214362,3.1770258,3.0490258,3.0916924,3.2328207,2.9243078,2.7273848,2.5600002,2.4713848,2.6518977,2.9243078,3.5314875,4.092718,4.5128207,4.95918,5.5072823,5.58277,5.097026,4.4767184,4.673641,4.516103,4.7261543,4.7524104,4.4832826,4.2502565,3.6562054,3.0916924,2.7831798,2.861949,3.3575387,3.5774362,3.757949,3.6693337,3.501949,3.8695388,3.0818465,2.8324106,2.6945643,2.5665643,2.6715899,2.6584618,2.8258464,2.8356924,2.546872,2.0118976,2.0578463,1.6804104,1.4572309,1.4769232,1.3259488,1.2832822,1.2504616,1.1126155,0.9419488,1.0010257,1.017436,0.9682052,0.955077,1.0075898,1.0765129,1.1158975,1.2832822,1.3915899,1.4441026,1.6344616,1.8740515,1.8642052,1.9659488,2.0775387,1.6049232,1.4802053,1.214359,1.0568206,1.1552821,1.585231,2.048,2.5304618,2.8849232,3.0424619,3.0030773,3.5183592,4.2863593,4.31918,3.6857438,3.511795,3.1409233,2.7831798,2.6026669,2.6453335,2.8225644,3.1245131,3.1671798,3.3312824,3.5511796,3.3247182,3.4691284,3.5282054,3.4166157,3.2262566,3.2229745,3.18359,3.2623591,3.1245131,2.8291285,2.8488207,3.515077,4.46359,5.1265645,5.405539,5.651693,6.009436,6.1046157,6.5870776,7.2205133,6.875898,5.792821,5.3202057,5.353026,5.5663595,5.4482055,4.7524104,5.2578464,5.674667,5.76,6.3179493,6.232616,6.2588725,6.2687182,6.51159,7.634052,7.9195905,8.004924,7.5191803,6.409847,4.9132314,4.8804107,6.232616,7.240206,7.200821,6.416411,7.4404106,8.224821,8.375795,7.821129,6.806975,6.498462,6.189949,6.1078978,6.482052,7.5520005,7.643898,8.14277,8.576,8.530052,7.6635904,7.752206,8.681026,8.490667,7.138462,6.498462,8.953437,9.872411,10.013539,10.115283,10.880001,9.846154,9.734565,9.888822,9.997129,10.098872,9.5606165,10.092308,11.2672825,12.570257,13.380924,13.22995,11.802258,10.049642,8.881231,9.170052,9.567181,9.777231,9.45559,8.851693,8.825437,10.594462,10.443488,10.203898,10.656821,11.526565,11.546257,11.437949,11.362462,11.047385,9.810052,9.580308,9.393231,9.380103,9.488411,9.4916935,9.035488,8.700719,8.667898,8.871386,8.996103,8.992821,8.871386,8.562873,8.218257,8.211693,1.9068719,2.1891284,2.3171284,2.5271797,2.8488207,3.1081028,3.1474874,2.8192823,2.7437952,3.121231,3.7284105,4.1878977,4.713026,5.3202057,5.5696416,4.588308,4.598154,4.7261543,5.0215387,5.35959,5.4416413,5.8945646,6.2687182,6.7577443,7.059693,6.373744,5.10359,6.3179493,7.5454364,7.4371285,5.7764106,5.431795,5.031385,4.6080003,4.3027697,4.388103,4.2502565,5.0182567,5.930667,6.5936418,6.9776416,6.5378466,6.4754877,6.931693,7.6274877,7.830975,7.2172313,6.8594875,6.449231,6.088206,6.2916927,5.930667,5.8420515,6.2720003,6.7872825,6.2720003,5.3070774,4.5554876,4.5095387,5.1265645,5.8157954,5.2512827,5.284103,5.612308,5.9602056,6.0750775,5.674667,5.8157954,6.426257,7.1023593,7.138462,7.3419495,7.00718,6.8266673,6.9776416,7.1056414,7.450257,7.637334,8.057437,8.999385,10.650257,11.648001,12.389745,12.612924,11.976206,10.049642,10.630565,11.204924,11.605334,11.956513,12.704822,12.973949,12.626052,12.314258,12.182976,11.861334,11.923694,10.57477,9.45559,9.248821,9.701744,8.999385,8.572719,7.9097443,7.1187696,6.9349747,6.7872825,6.4689236,6.2752824,6.235898,6.11118,5.730462,5.586052,5.4613338,5.293949,5.1659493,5.156103,5.356308,5.5762057,5.6976414,5.7009234,5.717334,5.720616,5.609026,5.4383593,5.412103,5.2545643,4.5522056,4.1156926,4.388103,5.435077,6.5936418,7.2336416,7.755488,8.251078,8.523488,9.540924,9.91836,10.712616,11.861334,12.202667,11.861334,13.059283,13.804309,13.856822,14.736411,14.54277,15.80636,16.807386,16.39713,14.017642,14.319591,14.158771,14.191591,14.598565,15.07118,13.935591,13.948719,14.473847,15.064616,15.451899,14.552616,14.519796,15.015386,15.392821,14.670771,14.500104,15.547078,17.10277,18.395899,18.609232,18.507488,17.706669,17.027283,16.357744,14.644514,14.647796,15.445334,16.489027,17.004309,15.980309,15.07118,14.867694,15.031796,15.05477,14.283488,13.846975,13.581129,13.298873,13.272616,14.234258,15.07118,16.147694,17.165129,17.99549,18.694565,18.386053,17.860924,17.024002,16.846771,19.373951,20.46359,19.029335,18.051283,18.031591,16.95836,16.31836,16.784412,18.136618,19.383797,18.747078,13.732103,11.894155,11.283693,10.587898,9.120821,7.9885135,8.211693,8.713847,9.147078,9.895386,9.475283,9.321027,9.478565,9.91836,10.528821,11.989334,11.352616,9.741129,8.178872,7.584821,7.030154,6.928411,7.204103,7.778462,8.5661545,8.385642,8.615385,8.904206,9.222565,9.869129,7.7718983,6.5050263,6.1768208,6.2490263,5.536821,4.089436,2.428718,1.6968206,1.723077,1.017436,0.77128214,1.2406155,2.4484105,3.4822567,2.4713848,2.353231,1.7920002,1.3686155,1.2800001,1.3751796,1.2898463,1.467077,3.3509746,5.5958977,4.082872,5.4416413,4.1878977,6.114462,11.227899,13.761642,8.973129,7.683283,10.210463,15.317334,20.187899,10.820924,5.0576415,2.665026,3.3444104,6.744616,5.9470773,5.549949,6.173539,7.75877,9.544206,7.3485136,8.283898,9.747693,9.764103,6.9710774,6.413129,5.536821,5.7042055,7.0137444,8.303591,6.820103,5.8256416,4.841026,3.636513,2.2055387,0.9419488,0.71548724,0.54482055,0.17723078,0.11158975,1.9528207,4.7917953,5.1200004,2.6715899,0.4201026,0.9878975,4.9952826,10.545232,13.515489,7.5585647,3.0687182,1.4178462,0.86974365,0.4955898,0.18379489,1.6443079,5.3103595,5.353026,1.8642052,0.8598975,2.8324106,2.9833848,3.751385,5.3924108,6.009436,3.9909747,3.7973337,2.8553848,0.92225647,0.06564103,1.0108719,1.5327181,2.1169233,2.789744,3.121231,5.412103,6.7085133,7.3386674,7.7325134,8.41518,8.576,9.186462,8.966565,8.03118,7.9097443,7.8080006,8.195283,8.78277,9.124104,8.63836,8.096821,7.210667,6.3310776,5.832206,6.117744,6.5772314,7.318975,8.293744,8.989539,8.4283085,9.130668,9.852718,10.115283,10.115283,10.738873,11.300103,10.79795,10.433641,10.354873,9.619693,8.687591,8.3593855,7.9885135,7.204103,5.914257,5.5269747,4.781949,4.240411,4.06318,3.9876926,4.069744,3.82359,3.7973337,4.1222568,4.5390773,4.7360005,4.95918,5.353026,5.586052,4.84759,4.348718,4.07959,3.7874875,3.4133337,3.0949745,3.121231,3.1442053,3.1409233,3.2131286,3.5741541,4.023795,4.3585644,4.535795,4.532513,4.33559,3.8662567,3.757949,3.5774362,3.1934361,2.7831798,2.1431797,2.0118976,2.0676925,2.100513,2.0151796,1.9003079,1.9429746,2.0020514,2.1300514,2.5895386,2.609231,2.537026,2.6223593,2.9604106,3.495385,3.7087183,4.086154,4.44718,4.7294364,4.9788723,5.1298466,5.35959,5.8420515,6.816821,8.612103,8.28718,7.13518,5.8125134,5.0838976,5.832206,4.2863593,3.6594875,3.826872,4.827898,6.8660517,5.7009234,4.210872,5.986462,8.973129,5.4547696,6.75118,9.504821,7.460103,2.0808206,2.5238976,3.3312824,3.895795,7.860513,13.37436,13.092104,8.4283085,6.7117953,10.056206,15.268104,13.869949,6.9743595,2.556718,5.172513,12.757335,16.62359,16.764719,12.314258,7.39118,4.414359,4.07959,2.2383592,3.0030773,4.6539493,5.786257,5.3169236,4.8804107,3.9089234,2.989949,2.5698464,2.9702566,2.7798977,2.2121027,2.0676925,2.409026,2.5764105,2.4451284,2.1989746,2.0906668,2.3335385,3.0982566,3.3542566,3.757949,4.3290257,4.9099493,5.172513,4.9329233,4.965744,4.588308,3.9154875,3.8596926,4.1485133,4.667077,4.7589746,4.33559,3.8728209,3.515077,2.92759,2.7634873,3.1540515,3.7218463,3.2853336,3.2918978,3.239385,3.0490258,3.0785644,2.7076926,2.5173335,2.4024618,2.4451284,2.9144619,2.7109745,2.6683078,2.540308,2.2121027,1.6902566,1.7099489,1.5983591,1.5163078,1.5524104,1.7394873,1.3784616,1.1946667,1.0404103,0.9321026,1.0305642,1.1520001,1.1158975,1.204513,1.4309745,1.5524104,1.4112822,1.5655385,1.7985642,1.9068719,1.6771283,1.6771283,1.9922053,2.1497438,2.03159,1.8740515,1.975795,1.5425643,1.204513,1.2077949,1.4276924,1.5491283,2.1234872,2.7011285,3.1113849,3.4592824,3.9187696,4.594872,4.565334,3.8432825,3.3903592,3.6693337,3.43959,3.1376412,2.9472823,2.7766156,3.3476925,3.9614363,4.5029745,4.6178465,3.6758976,3.2000003,3.2820516,3.3575387,3.2295387,3.0687182,3.05559,2.9702566,2.865231,2.8356924,3.0194874,3.3214362,4.1747694,4.84759,5.1298466,5.333334,5.366154,5.0609236,5.802667,7.171283,6.9382567,6.4722056,6.055385,6.2129235,6.636308,6.180103,5.362872,5.477744,5.586052,5.35959,5.077334,4.7524104,4.8311796,5.024821,5.4383593,6.554257,7.4765134,7.4732313,6.9842057,6.1440005,4.7589746,4.010667,4.7950773,5.651693,5.7796926,5.0576415,6.701949,7.4863596,7.712821,7.3780518,6.157129,5.9569235,6.0619493,6.1308722,6.422975,7.788308,7.2631803,8.021334,9.015796,9.383386,8.470975,7.936001,7.899898,7.312411,6.3310776,6.3179493,8.008205,9.225847,9.7903595,9.905231,10.177642,9.074872,9.163487,9.511385,9.764103,10.151385,10.6469755,11.247591,11.897437,12.501334,12.931283,13.170873,11.772718,10.029949,8.956718,9.258667,9.93477,10.138257,9.593436,8.795898,9.025641,10.423796,10.427077,10.407386,10.893129,11.562668,11.113027,10.735591,10.902975,11.204924,10.328616,10.043077,9.888822,9.9282055,9.93477,9.386667,8.960001,8.592411,8.41518,8.467693,8.681026,8.52677,8.293744,8.093539,7.955693,7.837539,2.1530259,2.103795,2.2646155,2.7700515,3.5249233,4.194462,4.0369234,3.7054362,3.4560003,3.373949,3.387077,3.9253337,4.644103,5.4514875,5.930667,5.356308,4.8672824,5.0116925,5.3727183,5.5991797,5.4153852,5.540103,6.4295387,7.4075904,7.899898,7.460103,5.789539,6.452513,7.2861543,7.27959,6.5444107,5.2512827,4.8738465,4.8738465,4.900103,4.7917953,4.7294364,4.926359,5.756718,6.9152827,7.4141545,7.427283,7.1023593,7.2237954,7.6964107,7.5388722,7.0990777,6.925129,6.8988724,6.87918,6.6822567,5.9995904,6.0849237,6.377026,6.491898,6.2096415,5.5893335,5.110154,5.0084105,5.156103,5.097026,5.402257,5.7632823,6.1538467,6.308103,5.720616,5.805949,6.0947695,6.308103,6.3442054,6.2720003,6.514872,5.6976414,5.58277,6.5050263,7.384616,7.5552826,8.211693,8.864821,9.380103,9.980719,11.113027,11.398565,11.634872,11.795693,11.001437,10.732308,11.204924,12.071385,12.911591,13.22995,13.5089245,13.443283,12.980514,12.337232,12.009027,11.336206,9.888822,8.874667,8.858257,9.750975,10.043077,9.373539,8.598975,7.896616,6.774154,6.5312824,6.416411,6.2063594,5.8420515,5.402257,5.2676926,5.2709746,5.2348723,5.1659493,5.2644105,4.972308,4.8147697,4.926359,5.35959,6.1046157,6.091488,5.970052,5.7796926,5.421949,4.6539493,3.7743592,3.3903592,3.4330258,3.7874875,4.2863593,4.9460516,5.7435904,6.6592827,7.4240007,7.522462,7.8145647,8.592411,9.504821,10.420513,11.460924,11.556104,10.896411,11.175385,12.649027,14.112822,13.627078,14.549335,15.908104,16.774565,16.249437,15.858873,15.094155,14.385232,14.106257,14.555899,14.165335,14.772514,15.573335,15.95077,15.488001,14.316309,14.244103,14.828309,15.891693,17.503181,17.08636,17.460514,18.392616,19.416616,19.80718,20.952618,20.808207,19.784206,18.454975,17.562258,16.502155,16.006565,16.567797,17.752617,18.202257,16.774565,15.776822,15.24513,15.113848,15.199181,15.465027,15.543797,15.084309,14.575591,15.320617,16.088617,16.738462,16.764719,16.853334,18.891489,19.157335,18.228514,17.460514,17.332514,17.457232,19.055592,18.786463,19.134361,19.984411,18.632206,17.824821,18.806156,21.691078,24.031181,20.79836,15.110565,13.174155,12.911591,12.698257,11.369026,9.025641,8.402052,8.63836,9.275078,10.240001,9.93477,9.682052,9.133949,8.697436,9.55077,11.529847,11.52,10.525539,9.147078,7.584821,6.669129,6.547693,6.7807183,7.3091288,8.467693,8.444718,9.26195,9.800206,9.760821,9.6754875,7.39118,6.6560006,6.4557953,6.0849237,5.156103,3.9253337,2.1431797,1.5458462,1.8215386,0.6268718,0.7220513,2.1858463,3.8137438,4.6933336,4.1813335,2.7044106,2.0676925,2.0873847,2.2055387,1.5097437,1.6082052,1.4309745,6.4295387,13.88636,12.908309,8.123077,5.674667,10.148104,17.742771,16.265848,9.45559,6.954667,11.592206,19.771078,21.4679,10.079181,3.8990772,2.0676925,3.1803079,5.280821,5.8289237,5.930667,7.450257,9.714872,9.504821,8.297027,7.3550773,8.3364105,9.974154,8.057437,7.4207187,6.6592827,6.928411,8.024616,8.375795,6.5706673,5.5958977,4.522667,3.121231,1.8773335,0.7778462,0.4397949,0.2855385,0.2100513,0.56451285,2.7733335,6.547693,7.9524107,5.6451287,0.88615394,2.0086155,2.0611284,4.6178465,8.254359,6.547693,5.142975,2.6584618,1.4998976,1.5491283,0.18379489,1.5753847,3.4527183,2.858667,0.50543594,0.761436,1.3850257,1.4966155,3.0096412,5.3005133,5.2020516,4.7392826,4.3027697,2.8455386,0.8008206,0.09189744,1.1520001,1.8871796,2.0939488,2.1464617,2.9768207,5.4908724,6.2916927,7.2270775,8.595693,9.170052,9.242257,10.066052,9.938052,8.618668,7.325539,7.397744,8.3134365,9.02236,9.176616,9.140513,8.674462,8.067283,7.0826674,6.0685134,5.937231,6.9120007,7.5421543,7.9195905,8.149334,8.329846,8.185436,8.533334,9.107693,9.77395,10.545232,11.057232,10.781539,10.368001,9.888822,8.851693,8.838565,9.009232,8.73354,7.7456417,6.1341543,5.32677,4.466872,4.1091285,4.269949,4.4406157,4.7950773,4.2863593,3.9023592,4.06318,4.6244106,4.7327185,4.532513,4.378257,4.394667,4.457026,4.5029745,4.414359,4.1058464,3.6430771,3.2656412,3.498667,3.4100516,3.4034874,3.5872824,3.767795,3.9154875,4.07959,4.020513,3.82359,3.9220517,3.761231,3.879385,4.0500517,3.892513,2.868513,2.2580514,1.8871796,1.8018463,1.9889232,2.3794873,2.3926156,2.2777438,2.1070771,1.9659488,1.9528207,2.4057438,2.1956925,2.1530259,2.553436,3.1277952,3.0293336,3.5183592,4.07959,4.650667,5.61559,5.579488,5.405539,5.733744,6.4754877,6.806975,7.0367184,6.6822567,6.1472826,5.989744,6.941539,7.026872,6.180103,4.916513,4.204308,5.4613338,5.586052,5.0116925,5.0609236,5.85518,6.3310776,3.8301542,3.892513,4.1780515,4.194462,5.293949,5.428513,3.4658465,5.146257,10.896411,15.839181,14.933334,8.254359,4.775385,7.79159,14.907078,6.4590774,2.3729234,4.1911798,10.240001,15.609437,19.98113,17.243898,13.223386,10.194052,6.9120007,3.3214362,3.0851285,5.037949,7.1581545,6.560821,6.232616,5.031385,3.879385,3.2131286,3.006359,2.6026669,2.0184617,1.6508719,1.6836925,2.0742567,2.4549747,1.9528207,1.7033848,2.0611284,2.609231,2.6223593,2.8521028,3.7809234,5.159385,6.0258465,4.634257,4.525949,4.342154,3.7874875,3.6168208,3.9811285,4.1485133,4.020513,3.7021542,3.495385,3.4691284,3.3903592,3.4133337,3.4921029,3.3575387,3.0752823,3.0326157,3.058872,2.993231,2.7011285,2.5042052,2.4746668,2.4385643,2.4516926,2.793026,2.8521028,2.2449234,1.6836925,1.5327181,1.8018463,1.654154,1.6278975,1.8215386,2.1431797,2.28759,1.8018463,1.5425643,1.4605129,1.4211283,1.1913847,1.1158975,1.1979488,1.4605129,1.8084104,2.028308,2.5435898,2.8816411,3.0030773,2.9472823,2.8389745,2.7766156,2.5862565,2.300718,1.9462565,1.5556924,2.0676925,1.913436,1.6311796,1.4539489,1.2832822,1.3554872,1.5195899,1.7690258,2.1989746,3.006359,4.1911798,5.0642056,4.903385,3.9384618,3.3411283,3.318154,3.5314875,3.5741541,3.4724104,3.692308,4.059898,4.4438977,4.381539,3.8367183,3.190154,2.993231,3.18359,3.511795,3.6332312,3.0818465,2.9604106,2.8914874,2.930872,3.1277952,3.5544617,3.895795,4.2830772,4.5456414,4.6276927,4.578462,4.4438977,4.007385,4.4701543,5.6451287,5.9503593,6.0980515,5.924103,5.861744,6.2030773,7.0957956,6.9743595,7.171283,7.200821,6.921847,6.5312824,5.687795,5.175795,4.827898,4.857436,5.858462,6.665847,6.8955903,7.02359,6.7610264,5.0510774,4.4898467,4.850872,5.1954875,5.1167183,4.775385,5.924103,6.3474874,6.633026,6.633026,5.4613338,5.280821,5.1331286,5.07077,5.5171285,7.2631803,7.6176414,7.5421543,8.182155,9.216001,8.851693,8.080411,8.182155,7.466667,6.0619493,5.8912826,7.062975,8.52677,9.803488,10.496001,10.299078,9.176616,8.484103,8.73354,9.527796,9.55077,10.236719,11.35918,12.25518,12.78359,13.321847,12.087796,10.515693,9.649232,9.7214365,10.161232,9.882257,9.619693,9.278359,8.904206,8.697436,9.770667,10.469745,10.7158985,10.817642,11.490462,10.807796,10.469745,10.417232,10.509129,10.55836,10.643693,10.226872,9.938052,9.754257,8.973129,8.690872,8.192,7.9228725,8.034462,8.375795,8.083693,7.965539,7.9885135,8.067283,8.057437,2.2613335,2.1234872,2.4681027,3.249231,4.06318,4.1583595,4.138667,3.7940516,3.370667,2.9604106,2.5337439,3.245949,4.1550775,5.1364107,5.901129,5.989744,5.7764106,5.8912826,6.170257,6.380308,6.235898,6.550975,7.171283,7.653744,7.6734366,7.0104623,5.865026,6.432821,7.0104623,6.820103,6.009436,5.536821,5.2020516,4.9132314,4.6933336,4.6802053,4.775385,5.2315903,6.173539,7.0531287,6.633026,7.2336416,6.928411,6.669129,6.7840004,6.9776416,6.8496413,6.7610264,6.7905645,6.9120007,7.000616,6.7085133,6.482052,6.242462,5.940513,5.549949,5.730462,5.6287184,5.658257,5.664821,4.9493337,4.893539,5.0838976,5.1167183,4.9493337,4.8804107,5.228308,5.536821,5.730462,5.85518,6.0652313,5.76,5.8256416,6.304821,6.8660517,6.8004107,6.7150774,7.427283,8.454565,9.711591,11.480617,13.046155,13.495796,13.24636,12.652308,12.015591,10.817642,11.264001,11.72677,11.782565,12.228924,12.324103,12.386462,12.028719,11.32636,10.811078,10.551796,9.77395,9.32759,9.43918,9.714872,9.488411,8.92718,8.28718,7.686565,7.0793853,6.8365135,6.442667,5.976616,5.536821,5.2414365,5.0018463,4.8836927,4.8016415,4.716308,4.630975,4.6966157,4.7556925,4.916513,5.1889234,5.504,5.4449234,5.435077,5.2611284,4.850872,4.2863593,3.6627696,3.318154,3.370667,3.7448208,4.164923,4.5817437,5.6976414,6.3540516,6.422975,6.803693,7.328821,8.687591,9.580308,9.783795,10.115283,10.029949,9.993847,10.28595,10.902975,11.588924,11.559385,12.3306675,14.024206,16.105026,17.398155,17.56554,15.031796,13.377642,13.525334,13.764924,13.410462,14.930053,16.321642,16.33477,14.473847,15.314053,14.959591,14.677335,15.07118,16.098463,16.981335,16.984617,17.316103,18.15631,18.635489,19.99754,20.867283,20.548925,19.18031,17.723078,15.908104,15.409232,15.763694,16.449642,16.873028,16.617027,15.809642,15.218873,15.153232,15.455181,15.78995,15.445334,14.539488,13.722258,14.171899,15.156514,16.298668,16.79754,16.922258,18.025026,19.590565,18.999796,17.946259,17.28,16.99118,18.57313,18.838976,18.405745,18.320412,20.069746,19.423182,20.184616,23.08595,25.77395,22.810259,17.417847,15.172924,14.418053,13.925745,12.918155,10.9456415,9.544206,8.743385,8.730257,9.8592825,9.819899,10.036513,9.55077,8.641642,8.832001,10.000411,10.781539,10.594462,9.386667,7.6701546,6.774154,6.4032826,6.088206,5.933949,6.626462,7.351795,8.79918,9.875693,10.112,9.626257,6.931693,6.088206,6.1538467,6.1374364,4.97559,4.06318,2.2449234,1.3718976,1.5261539,1.0043077,1.522872,3.045744,3.259077,2.038154,1.4473847,1.9331284,5.0116925,9.110975,12.140308,11.483898,10.253129,8.484103,9.186462,10.174359,4.073026,3.9844105,4.634257,7.1876926,10.010257,8.661334,6.0291286,3.9318976,6.7905645,13.433437,17.076513,6.301539,2.3762052,2.9538465,5.169231,5.658257,6.8430777,7.0432825,7.9950776,9.741129,10.617436,10.765129,8.329846,8.477539,10.66995,8.65477,6.409847,6.2030773,7.213949,8.224821,7.634052,6.442667,5.5204105,4.1550775,2.4910772,1.4998976,0.90912825,0.8992821,0.9419488,1.1552821,2.3105643,2.0086155,3.751385,5.1856413,4.5095387,0.46933338,0.93866676,2.5632823,5.3792825,7.680001,6.0225644,6.764308,3.2820516,2.3860514,4.0992823,1.6475899,1.0371283,1.9003079,1.8740515,1.0929232,2.1792822,3.4264617,3.4002054,3.8006158,4.348718,2.7864618,3.945026,3.0129232,1.8149745,1.2077949,1.0568206,1.8838975,2.3302567,2.9768207,3.6430771,3.3903592,4.9099493,5.937231,7.0531287,8.260923,9.012513,9.4457445,10.105436,10.072617,9.40636,9.117539,8.3823595,8.641642,8.973129,9.061745,9.199591,8.628513,8.300308,8.021334,7.686565,7.27959,8.303591,8.484103,8.027898,7.4240007,7.4404106,7.4896417,7.7390776,8.411898,9.432616,10.44677,10.528821,10.368001,10.299078,10.138257,9.16677,9.058462,8.946873,8.36595,7.253334,5.9634876,5.146257,4.322462,4.020513,4.279795,4.634257,4.5095387,4.2207184,4.138667,4.3027697,4.414359,4.71959,5.031385,4.778667,4.1583595,4.1025643,3.9253337,3.8104618,3.761231,3.8104618,3.9975388,4.414359,4.3585644,4.197744,4.086154,3.9778464,4.141949,4.027077,3.8038976,3.7251284,4.1058464,3.8104618,3.9056413,3.945026,3.6594875,2.9669745,2.425436,2.156308,2.0512822,2.028308,2.038154,2.2646155,2.0709746,2.0118976,2.0512822,1.5491283,1.9823592,2.481231,2.7503593,2.9046156,3.4691284,3.7054362,3.6758976,3.7284105,3.9680004,4.2469745,4.886975,4.785231,5.044513,5.8945646,6.6822567,5.937231,5.802667,5.9667697,6.229334,6.47877,6.9842057,7.1647186,6.8266673,6.157129,5.6943593,6.882462,6.9842057,7.062975,6.7544622,4.2830772,3.31159,3.882667,4.926359,5.76,6.0750775,5.3202057,4.381539,4.7327185,7.1581545,11.762873,22.038977,15.012104,6.5936418,4.9920006,10.722463,7.0990777,4.5423594,4.923077,6.813539,5.5138464,10.568206,12.517745,11.713642,8.5202055,3.31159,4.906667,5.7764106,7.5913854,10.210463,11.664412,11.218052,10.538668,9.31118,7.27959,4.2502565,2.5993848,1.8543591,1.5688206,1.5819489,2.0020514,2.3302567,2.0086155,4.0992823,7.1122055,5.0149746,2.92759,2.7798977,3.7087183,4.9296412,5.7468724,4.4438977,3.892513,3.515077,3.1967182,3.2984617,4.0369234,3.3214362,2.7175386,2.7536411,2.8947694,3.2820516,3.2754874,3.2656412,3.2361028,2.7602053,2.3991797,2.1924105,2.156308,2.2350771,2.2744617,2.284308,2.612513,2.7798977,2.6518977,2.425436,2.537026,2.0808206,1.595077,1.3489232,1.3259488,1.4309745,1.4473847,1.6672822,2.0053334,1.9954873,1.6935385,1.3981539,1.2865642,1.3718976,1.5195899,1.3883078,1.5786668,1.6902566,1.6640002,1.785436,1.8674873,1.9987694,2.044718,1.9856411,1.8871796,2.3827693,2.6453335,2.8127182,2.8160002,2.3860514,2.1267693,1.7657437,1.5130258,1.394872,1.2340513,1.3653334,1.7493335,1.9889232,2.2711797,3.3608208,4.71959,4.9920006,4.5390773,3.6857438,2.7076926,3.0162053,2.9538465,2.92759,3.1803079,3.7907696,3.9712822,3.826872,3.8367183,4.066462,4.1517954,3.8695388,3.7218463,3.5478978,3.2164104,2.6190772,2.789744,2.9210258,2.9768207,3.0162053,3.190154,3.9023592,4.44718,4.578462,4.384821,4.2962055,4.2601027,3.9811285,4.1156926,4.525949,4.2535386,4.3716927,4.5554876,5.031385,5.5762057,5.5204105,5.0576415,4.9854364,5.0477953,5.07077,4.9920006,5.146257,4.788513,4.5128207,4.7491283,5.7501545,5.4613338,5.8420515,6.5083084,6.810257,5.8453336,4.8344617,4.578462,4.7360005,4.8672824,4.457026,5.5269747,6.482052,6.9349747,6.5870776,5.2315903,5.077334,4.923077,4.9887185,5.4514875,6.445949,7.2205133,7.0367184,7.7357955,9.334154,10.023385,8.372514,7.8506675,7.387898,6.5706673,5.658257,6.7216415,8.123077,9.101129,9.563898,10.092308,9.143796,8.3364105,8.254359,8.779488,9.074872,9.544206,10.174359,10.748719,11.08677,11.0375395,10.489437,9.796924,9.921641,10.725744,10.981745,9.616411,9.366975,9.156924,8.546462,7.7325134,8.533334,9.156924,9.196308,9.042052,9.878975,9.977437,9.563898,9.416205,9.708308,10.023385,10.371283,10.115283,9.728001,9.42277,9.130668,9.084719,8.592411,8.4053335,8.677744,8.950154,8.618668,8.402052,8.503796,8.65477,8.1066675,2.1070771,2.4976413,3.2656412,3.8990772,4.1747694,4.1780515,4.3290257,3.882667,3.4625645,3.3411283,3.4264617,4.0008206,4.8640003,5.5729237,5.970052,6.166975,6.0783596,6.4295387,6.7971287,6.8529234,6.36718,6.957949,7.27959,7.387898,7.213949,6.557539,6.1078978,6.363898,6.6527185,6.4065647,5.159385,4.8705645,4.772103,4.6178465,4.384821,4.279795,4.6539493,5.0904617,5.8518977,6.685539,6.813539,7.0465646,6.482052,6.2884107,6.6625648,6.816821,6.629744,6.770872,6.744616,6.6592827,7.1909747,6.695385,6.626462,6.485334,6.166975,5.9634876,6.0061545,6.1768208,6.12759,5.7009234,4.9329233,4.71959,5.034667,5.169231,5.0084105,5.0543594,4.6933336,4.824616,4.926359,4.969026,5.425231,5.2053337,5.681231,6.370462,6.8529234,6.7807183,6.633026,7.253334,8.3823595,10.029949,12.458668,13.59754,13.66318,13.541744,13.466257,13.036308,11.946668,11.739899,11.762873,11.851488,12.327386,12.337232,12.235488,11.680821,10.771693,10.066052,9.95118,9.747693,9.803488,10.003693,9.796924,9.954462,9.419488,8.585847,7.709539,6.918565,6.6822567,6.196513,5.756718,5.4416413,5.1200004,4.8607183,4.7622566,4.6112823,4.3290257,3.9778464,3.892513,4.1058464,4.417641,4.644103,4.594872,4.535795,4.4110775,4.1485133,3.767795,3.370667,3.0884104,2.9538465,3.0424619,3.2886157,3.4592824,4.0303593,4.7491283,5.4449234,5.917539,5.943795,6.1997952,6.994052,7.7390776,8.3134365,9.058462,9.334154,9.603283,9.842873,10.276103,11.35918,11.047385,11.592206,12.934566,14.818462,16.768002,17.851078,16.072206,13.99795,12.895181,12.750771,12.737642,13.978257,15.428925,16.275694,15.940925,17.168411,16.840206,16.04595,15.514257,15.609437,17.851078,17.70995,17.539284,17.946259,17.801847,18.514053,18.773335,18.395899,17.522873,16.626873,15.195899,14.86113,14.844719,14.838155,14.976001,15.95077,16.114874,15.75713,15.209026,14.857847,14.87754,14.55918,13.751796,12.983796,13.472821,14.805334,15.91795,16.449642,16.617027,17.211079,18.67159,18.464823,17.792002,17.588514,18.5239,19.505232,19.43631,19.042463,19.18031,20.834463,20.663797,20.09272,20.217438,20.949335,21.008411,17.860924,16.370872,15.136822,13.699283,12.547283,11.516719,10.33518,9.5835905,9.521232,10.075898,10.144821,10.436924,10.043077,9.068309,8.625232,9.091283,9.7903595,10.006975,9.452309,8.257642,7.1122055,6.619898,6.265436,5.9602056,6.0356927,6.3376417,7.962257,9.409642,9.984001,9.777231,7.276308,6.048821,5.8847184,6.0619493,5.330052,4.5456414,2.8258464,1.7788719,1.6508719,1.3653334,2.8947694,3.2262566,2.4746668,1.2865642,0.8467693,3.9089234,9.337437,11.746463,10.932513,11.890873,9.603283,6.124308,4.420923,4.0992823,1.394872,1.8281027,2.6354873,4.4438977,6.242462,5.3760004,3.9286156,3.1671798,4.3749747,6.629744,6.8299494,2.4943593,2.4024618,4.5390773,6.810257,7.0432825,6.892308,7.1614366,8.441437,10.345026,11.506873,12.304411,10.06277,9.488411,10.70277,9.242257,6.2490263,6.294975,7.059693,7.4699492,7.702975,6.629744,5.35959,3.8564105,2.4024618,1.5786668,1.1224617,1.1126155,0.9747693,0.84348726,1.5392822,1.7952822,2.1989746,3.5872824,4.3027697,0.2100513,0.38400003,1.8806155,5.9602056,10.79795,11.464206,8.917334,3.9384618,2.2744617,3.892513,2.993231,0.94523084,1.4473847,1.8740515,1.9462565,3.7218463,3.4789746,3.0162053,2.8914874,3.1540515,3.370667,3.6660516,2.349949,1.4080001,1.3653334,1.2800001,2.3696413,2.8356924,3.373949,4.069744,4.4110775,5.9569235,6.6527185,7.3682055,8.231385,8.615385,9.3078985,9.586872,10.010257,10.522257,10.463181,9.3768215,9.061745,8.887795,8.756514,9.107693,8.362667,8.182155,8.385642,8.63836,8.448001,8.356103,7.7456417,7.351795,7.240206,6.813539,6.8529234,7.433847,8.4283085,9.537642,10.266257,9.91836,9.557334,9.672206,9.980719,9.393231,9.38995,9.409642,8.946873,7.837539,6.23918,5.0215387,4.056616,3.9286156,4.585026,5.353026,4.522667,4.493129,4.4800005,4.3552823,4.647385,4.6145644,4.6572313,4.4865646,4.128821,3.9023592,3.6791797,3.5544617,3.7284105,4.2305646,4.9132314,4.4045134,4.1550775,4.020513,3.948308,4.0008206,3.8564105,3.6135387,3.5774362,3.748103,3.8104618,3.69559,3.629949,3.5446157,3.2787695,2.5895386,2.172718,2.0906668,1.9167181,1.6640002,1.8051283,1.9856411,1.9167181,1.8773335,1.8970258,1.7526156,1.9593848,2.4418464,2.7634873,2.8816411,3.1343591,3.495385,3.5446157,3.5872824,3.6496413,3.495385,4.388103,4.5095387,4.4865646,4.827898,5.930667,5.789539,5.914257,6.0160003,6.166975,6.810257,6.9809237,7.02359,7.138462,7.0400004,5.937231,6.436103,6.882462,7.453539,7.9950776,8.008205,7.3550773,7.9917955,7.821129,6.6002054,5.924103,4.588308,4.522667,4.7589746,6.738052,14.322873,21.50072,15.274668,7.3386674,3.895795,5.654975,4.0369234,3.5052311,4.5390773,5.622154,3.255795,4.775385,6.957949,7.427283,5.9930263,4.6178465,5.7731285,6.373744,7.9294367,10.374565,12.071385,11.930258,12.491488,12.225642,10.893129,9.55077,9.284924,4.453744,1.3292309,1.4769232,1.7624617,2.0742567,1.8149745,3.0916924,5.034667,3.820308,5.874872,4.568616,3.629949,4.2174363,4.9362054,4.1517954,3.4789746,3.0884104,2.9965131,3.0654361,3.4921029,2.733949,2.1792822,2.3105643,2.7109745,2.9407182,2.9833848,2.8849232,2.5895386,1.9396925,1.847795,1.6311796,1.5491283,1.6705642,1.8642052,1.8674873,2.3926156,2.7569232,2.7241027,2.4910772,2.225231,2.0217438,1.7460514,1.4539489,1.4080001,1.4539489,1.5064616,1.7394873,2.0184617,1.8937438,1.7033848,1.6771283,1.595077,1.5425643,1.9035898,1.7427694,2.0250258,2.4320002,2.7273848,2.7667694,2.7667694,2.4681027,2.1136413,1.7985642,1.4736412,1.9200002,2.6223593,2.9604106,2.8127182,2.546872,2.2646155,2.1333334,1.9495386,1.6475899,1.3226668,1.5031796,1.8051283,2.0151796,2.300718,3.2196925,4.778667,5.0642056,4.5456414,3.6791797,2.9046156,3.2951798,3.1048207,2.986667,3.1934361,3.5478978,3.9614363,4.1091285,4.201026,4.20759,3.882667,4.0303593,3.9351797,3.6594875,3.2787695,2.858667,2.9801028,2.9538465,2.9768207,3.0949745,3.190154,3.620103,4.1813335,4.4701543,4.4865646,4.601436,4.588308,4.4701543,4.2994876,4.07959,3.7284105,3.495385,3.7054362,4.1682053,4.535795,4.2929235,3.9712822,4.2141542,4.70318,5.1856413,5.4875903,5.3103595,4.9132314,4.535795,4.378257,4.594872,4.4012313,4.6900516,5.3136415,5.927385,5.9963083,5.2381544,4.7360005,4.525949,4.44718,4.1222568,5.5171285,6.380308,6.62318,6.3277955,5.76,5.149539,4.768821,4.8705645,5.421949,6.0947695,7.2960005,7.8080006,8.477539,9.435898,10.095591,8.746667,7.958975,7.466667,7.00718,6.304821,7.0498466,8.086975,8.940309,9.409642,9.5835905,8.92718,8.507077,8.303591,8.3823595,8.910769,8.79918,8.937026,9.245539,9.531077,9.498257,9.403078,9.380103,9.662359,10.20718,10.673231,9.622975,9.245539,8.976411,8.425026,7.3714876,7.906462,7.9130263,7.6077952,7.3649235,7.709539,7.525744,7.4207187,7.755488,8.480822,9.137232,8.979693,8.763078,8.651488,8.684308,8.776206,8.2904625,7.79159,7.683283,7.939283,8.086975,8.162462,8.14277,8.546462,9.147078,8.969847,2.7766156,3.2361028,3.9023592,4.201026,4.082872,4.0303593,4.266667,3.9318976,3.7251284,3.879385,4.1583595,5.024821,5.6352825,5.9963083,6.045539,5.668103,5.72718,6.416411,7.1614366,7.381334,6.5017443,7.2237954,7.328821,7.194257,6.954667,6.5083084,6.3474874,6.2687182,6.183385,5.917539,5.21518,4.8771286,4.6966157,4.565334,4.378257,4.0402055,4.4701543,4.857436,5.4908724,6.3901544,7.3091288,7.1614366,6.6067696,6.3474874,6.4689236,6.432821,6.5247183,6.5837955,6.3901544,6.2523084,7.020308,6.76759,6.6034875,6.491898,6.409847,6.3540516,6.3310776,6.9054365,6.954667,6.245744,5.431795,4.84759,5.0215387,5.0838976,4.890257,5.0051284,4.7524104,4.8804107,4.821334,4.6080003,4.8640003,5.044513,5.4974365,6.157129,6.931693,7.6898465,8.109949,8.425026,9.074872,10.35159,12.373334,13.430155,13.715693,13.90277,14.122667,13.965129,13.361232,12.708103,12.005745,11.523283,11.808822,11.88759,11.59877,11.030975,10.361437,9.83959,9.8363085,9.829744,9.810052,9.780514,9.734565,10.04636,9.32759,8.231385,7.1647186,6.2884107,6.0028725,5.648411,5.4383593,5.3431797,5.0543594,4.6769233,4.4701543,4.1780515,3.7448208,3.3247182,3.1540515,3.2918978,3.4658465,3.5249233,3.442872,3.255795,3.0916924,2.9111798,2.7208207,2.5796926,2.3729234,2.3433847,2.3696413,2.3893335,2.4024618,3.2196925,3.6627696,4.20759,4.857436,5.1331286,5.169231,5.3924108,6.0980515,7.13518,7.896616,8.349539,8.884514,9.38995,9.911796,10.650257,10.794667,11.736616,12.662155,13.482668,14.8480015,15.796514,15.471591,14.368821,13.164309,12.721231,12.471796,13.161027,14.332719,16.02954,18.786463,20.256823,19.324718,17.637745,16.288822,15.799796,18.070976,17.78872,17.34236,17.490053,17.375181,17.211079,16.305231,15.776822,15.931078,16.272411,15.589745,15.461744,15.002257,14.313026,14.49354,15.701335,16.469334,16.377438,15.652103,15.1466675,14.552616,14.41477,13.912617,13.223386,13.499078,15.090873,15.8884115,15.960617,15.799796,16.295385,18.20554,19.03918,19.334566,19.56759,20.171488,21.090464,21.605745,21.513847,21.300514,22.14072,22.12431,20.197744,18.468103,17.913437,18.372925,17.289848,17.864206,16.692514,13.607386,11.697231,10.637129,10.282667,10.174359,10.246565,10.834052,11.136001,11.122872,10.630565,9.6984625,8.569437,8.635077,9.065026,9.396514,9.357129,8.881231,7.529026,7.200821,7.030154,6.695385,6.413129,6.196513,7.394462,8.79918,9.701744,9.911796,7.955693,6.5280004,6.166975,6.298257,5.2512827,4.562052,3.626667,2.8553848,2.5042052,2.665026,3.95159,3.1048207,2.6584618,3.1934361,3.3214362,7.315693,10.8996935,11.241027,9.048616,8.576,6.0356927,2.806154,1.4572309,1.8937438,1.3587693,1.2077949,1.401436,2.2547693,3.1967182,2.7700515,2.034872,2.0644104,2.2613335,2.0644104,0.93866676,1.148718,3.121231,5.8486156,8.113232,8.4972315,6.9087186,7.0957956,8.5202055,10.282667,11.113027,11.874462,10.633847,9.728001,9.708308,9.347282,7.00718,6.619898,6.518154,6.51159,7.893334,6.672411,5.0576415,3.495385,2.2744617,1.522872,0.98461545,0.86974365,0.764718,0.6301539,0.78769237,1.9593848,1.8051283,3.5544617,5.362872,0.29538465,0.22646156,1.0732309,4.332308,9.202872,12.58995,12.1698475,7.2172313,4.6834874,5.4482055,4.325744,1.4736412,1.6443079,1.8806155,1.782154,3.5216413,4.604718,3.0687182,1.9790771,2.8324106,5.543385,3.3542566,2.2744617,1.7558975,1.719795,2.546872,3.3969233,3.7185643,4.069744,4.768821,5.8978467,6.9152827,7.062975,7.6274877,8.621949,8.786052,9.524513,9.137232,9.403078,10.518975,11.099898,10.502565,9.990565,9.353847,8.835282,9.124104,8.155898,7.9819493,8.392206,8.904206,8.759795,8.119796,7.27959,6.99077,7.145026,6.741334,7.1122055,7.8145647,8.756514,9.6984625,10.243283,9.613129,9.337437,9.547488,9.921641,9.685334,9.458873,9.068309,8.533334,7.6307697,5.917539,5.100308,4.4898467,4.6211286,5.3103595,5.6451287,4.5128207,4.601436,4.6112823,4.3585644,4.7950773,4.453744,4.345436,4.2141542,4.0402055,4.0434875,3.8629746,3.8137438,4.0008206,4.466872,5.182359,4.2863593,4.0041027,3.8334363,3.7218463,4.056616,3.7120004,3.5282054,3.639795,3.8400004,3.5905645,3.7284105,3.6430771,3.4592824,3.1934361,2.740513,2.2416413,2.3204105,2.1497438,1.7263591,1.8674873,1.7526156,1.8904617,1.8937438,1.8346668,2.2219489,2.3072822,2.4484105,2.553436,2.605949,2.6453335,3.2262566,3.1934361,3.1376412,3.2853336,3.4822567,3.8301542,3.948308,3.9187696,4.07959,5.037949,5.5138464,6.0750775,6.3343596,6.416411,6.957949,7.056411,6.6592827,6.6067696,6.9152827,6.806975,6.987488,7.0957956,6.8594875,7.4929237,11.700514,11.894155,10.935796,9.609847,8.749949,9.235693,4.670359,5.159385,6.055385,7.3058467,13.456411,14.555899,11.408411,8.01477,5.6451287,2.8521028,2.2514873,2.5107694,3.7218463,4.84759,3.757949,2.9013336,4.4340515,5.3760004,4.9427695,4.5489235,4.4964104,5.674667,7.9524107,10.44677,11.52,9.229129,11.772718,14.519796,14.933334,12.544001,13.843694,6.4000006,1.2964103,1.401436,1.3357949,1.719795,1.5885129,1.8182565,2.540308,3.1113849,6.0061545,4.4110775,2.9243078,3.186872,3.8662567,3.6594875,3.0326157,2.737231,2.8717952,2.8816411,3.1081028,2.733949,2.3466668,2.2482052,2.4484105,2.4943593,2.5140514,2.3926156,2.0906668,1.6738462,1.4966155,1.2504616,1.214359,1.4309745,1.7165129,1.7296412,2.1070771,2.3893335,2.4320002,2.412308,2.15959,2.3040001,2.28759,2.0217438,1.913436,1.9659488,1.8904617,1.9593848,2.0808206,1.8149745,1.9462565,2.100513,1.9659488,1.7723079,2.2711797,2.281026,2.5107694,2.793026,3.0326157,3.1967182,3.495385,3.0851285,2.4976413,2.0151796,1.657436,1.9364104,2.6026669,2.8717952,2.6683078,2.6157951,2.356513,2.1891284,2.0053334,1.7788719,1.5425643,1.6672822,1.8313848,2.0184617,2.2613335,2.6289232,4.092718,4.578462,4.1714873,3.2787695,2.6354873,2.8455386,2.930872,3.0982566,3.3280003,3.4034874,3.761231,4.06318,4.1189747,3.8859491,3.4494362,3.7940516,3.8990772,3.7776413,3.5478978,3.446154,3.4330258,3.2853336,3.1967182,3.2361028,3.3411283,3.5446157,3.9844105,4.4274874,4.7261543,4.7917953,4.7261543,4.6933336,4.4012313,3.9318976,3.754667,3.6036925,4.013949,4.397949,4.4110775,3.945026,4.013949,4.069744,4.4012313,4.9854364,5.474462,5.221744,5.031385,4.667077,4.1156926,3.626667,4.2601027,4.5554876,4.713026,4.9920006,5.7107697,5.2644105,4.9526157,4.6769233,4.3716927,4.020513,5.0871797,5.865026,6.4065647,6.665847,6.491898,5.366154,4.9132314,5.0576415,5.540103,5.930667,7.2631803,8.333129,8.986258,9.31118,9.613129,8.881231,8.267488,7.8637953,7.6307697,7.397744,7.653744,8.283898,8.825437,8.960001,8.513641,8.001641,8.034462,8.129642,8.2215395,8.661334,8.352821,8.231385,8.310155,8.43159,8.2445135,8.5202055,8.818872,9.225847,9.69518,10.069334,9.271795,8.704,8.352821,7.962257,7.0367184,7.273026,6.7840004,6.2851286,6.157129,6.452513,6.0291286,5.61559,5.868308,6.705231,7.325539,7.0793853,7.0826674,7.394462,7.827693,7.958975,7.857231,7.5881033,7.3353853,7.1515903,6.921847,7.27959,7.643898,8.323282,9.120821,9.340718,3.889231,4.069744,4.332308,4.266667,3.9220517,3.820308,3.892513,3.9023592,4.07959,4.378257,4.466872,5.8486156,6.2096415,6.3245134,6.2227697,5.172513,5.3792825,6.2588725,7.318975,7.834257,6.8463597,7.3025646,7.3058467,7.02359,6.6822567,6.560821,6.340924,6.1013336,5.737026,5.5007186,5.986462,5.6320004,5.106872,4.775385,4.6244106,4.2535386,4.3651285,4.7917953,5.4908724,6.426257,7.571693,7.3353853,7.00718,6.5739493,6.12759,5.8847184,6.4754877,6.1505647,5.83877,6.0160003,6.7117953,7.1187696,6.6822567,6.3901544,6.51159,6.6002054,6.8496413,7.6635904,7.939283,7.3682055,6.432821,5.3037953,5.0510774,4.844308,4.535795,4.6605134,5.287385,5.5663595,5.3924108,4.955898,4.7524104,5.2480006,5.425231,5.943795,7.0859494,8.763078,10.069334,10.174359,10.256411,10.870154,11.949949,13.525334,14.628103,15.067899,14.989129,14.874257,14.358975,13.61395,12.370052,11.113027,11.113027,11.37559,11.073642,10.607591,10.249847,10.121847,10.148104,10.197334,9.846154,9.373539,9.77395,9.609847,8.5661545,7.2861543,6.2194877,5.602462,5.1298466,4.916513,4.916513,4.972308,4.8016415,4.2896414,3.876103,3.4133337,2.9111798,2.5271797,2.4451284,2.3893335,2.2711797,2.1464617,2.231795,1.9495386,1.9003079,1.9331284,1.975795,2.034872,1.719795,1.6705642,1.5392822,1.3259488,1.3620514,2.2055387,2.7011285,3.0030773,3.4330258,4.4832826,4.6276927,4.7589746,5.504,6.5870776,6.816821,7.1187696,7.765334,8.562873,9.147078,8.986258,10.226872,11.664412,12.304411,12.202667,12.498053,12.402873,13.069129,13.778052,14.017642,13.472821,12.658873,13.177437,13.988104,15.698052,20.54236,22.317951,20.854155,18.500925,16.754873,16.262566,17.355488,17.135592,16.850052,17.024002,17.460514,16.600616,14.818462,14.148924,15.067899,16.482462,16.538258,16.777847,16.170668,15.087591,15.31077,16.026258,16.617027,16.571077,16.042667,15.868719,14.867694,15.05477,15.0777445,14.611693,14.345847,15.714462,16.121437,15.671796,15.048206,15.514257,18.097233,20.263386,21.940514,22.774155,22.111181,22.839796,24.086977,24.04431,23.08595,23.785027,23.364925,20.841026,19.403488,19.163898,17.161848,16.646564,19.337847,18.884924,14.614976,11.539693,9.563898,9.898667,10.47959,10.774975,11.795693,12.452104,12.1698475,11.45436,10.433641,8.845129,8.779488,8.979693,9.291488,9.475283,9.216001,7.955693,7.9261546,7.9491286,7.6209235,7.328821,6.8693337,7.2172313,8.178872,9.330873,10.013539,8.730257,7.315693,6.8233852,6.7314878,4.9362054,4.210872,4.4077954,4.325744,4.020513,4.8049235,4.4340515,2.986667,3.6463592,6.449231,8.277334,11.021129,9.944616,9.061745,8.608821,5.044513,3.1048207,1.8904617,2.2219489,3.062154,1.5031796,1.6213335,1.4900514,1.1881026,0.82379496,0.5415385,0.7089231,0.7089231,0.58420515,0.6301539,1.401436,2.2383592,3.9876926,6.413129,8.615385,9.025641,7.3583593,7.565129,8.618668,9.590155,9.632821,10.072617,9.974154,9.3078985,8.55959,8.723693,7.968821,7.0859494,6.2063594,6.0225644,7.79159,6.3179493,4.6112823,3.045744,1.8806155,1.2471796,0.636718,0.4397949,0.6498462,1.0338463,1.1158975,2.0020514,2.2580514,5.228308,8.0377445,1.5983591,0.46276927,1.1618463,1.9331284,3.3345644,8.264206,14.532925,12.3536415,10.197334,9.540924,4.850872,2.1530259,1.847795,1.6508719,1.2931283,2.5173335,7.1581545,5.3366156,3.2131286,3.761231,6.76759,2.7831798,2.422154,2.5173335,2.5107694,4.4438977,4.571898,4.8147697,5.3431797,6.245744,7.5191803,7.3682055,7.171283,7.8703594,9.130668,9.340718,10.026668,9.051898,8.612103,9.4916935,11.063796,11.296822,10.9226675,10.043077,9.16677,9.193027,8.1066675,7.8834877,8.205129,8.562873,8.300308,8.086975,7.683283,7.322257,7.1614366,7.269744,8.024616,8.576,9.160206,9.816616,10.404103,9.731283,9.649232,9.711591,9.701744,9.642668,9.051898,8.001641,7.1876926,6.521436,5.169231,5.1298466,5.1659493,5.5105643,5.8420515,5.3070774,4.4800005,4.493129,4.535795,4.417641,4.585026,4.279795,4.325744,4.138667,3.8596926,4.325744,4.2371287,4.322462,4.332308,4.3552823,4.8344617,4.391385,4.2305646,3.9154875,3.5872824,3.9581542,3.764513,3.7710772,3.8728209,3.876103,3.508513,3.7185643,3.7120004,3.508513,3.239385,3.1540515,2.7076926,2.802872,2.5993848,2.0742567,2.0118976,1.6377437,1.910154,1.9889232,1.8904617,2.487795,2.681436,2.5173335,2.359795,2.3236926,2.284308,3.114667,2.8521028,2.674872,3.0720003,3.8662567,3.3575387,3.367385,3.6430771,4.076308,4.6769233,5.1265645,5.943795,6.6034875,6.8430777,6.672411,6.8955903,6.5247183,6.183385,6.3901544,7.5552826,8.080411,7.6964107,6.2687182,5.98318,11.332924,13.266052,10.883283,9.842873,11.533129,13.088821,6.5050263,6.994052,7.6996927,7.276308,9.905231,8.257642,8.100103,9.517949,9.724719,3.0752823,3.5413337,3.1343591,3.239385,3.9712822,4.1813335,3.6529233,5.034667,5.8420515,4.8804107,2.2449234,1.9856411,4.1025643,7.3091288,10.098872,10.752001,5.979898,10.049642,15.222155,16.30195,10.627283,12.104206,5.8814363,1.4441026,1.2996924,0.9682052,1.4276924,1.4736412,1.5655385,2.1464617,3.6463592,3.1245131,2.2547693,1.8806155,2.2383592,2.9735386,3.0982566,2.6683078,2.537026,2.8160002,2.8914874,3.186872,3.1113849,2.7864618,2.3991797,2.1989746,2.100513,2.0676925,2.034872,1.9823592,1.9364104,1.394872,1.0929232,1.1684103,1.5097437,1.7657437,1.975795,1.9626669,1.9462565,2.0512822,2.294154,2.3302567,2.809436,2.9801028,2.7175386,2.5206156,2.612513,2.3401027,2.1234872,2.03159,1.7690258,2.2646155,2.3696413,2.2153847,2.1234872,2.5961027,2.9111798,3.0391798,2.8947694,2.6978464,2.9833848,3.4494362,3.1442053,2.6157951,2.2186668,2.0873847,2.3433847,2.674872,2.8324106,2.8488207,3.0358977,2.7470772,2.1464617,1.8051283,1.847795,1.9495386,1.8510771,1.9364104,2.0709746,2.1070771,1.8773335,2.9505644,3.5282054,3.31159,2.5206156,1.8707694,1.7657437,2.2678976,2.9144619,3.3378465,3.2886157,3.3247182,3.4691284,3.4494362,3.2918978,3.3247182,3.5216413,3.7842054,3.8301542,3.7316926,3.9089234,3.876103,3.8038976,3.5872824,3.3542566,3.4494362,3.826872,4.1714873,4.598154,4.9788723,4.969026,4.788513,4.673641,4.3749747,3.9778464,3.892513,4.1124105,4.900103,5.412103,5.2414365,4.4274874,4.6769233,3.9876926,3.6529233,4.0303593,4.519385,4.906667,4.969026,4.640821,3.9876926,3.1967182,4.601436,5.221744,4.9132314,4.3651285,5.100308,4.900103,5.07077,5.0838976,4.7294364,4.1091285,4.1878977,5.0215387,6.173539,7.0334363,6.813539,5.6451287,5.293949,5.412103,5.684513,5.805949,6.9021544,7.9425645,8.635077,8.917334,8.966565,8.753231,8.549745,8.323282,8.169026,8.283898,8.14277,8.4283085,8.461129,7.958975,7.0367184,6.7282057,7.059693,7.571693,7.975385,8.182155,8.300308,8.211693,8.073847,7.8769236,7.4108725,7.8473854,8.093539,8.717129,9.494975,9.416205,8.369231,7.778462,7.4830775,7.1909747,6.482052,6.449231,5.927385,5.435077,5.3727183,6.0356927,5.914257,4.8344617,4.4012313,4.886975,5.2480006,5.5236926,5.8092313,6.3179493,6.8463597,6.806975,7.5881033,7.6898465,7.318975,6.685539,6.0061545,6.373744,7.1122055,7.8834877,8.457847,8.723693,3.570872,4.4242053,5.225026,4.841026,3.7349746,3.9680004,3.4560003,3.748103,4.394667,5.10359,5.737026,6.675693,7.177847,7.177847,6.7840004,6.2720003,6.4295387,6.9743595,7.460103,7.578257,7.125334,6.626462,6.6100516,6.2063594,5.536821,5.7074876,5.7796926,5.7435904,5.6385646,5.609026,5.8912826,5.681231,5.152821,4.6966157,4.594872,5.034667,4.5095387,5.0576415,5.9667697,6.7544622,7.1548724,6.803693,6.2555904,6.157129,6.3606157,5.920821,6.298257,5.7435904,5.720616,6.4557953,6.941539,7.322257,7.325539,7.056411,6.9054365,7.5520005,7.9195905,7.9917955,8.152616,8.228104,7.506052,6.1538467,5.7501545,5.622154,5.4153852,5.110154,5.5138464,5.677949,5.6352825,5.47118,5.32677,5.5565133,5.549949,5.8978467,6.806975,8.103385,9.554052,10.240001,10.9456415,11.9860525,13.184001,15.199181,16.534975,17.11918,16.938667,16.022976,14.276924,13.252924,12.855796,12.849232,12.849232,13.275898,13.262771,12.360206,11.063796,10.817642,10.453334,11.211488,11.382154,10.761847,10.666668,9.750975,8.487385,7.125334,6.0291286,5.674667,4.772103,4.2896414,4.1025643,4.0303593,3.8596926,3.5544617,3.1409233,2.6157951,1.9889232,1.2832822,1.1093334,1.1224617,1.2406155,1.339077,1.2668719,1.4244103,1.4998976,1.5392822,1.5097437,1.3259488,1.204513,1.2209232,1.014154,0.6892308,0.82379496,1.1913847,1.6475899,2.2777438,3.0916924,4.0434875,4.6178465,4.9788723,5.536821,6.232616,6.560821,6.8430777,6.9120007,7.0957956,7.53559,8.195283,9.511385,9.7673855,10.049642,10.630565,10.971898,10.604308,11.273847,12.672001,13.889642,13.413745,13.059283,14.188309,14.87754,15.232001,17.378464,18.441847,18.881643,18.028309,16.544823,16.433231,16.764719,17.42113,18.025026,18.326975,18.202257,16.994463,15.254975,13.984821,13.797745,14.907078,15.724309,16.836924,17.043694,16.200207,15.212309,16.298668,16.295385,15.78995,15.123693,14.404924,14.086565,15.051488,16.17395,16.640001,15.944206,15.993437,16.154257,16.02954,15.66195,15.504412,16.357744,18.776617,21.993027,25.002668,26.564924,24.549746,23.335386,22.600206,22.600206,24.139488,22.918566,21.028105,20.772104,21.362873,18.921026,16.981335,19.058874,19.692308,17.056822,12.954257,10.893129,10.7158985,11.441232,12.22236,12.343796,13.1872835,13.46954,12.780309,11.372309,10.161232,9.990565,9.747693,10.125129,10.535385,9.094564,8.39877,8.342975,8.4283085,8.388924,8.195283,7.4141545,7.00718,7.4207187,8.6580515,10.269539,9.573745,7.9885135,6.994052,6.678975,5.7534366,4.4832826,4.9526157,5.5138464,5.7829747,6.636308,4.7327185,3.1113849,3.8990772,7.6898465,13.548308,14.086565,11.126155,6.885744,3.383795,2.4582565,1.5524104,1.6213335,1.2307693,0.36758977,0.4266667,2.540308,2.297436,2.028308,2.2613335,1.723077,1.785436,1.8838975,1.6738462,1.4244103,1.9987694,3.2065644,4.7622566,6.294975,7.387898,7.584821,8.241231,9.212719,9.800206,9.6065645,8.546462,9.143796,9.8592825,10.092308,9.370257,7.3714876,7.637334,7.834257,7.315693,6.5837955,7.27959,5.533539,4.069744,2.5928206,1.3587693,1.1749744,0.80738467,0.56123084,0.9353847,1.7394873,2.1070771,1.1158975,3.058872,8.477539,12.672001,5.674667,1.2209232,3.117949,3.6693337,2.4910772,6.5312824,11.460924,15.238565,16.472616,13.200411,2.8980515,1.8609232,1.2077949,1.6902566,3.1409233,4.4701543,8.766359,10.656821,9.173334,5.58277,3.373949,2.0644104,2.1333334,2.878359,3.748103,4.332308,4.345436,5.5105643,6.9809237,8.165744,8.726975,8.214975,8.352821,8.720411,9.025641,9.110975,10.000411,9.32759,8.717129,9.097847,10.696206,10.745437,10.456616,9.705027,8.887795,8.910769,8.116513,7.9917955,7.9261546,7.788308,7.936001,8.192,8.218257,8.004924,7.817847,8.208411,8.27077,8.897642,9.563898,10.072617,10.57477,10.148104,9.373539,8.677744,8.300308,8.300308,8.116513,7.6767187,6.987488,6.157129,5.402257,4.414359,4.3749747,4.6276927,4.8082056,4.8672824,4.7327185,4.562052,4.57518,4.585026,3.9975388,4.1452312,4.1156926,3.9286156,3.8006158,4.164923,4.2141542,4.3651285,4.210872,4.027077,4.7622566,4.5522056,4.2830772,3.8531284,3.370667,3.1277952,3.4822567,3.6627696,3.748103,3.6562054,3.1442053,2.9735386,2.7831798,2.7109745,2.6551797,2.28759,2.9833848,2.8291285,2.2055387,1.6082052,1.6311796,1.5721027,1.7296412,1.8084104,1.7920002,1.9364104,2.425436,2.3204105,2.284308,2.3827693,2.0906668,2.7634873,2.930872,3.2820516,3.817026,3.8301542,3.5380516,3.9220517,4.4045134,4.8738465,5.691077,5.7403083,5.799385,6.1407185,6.5739493,6.439385,5.8518977,6.6133337,7.026872,6.6034875,6.042257,6.0685134,6.4295387,7.0400004,7.0104623,4.6539493,8.218257,9.465437,10.8767185,11.54954,7.2172313,10.525539,10.171078,7.003898,5.792821,15.228719,15.484719,12.3536415,12.645744,13.965129,4.699898,6.5312824,5.2676926,3.9614363,3.764513,3.9351797,4.132103,5.0510774,4.397949,2.4910772,2.2580514,1.4900514,1.7362052,3.4166157,5.8945646,7.4929237,7.076103,9.810052,10.476309,7.90318,4.97559,4.5489235,2.7208207,1.339077,1.0272821,1.1749744,1.467077,1.5688206,1.7591796,2.1825643,2.8521028,2.2908719,1.8313848,1.6836925,1.9954873,2.8389745,2.8389745,2.8750772,2.9669745,3.1376412,3.4166157,3.5774362,3.1113849,2.6847181,2.5665643,2.6387694,2.041436,2.038154,2.1924105,2.2055387,1.9364104,1.5589745,1.3456411,1.4736412,1.7558975,1.6311796,2.3401027,2.0775387,1.975795,2.3926156,2.930872,2.477949,3.062154,3.18359,2.678154,2.7175386,2.4484105,2.2514873,1.9298463,1.6475899,1.9528207,2.2219489,2.15959,2.3991797,2.8914874,2.9144619,3.367385,3.6529233,3.8465643,3.9253337,3.754667,3.1540515,2.4582565,2.0217438,1.9396925,2.0151796,2.4155898,2.930872,3.2787695,3.5380516,4.135385,4.2568207,3.2820516,2.5009232,2.4024618,2.6715899,2.1825643,2.1956925,2.1103592,1.7788719,1.5097437,2.1956925,2.5862565,2.5107694,2.1136413,1.847795,1.5655385,1.8346668,2.4188719,2.8980515,2.6551797,2.8258464,3.1540515,3.249231,3.1638978,3.370667,3.629949,3.8400004,3.754667,3.5183592,3.6758976,3.8498464,3.9745643,3.7776413,3.387077,3.3280003,4.2896414,4.8705645,5.0674877,5.225026,6.042257,5.723898,5.225026,4.7622566,4.3716927,3.9056413,3.7349746,4.571898,5.4613338,5.76,5.110154,4.647385,3.626667,3.2525132,3.7382567,4.2863593,5.3858466,4.8738465,4.164923,3.6758976,2.806154,3.7710772,5.139693,5.0609236,3.892513,4.197744,4.562052,5.139693,5.4580517,5.172513,4.073026,3.5249233,4.201026,4.9887185,5.4974365,6.058667,5.973334,5.540103,5.3366156,5.5007186,5.7074876,6.36718,6.8430777,7.5881033,8.392206,8.392206,8.648206,8.576,8.185436,7.8080006,8.103385,8.113232,8.080411,7.7325134,6.9382567,5.7074876,6.36718,6.8496413,7.0531287,7.145026,7.584821,8.474257,8.605539,8.2215395,7.7259493,7.6898465,7.7259493,7.581539,7.9819493,8.674462,8.392206,7.1483083,7.066257,7.131898,6.764308,5.799385,5.677949,5.618872,5.152821,4.5587697,4.850872,5.4613338,4.8738465,4.2141542,4.138667,4.821334,5.408821,5.5171285,5.4613338,5.4383593,5.5236926,5.5236926,5.723898,5.970052,5.970052,5.3103595,5.677949,6.482052,7.1122055,7.3583593,7.430565,3.9844105,4.089436,4.6572313,4.529231,3.892513,4.2601027,3.8465643,4.4340515,5.4843082,6.6527185,7.77518,8.188719,8.103385,7.6964107,7.24677,7.125334,7.2172313,7.2894363,7.3091288,7.384616,7.7718983,7.1844106,6.5312824,5.654975,5.031385,5.7796926,5.920821,6.114462,6.0947695,5.8814363,5.7796926,6.1013336,6.055385,5.733744,5.349744,5.2414365,5.3431797,5.4875903,6.0258465,6.6034875,6.166975,6.2227697,6.3212314,6.416411,6.4623594,6.432821,6.665847,6.058667,5.730462,5.933949,6.052103,6.8693337,7.1220517,7.174565,7.397744,8.152616,8.303591,8.1755905,7.9885135,7.7948723,7.496206,6.9021544,6.6592827,6.5706673,6.521436,6.47877,6.5870776,6.5050263,6.3310776,6.012718,5.349744,5.2676926,5.398975,6.117744,7.7292314,10.456616,11.07036,12.1238985,12.793437,13.131488,14.073437,14.683899,16.07877,17.083078,17.362053,17.414566,15.570052,14.309745,14.247386,14.762668,14.020925,14.457437,14.073437,13.371078,12.773745,12.635899,11.900719,11.936821,11.385437,10.085744,9.078155,7.8703594,7.0531287,6.121026,4.969026,3.882667,3.446154,3.4560003,3.3247182,2.9144619,2.5173335,2.2022567,1.8379488,1.5261539,1.2504616,0.8533334,0.88943595,0.9288206,1.0502565,1.1749744,1.0699488,1.1913847,1.273436,1.3587693,1.3554872,1.0338463,0.9419488,0.90584624,0.7417436,0.512,0.51856416,0.80738467,1.2898463,1.9232821,2.7634873,3.9712822,4.71959,5.221744,5.661539,6.0160003,6.0717955,6.235898,6.5706673,6.885744,7.243488,7.9491286,8.280616,8.700719,9.110975,9.5146675,10.029949,10.545232,11.067078,12.081232,13.423591,14.267078,14.322873,14.742975,14.201437,13.387488,14.998976,16.55795,17.80513,17.723078,16.571077,15.885129,17.201233,18.011898,18.04472,17.23077,15.714462,15.42236,14.454155,13.643488,13.571283,14.565744,15.481437,16.469334,17.483488,17.877335,16.410257,16.695797,16.213335,15.117129,13.991385,13.866668,13.433437,14.007796,15.156514,16.256,16.505438,16.869745,16.672821,16.262566,16.114874,16.833643,18.067694,19.528206,21.241438,23.023592,24.477541,25.238976,24.49395,23.72595,23.532309,23.61436,22.170258,21.169233,21.395695,22.025848,20.630976,18.202257,18.06113,18.592821,18.051283,14.552616,11.798975,11.175385,11.828514,13.092104,14.49354,14.592001,14.260514,13.653335,12.849232,11.835078,10.873437,10.417232,10.584617,10.778257,9.67877,8.349539,8.362667,8.503796,8.277334,7.9261546,7.719385,7.318975,7.427283,8.234667,9.416205,9.314463,8.018052,6.8627696,6.4689236,6.7544622,5.3760004,5.35959,5.933949,6.7117953,7.6767187,5.225026,3.7382567,3.3936412,4.466872,7.3485136,6.2063594,4.4242053,3.3345644,2.9833848,2.1136413,2.1202054,2.166154,2.1366155,2.3466668,3.5413337,3.8465643,2.6551797,1.654154,1.4441026,1.5425643,1.5130258,1.7657437,1.9593848,2.1530259,2.802872,3.6726158,4.8771286,6.2096415,7.0432825,6.3507695,7.890052,8.5891285,9.478565,10.128411,8.667898,8.553026,8.89436,9.212719,9.02236,7.821129,7.837539,8.208411,7.7292314,6.5444107,6.1538467,4.644103,3.3805132,2.1431797,1.1881026,1.2471796,0.8041026,0.6826667,0.8763078,1.3095386,1.8609232,2.0151796,1.9429746,3.623385,5.421949,2.100513,1.7362052,3.4789746,4.841026,5.1889234,5.723898,12.599796,15.596309,11.447796,4.0467696,4.4373336,1.7887181,1.785436,2.7142565,4.0434875,6.449231,8.411898,7.1844106,4.7524104,3.387077,5.6287184,3.5314875,3.4527183,4.1780515,4.893539,5.175795,5.3727183,6.695385,8.083693,8.812308,8.4972315,8.792616,8.986258,9.02236,8.996103,9.170052,8.900924,8.477539,8.608821,9.321027,9.95118,10.138257,9.882257,9.449026,9.078155,8.982975,8.592411,8.2445135,7.972103,7.8736415,8.116513,7.9261546,8.096821,8.356103,8.569437,8.746667,9.051898,9.229129,9.478565,9.764103,9.80677,9.622975,9.3768215,9.009232,8.493949,7.8506675,7.460103,6.925129,6.2818465,5.7074876,5.536821,5.3005133,5.208616,5.0674877,4.7950773,4.414359,3.8531284,3.8432825,4.1189747,4.2174363,3.4855387,3.564308,3.4592824,3.4264617,3.6496413,4.240411,4.201026,4.0402055,3.7316926,3.5413337,4.0402055,3.9220517,3.6332312,3.2853336,3.058872,3.2262566,3.4231799,3.5216413,3.5183592,3.4133337,3.2032824,3.442872,3.3280003,3.1113849,2.865231,2.4582565,2.8422565,2.6912823,2.1267693,1.5753847,1.7657437,1.8707694,2.0578463,1.9954873,1.785436,1.9495386,2.2219489,2.0709746,2.0742567,2.28759,2.2482052,2.8225644,3.3247182,3.8006158,3.9975388,3.3542566,3.1770258,3.6496413,4.07959,4.3618464,4.9952826,4.955898,5.3136415,5.8912826,6.5017443,6.9645133,6.4557953,6.6428723,6.6625648,6.518154,7.0793853,6.918565,6.3868723,6.5017443,7.138462,6.997334,7.4863596,6.806975,6.5083084,6.747898,6.2884107,10.535385,10.033232,8.395488,11.69395,28.471798,21.697643,10.453334,5.1298466,6.088206,3.636513,7.177847,5.681231,4.6211286,5.6320004,6.5378466,6.048821,5.8518977,4.525949,2.7798977,3.4560003,4.7655387,3.3936412,3.56759,6.0980515,8.372514,4.9493337,3.8564105,3.5052311,3.045744,2.3630772,1.6902566,1.1191796,0.88943595,0.98133343,1.1388719,1.2274873,1.4145643,1.5786668,1.7001027,1.8510771,1.6607181,1.3817437,1.4736412,1.975795,2.4976413,2.7602053,2.7733335,2.9538465,3.4166157,3.9778464,3.7874875,2.8553848,2.1792822,2.15959,2.6026669,1.975795,2.169436,2.4549747,2.3926156,1.8412309,1.7066668,1.7657437,1.7755898,1.6213335,1.3029745,2.0118976,2.3696413,2.6683078,2.9243078,2.9046156,3.2065644,3.4034874,3.387077,3.2918978,3.5347695,3.2262566,2.8160002,2.3302567,1.9790771,2.1366155,3.255795,3.2820516,3.767795,4.8640003,5.3202057,5.0477953,4.818052,4.667077,4.532513,4.2535386,4.604718,4.125539,3.0785644,1.9167181,1.3062565,1.7887181,2.8258464,3.4888208,3.6562054,4.0008206,4.2994876,3.9023592,3.2328207,2.6453335,2.425436,2.2416413,2.2514873,2.3466668,2.281026,1.6705642,1.719795,1.8773335,2.0086155,2.0775387,2.1530259,1.9593848,2.0939488,2.4943593,2.8455386,2.5829747,3.006359,3.2787695,3.2065644,2.9538465,3.05559,2.9604106,2.937436,2.793026,2.5993848,2.7011285,3.0096412,3.3214362,3.5282054,3.5544617,3.387077,3.8531284,4.315898,4.571898,4.7327185,5.2381544,4.95918,4.3651285,4.092718,4.1517954,3.9417439,3.692308,4.069744,4.781949,5.349744,5.110154,4.2174363,3.6529233,3.6463592,4.1846156,5.0084105,5.7829747,5.4843082,5.0116925,4.5817437,3.7349746,3.9975388,4.778667,4.6802053,3.7874875,3.6726158,3.8432825,4.4734364,5.077334,5.0838976,3.8301542,3.8662567,4.667077,4.9132314,4.6802053,5.4482055,6.045539,6.121026,5.98318,5.865026,5.927385,6.4000006,6.633026,7.059693,7.584821,7.574975,8.14277,8.083693,7.8736415,7.6931286,7.430565,7.394462,7.5454364,7.197539,6.262154,5.2545643,5.730462,5.8223596,6.196513,6.9087186,7.4240007,8.004924,7.9917955,7.643898,7.315693,7.433847,7.4404106,7.450257,7.5191803,7.568411,7.3682055,6.5805135,5.9963083,5.7731285,5.723898,5.346462,5.3891287,5.2578464,4.7491283,4.0467696,3.7054362,4.3749747,4.128821,3.5774362,3.370667,4.197744,4.667077,4.9099493,4.9526157,4.903385,4.9493337,5.0674877,5.408821,5.7403083,5.901129,5.799385,5.9503593,6.7610264,7.5946674,7.893334,7.174565,3.7152824,4.279795,4.44718,4.2568207,4.017231,4.2962055,4.332308,5.142975,6.2851286,7.4240007,8.329846,8.5891285,8.224821,7.906462,7.762052,7.384616,7.259898,7.384616,7.581539,7.768616,7.972103,7.4699492,6.9120007,6.114462,5.4416413,5.799385,6.0160003,5.861744,5.605744,5.353026,5.0576415,5.077334,5.395693,5.536821,5.5072823,5.789539,5.8256416,5.920821,6.245744,6.5378466,6.0947695,5.9536414,6.088206,6.2063594,6.2162056,6.232616,6.675693,6.2720003,6.1407185,6.2818465,5.58277,6.180103,6.413129,6.5969234,6.951385,7.578257,7.9885135,7.9195905,7.7259493,7.5388722,7.2631803,7.315693,7.4075904,7.522462,7.6767187,7.9195905,7.75877,7.1876926,6.5870776,6.058667,5.4580517,5.421949,6.1538467,7.4699492,9.281642,11.588924,12.225642,12.895181,13.351386,13.676309,14.260514,14.884104,16.46277,17.240616,16.70236,15.573335,14.864411,14.378668,14.198155,14.096412,13.53518,13.702565,13.302155,12.84595,12.465232,11.900719,10.962052,10.916103,10.220308,8.858257,8.342975,7.4436927,6.678975,5.8190775,4.8377438,3.9187696,3.7710772,3.7382567,3.3542566,2.5796926,1.8346668,1.332513,1.0108719,0.84348726,0.73517954,0.5284103,0.78769237,0.8369231,0.88287187,0.9517949,0.892718,0.88615394,0.94523084,0.95835906,0.8795898,0.7220513,0.7318975,0.57764107,0.42338464,0.36758977,0.4135385,0.74830776,1.2438976,1.910154,2.7175386,3.5774362,4.5390773,5.333334,5.930667,6.170257,5.7501545,5.6418467,5.914257,6.3901544,7.0465646,8.008205,7.9819493,8.129642,8.434873,8.891078,9.511385,9.974154,10.732308,11.644719,12.550565,13.252924,13.764924,14.119386,14.004514,13.686155,14.027489,14.454155,16.475899,17.45395,17.060104,17.27672,17.877335,18.038155,17.076513,15.218873,13.561437,13.472821,13.728822,14.04718,14.165335,13.850258,14.099693,15.176207,17.132309,18.71754,17.385027,16.584206,16.009848,15.018668,13.909334,13.925745,13.298873,13.354668,14.486976,16.288822,17.545847,18.051283,17.808413,17.30954,17.079796,17.706669,18.33354,19.767796,21.474463,22.757746,22.757746,24.612104,25.074873,24.82872,24.38236,24.07713,23.207386,23.765335,24.42831,24.208412,22.459078,20.90995,18.582975,17.801847,18.06113,16.042667,13.466257,12.557129,12.711386,13.75836,15.963899,16.712206,15.543797,14.178463,13.348104,12.793437,12.035283,11.0605135,10.476309,10.253129,9.718155,8.73354,8.421744,8.461129,8.41518,7.7390776,7.8473854,7.5881033,7.7423596,8.461129,9.265231,8.887795,7.827693,6.62318,5.989744,6.803693,6.2030773,6.1538467,6.636308,7.2894363,7.4207187,4.818052,3.9778464,3.767795,3.7874875,4.378257,4.164923,3.2032824,2.989949,3.4691284,3.05559,2.9440002,2.609231,2.546872,2.9210258,3.5872824,2.9472823,2.2449234,1.8609232,2.0184617,2.7602053,2.8127182,3.2000003,3.4494362,3.4921029,3.6660516,4.916513,5.8814363,6.2851286,6.2162056,6.1440005,7.1844106,7.8014364,8.992821,10.069334,8.661334,8.369231,8.500513,8.763078,8.960001,8.969847,8.474257,8.402052,7.827693,6.7249236,5.9569235,4.394667,2.9669745,1.9035898,1.3259488,1.2209232,0.88287187,0.90584624,0.95835906,1.1224617,1.910154,1.9528207,1.2471796,2.2416413,3.826872,1.2964103,1.7296412,4.4964104,5.9602056,5.5663595,5.8157954,13.689437,12.855796,7.8080006,4.164923,8.684308,3.515077,2.3269746,3.95159,6.675693,8.205129,7.1548724,5.5926156,4.4242053,4.089436,4.585026,3.8400004,3.6594875,4.3716927,5.4547696,5.5138464,7.0925136,7.506052,8.4053335,9.662359,9.380103,9.800206,9.449026,8.78277,8.346257,8.792616,8.214975,7.834257,8.3593855,9.449026,9.728001,9.888822,9.777231,9.508103,9.124104,8.598975,8.628513,8.182155,7.640616,7.4929237,8.310155,8.533334,8.661334,8.838565,9.101129,9.383386,9.984001,10.194052,10.194052,10.056206,9.741129,9.42277,9.232411,9.02236,8.661334,8.04759,7.6012316,7.00718,6.3179493,5.7764106,5.8157954,5.7764106,5.805949,5.6254363,5.100308,4.240411,3.639795,3.3903592,3.511795,3.6726158,3.1737437,3.1015387,3.3542566,3.5741541,3.7251284,4.1025643,3.8071797,3.5741541,3.4002054,3.3641028,3.6135387,3.7284105,3.6726158,3.501949,3.3444104,3.4133337,3.515077,3.515077,3.515077,3.4592824,3.1638978,3.43959,3.4034874,3.18359,2.917744,2.7667694,3.006359,2.7273848,2.1792822,1.7493335,1.9659488,1.8182565,1.910154,1.9626669,1.9200002,1.9429746,2.169436,2.2646155,2.356513,2.4976413,2.681436,2.8356924,3.0424619,3.6168208,4.089436,3.2262566,3.1376412,3.4264617,3.7973337,4.0467696,4.06318,4.7261543,5.3727183,5.8190775,6.2063594,7.02359,7.059693,7.6570263,7.604513,7.0498466,7.50277,7.4075904,6.2227697,5.9536414,6.7971287,7.1154876,8.116513,7.8441033,7.1515903,6.452513,5.72718,8.92718,9.921641,11.116308,16.180513,30.034054,21.88472,12.970668,8.743385,8.631796,6.0652313,8.457847,7.827693,6.8496413,6.7117953,7.131898,5.3169236,5.474462,5.464616,4.519385,3.239385,3.7185643,3.4494362,5.1167183,7.4797955,5.349744,2.6387694,1.7690258,1.6508719,1.6246156,1.4539489,0.8730257,0.6892308,0.827077,1.0732309,1.0666667,1.3226668,1.401436,1.3095386,1.1552821,1.1355898,1.148718,1.1093334,1.3226668,1.7427694,2.0086155,2.6157951,2.9538465,3.2262566,3.570872,4.0369234,3.9909747,3.006359,2.2482052,2.1497438,2.3926156,2.1891284,2.4910772,2.6026669,2.3827693,2.2646155,1.9561027,1.8609232,1.8576412,1.8609232,1.8149745,2.6256413,2.993231,3.2361028,3.436308,3.4297438,3.7940516,3.639795,3.692308,4.0303593,4.096,3.8432825,3.43959,3.0227695,2.9210258,3.6726158,4.059898,4.201026,5.0116925,6.445949,7.512616,8.759795,6.7117953,4.7327185,4.06318,3.8038976,4.6244106,5.2480006,5.549949,4.886975,2.0906668,1.7263591,2.4155898,3.3969233,4.0434875,3.8498464,4.138667,4.013949,3.442872,2.6584618,2.1530259,2.044718,2.0053334,2.15959,2.3236926,2.0020514,1.4375386,1.6935385,1.9659488,1.9954873,2.0808206,1.7558975,1.8051283,2.28759,2.8291285,2.6289232,2.6912823,3.0030773,2.9472823,2.546872,2.481231,2.4385643,2.4057438,2.2449234,2.1103592,2.4648206,2.674872,2.858667,3.121231,3.4756925,3.8596926,3.9811285,4.07959,4.309334,4.598154,4.650667,4.4406157,3.8564105,3.5872824,3.761231,3.9417439,3.6660516,3.8728209,4.4077954,4.9362054,4.955898,4.519385,4.3716927,4.4964104,4.781949,5.0510774,5.402257,5.546667,5.5302567,5.290667,4.6539493,4.893539,5.110154,4.7458467,4.013949,3.895795,3.639795,3.9023592,4.4865646,4.844308,4.069744,4.013949,4.571898,4.8607183,4.821334,5.2315903,5.5532312,6.048821,6.3934364,6.4722056,6.3934364,6.5345645,6.62318,6.872616,7.1680007,7.069539,7.210667,7.322257,7.204103,6.921847,6.7971287,6.9743595,6.872616,6.616616,6.2162056,5.5630774,5.579488,5.8912826,6.38359,6.820103,6.8365135,7.000616,6.6592827,6.2818465,6.2818465,7.0137444,7.318975,7.1089234,6.8955903,6.806975,6.5903597,6.0947695,5.3727183,4.8311796,4.644103,4.785231,4.8640003,4.713026,4.4800005,4.0303593,2.9505644,3.4166157,3.6069746,3.4756925,3.373949,4.069744,4.384821,4.598154,4.6933336,4.7261543,4.8049235,5.2742567,5.720616,5.910975,5.8847184,5.9667697,5.8223596,6.0947695,6.7085133,7.213949,6.7905645,4.348718,4.9920006,4.8311796,4.4865646,4.2863593,4.273231,4.7327185,5.412103,6.2162056,6.9776416,7.4765134,7.857231,7.9294367,8.109949,8.274052,7.752206,7.3682055,7.3682055,7.433847,7.433847,7.4469748,7.1909747,7.141744,6.7249236,6.0717955,6.0225644,6.0324106,5.4908724,5.0018463,4.778667,4.640821,4.529231,5.080616,5.4383593,5.5171285,5.98318,6.058667,6.121026,6.173539,6.12759,5.7764106,5.4514875,5.435077,5.3891287,5.290667,5.4613338,6.166975,6.1374364,6.0783596,6.0356927,5.428513,5.9602056,6.2785645,6.73477,7.3682055,7.9327188,8.411898,8.300308,8.113232,8.021334,7.8441033,7.9294367,8.073847,8.192,8.251078,8.28718,7.9491286,7.4043083,6.875898,6.5280004,6.4557953,6.692103,7.5388722,8.838565,10.262975,11.306667,11.85477,12.25518,12.58995,12.980514,13.594257,14.178463,15.707899,16.390566,15.497848,13.371078,13.5778475,13.564719,13.387488,13.078976,12.632616,12.3076935,12.045129,11.707078,11.195078,10.456616,10.381129,10.394258,9.911796,9.202872,9.412924,9.091283,8.0377445,6.7544622,5.5204105,4.388103,3.8596926,3.5347695,3.0490258,2.294154,1.4441026,0.83035904,0.5513847,0.47917953,0.45620516,0.30194873,0.53825647,0.60389745,0.6301539,0.6662565,0.67938465,0.5546667,0.5973334,0.6301539,0.60389745,0.55794877,0.574359,0.3708718,0.26256412,0.32820517,0.4266667,0.8336411,1.3784616,2.1300514,2.9571285,3.5347695,4.325744,5.1659493,5.8157954,6.012718,5.4941545,4.9132314,4.8147697,5.1200004,5.868308,7.2270775,7.2992826,7.171283,7.525744,8.251078,8.43159,8.858257,9.718155,10.482873,10.985026,11.398565,11.884309,12.773745,13.643488,14.240822,14.480412,14.178463,16.39713,18.057848,18.277744,18.392616,17.723078,17.601643,16.738462,14.976001,13.282462,12.58995,13.528616,14.5263605,14.41477,12.402873,13.000206,14.467283,16.416822,17.795284,16.902565,15.878566,15.510976,14.936617,14.168616,14.102976,13.827283,13.676309,14.562463,16.367592,17.946259,18.507488,18.405745,18.277744,18.25477,17.962667,18.185848,19.104822,20.476719,21.743591,22.029129,23.23036,24.231386,24.49067,24.182156,24.211695,23.42072,23.995079,24.402054,23.896618,22.537848,23.046566,20.04349,17.906874,17.578669,16.548103,15.120412,14.841437,14.5952835,14.598565,16.410257,17.96595,16.564514,14.578873,13.243078,12.658873,12.310975,11.825232,11.158976,10.440206,9.947898,9.412924,8.897642,8.65477,8.533334,7.9819493,7.972103,7.8802056,7.906462,8.310155,9.40636,8.89436,7.8506675,6.4754877,5.536821,6.3442054,6.3573337,6.452513,7.128616,7.7357955,6.5050263,4.450462,4.1025643,4.2601027,4.1583595,3.4691284,3.748103,3.4888208,3.4264617,3.5938463,3.3345644,3.4921029,3.2918978,3.3017437,3.5807183,3.6890259,3.31159,3.3444104,3.255795,3.249231,4.279795,4.0500517,4.46359,4.8016415,4.7294364,4.31918,5.720616,6.3606157,6.170257,5.76,6.4065647,6.75118,7.0334363,8.385642,9.931488,8.795898,8.720411,8.861539,8.999385,9.15036,9.5606165,8.753231,8.247795,7.4830775,6.5083084,5.9634876,4.273231,2.7798977,1.9200002,1.6082052,1.2438976,0.93866676,0.90912825,1.595077,2.7963078,3.6726158,1.8084104,0.92225647,3.2328207,6.5247183,4.1517954,2.2547693,4.709744,7.5913854,8.861539,8.36595,13.722258,10.28595,7.1089234,7.6964107,9.997129,4.4340515,2.6683078,5.1232824,8.677744,6.669129,5.536821,5.612308,5.428513,4.713026,4.3684106,4.9427695,5.037949,5.3398976,5.8256416,5.76,8.205129,8.257642,8.89436,10.276103,9.760821,10.433641,9.93477,8.779488,7.768616,7.968821,7.752206,7.515898,8.050873,9.179898,9.747693,9.636104,9.517949,9.399796,9.153642,8.52677,8.720411,8.441437,7.9097443,7.6603084,8.5661545,9.458873,9.432616,9.337437,9.603283,10.233437,10.683078,10.81436,10.692924,10.394258,10.010257,9.708308,9.235693,8.858257,8.595693,8.195283,7.5191803,6.928411,6.363898,5.910975,5.8157954,5.7698464,5.8125134,5.5991797,4.9788723,4.013949,3.5511796,2.989949,2.9801028,3.3411283,3.0523078,2.865231,3.2164104,3.498667,3.501949,3.4297438,3.1245131,3.0358977,3.05559,3.1409233,3.3017437,3.3542566,3.4330258,3.43959,3.4527183,3.7087183,3.626667,3.4921029,3.4921029,3.5314875,3.2262566,3.3345644,3.2754874,3.121231,2.9669745,2.92759,3.2196925,2.8914874,2.3926156,2.041436,2.038154,1.7887181,1.8510771,1.9889232,2.044718,1.9626669,2.2055387,2.3893335,2.537026,2.6551797,2.7437952,2.8488207,2.9210258,3.5774362,4.3618464,3.761231,3.5774362,3.5282054,3.757949,4.1025643,4.086154,4.525949,5.156103,5.7107697,6.189949,6.8693337,6.7216415,7.972103,8.2445135,7.2336416,6.7183595,7.1187696,6.038975,5.658257,6.2752824,6.298257,7.821129,8.027898,8.096821,8.01477,6.5444107,5.8420515,9.176616,12.704822,15.540514,19.728413,13.620514,10.410667,11.707078,14.464001,10.965334,9.212719,8.920616,8.129642,6.8299494,6.961231,5.07077,4.8705645,5.7632823,6.1046157,3.1803079,2.353231,2.4024618,4.027077,5.412103,2.225231,1.5753847,1.6410258,1.6968206,1.5688206,1.6311796,1.0469744,0.8598975,0.97805136,1.1815386,1.1126155,1.4441026,1.3817437,1.1093334,0.86646163,0.9714873,0.9911796,1.1126155,1.4900514,1.9232821,1.847795,2.7437952,3.1737437,3.501949,3.8137438,3.892513,3.639795,2.7667694,2.1989746,2.1858463,2.3072822,2.5862565,2.6715899,2.612513,2.546872,2.674872,2.3204105,2.300718,2.3401027,2.3663592,2.5009232,2.8225644,3.2262566,3.5478978,3.761231,3.9844105,4.2240005,3.9614363,4.0303593,4.4274874,4.3290257,4.414359,4.2174363,3.9909747,4.1124105,5.0904617,5.0018463,5.61559,6.7610264,8.937026,13.305437,16.978052,11.88759,6.314667,3.8695388,3.4855387,3.498667,4.161641,5.280821,6.042257,5.0149746,3.0326157,2.5698464,3.3641028,4.4701543,4.2207184,4.31918,4.073026,3.5840003,2.986667,2.428718,2.0118976,1.9396925,2.1300514,2.3204105,2.0644104,1.4834872,1.8051283,2.0676925,1.9790771,1.9298463,1.5097437,1.5786668,2.1103592,2.7503593,2.793026,2.353231,2.4746668,2.477949,2.2121027,2.048,2.3105643,2.4910772,2.3302567,2.0545642,2.3794873,2.5993848,2.7241027,2.930872,3.3378465,4.020513,4.0336413,4.1156926,4.2896414,4.466872,4.457026,4.420923,3.9614363,3.5478978,3.442872,3.7054362,3.4002054,3.4888208,3.757949,4.027077,4.1517954,4.5095387,4.7458467,5.0084105,5.2545643,5.2348723,5.074052,5.428513,5.756718,5.730462,5.2447186,5.543385,5.5269747,5.034667,4.378257,4.3290257,3.7251284,3.754667,4.2962055,4.772103,4.1452312,3.7251284,3.9351797,4.338872,4.70318,4.9920006,4.9821544,5.474462,6.1472826,6.669129,6.678975,6.5837955,6.5312824,6.5444107,6.5936418,6.5870776,6.36718,6.498462,6.488616,6.242462,6.0685134,6.4689236,6.380308,6.3868723,6.51159,6.2096415,5.8912826,6.163693,6.3212314,6.114462,5.756718,6.012718,5.7698464,5.3825645,5.395693,6.560821,7.0826674,6.616616,6.2687182,6.314667,6.2227697,5.85518,5.044513,4.138667,3.5511796,3.7973337,4.201026,4.2436924,4.0369234,3.5380516,2.537026,2.9111798,3.2918978,3.498667,3.623385,4.0336413,4.128821,4.20759,4.2568207,4.276513,4.2863593,4.8344617,5.3202057,5.4383593,5.3070774,5.4580517,5.412103,5.467898,5.868308,6.4065647,6.4295387,5.4908724,5.674667,5.5007186,5.146257,4.7425647,4.381539,4.8672824,5.2709746,5.622154,5.8945646,6.0061545,6.8004107,7.5881033,8.172308,8.36595,7.9852314,7.4863596,6.994052,6.49518,6.2162056,6.633026,6.547693,6.9382567,6.9087186,6.4032826,6.183385,5.72718,5.034667,4.562052,4.4734364,4.644103,4.7392826,5.3234878,5.586052,5.5204105,5.930667,6.3442054,6.173539,5.8486156,5.536821,5.142975,4.896821,4.8147697,4.663795,4.5062566,4.709744,5.425231,5.658257,5.4974365,5.2480006,5.4482055,6.12759,6.6560006,7.3682055,8.260923,8.976411,9.232411,9.061745,8.87795,8.825437,8.779488,8.516924,8.392206,8.260923,8.04759,7.752206,7.565129,7.584821,7.6143594,7.709539,8.152616,8.549745,8.92718,9.593436,10.345026,10.466462,10.532104,11.057232,11.431385,11.785847,13.019898,13.298873,14.336001,14.998976,14.54277,12.586668,12.593232,12.412719,12.373334,12.363488,11.835078,11.122872,10.919386,10.525539,9.862565,9.462154,10.761847,10.765129,10.6469755,10.981745,11.730052,11.867898,10.640411,8.982975,7.256616,5.2480006,4.06318,3.2984617,2.6617439,1.9692309,1.148718,0.6071795,0.3511795,0.30194873,0.31507695,0.17066668,0.19364104,0.2855385,0.3446154,0.36758977,0.446359,0.3052308,0.30851284,0.44964105,0.60389745,0.49887183,0.43651286,0.3052308,0.3117949,0.4594872,0.54482055,0.9911796,1.6114873,2.4582565,3.3509746,3.879385,4.138667,4.8016415,5.3924108,5.618872,5.3760004,4.2305646,3.69559,3.6562054,4.1878977,5.5532312,5.927385,5.805949,6.3573337,7.269744,6.738052,7.427283,8.123077,8.65477,9.061745,9.577026,9.833026,11.319796,12.747488,13.850258,15.38954,15.281232,16.918976,18.422155,18.858667,18.235079,16.774565,16.833643,16.86318,16.036104,14.250668,12.895181,13.696001,14.536206,13.988104,11.316514,13.095386,14.884104,15.875283,15.862155,15.24513,15.015386,15.081027,14.995693,14.634667,14.208001,14.513232,14.614976,15.182771,16.324924,17.59836,17.99549,18.17272,18.697847,19.10154,17.8839,18.20554,18.153027,18.432001,19.456001,21.369438,21.238155,21.956924,22.518156,22.715078,23.174566,22.245745,21.425232,20.926361,20.686771,20.36513,22.66913,21.211899,19.02277,17.562258,16.705643,16.518566,17.027283,16.649847,15.645539,16.134565,17.778873,17.030565,15.172924,13.223386,11.933539,11.657847,12.402873,12.5374365,11.631591,10.459898,10.177642,9.718155,9.216001,8.818872,8.67118,8.1755905,8.2904625,8.073847,7.88677,9.373539,9.268514,8.172308,6.6560006,5.579488,6.0685134,6.3245134,6.4000006,7.2369237,7.9130263,5.6385646,4.493129,3.9680004,3.9909747,4.086154,3.373949,3.2984617,3.5183592,3.6824617,3.6036925,3.2820516,3.9417439,4.1517954,4.5095387,5.0576415,5.3037953,5.4416413,5.546667,5.0018463,4.345436,5.284103,4.7589746,5.0543594,5.4514875,5.474462,4.896821,5.8125134,5.979898,5.85518,5.907693,6.619898,6.7610264,6.764308,8.041026,9.819899,9.160206,9.429334,9.472001,9.344001,9.186462,9.242257,8.4053335,7.7357955,6.8594875,5.9602056,5.7698464,4.1846156,2.809436,2.0906668,1.8609232,1.3259488,1.0108719,0.81066674,2.2186668,4.663795,5.5269747,1.8281027,0.8795898,4.1911798,9.051898,8.533334,4.128821,3.9680004,8.129642,13.377642,13.147899,11.723488,8.2215395,7.890052,9.77395,6.7282057,4.017231,3.5905645,6.2720003,8.707283,3.3575387,5.028103,6.7544622,6.514872,5.0904617,6.0750775,7.4896417,7.6077952,7.1844106,6.7150774,6.436103,8.149334,8.4972315,9.26195,10.210463,9.110975,10.226872,10.203898,9.160206,7.8441033,7.634052,7.9885135,7.8408213,7.9524107,8.641642,9.764103,9.32759,9.081436,9.058462,9.130668,8.999385,9.061745,9.081436,8.89436,8.687591,9.012513,10.30236,10.174359,9.957745,10.292514,11.1294365,10.8767185,10.709334,10.551796,10.371283,10.171078,10.108719,9.360411,8.713847,8.385642,8.03118,7.1056414,6.547693,6.121026,5.737026,5.4613338,5.4941545,5.3792825,5.024821,4.453744,3.7842054,3.436308,2.7536411,2.7109745,3.249231,3.2656412,3.0293336,3.0260515,3.0523078,2.934154,2.4943593,2.481231,2.5993848,2.7503593,2.9078977,3.1245131,2.92759,2.9636924,3.0752823,3.2984617,3.8596926,3.757949,3.564308,3.5511796,3.6463592,3.4297438,3.370667,3.2722054,3.2295387,3.2098465,3.0523078,3.4034874,3.1573336,2.7437952,2.3893335,2.103795,2.100513,2.1825643,2.2022567,2.1497438,2.1431797,2.3368206,2.3991797,2.556718,2.7241027,2.4943593,2.989949,3.2853336,3.945026,4.7360005,4.6539493,4.279795,3.9253337,3.8662567,4.161641,4.640821,4.2601027,4.6605134,5.435077,6.189949,6.547693,5.796103,7.269744,7.9458466,6.987488,5.733744,6.5969234,6.052103,5.7731285,6.0061545,5.546667,6.439385,6.3573337,7.3353853,8.891078,8.04759,2.8455386,7.755488,12.314258,12.885334,12.645744,8.011488,5.0871797,9.055181,16.269129,14.250668,8.411898,8.569437,8.12636,6.0061545,6.6592827,5.549949,4.2535386,5.139693,6.688821,3.4822567,2.2350771,1.2898463,0.8763078,0.8533334,0.7122052,1.7033848,2.044718,1.8904617,1.6640002,2.0742567,1.3981539,1.1979488,1.2209232,1.276718,1.2242053,1.4441026,1.2964103,1.0568206,0.96492314,1.2274873,1.1060513,1.1946667,1.8281027,2.537026,2.0709746,2.9111798,3.170462,3.5938463,4.2601027,4.59159,3.314872,2.3204105,1.9429746,2.1464617,2.5238976,3.0129232,2.6945643,2.6453335,2.9997952,2.937436,2.9571285,3.0982566,3.0687182,2.937436,3.1442053,2.6289232,3.170462,3.7120004,3.9122055,4.1714873,4.263385,4.2436924,4.352,4.5587697,4.5489235,4.916513,4.923077,4.9132314,5.1889234,6.0160003,5.9995904,7.0334363,8.172308,11.241027,20.818052,28.90831,20.217438,10.075898,5.2480006,3.9351797,2.1136413,2.0644104,2.8914874,4.647385,8.3364105,5.2414365,3.3444104,3.3608208,4.562052,4.772103,4.6276927,4.1682053,3.7940516,3.5840003,3.2820516,2.4451284,2.2678976,2.4057438,2.4713848,2.0151796,1.8937438,2.100513,2.1956925,2.0578463,1.8609232,1.4769232,1.6311796,2.0676925,2.5600002,2.9243078,2.3860514,2.1497438,2.0906668,2.0873847,2.0250258,2.5009232,2.7470772,2.5895386,2.228513,2.2580514,2.665026,2.9013336,3.121231,3.43959,3.9154875,3.9614363,4.3585644,4.453744,4.276513,4.525949,4.598154,4.2568207,3.6758976,3.1770258,3.2262566,2.9144619,2.8521028,2.8422565,2.878359,3.1409233,4.1124105,4.601436,5.0084105,5.431795,5.677949,5.0149746,5.2545643,5.723898,5.930667,5.5729237,5.802667,5.927385,5.4875903,4.6605134,4.2863593,3.7251284,3.9811285,4.6244106,4.9788723,4.125539,3.4100516,3.2853336,3.570872,4.073026,4.578462,4.6276927,4.893539,5.5532312,6.3507695,6.636308,6.5706673,6.370462,6.0816417,5.8847184,6.088206,5.874872,5.8092313,5.930667,6.0356927,5.674667,5.917539,5.9602056,6.2588725,6.692103,6.560821,6.1013336,5.9634876,5.7009234,5.2447186,4.893539,5.435077,5.6418467,5.330052,5.093744,6.265436,6.7840004,6.314667,6.045539,6.2588725,6.3245134,6.0849237,5.32677,4.1025643,2.9407182,2.8422565,3.6069746,3.7907696,3.4100516,2.7700515,2.4681027,2.878359,3.0916924,3.3805132,3.7448208,3.9089234,3.7710772,3.748103,3.7021542,3.5610259,3.314872,3.6758976,4.1452312,4.3684106,4.3585644,4.5128207,4.768821,5.093744,5.412103,5.677949,5.8486156,4.7458467,5.221744,5.605744,5.6352825,5.297231,4.821334,4.5522056,5.2545643,5.792821,5.7501545,5.431795,7.066257,7.5585647,7.50277,7.253334,6.9120007,6.705231,5.654975,4.8672824,5.0838976,6.6822567,6.2555904,6.3310776,6.363898,6.0717955,5.4613338,4.644103,4.073026,4.0303593,4.338872,4.3651285,4.352,4.6605134,4.9394875,5.3431797,6.514872,7.174565,6.47877,5.7764106,5.5072823,5.2020516,5.1922054,5.2414365,5.586052,5.832206,4.9887185,5.208616,5.0904617,5.182359,5.4843082,5.4482055,5.8125134,6.308103,6.6560006,7.0465646,8.132924,8.339693,8.612103,8.720411,8.55959,8.132924,8.083693,7.752206,7.384616,7.2861543,7.8112826,8.4972315,8.914052,9.147078,9.26195,9.324308,9.26195,9.357129,9.613129,10.102155,10.955488,10.541949,11.306667,11.776001,12.199386,14.555899,15.327181,15.363283,15.199181,14.867694,13.915898,12.245335,11.907283,11.585642,11.004719,10.955488,10.5780525,10.052924,9.527796,9.219283,9.416205,10.587898,10.587898,10.807796,11.792411,13.243078,13.243078,12.832822,12.068104,10.630565,7.8112826,6.9710774,5.549949,3.8301542,2.1497438,0.9156924,0.6104616,0.2855385,0.1148718,0.108307704,0.12143591,0.13456412,0.23958977,0.24287182,0.17723078,0.27569234,0.3117949,0.17394873,0.27897438,0.5218462,0.28882053,0.27897438,0.28225642,0.49230772,0.8041026,0.8402052,1.2537436,1.8970258,2.7634873,3.623385,4.013949,3.8432825,4.532513,5.362872,5.8289237,5.6451287,4.1189747,3.5446157,3.6693337,4.0402055,4.027077,4.578462,4.890257,5.3760004,5.8092313,5.3103595,6.163693,6.688821,7.1581545,7.7456417,8.513641,9.40636,10.561642,11.227899,11.995898,14.815181,14.815181,15.228719,15.491283,15.780104,17.014154,16.20677,15.898257,15.507693,14.76595,13.702565,13.164309,13.459693,13.633642,13.39077,13.121642,14.795488,16.000002,16.164104,15.343591,14.221129,14.966155,15.629129,16.000002,15.734155,14.342566,14.198155,14.8480015,15.537232,16.183796,17.378464,17.063385,17.706669,18.5239,18.858667,18.189129,18.530462,18.54359,17.926565,17.316103,18.281027,18.353231,19.104822,19.945026,20.502975,20.598156,21.172514,20.027079,18.707693,17.77559,16.800821,17.972515,20.214155,20.775387,19.462566,18.645334,17.94954,17.125746,16.699078,16.587488,16.098463,16.597334,17.115898,16.377438,14.299898,11.992617,11.162257,12.0549755,13.062565,12.911591,10.666668,10.725744,10.368001,10.085744,9.9282055,9.475283,8.41518,8.94359,9.042052,8.448001,8.667898,9.301334,8.546462,7.4469748,6.7544622,6.9120007,7.6931286,7.1844106,7.1220517,7.312411,5.61559,4.7622566,3.0260515,1.972513,2.0808206,2.7766156,3.7185643,3.751385,4.2436924,5.2447186,5.477744,5.172513,4.7392826,5.540103,7.318975,8.208411,6.892308,5.7468724,4.824616,4.457026,5.2480006,5.6385646,5.681231,5.61559,5.6418467,5.933949,5.861744,5.5138464,5.674667,6.2523084,6.301539,6.9120007,7.752206,8.684308,9.45559,9.6754875,9.990565,9.147078,8.395488,8.267488,8.55959,7.6931286,7.000616,6.4032826,5.8453336,5.293949,4.4406157,3.0720003,2.1956925,1.8904617,1.3259488,1.2537436,1.1815386,1.2832822,1.7558975,2.793026,1.6311796,0.9682052,1.4080001,3.8104618,9.278359,7.9097443,3.43959,3.817026,10.436924,18.12677,6.764308,4.086154,5.6418467,6.498462,1.2373334,3.8367183,6.810257,7.7948723,6.432821,4.394667,8.008205,8.326565,7.9294367,7.8834877,7.7357955,10.850462,9.091283,8.195283,9.147078,8.195283,7.0826674,6.997334,7.9852314,9.025641,8.011488,9.061745,9.596719,9.432616,9.065026,9.6754875,10.075898,9.353847,8.523488,8.39877,9.5835905,9.242257,9.025641,8.818872,8.851693,9.718155,9.537642,9.554052,9.8592825,10.171078,9.842873,10.817642,10.906258,11.024411,11.411694,11.641437,10.420513,10.108719,9.961026,9.744411,9.7214365,9.69518,9.248821,8.822155,8.448001,7.752206,7.1647186,6.5706673,5.733744,4.9493337,5.034667,5.4383593,5.1364107,4.6900516,4.332308,3.9680004,3.5511796,3.0916924,2.8291285,3.058872,4.1189747,3.876103,3.31159,2.793026,2.4451284,2.1530259,2.4320002,2.5206156,2.733949,3.0884104,3.2951798,3.3312824,3.3312824,3.4067695,3.495385,3.370667,4.0303593,4.1222568,4.128821,4.1025643,3.6627696,3.6627696,3.7907696,3.9187696,3.9187696,3.6627696,3.6627696,3.5347695,3.1803079,2.737231,2.5796926,3.006359,2.937436,2.6026669,2.3630772,2.7175386,2.6683078,2.7175386,2.8717952,2.9702566,2.7011285,3.4691284,3.945026,4.378257,4.788513,4.95918,4.6539493,4.2929235,3.757949,3.3247182,3.6758976,4.263385,4.6933336,4.926359,5.169231,5.8912826,5.927385,6.5936418,7.0531287,7.1023593,7.1876926,7.3452315,6.5903597,6.3507695,6.547693,5.586052,5.937231,5.3858466,5.533539,6.678975,7.827693,2.9078977,6.2194877,10.712616,18.162872,39.18113,29.696003,11.158976,2.6223593,6.5345645,8.743385,5.142975,8.78277,8.684308,4.450462,6.2555904,4.082872,3.0916924,4.4701543,6.193231,3.006359,2.481231,1.6804104,0.8566154,0.32164106,0.44307697,1.4933335,2.048,1.9561027,1.5753847,1.7690258,1.3686155,1.394872,1.4933335,1.4309745,1.1126155,1.332513,1.1520001,1.1520001,1.3850257,1.3718976,1.0568206,0.88615394,1.7755898,3.0227695,2.3040001,2.3040001,2.6617439,3.4067695,4.923077,7.9491286,4.7261543,2.8324106,2.0217438,2.1333334,3.0982566,3.255795,2.8750772,3.0227695,3.5971284,3.3411283,4.1583595,3.623385,3.1081028,3.2656412,3.9975388,3.4724104,3.7349746,4.066462,4.073026,3.7087183,3.4756925,4.0500517,4.6539493,5.037949,5.477744,5.208616,5.0149746,5.1298466,5.7829747,7.1876926,6.5280004,6.7840004,6.918565,9.856001,22.4919,40.484104,28.87877,15.0777445,9.452309,5.32677,1.9331284,3.006359,3.8006158,4.0402055,7.936001,6.616616,3.9975388,2.9538465,3.7973337,4.273231,4.076308,4.0369234,3.9089234,3.8071797,4.210872,3.5282054,2.934154,2.7109745,2.7602053,2.6256413,2.612513,2.5829747,2.428718,2.166154,1.9232821,1.6180514,1.7985642,2.041436,2.2646155,2.7175386,3.1081028,2.802872,2.356513,2.1858463,2.5632823,2.5993848,2.03159,1.8674873,2.2219489,2.3204105,2.8914874,3.2295387,3.6758976,4.194462,4.378257,4.31918,4.7228723,4.6933336,4.269949,4.4406157,4.1091285,3.626667,3.0687182,2.6518977,2.7011285,2.5173335,2.3269746,2.2514873,2.4943593,3.31159,4.2141542,4.650667,4.926359,5.2644105,5.8125134,4.8377438,4.893539,5.4580517,6.012718,6.0717955,6.2916927,6.7314878,6.2063594,4.6178465,2.9440002,3.1048207,4.141949,5.093744,5.3825645,4.821334,4.125539,3.629949,3.4724104,3.6627696,4.089436,4.578462,5.175795,5.6287184,5.940513,6.3934364,6.73477,6.4557953,5.973334,5.648411,5.7829747,5.733744,5.4482055,5.648411,6.294975,6.5772314,5.796103,5.0674877,5.3136415,6.121026,5.7665644,5.1331286,4.854154,5.228308,5.868308,5.720616,5.5138464,5.72718,5.648411,5.4843082,6.363898,6.803693,6.810257,6.885744,7.0432825,6.8365135,7.066257,6.997334,5.7107697,3.757949,3.1573336,3.3772311,2.993231,2.8914874,3.1048207,2.8225644,3.0194874,2.8488207,2.993231,3.495385,3.7382567,3.495385,3.5971284,3.5872824,3.2295387,2.5337439,2.9735386,3.4133337,3.8071797,4.0500517,3.95159,3.8662567,4.4045134,4.6178465,4.381539,4.394667,5.0871797,5.2709746,5.21518,5.1331286,5.07077,4.906667,5.1265645,5.861744,6.3507695,6.23918,5.579488,6.482052,7.250052,7.5421543,7.4075904,7.2894363,6.564103,5.7468724,5.182359,5.228308,6.232616,6.3606157,5.976616,5.543385,5.1659493,4.594872,4.197744,4.2240005,4.2436924,4.1714873,4.2535386,3.9286156,4.073026,4.8836927,5.933949,6.1505647,6.2227697,6.170257,5.8847184,5.5269747,5.543385,5.9930263,6.042257,6.1768208,6.23918,5.4153852,4.8640003,4.5390773,4.5817437,4.962462,5.47118,5.3103595,5.2644105,5.868308,7.02359,7.975385,8.280616,8.4512825,8.536616,8.470975,8.083693,8.113232,7.8080006,7.781744,8.316719,9.337437,9.856001,9.705027,8.979693,8.152616,8.067283,7.781744,7.8112826,8.198565,9.055181,10.564924,10.883283,11.516719,12.068104,12.888617,15.07118,16.003283,14.9628725,13.787898,13.164309,12.62277,10.597744,10.637129,11.434668,12.084514,12.0549755,11.392001,10.548513,9.593436,8.700719,8.132924,9.6754875,10.729027,11.58236,12.452104,13.476104,15.537232,15.963899,13.794462,9.957745,7.276308,5.622154,4.6080003,3.6135387,2.665026,2.4155898,1.4867693,0.64000005,0.18707694,0.1148718,0.098461546,0.098461546,0.15097436,0.16738462,0.15425642,0.21333335,0.18051283,0.23958977,0.37415388,0.4266667,0.108307704,0.15425642,0.26912823,0.41682056,0.6071795,0.88943595,1.2340513,2.0151796,2.8521028,3.4527183,3.6102567,4.1517954,4.4110775,4.699898,4.9788723,4.8640003,4.0041027,3.5807183,3.5741541,3.6824617,3.308308,4.06318,4.6900516,4.6802053,4.325744,4.7228723,5.3037953,5.658257,5.973334,6.445949,7.2927184,8.507077,9.796924,11.175385,12.337232,12.655591,12.996924,13.210258,13.302155,13.51877,14.352411,14.884104,16.262566,16.75159,15.458463,12.33395,12.1698475,12.448821,12.882052,13.453129,14.41477,15.455181,16.515284,16.610462,15.645539,14.418053,15.530668,16.059078,16.636719,17.152,16.73518,15.182771,14.54277,14.818462,15.835898,17.257027,18.198977,18.198977,18.25477,18.504206,18.212105,17.831387,17.59836,17.348925,17.174976,17.43754,16.866463,17.076513,18.57313,20.28308,19.561028,21.103592,21.215181,20.857437,20.079592,18.008617,16.994463,18.514053,19.557745,19.403488,19.610258,19.131079,18.402462,17.45395,16.597334,16.439796,16.28554,15.944206,15.241847,13.991385,12.018872,11.303386,11.464206,12.363488,13.138052,12.1928215,11.59877,11.10318,10.568206,9.938052,9.242257,9.002667,9.665642,9.819899,9.265231,8.996103,8.763078,8.461129,7.9524107,7.3386674,6.961231,7.8014364,7.6931286,6.6625648,5.3825645,5.1889234,5.0838976,3.6562054,2.4484105,2.162872,2.6551797,3.5544617,4.0500517,4.381539,4.7491283,5.284103,5.5729237,5.8157954,6.045539,6.6067696,8.172308,7.9294367,7.5421543,6.9152827,6.265436,6.1538467,5.7140517,5.540103,5.72718,6.038975,5.910975,5.612308,5.5105643,6.0652313,6.921847,6.9120007,8.070564,8.598975,9.330873,10.200616,10.236719,9.96759,10.387693,10.023385,8.940309,8.756514,8.231385,7.066257,6.2227697,5.789539,4.9788723,4.5029745,3.0785644,1.9790771,1.5655385,1.2800001,1.401436,1.3095386,1.0371283,0.96492314,1.8281027,1.2832822,0.9124103,1.2865642,2.6453335,4.8836927,6.9710774,3.43959,3.82359,8.753231,9.947898,6.4656415,6.1308722,8.205129,9.465437,4.2141542,5.5171285,7.8080006,7.834257,6.088206,6.8233852,5.8190775,5.7140517,6.36718,7.2894363,7.650462,9.163487,9.609847,9.110975,8.490667,9.317744,7.2205133,6.419693,6.557539,7.433847,8.986258,9.147078,8.825437,8.779488,9.137232,9.40636,9.5835905,8.628513,7.8506675,7.9228725,8.861539,8.881231,8.789334,8.467693,8.434873,9.816616,9.938052,10.19077,10.082462,9.642668,9.452309,10.115283,10.617436,11.083488,11.382154,11.1064625,10.400822,9.622975,8.930462,8.457847,8.316719,9.426052,9.409642,8.923898,8.277334,7.433847,7.0432825,6.6428723,6.0028725,5.2709746,4.9854364,4.706462,4.6211286,4.5817437,4.522667,4.4800005,4.493129,4.2962055,3.8859491,3.5478978,3.8400004,3.3017437,2.9440002,2.4385643,1.9626669,2.176,2.484513,3.0129232,3.3772311,3.4658465,3.4297438,3.1638978,3.3214362,3.5577438,3.636513,3.446154,3.820308,3.9220517,3.889231,3.7973337,3.6627696,3.370667,3.255795,3.31159,3.436308,3.4560003,3.629949,3.6496413,3.3936412,2.9538465,2.6387694,2.6190772,2.9440002,3.0129232,2.8882053,3.3017437,3.2722054,2.7208207,2.4451284,2.6486156,2.9571285,3.0818465,2.9636924,3.4855387,4.516103,4.9099493,4.6145644,4.493129,4.164923,3.5347695,2.7864618,4.076308,5.1364107,5.3005133,4.8705645,5.1331286,5.32677,5.5926156,5.861744,6.2818465,7.2369237,6.380308,5.7501545,5.7107697,5.835488,4.900103,5.5105643,5.3727183,5.677949,6.675693,7.6570263,5.2381544,9.156924,9.7903595,12.905026,39.696415,38.92185,18.12349,4.315898,4.8640003,7.4732313,5.7764106,8.963283,8.832001,5.297231,6.3901544,5.720616,4.066462,3.5052311,3.8006158,2.3696413,2.4713848,2.166154,1.4834872,0.8533334,1.1027694,2.169436,2.3072822,2.169436,2.2350771,2.7831798,2.3401027,2.1169233,2.0644104,2.0906668,2.0644104,1.6804104,1.3981539,1.339077,1.4309745,1.3981539,1.2668719,1.0108719,1.4375386,2.2153847,1.8773335,1.585231,1.6935385,2.4910772,3.5478978,3.7152824,2.8258464,2.5600002,2.2022567,2.034872,3.3411283,3.7054362,3.754667,3.6135387,3.5905645,4.1846156,4.3290257,4.135385,3.9253337,3.8104618,3.692308,3.5971284,3.8728209,3.9909747,4.023795,4.6244106,4.381539,4.578462,4.818052,5.034667,5.5138464,5.989744,5.861744,5.5269747,5.8256416,8.027898,7.4174366,7.762052,7.581539,8.625232,15.839181,24.536617,18.477951,11.044104,8.093539,7.962257,6.0816417,4.086154,3.1113849,3.8662567,6.629744,5.3398976,3.754667,2.9243078,3.0490258,3.4658465,4.06318,4.7261543,4.778667,4.4734364,4.9920006,4.640821,4.066462,3.8990772,3.9680004,3.2951798,2.8750772,2.7700515,2.422154,1.7788719,1.2996924,1.3653334,1.4769232,1.7362052,2.2121027,2.9472823,3.2984617,3.1671798,2.6256413,2.0020514,1.8937438,2.2908719,2.2088206,2.2350771,2.4681027,2.5271797,3.0720003,3.2984617,3.446154,3.6496413,3.9384618,4.082872,3.9909747,3.892513,3.892513,3.9647183,3.751385,3.442872,2.9702566,2.5238976,2.5435898,2.300718,2.166154,2.231795,2.5238976,3.0293336,3.639795,4.2896414,4.896821,5.4482055,6.009436,5.481026,5.110154,4.857436,4.824616,5.2545643,5.7009234,5.72718,5.5236926,4.9952826,3.761231,3.7743592,4.138667,4.2962055,4.092718,3.7842054,3.8400004,4.0467696,4.1813335,4.2141542,4.309334,4.630975,5.0838976,5.395693,5.579488,5.940513,6.4295387,6.669129,6.4590774,5.907693,5.4153852,5.349744,5.0871797,5.110154,5.4449234,5.6352825,5.7042055,5.609026,5.858462,6.265436,5.9503593,5.540103,5.474462,5.832206,6.3474874,6.4065647,5.691077,5.0215387,4.630975,4.906667,6.413129,6.8594875,7.1581545,7.2861543,7.1614366,6.6395903,7.496206,7.4732313,6.301539,4.588308,3.7940516,3.826872,3.6463592,3.5807183,3.5347695,2.9702566,2.674872,2.3893335,2.5238976,3.0752823,3.639795,3.4560003,3.501949,3.3969233,3.0227695,2.5206156,2.9604106,3.062154,3.0194874,2.9604106,2.9505644,3.3542566,3.8301542,4.092718,4.076308,3.9318976,4.896821,4.8607183,4.818052,4.906667,4.9329233,4.378257,5.2545643,6.232616,6.8397956,6.7971287,5.9995904,6.3179493,6.875898,7.066257,6.8594875,6.8004107,6.193231,5.986462,6.0717955,6.3212314,6.6133337,6.491898,5.9667697,5.366154,4.8082056,4.1878977,4.276513,4.4406157,4.391385,4.132103,3.9417439,3.5249233,4.023795,5.2709746,6.5444107,6.5706673,5.970052,5.8256416,5.7632823,5.723898,5.9602056,6.5378466,6.363898,6.038975,5.674667,4.900103,4.713026,4.7261543,4.9296412,5.297231,5.789539,5.182359,5.1626673,6.0849237,7.384616,7.5585647,7.755488,7.788308,7.821129,8.004924,8.474257,8.274052,7.8703594,7.817847,8.214975,8.704,8.717129,8.487385,7.9917955,7.322257,6.678975,6.6395903,7.0465646,7.9950776,9.265231,10.322052,11.444513,12.196103,12.356924,12.3536415,13.266052,13.787898,13.433437,12.708103,11.946668,11.300103,10.118565,10.338462,10.981745,11.447796,11.542975,11.067078,10.039796,8.996103,8.297027,8.14277,9.96759,11.457642,12.517745,13.725539,16.31836,18.835693,18.569847,15.90154,12.137027,9.501539,6.0225644,3.8629746,2.7076926,2.28759,2.3893335,1.2504616,0.7450257,0.49230772,0.29210258,0.128,0.10502565,0.13784617,0.15097436,0.13456412,0.1148718,0.08861539,0.16738462,0.21333335,0.16410258,0.04266667,0.08205129,0.17066668,0.28225642,0.43323082,0.67282057,1.2931283,2.2088206,3.062154,3.5938463,3.6463592,3.9122055,4.082872,4.2240005,4.3290257,4.312616,4.240411,3.8137438,3.5314875,3.4002054,2.937436,3.8596926,4.1813335,3.9581542,3.6758976,4.2469745,4.086154,4.4767184,4.854154,5.152821,5.8092313,7.2992826,8.605539,10.006975,11.122872,10.896411,11.67754,11.946668,11.989334,12.06154,12.416001,13.66318,14.79877,15.793232,15.872002,13.522053,13.213539,13.289026,13.952001,14.976001,15.675078,16.354464,17.024002,16.90913,16.059078,15.343591,16.25272,15.95077,15.977027,16.81395,17.900309,16.935387,15.724309,15.261539,15.698052,16.347898,17.6279,18.497643,19.058874,19.318155,19.18031,17.946259,17.079796,16.62359,16.682669,17.417847,16.613745,17.030565,18.313848,19.748104,20.263386,20.368412,20.404514,21.03795,21.766565,20.900105,18.95713,18.819284,18.904617,18.917746,19.85313,20.040207,20.007385,18.983387,17.444103,17.11918,16.633438,15.67836,14.729847,13.797745,12.416001,11.398565,12.12718,13.1872835,13.702565,13.341539,11.808822,11.0375395,10.384411,9.793642,9.800206,9.747693,9.747693,9.40636,8.89436,8.940309,8.241231,8.096821,7.857231,7.2270775,6.2588725,6.87918,7.430565,6.3934364,4.4045134,4.266667,5.0116925,4.082872,2.9144619,2.4451284,3.117949,4.141949,4.8804107,5.110154,5.10359,5.618872,6.2916927,6.8233852,6.9021544,7.00718,8.418462,8.598975,8.346257,7.328821,6.045539,5.865026,5.4383593,5.3234878,5.4514875,5.661539,5.684513,5.5663595,6.0652313,6.9054365,7.6964107,7.936001,8.87795,9.521232,10.417232,11.303386,11.099898,10.492719,10.729027,10.492719,9.622975,9.097847,8.329846,6.8988724,6.2194877,6.170257,5.100308,4.7360005,3.31159,2.2186668,1.8149745,1.4145643,1.4441026,1.3489232,1.3489232,1.585231,2.1169233,1.6114873,1.1060513,1.1815386,1.847795,2.556718,6.2063594,4.0336413,4.276513,7.4404106,6.265436,5.602462,5.8190775,7.8670774,9.6295395,5.9470773,5.431795,5.7501545,6.114462,6.6560006,8.418462,5.9963083,5.349744,5.5729237,6.0750775,6.5870776,7.1614366,8.280616,8.503796,7.906462,8.077128,6.7150774,5.8486156,5.4875903,5.858462,7.4174366,8.572719,8.621949,8.470975,8.477539,8.43159,8.4283085,7.9130263,7.683283,7.9885135,8.507077,8.612103,8.628513,8.349539,8.195283,9.209436,9.229129,9.40636,9.163487,8.707283,9.025641,8.848411,9.42277,10.108719,10.492719,10.374565,10.35159,9.688616,9.015796,8.684308,8.763078,9.67877,9.777231,9.40636,8.786052,7.9852314,7.322257,6.705231,6.1997952,5.7435904,5.139693,4.33559,4.3290257,4.598154,4.7983594,4.7556925,4.568616,4.3684106,4.07959,3.7809234,3.69559,3.1507695,2.9472823,2.740513,2.553436,2.7864618,3.1048207,3.4888208,3.7021542,3.7152824,3.7185643,3.3476925,3.249231,3.373949,3.5840003,3.6463592,3.8564105,3.892513,3.764513,3.623385,3.7448208,3.5544617,3.2196925,3.1376412,3.3214362,3.4297438,3.495385,3.3903592,3.0752823,2.7044106,2.6289232,2.9243078,3.0720003,3.0949745,3.0818465,3.2000003,3.0752823,2.7208207,2.5074873,2.6223593,3.058872,3.6660516,3.3476925,3.4724104,4.1714873,4.322462,4.5128207,4.772103,4.420923,3.6069746,3.314872,4.604718,5.4514875,5.622154,5.3169236,5.1922054,4.9985647,4.9952826,5.139693,5.5663595,6.560821,6.0061545,6.0028725,6.2851286,6.2555904,5.0051284,5.293949,4.9920006,5.159385,6.0291286,6.99077,5.35959,10.033232,11.707078,11.61518,21.526976,28.340515,14.404924,3.7940516,4.6112823,8.969847,6.8627696,8.320001,7.9950776,5.6254363,6.0225644,7.7948723,5.1856413,3.4067695,3.5807183,2.7602053,2.4976413,2.2613335,1.8937438,1.5425643,1.6771283,2.1464617,2.0217438,2.0578463,2.5304618,3.2754874,3.2032824,2.9997952,2.8816411,2.8980515,2.9538465,2.3729234,1.723077,1.3357949,1.2471796,1.211077,1.595077,1.4900514,1.7952822,2.4352822,2.3368206,1.972513,1.7755898,2.1234872,2.678154,2.409026,2.103795,1.9659488,1.8642052,2.0906668,3.367385,3.757949,4.391385,4.210872,3.5544617,4.1550775,3.8596926,4.017231,4.417641,4.6572313,4.128821,4.0303593,4.2601027,4.312616,4.2830772,4.8607183,4.457026,4.713026,5.024821,5.142975,5.175795,5.8847184,5.431795,4.916513,5.028103,6.0324106,5.83877,9.140513,9.944616,8.251078,10.072617,14.01436,13.010053,11.447796,12.681848,19.058874,25.96431,15.419078,5.3366156,2.8980515,4.562052,5.0018463,3.7185643,3.0030773,3.2918978,3.1737437,4.312616,5.175795,5.2545643,4.9329233,5.481026,5.474462,4.857436,4.460308,4.3618464,3.8564105,3.0982566,2.737231,2.2580514,1.6246156,1.2635899,1.2307693,1.4375386,1.7329233,2.038154,2.3368206,2.9210258,2.8882053,2.4943593,2.1169233,2.228513,2.4746668,2.6551797,2.8914874,3.0916924,2.9636924,3.1474874,3.318154,3.570872,3.7152824,3.2722054,3.7218463,3.442872,3.1803079,3.2722054,3.6332312,3.2328207,3.1737437,2.930872,2.4746668,2.2744617,2.3236926,2.1792822,2.2646155,2.6256413,2.9144619,3.4133337,4.1747694,4.8049235,5.2545643,5.802667,5.2611284,4.516103,4.2896414,4.709744,5.3169236,5.4416413,5.2020516,5.0674877,4.9854364,4.352,3.8367183,4.023795,4.1025643,3.8728209,3.7448208,3.8334363,4.1222568,4.342154,4.460308,4.6834874,4.824616,5.1889234,5.395693,5.4547696,5.7468724,6.1768208,6.445949,6.445949,6.1013336,5.353026,4.781949,4.8082056,4.9329233,5.0510774,5.4580517,5.6418467,5.8814363,6.166975,6.2752824,5.786257,5.4383593,5.7009234,5.9634876,5.940513,5.671385,5.208616,4.397949,4.141949,4.6834874,5.6287184,5.858462,6.482052,6.770872,6.6395903,6.619898,6.5772314,5.973334,5.2545643,4.604718,3.9154875,3.9023592,4.020513,4.138667,4.073026,3.5544617,3.242667,2.5042052,2.2186668,2.5895386,3.1409233,3.190154,3.1770258,3.1245131,2.9997952,2.7011285,2.7241027,2.6322052,2.5764105,2.609231,2.674872,3.0523078,3.3280003,3.4560003,3.4592824,3.4297438,5.464616,5.110154,5.0609236,5.0674877,4.7524104,3.6036925,5.4383593,6.5411286,7.2172313,7.3452315,6.38359,6.452513,6.564103,6.521436,6.308103,6.091488,5.914257,6.3212314,6.9382567,7.3419495,7.0531287,6.488616,5.937231,5.412103,4.919795,4.4373336,4.5390773,4.4045134,4.1583595,3.892513,3.6496413,3.3969233,4.2141542,5.5236926,6.6592827,6.8332314,5.9503593,5.677949,5.7403083,5.940513,6.1505647,6.7905645,6.6428723,6.2851286,5.8814363,5.1954875,5.356308,5.756718,6.193231,6.3474874,5.7764106,5.2020516,5.6418467,6.567385,7.4010262,7.50277,7.778462,7.509334,7.2172313,7.276308,7.906462,7.6734366,7.0990777,6.8332314,7.017026,7.276308,7.256616,7.2270775,7.062975,6.6395903,5.8256416,5.648411,5.98318,6.951385,8.251078,9.16677,10.47959,11.017847,10.840616,10.41395,10.604308,10.725744,10.981745,10.952206,10.65354,10.532104,10.069334,10.197334,10.5780525,10.909539,10.948924,10.262975,9.403078,8.736821,8.441437,8.4972315,10.489437,11.641437,12.885334,15.048206,18.852104,21.270975,20.427488,18.81272,16.784412,12.57354,7.0793853,3.370667,1.6344616,1.4145643,1.6082052,0.7187693,0.55794877,0.5152821,0.3511795,0.190359,0.13784617,0.14441027,0.13456412,0.0951795,0.049230773,0.036102567,0.072205134,0.06235898,0.01969231,0.049230773,0.068923086,0.13128206,0.23630771,0.40369233,0.6465641,1.4736412,2.3433847,2.9538465,3.2787695,3.5446157,3.3608208,3.5511796,3.748103,3.820308,3.8662567,3.9975388,3.7415388,3.43959,3.259077,3.1671798,3.7940516,3.7940516,3.6168208,3.5544617,3.761231,3.1803079,3.4166157,3.9154875,4.4373336,5.0576415,5.904411,7.253334,8.910769,10.161232,9.780514,10.203898,10.331899,10.266257,10.226872,10.551796,12.649027,13.801026,14.772514,15.451899,14.8709755,14.529642,14.670771,15.43877,16.341335,16.25272,16.95836,17.168411,16.68595,15.908104,15.832617,16.219898,15.675078,15.570052,16.46277,18.07754,18.133335,17.083078,16.049232,15.520822,15.340309,16.338053,17.749334,18.934155,19.636515,19.990976,18.23836,16.794258,15.977027,16.019693,17.060104,16.794258,17.355488,18.294155,19.334566,20.374975,19.91549,19.866259,20.647387,21.697643,21.4679,21.014977,20.187899,19.19672,18.582975,19.22954,19.843283,19.856411,19.206566,18.290873,17.992207,17.444103,15.91795,14.49354,13.627078,13.138052,11.83836,12.668719,13.791181,14.244103,13.965129,12.301129,10.886565,9.878975,9.5835905,10.453334,10.473026,9.626257,8.848411,8.598975,8.845129,8.425026,8.024616,7.5487185,6.87918,5.8486156,6.055385,6.698667,6.1374364,4.535795,3.892513,4.5029745,3.8662567,2.8816411,2.356513,2.989949,4.378257,5.297231,5.756718,5.917539,6.1013336,6.4000006,7.4436927,7.8539495,7.6931286,8.467693,8.621949,8.260923,7.259898,6.0619493,5.651693,5.477744,5.4153852,5.428513,5.5991797,6.11118,5.8223596,6.5083084,7.3649235,8.162462,9.278359,9.544206,10.417232,11.526565,12.35036,12.22236,11.861334,11.382154,10.617436,9.639385,8.736821,7.5618467,6.3343596,5.9536414,6.091488,5.1987696,4.5390773,3.570872,2.4943593,1.654154,1.5524104,1.3850257,1.0765129,1.6443079,2.8717952,3.3312824,1.9298463,1.0929232,0.9353847,1.2471796,1.4900514,5.6385646,5.677949,5.6418467,6.1768208,4.5456414,5.609026,5.723898,6.7544622,7.8834877,5.618872,6.380308,5.333334,5.431795,7.253334,9.025641,6.242462,5.0477953,4.8672824,5.277539,6.0061545,5.9470773,6.3901544,6.5936418,6.550975,6.9677954,6.226052,5.5236926,4.9854364,4.850872,5.477744,7.020308,7.7292314,7.7325134,7.4404106,7.5454364,7.6767187,7.4929237,7.568411,7.9950776,8.39877,8.569437,8.490667,8.1755905,7.939283,8.379078,7.9885135,7.827693,7.6012316,7.525744,8.2904625,7.9885135,8.55959,9.31118,9.714872,9.412924,9.993847,9.77395,9.429334,9.32759,9.544206,9.764103,9.895386,9.701744,9.127385,8.2904625,7.509334,6.7905645,6.311385,5.937231,5.2053337,4.2207184,4.1091285,4.519385,5.028103,5.139693,4.6080003,4.1714873,3.9614363,3.9680004,4.020513,3.5971284,3.5282054,3.5872824,3.639795,3.6463592,3.7021542,3.6693337,3.764513,3.9811285,4.092718,3.6824617,3.367385,3.3050258,3.4494362,3.5610259,3.6004105,3.7120004,3.7776413,3.7907696,3.8596926,3.7874875,3.3575387,3.1048207,3.1245131,3.0687182,3.1606157,3.2623591,3.0818465,2.7044106,2.6026669,3.1737437,3.2131286,3.058872,2.9144619,2.8521028,2.8127182,2.7536411,2.6978464,2.7864618,3.2787695,4.4274874,4.1156926,3.8596926,4.069744,4.0336413,4.6112823,4.972308,4.44718,3.5840003,4.1189747,5.3005133,5.5236926,5.4613338,5.431795,5.412103,4.7622566,4.6276927,4.673641,4.84759,5.3727183,5.579488,5.917539,6.232616,6.166975,5.156103,4.9985647,4.667077,4.7360005,5.5204105,7.076103,5.2742567,8.556309,11.008,10.187488,7.145026,13.013334,7.571693,3.9056413,5.7764106,7.6143594,6.7577443,7.0400004,6.816821,6.1505647,6.820103,8.402052,5.602462,3.623385,3.7152824,3.1540515,2.3236926,1.9396925,1.8018463,1.7788719,1.8313848,1.8970258,1.6869745,1.785436,2.3466668,3.0851285,3.4888208,3.6529233,3.754667,3.8038976,3.6496413,3.0687182,2.2482052,1.6049232,1.3062565,1.2832822,1.9167181,2.0939488,2.4516926,2.92759,2.7470772,2.477949,2.3138463,2.4320002,2.6584618,2.4582565,1.8838975,1.5524104,1.6836925,2.28759,3.1540515,3.31159,4.397949,4.378257,3.4560003,4.0467696,3.9187696,3.9975388,4.4701543,4.919795,4.3290257,4.3060517,4.3585644,4.4110775,4.516103,4.8607183,4.5062566,4.713026,5.0182567,5.0149746,4.3651285,5.3202057,4.788513,4.3585644,4.345436,3.817026,5.720616,11.1983595,12.763899,9.908514,9.097847,11.464206,14.815181,17.027283,20.627693,32.784412,51.521645,33.16513,11.72677,2.7733335,3.4100516,4.9132314,3.761231,3.242667,3.9253337,3.6627696,4.6276927,5.21518,5.293949,5.2348723,5.920821,5.730462,5.1889234,4.7491283,4.5456414,4.3749747,3.508513,3.062154,2.3696413,1.5195899,1.3423591,1.3292309,1.4834872,1.6311796,1.7132308,1.7690258,2.4057438,2.3958976,2.2580514,2.3630772,2.9243078,2.9210258,3.18359,3.4789746,3.5807183,3.2623591,3.5314875,3.623385,3.8301542,3.9318976,3.2098465,3.5249233,3.0949745,2.5665643,2.4320002,3.0227695,2.605949,2.8882053,2.9472823,2.6551797,2.6715899,2.7076926,2.5928206,2.6617439,2.930872,3.121231,3.446154,3.9811285,4.2601027,4.4077954,5.156103,4.7556925,3.9581542,3.8367183,4.5456414,5.3037953,5.175795,4.841026,4.630975,4.5554876,4.279795,3.754667,3.8564105,4.017231,4.0434875,4.1156926,4.086154,4.197744,4.3618464,4.598154,5.024821,5.1626673,5.395693,5.4941545,5.4449234,5.4547696,5.8289237,6.1505647,6.2752824,6.121026,5.671385,4.6244106,4.59159,4.7360005,4.893539,5.5532312,5.5236926,5.85518,6.0685134,5.8880005,5.218462,5.1200004,5.7107697,5.8453336,5.3103595,4.827898,4.8311796,4.135385,4.020513,4.6145644,4.9132314,4.916513,5.330052,5.579488,5.737026,6.521436,5.7435904,4.955898,4.598154,4.4800005,3.7874875,4.1452312,4.125539,4.0041027,3.9318976,3.9220517,3.8334363,3.0129232,2.4024618,2.3827693,2.7437952,3.006359,2.937436,2.802872,2.7044106,2.5796926,2.425436,2.4188719,2.4976413,2.5731285,2.5140514,2.6683078,2.8455386,2.9538465,2.9702566,2.9111798,6.409847,5.8223596,5.789539,5.4416413,4.493129,3.2229745,5.6943593,6.7249236,7.4404106,7.830975,6.7610264,6.5936418,6.3573337,6.2227697,6.1013336,5.668103,6.009436,6.7183595,7.381334,7.64718,7.2205133,6.49518,5.98318,5.687795,5.481026,5.110154,4.6769233,4.0500517,3.639795,3.5347695,3.5052311,3.6791797,4.565334,5.609026,6.3606157,6.4722056,5.858462,5.730462,5.904411,6.157129,6.2063594,6.9120007,7.0925136,7.062975,6.9021544,6.4557953,6.669129,7.4010262,7.972103,7.6767187,5.7632823,5.3234878,6.114462,6.688821,6.8004107,7.4207187,7.8441033,7.39118,6.872616,6.6034875,6.4000006,6.298257,5.6976414,5.3891287,5.6254363,6.124308,6.4295387,6.688821,6.619898,6.196513,5.6451287,5.0051284,4.84759,5.280821,6.2194877,7.4141545,8.280616,8.277334,7.9917955,7.830975,8.041026,8.04759,8.418462,9.019077,9.728001,10.423796,10.144821,9.977437,10.266257,10.692924,10.30236,9.088,8.736821,8.736821,8.766359,8.694155,10.689642,11.339488,12.937847,16.108309,19.784206,21.796104,21.064207,20.94277,20.673643,15.369847,8.155898,3.2689233,0.92553854,0.53825647,0.69251287,0.35446155,0.28882053,0.31507695,0.3446154,0.3708718,0.30851284,0.20348719,0.11158975,0.055794876,0.036102567,0.016410258,0.013128206,0.01969231,0.04266667,0.08205129,0.128,0.2297436,0.36758977,0.57764107,0.9353847,1.7723079,2.3827693,2.553436,2.5173335,2.9636924,2.674872,2.9505644,3.245949,3.3542566,3.4002054,3.4100516,3.4560003,3.3903592,3.3280003,3.6791797,3.6791797,3.5183592,3.4789746,3.515077,3.239385,2.7798977,2.7667694,3.3017437,4.1747694,4.857436,4.667077,6.0192823,7.9852314,9.344001,8.592411,8.267488,8.15918,8.100103,8.254359,9.114257,11.785847,13.653335,14.444309,14.552616,15.028514,14.752822,15.228719,15.95077,16.288822,15.497848,16.393847,16.505438,15.996719,15.474873,15.96718,16.082052,16.009848,16.193642,16.7319,17.381744,17.811693,17.473642,16.534975,15.442053,14.920206,15.589745,16.617027,17.818258,19.003078,19.984411,18.36308,16.676104,15.707899,15.691488,16.31836,16.928822,17.306257,18.008617,18.947283,19.419899,20.155079,20.457027,20.601437,20.466873,19.515078,21.454771,21.592617,20.565334,19.22954,18.635489,18.714258,18.330257,18.277744,18.599386,18.592821,18.336823,16.361027,14.401642,13.466257,13.846975,12.829539,12.793437,13.617231,14.536206,14.112822,13.02318,11.073642,9.787078,9.7903595,10.811078,10.925949,9.468719,8.579283,8.809027,9.107693,9.350565,8.503796,7.4797955,6.695385,6.0750775,5.9602056,6.196513,6.0816417,5.356308,4.2207184,4.132103,3.5314875,2.6420515,1.9987694,2.422154,4.066462,5.0543594,5.874872,6.498462,6.370462,5.8125134,7.4207187,8.411898,8.201847,8.411898,8.490667,8.214975,7.6931286,6.9054365,5.717334,5.7042055,5.723898,5.76,6.0291286,6.9710774,6.294975,6.6494365,7.325539,8.3134365,10.295795,10.427077,11.644719,12.76718,13.269335,13.266052,13.403898,12.3995905,10.788103,9.153642,8.155898,6.564103,5.8453336,5.5762057,5.431795,5.182359,3.9318976,3.4560003,2.4352822,1.1454359,1.4703591,1.1552821,0.8041026,1.8576412,3.8104618,4.1911798,3.2065644,2.0676925,1.4605129,1.4309745,1.4080001,5.4613338,7.9163084,7.430565,4.9132314,3.508513,6.6822567,6.301539,5.5958977,5.5663595,4.97559,7.9195905,6.8266673,6.193231,7.3747697,8.592411,5.8814363,4.3684106,4.1846156,4.9821544,5.943795,5.428513,4.9493337,4.630975,4.8804107,6.377026,5.901129,5.405539,4.896821,4.460308,4.2535386,4.9394875,6.0225644,6.491898,6.432821,7.0137444,7.4075904,7.269744,7.259898,7.6274877,8.192,8.507077,8.211693,7.8112826,7.6209235,7.762052,7.13518,6.636308,6.4623594,6.738052,7.4896417,7.8670774,8.553026,9.248821,9.508103,8.730257,9.475283,9.668923,9.665642,9.685334,9.810052,9.337437,9.435898,9.363693,8.818872,7.9228725,7.2172313,6.6560006,6.1308722,5.5696416,4.9362054,4.2502565,3.9876926,4.2994876,4.9427695,5.280821,4.7655387,4.1911798,3.9581542,4.1517954,4.5489235,4.194462,4.135385,4.269949,4.4012313,4.2535386,4.0402055,3.757949,3.879385,4.2962055,4.2994876,3.882667,3.5774362,3.3641028,3.2361028,3.18359,3.1277952,3.4002054,3.767795,4.0041027,3.876103,3.7842054,3.4002054,3.05559,2.809436,2.4681027,2.681436,3.2065644,3.308308,2.8882053,2.484513,2.9078977,3.1376412,3.0030773,2.6683078,2.6322052,2.9013336,2.8488207,2.7733335,2.9636924,3.692308,4.95918,4.7228723,4.325744,4.2929235,4.315898,4.785231,4.9427695,4.391385,3.7743592,4.775385,5.8190775,5.435077,4.9460516,4.9362054,5.277539,4.578462,4.457026,4.4832826,4.460308,4.457026,5.175795,5.467898,5.5630774,5.4908724,5.0609236,4.5423594,4.5029745,4.713026,5.425231,7.3747697,6.0750775,6.4623594,7.4436927,7.433847,4.338872,5.080616,4.634257,5.5696416,6.875898,3.9351797,6.413129,6.2588725,5.796103,6.2063594,7.5388722,6.514872,4.647385,3.5380516,3.4100516,3.0818465,2.0841026,1.5622566,1.4933335,1.6804104,1.7362052,1.847795,1.654154,1.6180514,1.9331284,2.5206156,3.259077,3.945026,4.4274874,4.5423594,4.1124105,3.5774362,2.8717952,2.1956925,1.7427694,1.6902566,2.0709746,2.5632823,3.045744,3.242667,2.7142565,2.6289232,2.7208207,2.9111798,2.9997952,2.6551797,1.7657437,1.4309745,1.7033848,2.300718,2.5961027,2.553436,3.8071797,4.138667,3.6890259,4.9526157,4.598154,4.128821,4.1747694,4.571898,4.3716927,4.3651285,4.125539,4.1813335,4.5554876,4.7622566,4.818052,4.772103,4.7983594,4.673641,3.7448208,4.818052,4.598154,4.4340515,4.2896414,2.7175386,7.6931286,12.452104,13.4859495,11.434668,11.07036,14.339283,20.65067,24.041027,28.274874,46.85785,71.634056,47.379696,17.58195,3.3378465,3.3411283,4.4045134,3.6857438,3.501949,4.2305646,4.322462,4.778667,4.709744,4.841026,5.421949,6.2227697,5.4580517,5.0904617,4.8738465,4.7491283,4.8640003,4.059898,3.6529233,2.7503593,1.5721027,1.4375386,1.5983591,1.5786668,1.4703591,1.3915899,1.5064616,1.9298463,1.9856411,2.1366155,2.6157951,3.4330258,3.3641028,3.508513,3.7120004,3.751385,3.3214362,3.9220517,3.8301542,3.7415388,3.7874875,3.5380516,3.318154,2.809436,2.166154,1.7493335,2.1103592,2.0053334,2.5928206,2.9735386,3.0293336,3.4067695,3.1967182,3.114667,3.114667,3.1671798,3.2853336,3.3509746,3.5577438,3.4592824,3.373949,4.381539,4.273231,3.7021542,3.5446157,4.086154,5.041231,4.969026,4.644103,4.2535386,3.945026,3.82359,3.7284105,3.6332312,3.7874875,4.161641,4.460308,4.4307694,4.352,4.4045134,4.6867695,5.221744,5.435077,5.5762057,5.605744,5.4908724,5.1954875,5.5236926,6.0028725,6.1046157,5.8847184,5.9667697,5.031385,4.6145644,4.5489235,4.7983594,5.467898,5.2742567,5.58277,5.6287184,5.182359,4.5554876,4.896821,5.5565133,5.5565133,4.919795,4.673641,4.778667,4.2929235,4.1747694,4.519385,4.562052,4.670359,4.4865646,4.453744,4.923077,6.173539,5.5663595,5.093744,4.7983594,4.522667,3.9187696,4.6605134,4.1813335,3.5741541,3.4527183,3.9384618,4.023795,3.4330258,2.733949,2.3335385,2.481231,2.7536411,2.740513,2.5206156,2.28759,2.3368206,2.3236926,2.5435898,2.6715899,2.5829747,2.3729234,2.3827693,2.5206156,2.6715899,2.6912823,2.428718,5.677949,5.481026,6.0717955,5.586052,4.197744,4.1517954,5.5663595,6.488616,7.4699492,8.201847,7.506052,6.2752824,6.2030773,6.3507695,6.242462,5.874872,6.705231,7.177847,7.177847,6.9776416,7.2336416,6.9776416,6.692103,6.626462,6.5017443,5.540103,4.391385,3.564308,3.3378465,3.5446157,3.5544617,4.3716927,5.2381544,6.012718,6.314667,5.5072823,5.5565133,5.7698464,6.11118,6.4623594,6.62318,7.256616,7.709539,7.5618467,7.0892315,7.24677,7.785026,9.107693,9.504821,8.536616,7.0334363,5.654975,5.76,5.910975,5.737026,5.920821,5.933949,6.11118,6.452513,6.5083084,5.3858466,5.0215387,4.9099493,5.2512827,5.832206,6.0258465,5.989744,6.419693,6.616616,6.3277955,5.7665644,5.290667,5.1987696,5.474462,6.0324106,6.7282057,7.1548724,6.9054365,6.547693,6.294975,6.0258465,6.160411,7.1483083,8.910769,10.607591,10.620719,10.486155,10.049642,9.77395,9.435898,8.116513,7.069539,7.3714876,7.837539,8.109949,8.681026,10.453334,11.792411,13.909334,16.843489,19.456001,20.187899,19.75795,18.720821,17.736206,17.578669,9.058462,3.767795,1.1191796,0.26584616,0.108307704,0.26584616,0.40697438,0.5152821,0.64000005,0.88615394,0.8598975,0.45292312,0.13456412,0.06235898,0.06235898,0.013128206,0.0,0.01969231,0.059076928,0.108307704,0.28882053,0.48246157,0.6892308,0.94523084,1.3128207,2.1431797,2.4057438,2.3269746,2.0841026,1.8149745,1.9856411,2.5600002,2.865231,2.789744,2.7766156,3.5577438,3.6529233,3.629949,3.6693337,3.570872,3.314872,2.8947694,2.802872,2.9702566,2.7634873,2.6289232,2.8324106,3.186872,3.5511796,3.8465643,4.1517954,5.1889234,6.2490263,6.636308,5.661539,5.904411,6.157129,6.738052,7.821129,9.4457445,10.837335,12.813129,14.188309,14.431181,13.686155,12.931283,13.538463,14.116103,13.899488,12.724514,13.459693,14.49354,15.323898,15.990155,17.089642,18.054565,18.15631,17.828104,17.138874,15.809642,15.356719,15.911386,16.229744,15.983591,15.763694,16.922258,17.293129,17.59836,18.166155,18.937437,18.241642,16.784412,16.193642,16.52513,16.282257,16.843489,17.02072,17.319386,17.942976,18.799591,20.95918,21.609028,21.333336,20.38154,18.661745,19.712002,21.897848,22.87918,21.943796,20.004105,17.85436,18.261335,18.579693,18.113642,18.12677,18.763489,16.833643,14.549335,13.35795,13.932309,14.372104,13.289026,13.321847,14.454155,14.037334,12.937847,11.720206,11.221334,11.286975,10.788103,10.765129,9.193027,8.41518,9.094564,10.194052,10.387693,9.485129,8.149334,6.99077,6.5772314,6.73477,7.003898,6.7840004,5.8814363,4.4996924,5.0871797,4.565334,3.2525132,2.1431797,2.8980515,3.889231,4.601436,5.2676926,5.85518,6.088206,5.3070774,6.567385,7.860513,8.457847,8.910769,9.458873,9.990565,9.373539,7.4863596,5.2020516,5.1922054,5.674667,6.0028725,6.1997952,6.957949,6.7150774,6.764308,7.384616,8.52677,9.796924,12.018872,14.020925,14.78236,14.303181,13.594257,13.499078,12.685129,10.965334,9.170052,9.170052,7.0104623,6.514872,5.8125134,4.841026,5.3398976,3.5347695,2.3401027,1.723077,1.4112822,0.88615394,0.6301539,1.3522053,2.4320002,3.1048207,2.4582565,8.034462,6.875898,4.709744,3.7251284,2.5796926,6.058667,9.370257,8.218257,3.8629746,3.1442053,7.768616,5.8781543,3.698872,4.450462,8.329846,6.3540516,6.052103,6.422975,6.8693337,7.1876926,5.85518,4.634257,4.0992823,4.345436,5.0051284,4.322462,4.71959,4.9132314,4.630975,4.6080003,5.402257,5.179077,4.6834874,4.240411,3.754667,3.570872,4.4865646,5.3727183,5.901129,6.560821,6.7314878,6.7577443,6.738052,6.8496413,7.325539,7.77518,7.522462,7.259898,7.3321033,7.7357955,7.9327188,7.578257,7.3747697,7.453539,7.3550773,8.172308,9.199591,9.82318,9.829744,9.416205,9.3768215,9.468719,9.504821,9.4457445,9.383386,8.3823595,8.188719,8.077128,7.716103,7.141744,6.1538467,5.7764106,5.2512827,4.4964104,4.1058464,4.2994876,4.1485133,4.066462,4.1452312,4.1189747,4.522667,4.5587697,4.3716927,4.20759,4.4406157,3.879385,3.4560003,3.4592824,3.7907696,3.9351797,4.240411,4.44718,4.6178465,4.5817437,3.9220517,3.5905645,3.4166157,3.1442053,2.8422565,2.9144619,3.1343591,3.3345644,3.4133337,3.4231799,3.570872,3.4002054,3.1376412,2.9472823,2.7733335,2.3335385,2.2744617,2.605949,2.7044106,2.412308,2.044718,1.9593848,2.4976413,2.8980515,2.92759,2.8521028,3.4133337,3.0227695,2.6289232,2.8882053,4.1813335,5.2414365,5.041231,4.699898,4.6933336,4.850872,4.522667,4.5587697,4.6080003,4.7622566,5.5696416,5.9963083,5.4908724,4.768821,4.325744,4.4110775,4.532513,4.5817437,4.818052,5.1659493,5.2020516,5.618872,6.0619493,6.12759,5.681231,4.850872,4.069744,4.2863593,4.9460516,5.5302567,5.5532312,7.958975,7.499488,5.98318,5.0609236,6.196513,13.761642,12.048411,7.8014364,4.9493337,4.6080003,9.380103,8.057437,5.297231,3.7415388,3.9975388,1.9593848,1.8445129,2.4582565,2.9243078,2.6551797,2.300718,1.8740515,1.8313848,2.103795,2.0906668,2.359795,2.1530259,1.8937438,1.8970258,2.349949,3.1081028,4.020513,4.57518,4.6276927,4.394667,3.8564105,3.2820516,2.7700515,2.3729234,2.1070771,1.8609232,2.605949,3.2656412,3.239385,2.3958976,2.4582565,2.4155898,2.3991797,2.3729234,2.166154,1.6311796,1.339077,1.332513,1.4867693,1.5097437,1.975795,3.062154,3.9384618,5.0871797,8.283898,4.9526157,3.7907696,3.8137438,4.420923,5.3858466,4.568616,4.017231,4.023795,4.384821,4.4110775,5.1659493,4.9788723,4.6145644,4.5029745,4.7458467,5.037949,5.110154,5.2578464,4.9362054,2.7766156,9.065026,9.6754875,8.228104,7.2992826,8.421744,14.989129,21.704206,24.247797,30.903797,62.546055,74.10544,42.023388,12.232206,2.6223593,3.0358977,2.8291285,3.242667,3.446154,3.3575387,3.6627696,4.4800005,3.5577438,3.8498464,5.5269747,5.9667697,5.074052,4.7425647,4.699898,4.850872,5.280821,4.4373336,3.7316926,2.9571285,2.1956925,1.8149745,1.7920002,1.8576412,1.7165129,1.3850257,1.1913847,1.3981539,1.8248206,2.3072822,2.7864618,3.31159,3.5052311,3.2623591,3.3772311,3.7349746,3.2951798,3.3312824,2.8553848,2.5764105,2.7076926,2.9768207,2.4746668,2.3040001,2.2121027,1.9528207,1.2832822,1.6344616,2.2547693,2.9440002,3.370667,3.0523078,3.1737437,2.9210258,2.7142565,2.6486156,2.5009232,2.4418464,2.9111798,3.2032824,3.3575387,4.1517954,3.8465643,3.43959,3.4034874,3.9680004,5.1265645,5.297231,4.9460516,4.240411,3.6529233,3.9811285,3.7021542,3.31159,3.4133337,4.010667,4.4865646,4.585026,4.4242053,4.388103,4.6605134,5.2348723,5.2348723,5.5532312,5.7074876,5.609026,5.586052,5.671385,6.058667,5.910975,5.330052,5.356308,5.7107697,5.2578464,4.781949,4.637539,4.7622566,4.8082056,5.225026,5.1331286,4.568616,4.4701543,5.093744,5.156103,5.034667,5.0510774,5.477744,4.7458467,4.709744,4.5817437,4.2436924,4.2568207,5.284103,4.972308,4.6539493,4.893539,5.477744,5.76,5.2611284,4.7622566,4.673641,5.0642056,5.113436,4.6244106,4.2272825,4.1091285,4.013949,3.8432825,2.9768207,2.1956925,1.8576412,1.9068719,1.7985642,2.172718,2.428718,2.4976413,2.8389745,2.7634873,2.9571285,2.8521028,2.5206156,2.6551797,2.8488207,2.6978464,2.5140514,2.3696413,2.0742567,5.1987696,5.658257,6.1078978,5.927385,5.4416413,5.920821,6.62318,7.3452315,8.077128,8.493949,7.936001,7.512616,7.059693,6.5837955,6.2227697,6.2162056,6.3934364,7.0104623,7.4765134,7.5881033,7.512616,7.2664623,6.8693337,6.445949,5.943795,5.1364107,4.7983594,4.525949,4.2962055,4.141949,4.1517954,4.0041027,4.2896414,4.923077,5.428513,4.9362054,5.2578464,5.671385,6.042257,6.3934364,6.9021544,6.3967185,6.76759,7.069539,7.1056414,7.430565,7.3616414,7.4896417,7.6274877,7.6242056,7.3649235,6.931693,6.5247183,6.0324106,5.4580517,4.919795,5.106872,6.0028725,6.8365135,7.24677,7.2664623,6.2752824,5.4974365,5.1987696,5.356308,5.648411,6.160411,6.747898,7.1056414,7.177847,7.1844106,6.432821,6.4065647,6.514872,6.554257,6.692103,6.3474874,5.435077,5.0609236,5.543385,6.416411,7.020308,7.6701546,8.707283,9.77395,9.826463,9.127385,8.533334,7.8670774,7.1844106,6.764308,6.3967185,6.9743595,7.525744,7.8080006,8.303591,8.490667,9.833026,12.619488,15.82277,17.08636,18.034874,16.705643,15.747283,15.904821,16.039387,8.467693,4.023795,1.5064616,0.23630771,0.059076928,0.15753847,0.32164106,0.42994875,0.47589746,0.54482055,0.8008206,1.1749744,0.86646163,0.08533334,0.036102567,0.026256412,0.009846155,0.009846155,0.029538464,0.059076928,0.39712822,0.58420515,0.73517954,0.86646163,0.92225647,1.1060513,1.1716924,1.3357949,1.591795,1.6935385,1.6016412,1.7788719,1.9922053,2.1333334,2.228513,2.550154,2.865231,3.239385,3.5774362,3.6562054,3.8498464,3.4756925,3.0030773,2.7470772,2.8717952,3.2656412,3.117949,2.9505644,3.0523078,3.4921029,3.5905645,4.460308,5.287385,5.5597954,5.0510774,4.788513,5.1200004,5.9963083,7.253334,8.602257,9.993847,12.347078,14.076719,14.598565,14.322873,13.574565,12.786873,12.570257,12.813129,12.678565,13.906053,14.700309,14.959591,15.159796,16.344616,16.968206,16.357744,15.816206,15.432206,14.063591,13.8075905,14.555899,15.688207,16.846771,17.93641,18.576412,18.294155,17.611488,17.063385,17.178257,17.204514,17.257027,17.283283,17.171694,16.7319,16.091898,15.983591,16.338053,16.768002,16.577642,18.582975,20.329027,21.221745,20.97231,19.61354,20.555489,22.104616,23.18113,23.138464,21.77313,18.924309,18.22195,18.261335,18.018463,16.869745,17.289848,16.823795,15.484719,14.168616,14.6642065,14.713437,14.326155,13.833847,13.4859495,13.453129,13.115078,11.874462,10.866873,10.620719,11.057232,12.182976,10.834052,9.357129,8.887795,9.363693,9.77395,9.524513,8.635077,7.4732313,6.73477,6.5017443,6.557539,6.426257,5.7764106,4.414359,4.778667,4.6178465,3.4494362,2.0775387,2.5698464,3.0326157,4.322462,5.4416413,5.976616,6.1013336,6.675693,7.719385,8.477539,8.743385,8.861539,10.154668,10.108719,9.078155,7.4732313,5.7764106,5.930667,6.2194877,6.452513,6.7840004,7.7259493,8.516924,8.421744,8.044309,7.975385,8.795898,11.503591,14.040616,15.202463,15.159796,15.43877,13.817437,13.00677,11.82195,10.033232,8.36595,6.6527185,6.1407185,5.8092313,5.1659493,4.2305646,3.8695388,2.6847181,1.8379488,1.5786668,1.2406155,1.020718,1.3883078,2.2547693,2.986667,2.409026,4.010667,3.8137438,4.089436,5.1265645,5.2381544,5.937231,8.011488,8.2215395,6.73477,7.1483083,6.2162056,4.699898,4.059898,4.6276927,5.609026,6.1505647,5.8256416,5.5991797,6.052103,7.394462,6.806975,6.114462,5.5696416,5.182359,4.7491283,5.618872,4.6802053,3.9351797,4.197744,5.1200004,4.955898,4.818052,4.4898467,4.023795,3.7284105,3.3805132,3.8301542,4.6080003,5.4514875,6.3179493,6.4689236,7.059693,7.207385,6.944821,7.213949,7.4010262,7.522462,7.4896417,7.394462,7.50277,7.269744,7.1614366,7.2894363,7.5881033,7.781744,8.776206,10.010257,10.420513,10.033232,9.938052,10.148104,9.905231,9.393231,8.828718,8.457847,8.139488,8.113232,8.1755905,8.12636,7.77518,6.7085133,5.927385,5.1265645,4.33559,3.8859491,4.3716927,4.519385,4.325744,3.9811285,3.889231,3.4133337,3.5282054,3.754667,3.8334363,3.7316926,3.6496413,3.754667,4.1550775,4.7261543,5.110154,4.818052,4.844308,4.7524104,4.4373336,4.128821,3.7316926,3.4297438,3.1442053,2.9013336,2.8291285,3.2623591,3.2984617,3.186872,3.0884104,3.0687182,2.8127182,2.8258464,2.8488207,2.7995899,2.809436,2.9144619,3.0391798,3.05559,2.9013336,2.5928206,2.048,2.281026,2.5271797,2.5107694,2.4385643,2.9801028,2.8849232,3.1540515,3.9745643,4.7294364,4.8147697,4.5390773,4.312616,4.3552823,4.6802053,4.6539493,4.5390773,4.6769233,5.297231,6.521436,6.422975,5.8945646,4.9952826,4.1583595,4.164923,4.2568207,4.1911798,4.5390773,5.031385,4.519385,4.6900516,5.225026,5.6287184,5.76,5.8289237,4.8607183,5.0609236,5.362872,5.3431797,5.211898,6.173539,7.3419495,7.3649235,5.861744,3.4231799,4.5390773,5.2381544,4.6211286,3.748103,5.6320004,5.1331286,4.138667,3.446154,3.0391798,2.1070771,1.9232821,2.4320002,2.9111798,2.9702566,2.5435898,2.1825643,2.03159,2.1956925,2.5337439,2.6289232,3.0227695,2.612513,2.297436,2.4713848,3.0227695,3.7087183,5.287385,5.914257,5.277539,4.578462,4.5489235,4.056616,3.2951798,2.553436,2.2153847,2.3926156,2.733949,3.0818465,3.2032824,2.809436,2.3433847,2.0250258,1.9068719,1.8642052,1.6180514,1.7066668,1.7099489,1.7920002,2.0118976,2.3269746,3.3280003,3.0785644,3.1409233,4.493129,7.515898,4.9460516,3.3641028,3.0916924,3.7809234,4.4340515,4.59159,4.644103,4.6112823,4.535795,4.4832826,4.850872,5.4449234,5.5663595,5.330052,5.674667,4.8738465,4.33559,4.453744,4.598154,3.131077,4.3585644,4.4964104,4.4996924,4.9526157,6.0685134,9.101129,14.834873,18.176,22.692104,40.621952,51.22626,27.050669,6.229334,2.1825643,3.5741541,2.9669745,3.692308,4.0303593,4.0533338,5.6287184,4.7655387,3.8400004,3.945026,5.044513,5.989744,5.549949,4.962462,4.699898,4.8377438,5.0609236,4.384821,3.7874875,3.255795,2.7766156,2.3401027,2.228513,2.03159,1.8215386,1.7001027,1.7887181,1.7033848,1.9528207,2.162872,2.359795,2.9801028,3.4297438,3.0654361,2.8422565,2.8914874,2.540308,2.7503593,2.612513,2.428718,2.4451284,2.8422565,2.612513,2.2777438,2.048,1.9200002,1.6607181,1.8773335,2.1464617,2.6387694,3.062154,2.6847181,2.740513,2.5271797,2.422154,2.5304618,2.6978464,2.7044106,2.8914874,3.2000003,3.4625645,3.4067695,3.0720003,2.665026,2.681436,3.3608208,4.6769233,5.139693,5.4186673,4.896821,3.8695388,3.5544617,3.6168208,3.56759,3.7021542,4.0303593,4.3027697,4.4406157,4.466872,4.6605134,5.225026,6.308103,5.605744,5.1922054,5.169231,5.47118,5.865026,5.549949,5.5958977,5.405539,5.0642056,5.330052,5.6451287,5.425231,5.110154,5.031385,5.408821,4.9394875,5.4153852,5.917539,5.973334,5.533539,5.920821,5.6320004,5.2381544,5.208616,5.930667,5.2644105,5.024821,4.46359,3.8006158,4.2338467,4.778667,4.4800005,4.6112823,5.3202057,5.612308,5.149539,5.3694363,5.7698464,6.0192823,5.933949,5.2381544,4.6211286,4.1222568,3.8104618,3.7809234,3.249231,3.0096412,2.9407182,2.8488207,2.4582565,1.6049232,1.7591796,1.9889232,2.0906668,2.5698464,2.4582565,2.4352822,2.477949,2.6453335,3.0818465,3.3641028,2.9997952,2.6354873,2.4910772,2.3433847,5.586052,5.7009234,5.920821,6.183385,6.5280004,7.0957956,7.282872,7.3747697,7.433847,7.394462,7.0892315,7.397744,7.030154,6.514872,6.2096415,6.301539,6.2490263,6.518154,7.128616,7.830975,8.096821,7.7948723,7.1647186,6.6560006,6.2030773,5.2381544,5.1232824,5.142975,4.7556925,4.161641,4.312616,4.1780515,4.20759,4.571898,5.100308,5.284103,5.543385,5.464616,5.579488,6.0685134,6.7544622,6.5247183,6.8004107,6.885744,6.672411,6.6428723,6.3442054,6.193231,6.2162056,6.311385,6.265436,6.157129,6.012718,5.76,5.4482055,5.2644105,5.5762057,6.3868723,7.3058467,8.169026,9.009232,7.3714876,6.042257,5.293949,5.080616,5.0674877,5.540103,6.2063594,6.7314878,7.00718,7.1548724,6.8496413,6.7938466,6.744616,6.675693,6.7840004,6.340924,5.5565133,5.093744,5.2709746,6.048821,6.8430777,7.6603084,8.43159,8.900924,8.63836,7.6274877,7.0859494,6.4689236,5.799385,5.664821,5.2578464,5.6320004,5.8814363,5.979898,6.764308,7.1548724,9.31118,12.11077,14.683899,16.393847,17.056822,15.904821,16.827078,18.901335,16.370872,9.193027,4.2535386,1.782154,1.2570257,1.4178462,0.83035904,0.51856416,0.7811283,1.6902566,3.0851285,4.007385,3.8301542,2.300718,0.3708718,0.17723078,0.14769232,0.08861539,0.036102567,0.07548718,0.34789747,0.49887183,0.46276927,0.45292312,0.4955898,0.45620516,0.4955898,0.90584624,1.270154,1.404718,1.3423591,1.463795,1.5721027,1.8379488,2.1300514,2.0184617,2.3696413,2.553436,2.9604106,3.4264617,3.255795,3.7382567,3.5216413,3.0785644,2.7798977,2.8980515,2.9997952,2.9768207,2.989949,3.0752823,3.1540515,3.4166157,4.082872,4.532513,4.5554876,4.348718,4.381539,5.097026,6.2227697,7.640616,9.38995,10.948924,12.4685135,13.190565,13.144616,13.161027,12.688411,11.913847,11.625027,11.871181,11.9860525,12.727796,13.991385,14.8480015,15.268104,16.141129,16.472616,16.328207,15.986873,15.37313,14.066873,13.98154,14.63795,15.993437,17.851078,19.859694,19.984411,18.97354,17.473642,16.370872,16.774565,17.509745,17.93641,17.795284,17.115898,16.233027,15.16636,14.923489,15.327181,15.82277,15.471591,16.082052,17.621334,19.305027,20.319181,19.833437,20.155079,21.238155,22.344208,22.678976,21.382566,17.910154,17.273438,17.716515,17.808413,16.426668,16.866463,16.850052,15.908104,14.697027,15.012104,14.605129,14.41477,14.043899,13.5778475,13.617231,13.6008215,12.314258,10.896411,10.236719,10.95877,12.763899,12.484924,11.474052,10.614155,10.31877,9.412924,9.373539,9.127385,8.310155,7.27959,6.6494365,6.370462,6.1505647,5.671385,4.594872,3.9548721,3.7152824,3.114667,2.3663592,2.6715899,2.7208207,3.6890259,4.926359,5.927385,6.3310776,6.675693,7.2960005,7.965539,8.461129,8.585847,10.06277,10.000411,9.386667,8.438154,6.5805135,6.232616,6.180103,6.5772314,7.2960005,7.9097443,9.068309,9.170052,8.687591,8.385642,9.304616,10.86359,12.557129,14.660924,16.672821,17.335796,13.351386,12.301129,12.166565,11.18195,7.8441033,6.99077,6.311385,5.924103,5.612308,4.8311796,4.194462,3.0194874,2.1333334,1.7591796,1.5097437,1.273436,1.3522053,1.8642052,2.5173335,2.605949,3.0129232,3.7284105,4.7261543,5.605744,5.5926156,7.2270775,7.8769236,7.7456417,7.748924,9.485129,7.276308,4.4865646,3.314872,4.089436,5.277539,5.4514875,5.477744,5.7074876,6.2523084,6.9809237,8.41518,7.821129,6.629744,5.648411,5.0510774,5.7796926,5.3858466,4.8147697,4.673641,5.211898,4.903385,5.142975,4.962462,4.352,4.263385,4.020513,4.2830772,4.775385,5.2315903,5.421949,5.8190775,6.4590774,6.6461544,6.419693,6.5739493,6.5772314,6.76759,6.770872,6.62318,6.76759,6.8233852,6.8988724,6.9842057,7.1581545,7.5946674,8.464411,9.42277,9.616411,9.229129,9.465437,9.888822,9.67877,9.088,8.4053335,7.9327188,8.260923,8.303591,8.021334,7.496206,6.954667,6.088206,5.284103,4.601436,4.1189747,3.9384618,4.06318,4.197744,4.059898,3.7251284,3.636513,3.498667,3.6660516,3.8564105,3.9056413,3.764513,4.2207184,5.028103,5.477744,5.467898,5.5204105,4.781949,4.562052,4.276513,3.8662567,3.7874875,3.636513,3.446154,3.3050258,3.2065644,3.045744,3.314872,3.242667,3.1015387,3.0162053,2.9636924,2.806154,2.7536411,2.6322052,2.4976413,2.6190772,2.8455386,3.0326157,3.0326157,2.7864618,2.3204105,1.8346668,2.1825643,2.477949,2.5271797,2.8291285,3.249231,3.3017437,3.7152824,4.4800005,4.8771286,4.571898,4.529231,4.332308,3.9680004,3.8432825,4.493129,4.417641,4.2601027,4.588308,5.8912826,6.301539,5.8486156,5.2611284,4.9394875,4.919795,5.0642056,4.7556925,4.8836927,5.2545643,4.578462,4.4012313,4.97559,5.405539,5.536821,5.9536414,5.3727183,5.0018463,4.857436,5.0051284,5.540103,5.976616,6.5903597,7.0367184,6.8562055,5.4875903,4.7524104,6.4689236,6.498462,4.821334,5.543385,4.388103,3.8071797,3.045744,2.0841026,1.6508719,2.481231,3.114667,3.5511796,3.629949,3.0227695,2.6026669,2.5238976,2.7142565,2.917744,2.678154,3.114667,2.7044106,2.4713848,2.986667,4.388103,4.634257,5.920821,6.3868723,5.756718,5.3202057,5.1298466,4.706462,3.9154875,2.9997952,2.5731285,2.6551797,2.878359,3.0358977,3.0326157,2.878359,2.3302567,2.0053334,2.0086155,2.1103592,1.7460514,2.0545642,2.0906668,2.2908719,2.7273848,3.1081028,3.7973337,3.6332312,3.6069746,4.1911798,5.346462,4.6933336,3.5314875,3.4658465,4.273231,3.892513,3.8728209,3.945026,3.9712822,4.076308,4.637539,4.4964104,5.1200004,5.5532312,5.5663595,5.6385646,5.225026,4.4307694,4.332308,4.604718,3.5216413,3.6824617,3.0851285,2.7733335,3.2000003,4.2240005,6.9809237,10.502565,13.705847,17.371899,24.146053,25.823181,13.958565,4.965744,3.6004105,2.9669745,4.273231,4.821334,4.276513,3.82359,6.1538467,6.6592827,7.253334,6.6592827,5.7107697,7.3321033,6.432821,5.4153852,5.044513,5.2020516,4.8672824,4.378257,3.7907696,3.2656412,2.9013336,2.7175386,2.5862565,2.2383592,1.8773335,1.8182565,2.5042052,2.103795,2.1464617,2.2711797,2.3466668,2.487795,2.868513,2.5337439,2.3171284,2.3958976,2.284308,2.300718,2.3729234,2.294154,2.1924105,2.5238976,2.612513,2.225231,1.8674873,1.782154,1.9462565,2.028308,2.162872,2.422154,2.6847181,2.6322052,2.425436,2.6354873,2.8225644,2.8816411,3.0391798,3.1081028,3.0851285,3.2820516,3.56759,3.3936412,3.1474874,2.9669745,2.8553848,3.1442053,4.5062566,5.0215387,5.3924108,5.156103,4.31918,3.367385,3.6004105,3.9286156,4.2305646,4.394667,4.322462,4.4077954,4.9460516,5.5204105,5.9995904,6.51159,6.0356927,5.146257,4.6605134,4.8804107,5.579488,5.786257,5.671385,5.4383593,5.330052,5.6352825,5.7501545,5.651693,5.549949,5.5171285,5.4875903,4.9394875,5.2480006,5.8289237,5.973334,4.818052,5.7403083,5.146257,4.4734364,4.6145644,5.914257,4.7983594,4.585026,4.4373336,4.2436924,4.6211286,4.453744,4.6211286,5.284103,5.933949,5.3727183,4.857436,5.3037953,5.8847184,6.170257,6.1308722,5.3037953,4.601436,4.092718,3.7940516,3.6496413,3.2984617,3.117949,3.0523078,3.0916924,3.2722054,2.2482052,2.0250258,2.0053334,1.975795,2.1103592,2.0020514,1.9790771,2.2514873,2.7963078,3.3444104,3.446154,3.1507695,2.865231,2.7634873,2.7766156,5.7074876,5.618872,6.055385,6.6560006,7.2664623,7.9261546,7.860513,7.653744,7.2369237,6.75118,6.557539,6.8266673,6.7150774,6.4656415,6.2687182,6.265436,6.449231,6.442667,6.8496413,7.64718,8.155898,7.9130263,7.3714876,6.987488,6.619898,5.5302567,5.182359,5.2020516,4.8705645,4.2994876,4.453744,4.2601027,4.2371287,4.4438977,4.850872,5.330052,5.671385,5.4153852,5.3234878,5.6320004,6.058667,6.669129,6.7807183,6.521436,6.0849237,5.76,5.536821,5.5204105,5.5762057,5.609026,5.5565133,5.4843082,5.72718,5.917539,6.045539,6.4656415,6.5739493,6.9842057,7.8441033,8.946873,9.7214365,8.664616,7.322257,6.2555904,5.684513,5.4974365,5.6451287,5.989744,6.432821,6.8299494,6.9809237,7.0432825,6.9710774,6.7774363,6.5706673,6.564103,6.229334,5.7403083,5.3202057,5.2053337,5.658257,6.3474874,6.885744,7.2861543,7.4010262,6.925129,6.088206,5.579488,5.077334,4.588308,4.460308,4.0008206,4.089436,4.0402055,4.007385,5.0182567,5.786257,8.94359,12.018872,14.188309,16.272411,15.819489,15.812924,18.678156,21.62872,16.676104,10.604308,4.969026,1.8674873,1.3981539,1.6640002,2.612513,2.7831798,2.917744,3.9384618,6.954667,7.6734366,7.3714876,4.5554876,0.69579494,0.23958977,0.190359,0.10502565,0.032820515,0.08205129,0.41025645,0.3446154,0.25928208,0.3052308,0.46276927,0.56123084,0.39712822,0.86646163,1.1355898,1.020718,1.020718,1.4473847,1.5261539,1.7362052,1.9856411,1.6213335,2.2514873,2.681436,3.05559,3.2754874,3.006359,3.2032824,3.186872,2.9735386,2.793026,3.058872,2.8488207,2.989949,3.2525132,3.4527183,3.4297438,3.9023592,4.194462,4.2535386,4.1682053,4.1714873,4.568616,5.5926156,6.8233852,8.208411,10.092308,11.441232,12.163283,12.245335,12.012309,12.107488,11.926975,11.30995,10.834052,10.712616,10.778257,11.621744,13.610668,15.415796,16.275694,16.006565,15.937642,15.911386,15.737437,15.254975,14.316309,14.720001,15.07118,16.114874,17.992207,20.22072,20.197744,19.222977,17.660719,16.370872,16.70236,17.831387,18.359797,18.011898,16.827078,15.133539,14.244103,13.801026,13.869949,14.290052,14.641232,14.6182575,15.317334,16.659693,18.080822,18.520617,18.668308,19.941746,21.169233,21.35959,19.72513,17.010874,16.607182,17.398155,18.162872,17.588514,17.624617,17.283283,16.630156,15.944206,15.707899,15.366566,14.880821,14.431181,14.093129,13.843694,13.984821,12.918155,11.602052,10.95877,11.867898,13.607386,14.54277,14.043899,12.491488,11.277129,9.852718,9.380103,9.278359,8.966565,7.8769236,7.0990777,6.36718,5.901129,5.5204105,4.637539,3.387077,3.0391798,2.802872,2.5304618,2.7306669,2.6617439,3.058872,4.1747694,5.6418467,6.4722056,6.518154,6.925129,7.788308,8.6580515,8.54318,9.885539,9.96759,9.649232,8.94359,6.987488,6.5247183,6.5411286,7.1056414,7.8670774,8.064001,9.4457445,9.869129,9.452309,8.94359,9.737847,10.364718,11.316514,13.571283,16.341335,17.073233,13.312001,12.012309,12.028719,11.562668,8.152616,7.466667,6.62318,6.3310776,6.370462,5.5762057,4.4800005,3.7284105,2.8455386,1.9167181,1.5655385,1.4605129,1.9462565,2.2186668,2.2908719,2.9965131,3.1081028,3.9384618,5.100308,6.042257,6.045539,6.3277955,6.3179493,6.242462,6.701949,8.674462,6.816821,4.197744,3.1507695,4.0402055,5.277539,5.2414365,5.5893335,5.85518,5.98318,6.3212314,8.362667,7.8047185,6.4557953,5.47118,5.362872,5.5597954,5.586052,5.3202057,4.84759,4.493129,4.7261543,5.106872,5.0018463,4.601436,4.923077,4.6211286,4.673641,4.890257,5.0116925,4.716308,5.037949,5.5171285,5.7435904,5.7140517,5.835488,5.654975,5.7042055,5.668103,5.618872,5.9930263,6.705231,6.918565,6.8693337,6.9120007,7.5421543,8.2445135,8.67118,8.681026,8.539898,8.930462,9.078155,8.874667,8.4512825,7.962257,7.5946674,7.6603084,7.515898,6.9776416,6.189949,5.618872,4.9952826,4.457026,4.056616,3.8629746,3.9581542,3.9778464,4.017231,3.882667,3.639795,3.620103,3.817026,3.9548721,4.1747694,4.4373336,4.516103,5.156103,6.449231,6.9120007,6.2916927,5.5565133,4.670359,4.2601027,3.9089234,3.5840003,3.6332312,3.6529233,3.620103,3.6168208,3.5774362,3.2951798,3.2820516,3.0785644,2.8914874,2.8160002,2.8521028,2.8521028,2.8225644,2.678154,2.550154,2.789744,2.9243078,3.1442053,3.062154,2.5731285,1.8871796,1.5819489,1.9495386,2.349949,2.605949,3.0194874,3.1507695,3.31159,3.7382567,4.315898,4.588308,4.5029745,4.7425647,4.460308,3.636513,3.0424619,3.895795,4.1222568,3.9614363,3.9811285,5.077334,6.0717955,5.7698464,5.5105643,5.5565133,5.077334,5.1298466,4.9460516,5.0871797,5.3891287,4.969026,4.5095387,5.034667,5.5532312,5.7074876,5.7764106,5.937231,5.3234878,4.6867695,4.6244106,5.5762057,6.3343596,6.4754877,6.7577443,7.2336416,7.256616,6.7216415,7.958975,7.4765134,5.3727183,5.3169236,5.3169236,4.6178465,3.1638978,1.7624617,2.0611284,3.255795,3.7940516,4.0467696,4.0303593,3.4133337,3.0785644,3.006359,3.3017437,3.5840003,2.9735386,3.1967182,2.809436,2.678154,3.370667,5.1265645,5.349744,6.2916927,6.550975,6.0324106,5.937231,5.61559,5.110154,4.384821,3.5905645,3.0654361,2.8488207,3.0391798,3.1934361,3.1540515,3.0358977,2.7175386,2.425436,2.3729234,2.4681027,2.3072822,2.7241027,2.6518977,2.809436,3.3247182,3.7251284,3.7448208,3.748103,3.7021542,3.8006158,4.466872,4.197744,3.6726158,3.9942567,4.8082056,4.332308,4.20759,4.135385,4.017231,4.082872,4.900103,4.6178465,5.028103,5.431795,5.5269747,5.4153852,5.609026,5.0051284,4.6112823,4.6178465,4.4077954,4.1222568,2.986667,2.097231,2.1366155,3.373949,6.498462,8.917334,11.405129,13.722258,14.6182575,11.47077,13.197129,13.37436,9.432616,2.6683078,7.2205133,7.276308,5.717334,4.8016415,6.1538467,7.4240007,9.537642,8.845129,6.4689236,8.329846,6.5378466,6.0028725,6.0028725,5.802667,4.6539493,4.4406157,3.895795,3.3050258,2.9046156,2.8849232,2.7044106,2.3466668,1.910154,1.7788719,2.6289232,2.231795,2.1891284,2.353231,2.4320002,1.975795,2.1989746,2.0841026,1.9561027,1.9790771,2.1267693,2.0644104,2.2383592,2.2482052,2.0644104,2.028308,2.2186668,2.0250258,1.8018463,1.7460514,1.9298463,1.9495386,2.1169233,2.1366155,2.1267693,2.5993848,2.5074873,2.806154,3.0030773,2.993231,3.0523078,3.0260515,3.1770258,3.4100516,3.564308,3.4067695,3.1934361,3.259077,3.1967182,3.255795,4.3290257,4.7589746,5.2480006,5.297231,4.7524104,3.8301542,3.889231,4.2371287,4.5062566,4.585026,4.644103,4.9526157,5.671385,6.2851286,6.557539,6.5444107,6.4656415,5.609026,5.0051284,5.080616,5.6320004,6.0619493,5.8945646,5.6320004,5.546667,5.6976414,5.58277,5.612308,5.658257,5.605744,5.353026,5.353026,5.609026,5.9470773,5.917539,4.781949,5.3103595,4.2207184,3.7710772,4.601436,5.720616,4.5095387,4.588308,4.673641,4.4242053,4.414359,4.076308,4.9460516,5.9634876,6.226052,4.962462,4.9788723,5.543385,5.924103,5.901129,5.7632823,5.2578464,4.775385,4.2568207,3.767795,3.498667,3.318154,3.1540515,3.0654361,3.1245131,3.442872,2.737231,2.5304618,2.5009232,2.422154,2.156308,1.8346668,1.6443079,1.8707694,2.4910772,3.186872,3.1343591,3.1015387,3.0752823,3.1015387,3.2722054,5.4974365,5.602462,6.3442054,6.9776416,7.4404106,8.316719,8.297027,8.2904625,7.817847,7.0104623,6.6034875,6.308103,6.449231,6.554257,6.4590774,6.3310776,6.8627696,6.8660517,6.8955903,7.174565,7.5913854,7.50277,7.325539,7.066257,6.633026,5.8518977,5.284103,5.1889234,5.024821,4.6933336,4.5423594,4.128821,4.210872,4.391385,4.59159,5.0576415,5.5236926,5.622154,5.5630774,5.4580517,5.3431797,6.521436,6.436103,6.052103,5.7829747,5.5007186,5.4974365,5.7534366,5.970052,6.0783596,6.262154,6.1341543,6.432821,6.7938466,7.177847,7.90318,7.653744,7.7292314,8.477539,9.4916935,9.639385,9.869129,9.019077,7.899898,7.0957956,6.9776416,6.7872825,6.5706673,6.669129,7.0367184,7.204103,7.3091288,7.2369237,6.9645133,6.5706673,6.2490263,5.976616,5.533539,5.1265645,4.955898,5.2020516,5.543385,5.431795,5.353026,5.3037953,4.7983594,4.4274874,3.9745643,3.6135387,3.3936412,3.2295387,2.8947694,2.7864618,2.605949,2.6026669,3.5478978,4.2535386,7.972103,11.480617,13.692719,15.688207,14.080001,15.852309,19.232822,20.883694,15.898257,11.625027,5.8289237,1.8018463,0.5349744,0.7056411,4.388103,5.7632823,5.668103,5.865026,9.058462,8.687591,9.842873,6.8430777,0.9321026,0.26584616,0.2297436,0.16738462,0.22646156,0.36102566,0.30851284,0.35446155,0.29538465,0.39056414,0.6662565,0.9321026,0.5546667,0.7844103,0.78769237,0.5677949,0.9714873,1.3751796,1.3193847,1.3981539,1.5688206,1.1684103,2.041436,2.9505644,3.3017437,3.1409233,3.1277952,2.806154,2.8455386,2.806154,2.7503593,3.2295387,3.2262566,3.4494362,3.7809234,4.164923,4.630975,5.1232824,4.8082056,4.5062566,4.535795,4.716308,5.1922054,6.245744,7.381334,8.579283,10.262975,10.840616,11.296822,11.602052,11.74318,11.730052,11.467488,10.794667,10.075898,9.691898,10.036513,11.667693,14.063591,16.311796,17.352207,15.9573345,15.382976,14.851283,14.562463,14.50995,14.519796,15.763694,15.940925,16.41354,17.683693,19.370668,19.140924,18.809437,17.900309,16.754873,16.521847,17.631182,18.281027,18.07754,16.800821,14.418053,14.04718,13.279181,12.675283,12.698257,13.702565,14.04718,14.116103,14.473847,15.353437,16.672821,16.948515,18.527182,19.86954,19.941746,18.20554,16.971489,16.758156,17.59836,18.914463,19.505232,19.009642,18.116924,17.713232,17.703386,17.024002,17.132309,16.049232,15.015386,14.444309,13.929027,14.306462,13.879796,13.128206,12.800001,13.88636,15.041642,16.423386,15.327181,12.278154,11.040821,11.017847,9.93477,9.3768215,9.366975,8.36595,7.6898465,6.6560006,5.933949,5.4514875,4.388103,3.2722054,2.9604106,2.7569232,2.5206156,2.665026,2.5895386,2.6584618,3.623385,5.2480006,6.2851286,6.445949,6.931693,8.060719,9.212719,8.851693,9.970873,10.043077,9.573745,8.720411,7.2960005,7.177847,7.430565,7.8834877,8.280616,8.280616,9.96759,10.768411,10.197334,9.094564,9.619693,10.125129,10.752001,12.294565,14.536206,16.239592,14.171899,12.511181,11.703795,11.122872,9.110975,7.8703594,7.056411,6.994052,7.059693,5.6385646,4.562052,4.2535386,3.4067695,2.0250258,1.4342566,1.972513,3.255795,3.3476925,2.4910772,3.1048207,3.751385,4.0402055,4.7556925,5.8814363,6.5870776,3.9614363,3.9089234,4.309334,4.5423594,5.4843082,4.345436,3.629949,3.889231,4.7917953,5.1265645,5.6943593,5.858462,5.668103,5.395693,5.533539,6.413129,5.8223596,5.097026,4.886975,5.1364107,5.0149746,4.9821544,4.893539,4.5554876,3.7185643,4.384821,4.594872,4.5456414,4.598154,5.2742567,4.6834874,4.450462,4.4406157,4.44718,4.210872,4.2863593,4.6867695,5.0182567,5.169231,5.3202057,4.919795,4.8049235,4.8082056,5.0084105,5.7074876,6.813539,6.928411,6.747898,6.8004107,7.4699492,8.03118,8.1066675,8.041026,8.021334,8.083693,7.571693,7.4010262,7.3058467,7.1483083,6.925129,6.117744,5.861744,5.543385,5.041231,4.7392826,4.332308,4.086154,3.876103,3.748103,3.9056413,4.1780515,4.1583595,3.9384618,3.7382567,3.892513,4.023795,4.0336413,4.3552823,4.9952826,5.504,6.180103,7.3649235,7.643898,6.6822567,5.2381544,4.4898467,4.027077,3.7185643,3.5511796,3.6135387,3.6004105,3.6332312,3.6660516,3.5971284,3.2722054,3.0490258,2.7470772,2.5140514,2.4516926,2.6157951,2.6584618,2.7995899,2.8225644,2.8324106,3.2164104,3.1343591,3.2623591,3.0523078,2.4057438,1.6836925,1.4112822,1.5491283,2.041436,2.6223593,2.8127182,2.7208207,3.0326157,3.4560003,3.8367183,4.161641,4.4800005,4.644103,4.1813335,3.2623591,2.6945643,3.2164104,3.757949,3.8432825,3.7316926,4.4274874,5.7829747,5.8157954,5.8223596,5.8945646,4.919795,4.6834874,4.699898,4.926359,5.225026,5.3694363,4.821334,5.175795,5.8847184,6.3277955,5.8092313,6.373744,6.038975,5.179077,4.535795,5.2315903,6.3540516,6.688821,6.7577443,6.8660517,7.0826674,7.4108725,7.322257,6.1505647,4.71959,5.362872,5.671385,4.4406157,2.9013336,2.0250258,2.5238976,3.8728209,4.2896414,4.240411,3.9614363,3.4724104,3.308308,3.2164104,3.7349746,4.394667,3.7087183,3.4658465,3.1015387,3.058872,3.639795,4.9854364,5.5893335,6.38359,6.4656415,5.989744,6.163693,5.989744,5.280821,4.529231,3.9712822,3.5872824,3.1245131,3.190154,3.4855387,3.7185643,3.5905645,3.639795,3.308308,2.9833848,2.9440002,3.3542566,3.757949,3.4527183,3.367385,3.7415388,4.1189747,3.8465643,3.626667,3.318154,3.4756925,5.349744,3.69559,3.3641028,4.0041027,5.0084105,5.5269747,5.398975,5.1659493,4.7589746,4.44718,4.827898,5.0149746,5.3234878,5.4383593,5.398975,5.586052,5.832206,5.7435904,5.3431797,4.9952826,5.402257,4.1911798,2.9735386,2.2219489,2.3958976,3.948308,6.813539,8.835282,10.217027,11.076924,11.457642,12.1928215,21.717335,24.6679,16.423386,3.121231,11.657847,10.748719,7.899898,6.6560006,6.5837955,7.384616,10.965334,10.712616,7.256616,8.480822,5.664821,6.23918,6.918565,6.235898,4.5128207,4.4274874,4.056616,3.5347695,3.062154,2.92759,2.612513,2.2449234,1.8445129,1.6738462,2.2482052,2.0250258,2.0184617,2.2153847,2.294154,1.6246156,1.7099489,1.8576412,1.7657437,1.5524104,1.7526156,1.8313848,1.9987694,2.0709746,1.9593848,1.654154,1.6607181,1.7788719,1.8149745,1.7460514,1.7033848,1.7887181,2.0512822,1.9298463,1.6968206,2.4582565,2.737231,2.7831798,2.806154,2.861949,2.8389745,2.612513,3.0687182,3.4330258,3.3969233,3.1277952,2.8849232,3.0523078,3.242667,3.4658465,4.1025643,4.2896414,4.9394875,5.1659493,4.8672824,4.7458467,4.378257,4.4373336,4.598154,4.8147697,5.32677,5.9995904,6.432821,6.7183595,6.8397956,6.669129,6.76759,6.3606157,6.055385,6.0685134,6.226052,6.370462,6.1505647,5.8420515,5.618872,5.5696416,5.353026,5.428513,5.5105643,5.5007186,5.464616,6.0061545,6.4689236,6.560821,6.298257,5.976616,5.1659493,3.7448208,3.9253337,5.366154,5.172513,4.519385,5.0116925,4.919795,4.0303593,3.6529233,3.757949,5.179077,6.2523084,6.117744,4.6900516,5.402257,6.0028725,6.0849237,5.6418467,5.077334,5.0543594,4.965744,4.4110775,3.6069746,3.4067695,3.2000003,3.0785644,3.0916924,3.1737437,3.1540515,2.92759,2.9997952,3.0818465,2.9505644,2.4451284,1.9068719,1.5392822,1.4933335,1.8609232,2.674872,2.6354873,2.9078977,3.18359,3.3608208,3.5314875,5.937231,6.0324106,5.920821,6.121026,6.813539,7.827693,8.169026,8.4283085,8.123077,7.2270775,6.163693,5.9569235,6.2884107,6.6560006,6.820103,6.820103,7.026872,7.207385,7.0432825,6.738052,7.020308,6.957949,6.9054365,6.413129,5.805949,6.196513,6.232616,6.294975,5.83877,4.893539,4.089436,4.1747694,4.5456414,4.6178465,4.640821,5.691077,5.6320004,6.009436,6.265436,6.160411,5.7829747,6.442667,6.2588725,6.1440005,6.340924,6.439385,6.5247183,7.177847,7.6176414,7.837539,8.605539,8.39877,8.182155,8.146052,8.369231,8.818872,8.684308,8.769642,9.278359,9.957745,10.115283,10.029949,9.724719,9.133949,8.500513,8.392206,8.086975,7.6996927,7.4240007,7.3747697,7.584821,7.706257,7.581539,7.39118,7.1548724,6.7150774,6.419693,5.579488,4.644103,3.9811285,3.8596926,3.7021542,3.7087183,3.6036925,3.245949,2.6256413,2.3794873,2.3204105,2.4484105,2.605949,2.4713848,2.1169233,1.8281027,1.6705642,1.7788719,2.3663592,2.9505644,6.173539,9.127385,11.122872,13.686155,12.819694,16.41354,17.664001,15.350155,13.824001,10.761847,5.654975,1.7362052,0.33805132,0.8992821,3.5872824,4.962462,5.333334,5.10359,4.7622566,3.636513,8.356103,7.4765134,1.0469744,0.5940513,0.62030774,0.63343596,1.1290257,1.6377437,0.74830776,1.6147693,1.079795,0.45292312,0.27241027,0.32164106,0.39384618,0.8598975,0.94523084,0.78769237,1.4342566,1.020718,0.71548724,0.90256417,1.401436,1.4506668,2.2055387,2.7995899,2.9997952,3.006359,3.4330258,3.4330258,3.1113849,2.8750772,2.861949,2.9604106,3.9253337,4.3749747,4.706462,5.353026,6.803693,6.9645133,5.805949,5.1265645,5.398975,5.7534366,6.0947695,6.8496413,7.6767187,8.749949,10.725744,10.154668,10.650257,11.2672825,11.500309,11.290257,10.023385,9.639385,9.537642,9.878975,11.611898,13.321847,15.110565,16.400412,16.873028,16.49559,15.468308,14.828309,14.027489,13.689437,15.593027,17.7559,18.504206,18.635489,18.760206,19.331284,17.59836,17.375181,17.18154,16.62031,16.387283,17.145437,17.700104,17.969233,17.545847,15.701335,15.835898,14.7331295,13.581129,12.934566,12.724514,12.934566,13.59754,14.037334,14.680616,17.073233,16.561232,16.984617,18.100513,19.134361,18.766771,17.083078,17.578669,18.46154,19.03918,19.698874,19.771078,18.983387,18.471386,18.563284,18.78318,18.83241,17.250463,15.353437,14.112822,14.158771,15.074463,15.698052,15.465027,14.946463,15.839181,16.594053,16.528412,12.553847,7.282872,9.002667,12.199386,11.460924,10.331899,9.892103,8.743385,8.146052,7.5191803,6.816821,5.7796926,3.9351797,3.239385,3.0490258,2.9078977,2.7241027,2.7602053,2.297436,2.5665643,3.6660516,5.0642056,5.5991797,5.733744,6.3442054,7.53559,8.851693,9.278359,10.289231,9.977437,9.212719,8.651488,8.713847,8.503796,8.113232,7.890052,7.9491286,8.195283,10.197334,11.483898,10.505847,8.5202055,9.5835905,10.108719,9.990565,11.119591,14.496821,20.233849,15.642258,13.111795,11.746463,10.817642,9.780514,8.329846,7.9917955,7.6701546,6.7150774,4.9427695,4.138667,3.0851285,2.4155898,2.0676925,1.3128207,3.5216413,4.7524104,4.3552823,2.8717952,2.028308,5.7632823,5.8912826,4.2994876,3.131077,4.7917953,5.1954875,4.4242053,3.692308,3.3608208,2.9440002,3.0194874,3.4034874,4.4767184,5.7632823,5.920821,6.1768208,5.097026,5.290667,6.2785645,4.4701543,4.4340515,3.3280003,3.4921029,4.634257,3.8301542,3.511795,4.194462,4.6867695,4.6933336,4.7917953,4.325744,4.450462,4.594872,4.637539,4.8836927,4.089436,3.7185643,3.387077,3.0752823,3.1113849,3.626667,4.312616,4.8016415,5.024821,5.2348723,4.6112823,4.585026,4.8771286,5.4514875,6.5017443,6.806975,6.232616,5.835488,5.979898,6.3474874,6.6527185,7.1876926,7.273026,6.6560006,5.5072823,4.604718,4.97559,5.4449234,5.4613338,5.080616,4.276513,4.824616,5.349744,5.3727183,5.32677,5.1922054,4.8738465,4.46359,4.1124105,4.027077,4.161641,4.1222568,3.9089234,3.7940516,4.31918,4.4045134,4.1878977,4.194462,4.713026,5.799385,7.177847,7.322257,6.557539,5.333334,4.210872,3.698872,3.3608208,3.1409233,2.989949,2.868513,2.7602053,2.6847181,2.6256413,2.5895386,2.6256413,2.3926156,2.2055387,2.162872,2.2613335,2.3958976,2.176,2.284308,2.3663592,2.3860514,2.6551797,2.5829747,2.5829747,2.412308,2.0742567,1.8313848,1.2931283,1.1585642,1.7624617,2.7044106,2.8389745,3.1081028,3.6758976,3.9089234,3.8465643,4.210872,4.2371287,3.4625645,2.737231,2.5238976,2.9144619,3.2820516,3.5905645,3.4264617,3.0129232,3.2196925,5.113436,5.8781543,6.4032826,6.8365135,6.5903597,6.0061545,5.2447186,4.7327185,4.768821,5.540103,5.1954875,5.221744,5.937231,6.8233852,6.5312824,5.979898,5.9536414,5.7468724,5.3169236,5.280821,5.280821,5.362872,5.717334,6.2884107,6.7905645,8.425026,7.5913854,5.654975,4.2994876,5.5072823,2.7995899,1.4900514,1.3915899,1.9003079,1.9987694,3.95159,4.3290257,4.1550775,3.876103,3.387077,3.1934361,3.006359,3.6529233,4.71959,4.562052,3.7448208,3.5478978,3.6102567,3.9122055,4.7917953,5.366154,5.792821,5.687795,5.431795,6.163693,6.2129235,5.356308,4.240411,3.5478978,4.013949,3.6102567,3.2820516,3.7152824,4.6178465,4.716308,5.044513,4.6244106,4.1517954,4.20759,5.2348723,5.1954875,4.44718,4.023795,4.1682053,4.3027697,5.0838976,4.667077,3.8859491,3.9089234,6.23918,3.6758976,2.349949,3.0818465,5.1856413,6.4557953,5.2348723,4.71959,4.322462,3.8498464,3.508513,4.7917953,5.277539,5.1922054,5.2348723,6.5772314,5.989744,6.413129,6.931693,6.76759,5.280821,3.8137438,3.045744,3.6069746,5.146257,6.3179493,8.379078,7.5585647,7.456821,9.3078985,11.992617,22.465643,22.971079,20.30277,15.488001,3.767795,16.807386,13.968411,8.402052,6.6067696,8.438154,9.95118,16.33477,15.845745,8.979693,8.467693,4.598154,5.2512827,6.242462,5.8190775,4.6834874,4.06318,4.023795,3.945026,3.5872824,3.0982566,2.5009232,1.8642052,1.5163078,1.6377437,2.2744617,1.7362052,1.7493335,1.7296412,1.5753847,1.6475899,1.5885129,1.7263591,1.6114873,1.214359,0.94523084,1.0929232,1.1027694,1.2307693,1.5556924,1.9823592,1.6771283,1.8116925,1.7329233,1.4572309,1.6771283,1.9593848,2.2482052,2.281026,2.1267693,2.2121027,2.3466668,2.5074873,2.8488207,3.2032824,3.0818465,2.789744,2.8980515,3.0752823,3.05559,2.6387694,2.4582565,2.4746668,2.806154,3.3936412,4.027077,3.698872,4.0008206,4.1714873,4.2929235,5.293949,4.6244106,4.5554876,5.142975,6.012718,6.377026,6.951385,6.994052,7.062975,7.1548724,6.7282057,6.741334,6.770872,6.685539,6.5903597,6.8365135,7.020308,6.5969234,6.1472826,5.937231,5.937231,5.924103,5.654975,5.684513,6.0750775,6.3934364,6.0258465,6.8594875,7.1581545,6.7577443,7.0498466,5.6451287,4.9821544,5.4908724,5.979898,3.6463592,3.892513,4.601436,4.4865646,3.6168208,3.4330258,3.9581542,5.1987696,6.058667,5.98318,4.95918,5.789539,6.0160003,5.904411,5.467898,4.457026,4.6276927,4.594872,4.0402055,3.3575387,3.6627696,3.4166157,2.9735386,2.8324106,3.1442053,3.692308,3.5216413,3.3247182,2.934154,2.3466668,1.723077,1.6738462,1.8084104,1.7493335,1.6508719,2.2121027,2.297436,2.740513,3.1803079,3.3476925,3.0654361,7.315693,7.207385,7.0793853,7.056411,7.2894363,7.962257,8.3823595,8.874667,8.825437,8.1066675,7.0432825,6.875898,6.806975,7.003898,7.3583593,7.50277,7.273026,7.0498466,6.7905645,6.5345645,6.38359,6.6560006,6.8397956,6.688821,6.2523084,5.8912826,5.858462,5.7074876,5.297231,4.6834874,4.1124105,3.6726158,3.8006158,4.1747694,4.706462,5.5204105,6.2687182,6.813539,7.1089234,7.1581545,7.003898,7.4863596,7.817847,7.975385,7.9491286,7.7456417,8.162462,8.553026,8.887795,9.055181,8.887795,8.553026,8.090257,7.893334,8.103385,8.612103,9.570462,9.90195,9.96759,10.131693,10.738873,9.803488,9.229129,8.743385,8.2445135,7.7948723,7.5585647,7.4732313,7.2369237,6.9152827,6.9382567,6.9021544,7.059693,7.0137444,6.672411,6.262154,5.47118,4.637539,3.9712822,3.511795,3.114667,2.917744,2.7766156,2.5993848,2.300718,1.7952822,1.6377437,1.5327181,1.4703591,1.4178462,1.3128207,1.2800001,1.1881026,1.1224617,1.1749744,1.4506668,1.8412309,4.71959,8.467693,11.680821,13.200411,13.6697445,14.490257,13.627078,11.18195,9.380103,7.207385,3.8006158,1.2274873,0.21989745,0.20348719,0.761436,1.1158975,1.3587693,1.5589745,1.7460514,1.1881026,2.5271797,2.281026,0.52512825,0.86317956,0.56451285,0.43323082,0.78769237,1.1290257,0.15097436,0.32164106,0.21661541,0.09189744,0.24287182,1.0043077,0.82379496,1.0075898,0.92225647,0.69579494,1.2274873,0.9288206,1.3062565,1.7526156,1.9790771,1.9987694,2.6387694,3.0490258,3.186872,3.2131286,3.495385,3.1540515,3.062154,3.0884104,3.2984617,3.9614363,4.604718,5.0609236,5.3136415,5.605744,6.4623594,6.8562055,5.786257,4.8147697,4.7294364,5.533539,6.157129,7.1876926,8.251078,9.314463,10.676514,9.810052,9.393231,9.432616,9.750975,9.974154,9.777231,9.875693,10.292514,11.21477,13.026463,13.751796,14.8480015,16.02954,16.925539,17.106052,16.108309,16.443079,16.722052,16.66954,17.109335,17.09949,17.808413,18.409027,18.58954,18.527182,16.91241,16.433231,16.823795,17.56882,17.913437,18.271181,18.448412,18.057848,17.335796,17.155283,17.23077,16.354464,14.887385,13.643488,13.88636,13.495796,13.938873,14.375385,14.788924,16.000002,16.902565,17.217642,17.591797,18.146463,18.46154,17.929848,17.270155,17.51959,18.615797,19.380514,18.546873,17.77559,17.430975,17.45395,17.332514,16.86318,16.820515,16.256,15.396104,15.648822,15.911386,16.098463,15.855591,15.409232,15.556924,16.433231,13.223386,8.759795,6.11118,8.562873,11.585642,12.209231,11.890873,11.1294365,9.462154,7.965539,7.525744,6.738052,5.2578464,3.8137438,3.3050258,3.239385,3.367385,3.4855387,3.446154,2.8258464,2.9440002,3.692308,4.7327185,5.5138464,5.149539,6.235898,7.6176414,8.5661545,8.789334,9.383386,9.9282055,9.787078,9.248821,9.544206,8.192,7.515898,7.9983597,9.012513,8.815591,9.462154,10.686359,10.706052,9.944616,11.034257,10.985026,10.407386,10.771693,13.029744,17.64431,16.902565,13.5548725,11.434668,11.211488,10.377847,8.116513,7.8769236,7.584821,6.380308,4.650667,4.1189747,4.775385,5.5236926,5.3858466,3.498667,2.7175386,4.5423594,4.900103,3.3280003,2.9440002,4.092718,3.764513,2.989949,3.006359,5.2414365,6.377026,5.47118,3.882667,2.7175386,2.809436,2.6584618,3.9548721,4.886975,5.152821,5.943795,6.9152827,6.7872825,6.2851286,5.5236926,4.020513,3.8859491,4.204308,4.4898467,4.4242053,3.8531284,3.751385,3.8695388,3.9318976,3.9220517,4.1091285,3.5282054,3.620103,4.0402055,4.388103,4.210872,4.06318,4.269949,4.1452312,3.6758976,3.515077,3.570872,4.1714873,4.4307694,4.342154,4.7950773,5.149539,5.1232824,5.0543594,5.169231,5.586052,5.7435904,5.609026,5.622154,5.865026,6.055385,5.3924108,5.356308,5.402257,5.211898,4.6900516,4.450462,4.699898,4.9526157,4.926359,4.5554876,4.8049235,5.786257,6.0980515,5.5204105,5.031385,4.450462,4.135385,3.9384618,3.8564105,4.0533338,4.069744,4.089436,4.0008206,3.892513,4.0369234,4.31918,4.4373336,4.588308,4.850872,5.175795,6.4000006,5.930667,4.8377438,3.8859491,3.564308,3.6168208,3.5971284,3.5347695,3.4067695,3.1507695,2.6880002,2.3729234,2.2744617,2.3696413,2.5632823,2.3696413,2.231795,2.1300514,2.1202054,2.3236926,2.3958976,2.5271797,2.4451284,2.2777438,2.556718,2.4549747,2.2055387,1.7558975,1.276718,1.1585642,1.3161026,1.5753847,1.8707694,2.1103592,2.166154,2.4451284,2.9078977,3.2951798,3.4921029,3.515077,4.096,3.8006158,3.1967182,2.7536411,2.8422565,3.2951798,3.6562054,3.3214362,2.678154,3.1113849,4.3585644,5.1232824,5.6287184,5.901129,5.7731285,5.8420515,5.5532312,5.330052,5.293949,5.2709746,5.0642056,5.159385,5.802667,6.7905645,7.4830775,6.3376417,4.785231,3.9220517,4.07959,4.8147697,5.07077,5.280821,5.622154,6.012718,6.1308722,7.4043083,7.643898,7.02359,6.3277955,6.961231,6.4590774,5.5893335,4.3585644,3.2262566,3.1081028,3.9975388,4.2502565,4.1222568,3.8301542,3.5577438,3.6463592,3.3476925,3.511795,4.1124105,4.2568207,3.948308,3.7251284,3.4724104,3.5052311,4.5587697,5.405539,5.5958977,5.113436,4.630975,5.481026,5.6287184,4.706462,3.8038976,3.511795,3.9286156,4.0041027,3.7940516,4.2469745,5.3136415,5.9470773,5.477744,5.5007186,5.477744,5.32677,5.405539,4.8311796,4.4964104,4.4438977,4.585026,4.670359,4.923077,4.601436,4.1222568,4.565334,7.6701546,5.83877,4.59159,3.7940516,3.764513,5.2578464,4.535795,4.069744,4.2994876,4.9788723,5.1954875,6.1538467,6.3179493,6.3179493,6.619898,7.50277,7.00718,7.765334,8.254359,7.9983597,7.574975,4.896821,4.2896414,4.6900516,5.4908724,6.5378466,11.247591,11.723488,12.337232,13.896206,13.653335,20.279797,20.004105,16.879591,12.547283,6.245744,15.770258,11.904001,7.197539,6.882462,8.891078,9.757539,11.565949,10.745437,8.4512825,10.555078,6.373744,6.370462,6.3540516,5.106872,4.391385,4.1682053,4.1517954,4.0303593,3.636513,2.9636924,2.8127182,2.176,1.7690258,1.7690258,1.7985642,1.8576412,1.6935385,1.5491283,1.657436,2.2580514,1.6016412,1.211077,1.1060513,1.1454359,1.0305642,1.079795,1.0272821,0.9321026,0.88287187,1.0075898,1.2570257,1.5097437,1.6804104,1.723077,1.6311796,1.8215386,1.8412309,1.9068719,2.1300514,2.5173335,2.5632823,2.3072822,2.3072822,2.674872,3.0687182,2.4746668,2.477949,2.5042052,2.428718,2.5796926,2.9144619,2.861949,2.8127182,2.9604106,3.3214362,3.5183592,3.6726158,3.879385,4.2830772,5.0871797,4.854154,5.287385,6.363898,7.509334,7.574975,7.141744,6.9710774,7.194257,7.351795,6.3868723,7.0826674,7.3419495,7.3353853,7.1089234,6.5903597,6.3245134,5.8157954,5.5138464,5.7796926,6.8627696,5.874872,6.048821,6.436103,6.3474874,5.356308,5.907693,6.0619493,5.7009234,5.3825645,6.3277955,5.287385,4.1813335,4.384821,5.2742567,4.2207184,4.7392826,4.5128207,3.9581542,3.5446157,3.8104618,4.775385,5.7731285,6.2490263,5.9536414,4.95918,5.7698464,5.8945646,5.920821,5.8486156,5.0904617,4.7327185,4.279795,3.9811285,3.7087183,2.930872,3.1245131,3.2131286,2.9669745,2.540308,2.484513,2.5764105,2.4451284,2.294154,2.228513,2.2613335,2.2022567,1.7985642,1.4834872,1.5491283,2.1398976,2.284308,2.425436,2.537026,2.5304618,2.2482052,7.8703594,7.9097443,7.683283,7.450257,7.39118,7.6110773,8.116513,8.648206,8.769642,8.395488,7.7948723,7.453539,7.256616,7.3616414,7.6767187,7.8670774,7.50277,7.2303596,6.8594875,6.409847,6.088206,6.514872,6.688821,6.567385,6.242462,5.940513,5.8125134,5.648411,5.3202057,4.818052,4.240411,3.892513,3.8564105,4.194462,4.9394875,6.1013336,6.8562055,7.397744,7.817847,8.169026,8.454565,8.746667,9.179898,9.399796,9.301334,9.005949,9.248821,9.632821,9.91836,9.915077,9.458873,8.667898,7.9983597,7.680001,7.785026,8.231385,9.366975,9.626257,9.412924,9.229129,9.639385,9.255385,9.048616,8.766359,8.346257,7.9195905,7.574975,7.463385,7.3353853,7.145026,7.030154,6.665847,6.4754877,6.0947695,5.4908724,4.9493337,4.0041027,3.367385,2.92759,2.5895386,2.2711797,2.048,1.8379488,1.6246156,1.3883078,1.1027694,0.94523084,0.8172308,0.7318975,0.67610264,0.636718,0.6662565,0.6268718,0.60389745,0.65969235,0.86317956,1.1027694,3.442872,6.1013336,8.576,11.657847,11.69395,11.59877,10.597744,8.661334,6.485334,4.9493337,2.7470772,1.0568206,0.28882053,0.059076928,0.03938462,0.068923086,0.16082053,0.28882053,0.4135385,0.57764107,1.0896411,0.98133343,0.380718,0.5021539,0.26912823,0.16410258,0.28225642,0.40369233,0.01969231,0.0032820515,0.0,0.14441027,0.5316923,1.2307693,0.6498462,0.5415385,0.5513847,0.6498462,1.1290257,1.1979488,1.5819489,1.8510771,1.910154,1.9889232,2.5993848,2.9571285,2.9833848,2.8422565,2.9243078,3.0982566,3.2065644,3.4198978,3.895795,4.788513,5.1232824,5.284103,5.159385,4.9329233,5.106872,5.4186673,4.706462,4.2535386,4.601436,5.5597954,6.0061545,6.6494365,7.702975,8.910769,9.540924,8.907488,8.448001,8.490667,9.02236,9.688616,10.075898,10.781539,11.467488,12.370052,14.28677,15.363283,15.891693,16.659693,17.624617,17.897026,18.051283,18.924309,19.541334,19.452719,18.740515,17.365335,17.463797,17.946259,18.139898,17.80513,16.479181,15.849027,16.02954,16.715488,17.19795,17.188105,17.496616,17.378464,16.866463,16.784412,16.955078,16.649847,15.58318,14.424617,14.769232,14.388514,14.818462,15.209026,15.435489,16.12472,17.125746,17.32595,17.220924,17.263592,17.893745,18.169437,18.448412,18.704412,18.852104,18.743795,18.267899,18.17272,17.900309,17.237335,16.31836,15.681643,16.787693,17.424412,17.089642,16.99118,16.07877,15.724309,15.501129,15.248411,15.067899,15.323898,12.47836,8.930462,7.0892315,9.360411,11.503591,12.740924,12.711386,11.483898,9.580308,8.224821,7.8769236,6.987488,5.3792825,4.269949,4.076308,3.8071797,3.5577438,3.3969233,3.3772311,2.9768207,3.0490258,3.5807183,4.453744,5.464616,5.2709746,6.170257,7.433847,8.421744,8.585847,8.92718,10.125129,10.28595,9.412924,9.393231,8.241231,7.6964107,8.362667,9.642668,9.731283,9.3768215,10.390975,11.1294365,11.155693,11.250873,11.336206,11.861334,11.900719,11.808822,13.236514,13.791181,12.186257,11.047385,11.113027,11.224616,8.868103,7.7981544,6.7150774,5.356308,4.4865646,3.7284105,4.092718,5.8781543,7.210667,4.0336413,1.7394873,3.1606157,4.128821,3.5052311,3.2000003,2.9407182,2.6256413,2.92759,4.1747694,6.370462,7.64718,6.242462,4.273231,3.0982566,3.3280003,3.249231,4.082872,4.890257,5.421949,6.0980515,6.4623594,6.8562055,6.688821,5.9536414,5.2414365,4.716308,4.338872,3.95159,3.7448208,4.263385,4.2371287,4.2863593,4.06318,3.629949,3.4691284,3.2032824,3.4756925,3.9581542,4.194462,3.5774362,3.817026,3.9811285,3.8564105,3.5413337,3.4527183,3.5971284,3.9614363,4.263385,4.450462,4.71959,5.3792825,5.47118,5.2545643,4.8607183,4.312616,4.059898,4.2240005,4.571898,4.9132314,5.074052,4.5456414,4.5029745,4.706462,4.9394875,4.9887185,4.8344617,5.034667,5.07077,4.841026,4.6802053,4.9821544,5.7534366,6.0192823,5.5729237,5.0051284,4.397949,3.9417439,3.6693337,3.570872,3.629949,3.9975388,4.2535386,4.276513,4.0992823,3.8859491,4.059898,4.397949,4.6112823,4.650667,4.7261543,5.1626673,4.6276927,3.9187696,3.4888208,3.43959,3.387077,3.255795,3.2098465,3.2262566,3.1113849,2.612513,2.294154,2.103795,2.0184617,2.044718,1.9364104,1.9396925,1.9626669,1.9987694,2.1398976,2.1989746,2.2580514,2.166154,2.03159,2.231795,2.1858463,2.0086155,1.5885129,1.1224617,1.1093334,1.4178462,1.8018463,1.8937438,1.7887181,2.0545642,2.3991797,2.665026,3.0293336,3.3444104,3.1671798,3.6693337,3.5282054,3.2262566,3.0162053,2.934154,3.114667,3.6857438,3.820308,3.4855387,3.43959,4.013949,4.644103,5.366154,5.917539,5.7632823,5.7009234,5.5991797,5.7534366,5.9602056,5.504,4.893539,5.0674877,5.76,6.744616,7.830975,6.5280004,4.893539,3.879385,3.751385,4.086154,4.4996924,4.8607183,5.398975,6.0783596,6.6067696,7.174565,6.9842057,6.954667,7.2336416,7.1876926,7.637334,7.785026,6.5083084,4.5522056,4.5029745,4.8049235,4.9394875,4.6244106,4.1189747,4.2141542,4.44718,4.076308,4.073026,4.46359,4.3552823,4.20759,4.1878977,4.010667,3.8662567,4.4110775,5.3924108,5.7435904,5.293949,4.6145644,5.024821,5.402257,4.6867695,4.0467696,4.007385,4.44718,4.5456414,4.6276927,5.0116925,5.61559,5.9536414,5.7435904,5.58277,5.6418467,5.8420515,5.858462,5.504,5.1954875,5.0477953,5.07077,5.182359,4.8705645,4.9362054,4.8640003,5.146257,7.2861543,4.57518,3.748103,3.56759,3.9384618,5.8847184,5.543385,5.0510774,5.031385,5.4843082,5.7698464,6.6494365,7.3682055,7.8112826,8.034462,8.277334,8.326565,9.209436,9.6,9.458873,10.023385,9.403078,8.172308,8.553026,10.70277,12.698257,15.140103,13.062565,13.167591,16.600616,18.947283,22.744617,29.952002,33.7198,30.542772,20.26995,16.613745,11.480617,8.868103,9.498257,10.81436,10.079181,9.229129,8.976411,9.330873,9.586872,5.2020516,5.431795,5.330052,3.8695388,3.9253337,3.82359,3.8137438,3.7874875,3.5840003,2.9669745,2.8849232,2.3696413,2.028308,1.9035898,1.5031796,1.7788719,1.7887181,1.585231,1.3915899,1.595077,1.2668719,0.9682052,0.8467693,0.86317956,0.8041026,0.79425645,0.8041026,0.7844103,0.7384616,0.73517954,0.892718,1.1355898,1.3718976,1.5655385,1.7558975,1.9626669,1.8838975,1.975795,2.3040001,2.546872,2.5009232,2.3072822,2.225231,2.3926156,2.8389745,2.3926156,2.4188719,2.297436,2.03159,2.2514873,2.7536411,2.6223593,2.356513,2.3072822,2.7044106,3.1737437,3.511795,3.8367183,4.2535386,4.8705645,5.3037953,6.091488,7.1154876,7.9294367,7.755488,6.9382567,6.547693,6.875898,7.2664623,6.1013336,6.7610264,7.450257,7.5618467,6.994052,6.1538467,5.98318,5.868308,5.7435904,6.2523084,8.743385,6.7774363,6.491898,6.3442054,5.83877,5.5072823,6.055385,6.2851286,5.904411,5.156103,4.7950773,4.919795,4.57518,4.640821,5.077334,4.9329233,5.093744,4.096,3.3805132,3.4592824,3.889231,4.7491283,5.5171285,5.6943593,5.3070774,4.903385,5.474462,5.4613338,5.405539,5.2578464,4.3716927,3.8006158,3.4625645,3.4789746,3.6069746,3.2328207,2.7831798,2.7109745,2.4648206,2.0151796,1.8904617,2.3335385,2.3335385,2.2449234,2.1825643,2.0118976,2.1103592,1.7887181,1.5556924,1.6147693,1.8838975,1.8215386,1.8904617,2.0086155,2.0217438,1.6968206,8.283898,8.231385,7.8080006,7.3682055,7.069539,6.87918,7.4732313,8.1755905,8.5891285,8.65477,8.648206,7.90318,7.463385,7.466667,7.706257,7.640616,7.1515903,7.020308,6.7971287,6.4590774,6.4000006,6.918565,6.8988724,6.678975,6.449231,6.2162056,5.87159,5.671385,5.4580517,5.097026,4.4832826,4.325744,4.493129,4.84759,5.5007186,6.806975,7.6110773,8.139488,8.710565,9.353847,9.803488,9.642668,9.921641,10.079181,9.915077,9.609847,9.842873,10.220308,10.282667,9.90195,9.271795,8.592411,8.169026,7.965539,7.9819493,8.231385,9.18318,9.452309,9.163487,8.720411,8.786052,8.838565,8.835282,8.592411,8.169026,7.857231,7.5388722,7.3353853,7.1844106,7.0334363,6.816821,6.163693,5.477744,4.775385,4.1091285,3.5511796,2.8422565,2.3991797,2.103795,1.8510771,1.5392822,1.3062565,1.0896411,0.8763078,0.6826667,0.5415385,0.42338464,0.32820517,0.27241027,0.25271797,0.25271797,0.256,0.23302566,0.23302566,0.29538465,0.44964105,0.56123084,2.3696413,4.096,5.9536414,10.144821,9.590155,9.442462,8.953437,7.6242056,5.21518,4.8672824,3.9351797,2.356513,0.6892308,0.13128206,0.059076928,0.032820515,0.03938462,0.068923086,0.10502565,0.64000005,1.0601027,0.9288206,0.38728207,0.15753847,0.059076928,0.013128206,0.0,0.0032820515,0.02297436,0.0032820515,0.0,0.2100513,0.5940513,0.8763078,0.4660513,0.50543594,0.69251287,0.93866676,1.3784616,1.3292309,1.6147693,1.8576412,1.9298463,1.9593848,2.5009232,2.6912823,2.6715899,2.6256413,2.7831798,3.2098465,3.4592824,3.8301542,4.414359,5.093744,5.0116925,4.9460516,4.673641,4.2305646,3.9154875,4.1452312,3.9778464,4.2469745,5.0904617,5.933949,6.2818465,6.6100516,7.50277,8.720411,9.179898,8.726975,8.582564,8.736821,9.222565,10.128411,10.692924,11.851488,12.829539,13.682873,15.284514,16.886156,17.673847,18.533745,19.403488,19.242668,19.86954,20.407797,20.719591,20.480001,19.167181,17.312822,16.97477,17.05354,17.02072,16.91241,15.970463,15.2155905,14.995693,15.29436,15.724309,16.019693,16.544823,16.613745,16.137848,15.599591,15.996719,15.960617,15.461744,14.923489,15.235283,15.560206,15.763694,15.812924,15.904821,16.485744,17.207796,17.529438,17.562258,17.683693,18.54031,18.60595,19.124514,19.026052,18.323694,18.133335,18.25477,18.60595,18.67159,18.120207,16.836924,16.02954,17.782156,18.84554,18.277744,17.417847,15.593027,14.713437,14.388514,14.345847,14.424617,13.659899,11.815386,9.731283,8.78277,10.866873,11.789129,12.793437,12.484924,10.807796,9.028924,8.408616,8.086975,7.269744,5.973334,5.024821,4.8147697,4.391385,3.8662567,3.4264617,3.3411283,3.1737437,3.3542566,3.8990772,4.716308,5.6320004,5.464616,5.7829747,6.8365135,8.100103,8.254359,8.530052,9.852718,10.079181,9.170052,9.209436,8.474257,7.653744,7.9491286,9.255385,10.171078,9.6065645,10.000411,10.712616,11.21477,11.1064625,11.52,13.679591,14.076719,12.068104,9.892103,11.1983595,11.769437,11.211488,10.19077,10.423796,9.222565,7.5421543,5.58277,3.9647183,3.7185643,3.0096412,3.5216413,5.658257,7.4240007,4.417641,1.9396925,2.5764105,3.5741541,3.8006158,3.7743592,2.605949,2.2482052,3.0358977,4.8311796,7.020308,8.6580515,7.056411,4.84759,3.639795,4.010667,3.9253337,4.1714873,4.713026,5.4416413,6.170257,6.1341543,6.619898,6.688821,6.2523084,6.048821,5.2644105,4.338872,3.5938463,3.3312824,3.8104618,3.6332312,3.8006158,3.7054362,3.2787695,2.9702566,3.0391798,3.259077,3.5807183,3.7185643,3.1442053,3.3050258,3.1770258,2.9407182,2.7569232,2.7569232,3.0654361,3.3641028,3.754667,4.1485133,4.2863593,4.857436,5.041231,4.768821,4.059898,3.0358977,2.6978464,3.062154,3.570872,3.892513,3.895795,3.7251284,3.9187696,4.3290257,4.7917953,5.152821,5.1922054,5.428513,5.474462,5.3825645,5.6451287,5.677949,5.8912826,5.87159,5.474462,4.857436,4.2830772,3.7940516,3.501949,3.3903592,3.3345644,3.8400004,4.1058464,4.0500517,3.8071797,3.7087183,3.8990772,4.2436924,4.325744,4.138667,4.092718,3.9548721,3.5577438,3.2754874,3.249231,3.3969233,3.249231,2.9144619,2.7142565,2.6945643,2.6289232,2.349949,2.172718,2.0020514,1.8379488,1.7755898,1.6771283,1.719795,1.8149745,1.9003079,1.9495386,1.8806155,1.8674873,1.8871796,1.9462565,2.0611284,1.9035898,1.719795,1.394872,1.0666667,1.0929232,1.3423591,1.8313848,1.9659488,1.7920002,2.0184617,2.294154,2.5271797,2.7667694,2.9505644,2.9046156,3.0851285,3.0030773,2.9801028,3.0785644,3.1048207,2.9243078,3.3509746,3.8071797,3.9614363,3.751385,3.8662567,4.3585644,5.093744,5.7468724,5.8092313,6.0291286,6.1472826,6.452513,6.744616,6.3277955,5.293949,5.3070774,5.970052,6.882462,7.64718,6.1472826,5.0477953,4.4012313,4.1485133,4.1156926,4.4996924,4.71959,5.074052,5.684513,6.47877,6.8430777,6.5706673,6.7282057,7.1647186,6.498462,7.1483083,7.243488,6.121026,4.6211286,5.07077,5.4908724,5.605744,5.1167183,4.4045134,4.519385,4.854154,4.6112823,4.630975,4.9099493,4.598154,4.525949,4.6539493,4.601436,4.397949,4.4701543,5.3070774,5.7468724,5.4153852,4.71959,4.854154,5.2053337,4.8836927,4.673641,4.8705645,5.293949,5.2381544,5.4153852,5.681231,5.874872,5.8256416,5.7468724,5.3825645,5.402257,5.901129,6.3967185,6.4000006,6.114462,5.835488,5.789539,6.1078978,5.5269747,5.8486156,5.8157954,5.5105643,6.373744,3.1967182,2.605949,3.5872824,5.1331286,6.23918,6.49518,6.3967185,6.3474874,6.616616,7.3452315,7.6570263,8.195283,8.356103,8.267488,8.776206,9.800206,11.421539,11.674257,10.988309,12.209231,14.358975,12.406155,11.930258,14.214565,16.269129,17.050259,13.407181,13.633642,18.835693,22.921848,27.795694,43.490463,50.898056,43.651287,28.107489,20.896822,17.371899,14.516514,11.588924,10.118565,8.5661545,6.6592827,7.2205133,9.265231,7.9852314,3.7087183,4.315898,4.673641,3.5446157,3.6004105,3.6069746,3.5347695,3.4888208,3.3641028,2.8389745,2.5829747,2.2744617,2.0742567,1.9495386,1.7066668,1.6475899,1.7329233,1.591795,1.2340513,1.0272821,0.88287187,0.81394875,0.7811283,0.764718,0.77456415,0.7384616,0.761436,0.7811283,0.74830776,0.6432821,0.65312827,0.92553854,1.2012309,1.3751796,1.5031796,1.8084104,1.847795,2.0808206,2.5042052,2.6518977,2.409026,2.3171284,2.2416413,2.2646155,2.7044106,2.3663592,2.3040001,2.2350771,2.1103592,2.100513,2.4385643,2.3368206,2.0611284,1.9396925,2.356513,2.9013336,3.5380516,4.020513,4.3749747,4.893539,5.58277,6.193231,6.9087186,7.522462,7.4436927,6.9809237,6.672411,6.987488,7.3550773,6.1538467,6.232616,6.961231,7.213949,6.672411,5.83877,5.865026,6.058667,6.0258465,6.672411,10.20718,8.080411,6.941539,6.157129,5.72718,6.2884107,6.2752824,6.380308,6.157129,5.5532312,4.923077,5.421949,5.395693,5.0642056,4.8114877,5.1889234,4.6276927,3.5380516,3.1770258,3.6529233,3.9614363,4.378257,4.8672824,4.955898,4.6966157,4.6900516,4.9394875,4.630975,4.46359,4.4274874,3.7842054,3.387077,3.1573336,3.1113849,3.2065644,3.3411283,2.7306669,2.4516926,2.231795,2.0053334,1.9003079,2.4057438,2.425436,2.3401027,2.2678976,2.0775387,2.162872,2.0118976,1.9035898,1.8904617,1.8051283,1.595077,1.5786668,1.6738462,1.7132308,1.4539489,8.513641,8.12636,7.532308,6.9842057,6.560821,6.1538467,6.744616,7.581539,8.36595,8.960001,9.380103,8.264206,7.4043083,7.1220517,7.177847,6.7577443,6.196513,6.304821,6.5083084,6.6461544,6.9809237,7.397744,7.177847,6.875898,6.6527185,6.2884107,5.668103,5.362872,5.2447186,5.10359,4.637539,4.601436,5.0642056,5.5729237,6.1013336,7.076103,8.152616,8.684308,9.366975,10.187488,10.417232,9.833026,10.000411,10.233437,10.184206,9.869129,10.148104,10.31877,10.125129,9.504821,8.595693,8.480822,8.585847,8.664616,8.648206,8.635077,9.265231,9.701744,9.5835905,9.07159,8.848411,8.700719,8.411898,7.965539,7.525744,7.463385,7.3452315,7.0432825,6.6494365,6.242462,5.861744,5.100308,4.1550775,3.3936412,2.9013336,2.4582565,2.1431797,1.7985642,1.5556924,1.3620514,0.97805136,0.761436,0.58092314,0.4135385,0.25928208,0.15425642,0.12143591,0.09189744,0.06564103,0.052512825,0.052512825,0.03938462,0.036102567,0.052512825,0.08861539,0.15097436,0.19364104,1.5360001,3.0490258,4.8377438,8.251078,8.113232,8.198565,8.041026,7.1647186,5.0838976,6.1308722,5.796103,3.7218463,1.0010257,0.17066668,0.08533334,0.049230773,0.06235898,0.12471796,0.23302566,0.7253334,0.99774367,0.83035904,0.35774362,0.068923086,0.04594872,0.036102567,0.02297436,0.009846155,0.016410258,0.006564103,0.0032820515,0.15097436,0.39056414,0.446359,0.5677949,0.86646163,1.0732309,1.2406155,1.7394873,1.3784616,1.7591796,2.162872,2.2449234,2.038154,2.5009232,2.4648206,2.4484105,2.6912823,3.1343591,3.2525132,3.570872,4.089436,4.630975,4.850872,4.562052,4.493129,4.2830772,3.892513,3.6135387,3.8564105,4.2469745,5.031385,5.9995904,6.482052,6.954667,7.194257,7.8670774,8.973129,9.852718,9.488411,9.642668,9.80677,10.115283,11.369026,11.753027,12.691693,13.794462,14.838155,15.799796,17.703386,19.006361,20.030361,20.578463,19.931898,20.102566,20.033642,19.977848,19.67918,18.353231,16.899282,16.354464,16.042667,15.819489,16.065641,15.67836,14.857847,14.395078,14.496821,14.79877,15.645539,16.147694,15.983591,15.192616,14.152206,14.818462,14.641232,14.427898,14.598565,15.163078,16.423386,16.479181,16.292105,16.393847,16.90913,17.447386,18.008617,18.635489,19.410053,20.4439,19.48554,19.01949,18.182566,17.211079,17.427694,17.93313,18.520617,19.15077,19.367386,18.320412,17.322668,19.032618,19.662771,18.267899,16.761436,14.857847,13.640206,13.10195,13.157744,13.633642,12.012309,10.548513,9.865847,10.397539,12.393026,12.265027,12.530872,11.67754,9.731283,8.251078,8.448001,8.116513,7.4699492,6.672411,5.858462,5.353026,4.8804107,4.342154,3.8334363,3.6430771,3.511795,3.7874875,4.4438977,5.2545643,5.7698464,5.290667,5.1298466,6.1538467,7.755488,7.8506675,7.965539,9.025641,9.225847,8.625232,9.170052,8.746667,7.532308,7.2861543,8.477539,10.269539,10.112,9.603283,9.711591,10.515693,11.195078,11.382154,14.539488,16.114874,14.057027,8.79918,10.397539,12.406155,11.746463,9.019077,8.493949,8.667898,6.7774363,4.381539,2.8521028,3.4034874,2.4516926,4.082872,5.910975,6.5312824,5.5007186,3.1507695,2.8947694,3.3280003,3.7218463,4.027077,2.5764105,2.422154,3.2262566,4.7622566,6.9152827,8.835282,7.8145647,5.7501545,4.2305646,4.529231,4.31918,4.2601027,4.4734364,5.0576415,6.114462,6.2588725,6.5805135,6.5378466,6.170257,6.1046157,5.093744,4.46359,3.9056413,3.3017437,2.7208207,2.4516926,2.5928206,2.7634873,2.809436,2.806154,2.8717952,2.802872,2.878359,3.0358977,2.868513,2.7437952,2.3401027,1.9659488,1.7952822,1.847795,2.0742567,2.425436,2.7798977,3.058872,3.2262566,3.6036925,3.7973337,3.5380516,2.8553848,2.0676925,2.041436,2.4516926,2.8980515,3.131077,3.0654361,3.0293336,3.387077,3.8990772,4.4340515,4.965744,5.5204105,5.789539,5.901129,6.0816417,6.6560006,6.564103,6.2720003,5.7501545,5.0642056,4.378257,3.8596926,3.4494362,3.2000003,3.1015387,3.0687182,3.318154,3.3969233,3.2656412,3.1442053,3.4822567,3.761231,3.9811285,3.8859491,3.5610259,3.446154,3.239385,3.0916924,3.045744,3.121231,3.318154,3.1934361,2.737231,2.349949,2.1431797,1.9429746,1.975795,1.9331284,1.8674873,1.8149745,1.7920002,1.6147693,1.591795,1.6771283,1.785436,1.8084104,1.7362052,1.719795,1.8904617,2.169436,2.2613335,1.9232821,1.5524104,1.204513,0.96492314,0.9353847,1.1979488,1.7920002,2.0512822,1.9331284,1.9922053,2.0906668,2.3696413,2.4451284,2.3302567,2.4385643,2.297436,2.3040001,2.5238976,2.8980515,3.2787695,3.045744,2.9801028,3.2065644,3.6168208,3.8564105,3.8728209,4.2962055,4.709744,5.041231,5.5696416,6.482052,6.961231,7.145026,7.131898,6.9677954,5.933949,5.72718,6.196513,6.8332314,6.764308,5.1954875,4.7622566,4.6900516,4.6244106,4.630975,5.0149746,5.0215387,4.890257,4.9296412,5.540103,6.117744,6.436103,6.698667,6.692103,5.796103,6.045539,5.182359,4.1485133,3.7743592,4.8082056,5.648411,5.8157954,5.3103595,4.5554876,4.388103,4.7294364,4.7491283,4.8705645,5.07077,4.903385,4.916513,5.0477953,5.028103,4.8147697,4.601436,5.028103,5.346462,5.159385,4.7294364,4.9854364,5.10359,5.1298466,5.3398976,5.7107697,5.917539,5.691077,5.6976414,5.8518977,6.0028725,5.9503593,5.622154,5.2611284,5.2414365,5.7501545,6.764308,7.1122055,7.076103,6.921847,6.951385,7.4797955,6.8627696,7.0465646,6.806975,6.160411,6.3573337,3.5183592,2.6912823,4.1485133,6.445949,6.4065647,8.096821,7.939283,7.6077952,8.323282,10.837335,9.409642,8.723693,8.717129,9.366975,10.696206,12.740924,15.432206,15.258258,12.763899,12.547283,16.436514,15.012104,13.216822,13.843694,17.506462,16.354464,12.652308,13.984821,20.079592,22.826668,29.367798,46.486977,51.091698,39.246773,26.190771,32.495594,37.651695,30.972721,15.366566,7.325539,6.0849237,4.348718,5.208616,7.8441033,7.53559,3.442872,3.95159,4.7425647,4.1780515,3.31159,3.4625645,3.3444104,3.2262566,3.0720003,2.537026,2.1366155,2.0250258,1.9692309,1.9561027,2.169436,1.6410258,1.5327181,1.4834872,1.3095386,0.9878975,0.67938465,0.7056411,0.79097444,0.827077,0.8795898,0.84348726,0.82379496,0.7778462,0.6826667,0.5349744,0.5349744,0.8763078,1.204513,1.2996924,1.0699488,1.3620514,1.5721027,1.9593848,2.4615386,2.7011285,2.284308,2.2383592,2.2088206,2.2055387,2.6354873,2.2449234,2.034872,2.1891284,2.4549747,2.1398976,2.2186668,2.231795,2.1202054,2.0611284,2.4746668,2.9669745,3.7185643,4.2305646,4.46359,4.850872,5.2512827,5.536821,6.0685134,6.738052,6.9743595,7.1876926,7.325539,7.64718,7.765334,6.6428723,5.9634876,6.38359,6.8332314,6.7183595,5.930667,5.865026,5.87159,5.802667,6.567385,10.115283,9.068309,7.2992826,6.183385,6.183385,6.8496413,6.294975,5.937231,5.874872,6.1341543,6.6592827,6.49518,6.1013336,5.421949,4.8147697,5.0674877,3.9647183,3.3903592,3.4888208,3.9647183,4.066462,4.027077,4.2994876,4.4767184,4.4340515,4.31918,4.3027697,3.757949,3.620103,3.9384618,3.882667,3.757949,3.5314875,3.1770258,2.8750772,3.0194874,3.0096412,2.7963078,2.5796926,2.4320002,2.2777438,2.5698464,2.4516926,2.3368206,2.3762052,2.4582565,2.3663592,2.2678976,2.2416413,2.225231,2.0250258,1.7985642,1.5819489,1.4834872,1.4703591,1.3751796,7.781744,7.4043083,6.941539,6.6002054,6.38359,6.1046157,6.432821,6.698667,7.6209235,8.917334,9.3078985,8.41518,7.1876926,6.1997952,5.6451287,5.3398976,5.169231,5.5762057,6.245744,6.820103,6.882462,6.626462,6.514872,6.2227697,5.7534366,5.4482055,4.6769233,4.322462,4.204308,4.210872,4.273231,4.4800005,4.5128207,5.0674877,6.0160003,6.3934364,7.4797955,7.9163084,8.625232,9.488411,9.353847,9.219283,9.734565,10.643693,11.372309,11.017847,10.502565,10.112,10.164514,10.220308,9.048616,8.815591,8.940309,9.117539,9.15036,8.940309,9.015796,9.508103,9.846154,9.737847,9.199591,8.664616,7.788308,6.9809237,6.6822567,7.3550773,7.39118,6.8430777,6.0061545,5.1167183,4.348718,3.7152824,3.0326157,2.5074873,2.1300514,1.6771283,1.4112822,1.0765129,0.7975385,0.6104616,0.48902568,0.34133336,0.2231795,0.13128206,0.068923086,0.04594872,0.02297436,0.016410258,0.016410258,0.016410258,0.016410258,0.0032820515,0.0,0.0,0.006564103,0.029538464,0.14112821,1.0108719,2.103795,3.1376412,4.089436,6.0783596,6.4754877,6.1538467,5.622154,5.034667,6.2194877,3.7152824,1.2307693,0.24287182,0.0,0.013128206,0.006564103,0.02297436,0.108307704,0.3052308,0.7187693,0.97805136,0.72861546,0.16738462,0.04594872,0.118153855,0.15425642,0.118153855,0.03938462,0.016410258,0.026256412,0.013128206,0.098461546,0.41025645,1.0666667,0.94523084,0.4955898,0.2855385,0.6170257,1.4966155,1.9331284,2.6387694,2.9013336,2.550154,1.9528207,2.5009232,2.540308,2.4484105,2.537026,3.0358977,2.793026,3.1606157,3.8038976,4.33559,4.348718,4.8114877,4.919795,4.4077954,3.8071797,4.457026,4.699898,5.4186673,6.2687182,6.8594875,6.774154,7.3353853,7.276308,7.7259493,8.92718,10.20718,10.328616,10.535385,10.663385,11.323078,13.88636,13.7386675,13.026463,13.426873,14.8709755,15.51754,17.860924,18.080822,17.660719,17.355488,17.19795,17.270155,17.975796,18.537027,18.464823,17.54913,17.253744,16.137848,15.727591,16.114874,15.931078,16.54154,15.858873,15.37313,15.481437,15.51754,15.701335,15.727591,15.241847,14.12595,12.527591,13.371078,13.029744,12.511181,12.724514,14.480412,15.849027,16.840206,17.578669,18.031591,18.021746,18.46154,18.907898,19.90236,21.287386,22.199797,20.480001,19.5479,18.569847,17.293129,16.036104,16.853334,18.376207,19.34113,19.285336,18.54031,17.64759,18.369642,18.14318,16.577642,15.442053,14.674052,13.5089245,12.819694,12.727796,12.619488,11.16554,9.787078,10.056206,11.795693,13.075693,12.73436,12.547283,11.503591,9.668923,8.178872,8.717129,8.3823595,7.6307697,6.8955903,6.5903597,6.114462,5.428513,4.6900516,4.1452312,4.1189747,3.754667,3.7349746,4.266667,5.037949,5.2348723,4.4898467,4.6966157,6.180103,7.9852314,7.890052,7.181129,8.1755905,8.487385,7.962257,8.681026,8.950154,8.605539,8.457847,9.133949,11.063796,11.158976,9.96759,9.705027,10.791386,11.841642,10.243283,12.461949,16.098463,17.03713,9.4457445,9.042052,11.533129,11.654565,9.068309,8.346257,7.5520005,5.0576415,2.9801028,3.0129232,6.3934364,3.0129232,5.3070774,6.521436,5.658257,7.4765134,3.692308,2.353231,2.0250258,1.8773335,1.6935385,1.522872,2.9735386,4.381539,5.3398976,6.6822567,7.3550773,7.9885135,7.2631803,5.504,4.699898,4.578462,4.0434875,4.1714873,5.10359,6.042257,6.163693,6.432821,6.5378466,6.5312824,6.8365135,5.0051284,4.637539,4.1189747,3.1376412,2.6847181,3.0391798,2.678154,2.412308,2.6223593,3.2820516,2.6945643,2.5107694,2.5731285,2.6617439,2.5009232,2.612513,2.1267693,1.657436,1.5163078,1.723077,1.4572309,1.5721027,1.6508719,1.6147693,1.723077,2.103795,2.2416413,2.1464617,1.8970258,1.6771283,1.9364104,2.0709746,2.2186668,2.5304618,3.190154,3.0424619,3.1606157,3.5577438,4.2436924,5.2348723,6.3934364,6.5017443,6.157129,5.8486156,5.937231,6.1078978,5.874872,5.093744,4.06318,3.5249233,3.367385,2.9144619,2.4582565,2.1530259,2.028308,1.9692309,2.1366155,2.5140514,2.9801028,3.31159,3.239385,3.4592824,3.5183592,3.3969233,3.495385,3.495385,3.8137438,4.020513,3.892513,3.4034874,2.92759,2.487795,2.1825643,1.9692309,1.6640002,1.8215386,1.6869745,1.6016412,1.6082052,1.4506668,1.1946667,1.211077,1.3883078,1.6016412,1.723077,2.041436,2.166154,2.3696413,2.674872,2.8849232,2.7602053,2.2088206,1.5688206,1.083077,0.8992821,1.4736412,1.9462565,1.9593848,1.785436,2.3335385,2.3827693,2.3860514,2.2777438,1.9856411,1.4506668,1.083077,1.2471796,1.8215386,2.6190772,3.387077,3.9351797,3.5511796,3.0096412,2.9407182,3.8465643,4.161641,4.6276927,4.5423594,4.240411,5.080616,5.937231,6.806975,6.8266673,6.11118,5.7829747,5.549949,5.674667,5.8289237,5.654975,4.775385,4.1058464,4.322462,4.3749747,4.069744,4.059898,4.9854364,5.474462,5.280821,4.8049235,5.110154,5.3202057,5.691077,6.294975,6.820103,6.5772314,5.6254363,4.8738465,4.20759,3.9417439,4.821334,5.346462,5.4974365,5.172513,4.630975,4.4865646,4.522667,4.6966157,4.8804107,5.0642056,5.356308,5.4153852,5.4974365,5.464616,5.1626673,4.394667,4.322462,4.522667,4.713026,4.900103,5.402257,5.546667,5.4941545,5.664821,5.904411,5.477744,5.1232824,4.916513,5.044513,5.4875903,6.012718,5.7435904,5.402257,5.333334,5.7403083,6.669129,7.6209235,8.152616,8.51036,8.822155,9.078155,8.237949,7.778462,7.8080006,8.237949,8.772923,5.868308,4.2535386,4.6572313,6.6494365,8.651488,13.499078,10.59118,7.719385,9.225847,15.977027,10.981745,9.048616,11.72677,16.65313,17.532719,19.93518,22.616617,21.218464,15.291079,8.28718,11.972924,14.303181,12.491488,11.782565,25.465437,14.808617,8.740103,11.004719,17.870771,18.12677,17.371899,20.010668,19.59713,17.939693,25.11754,57.62298,83.81047,70.803696,28.100925,7.568411,6.738052,5.9634876,5.717334,6.6067696,9.353847,4.8607183,4.2962055,4.7556925,4.4110775,2.5173335,2.6880002,2.7602053,2.9243078,2.9636924,2.2416413,2.156308,2.0644104,2.0644104,2.1333334,2.1202054,1.9626669,1.4933335,1.332513,1.4145643,0.97805136,0.79425645,0.7187693,0.6826667,0.6235898,0.48902568,0.46276927,0.5021539,0.49230772,0.44964105,0.5349744,0.44964105,0.72861546,1.0469744,1.2537436,1.3883078,1.1815386,1.276718,1.4998976,1.7723079,2.0906668,1.8576412,2.0644104,2.1989746,2.15959,2.2580514,1.9035898,1.8051283,2.0939488,2.4188719,1.9692309,2.1136413,2.1956925,2.294154,2.5731285,3.2820516,3.6332312,3.9876926,4.1058464,3.9844105,3.876103,3.826872,4.8114877,5.733744,6.193231,6.485334,6.7774363,7.5191803,8.201847,8.339693,7.460103,6.4590774,6.889026,7.6635904,7.857231,6.698667,5.8912826,4.9493337,4.7556925,5.674667,7.5520005,8.858257,7.39118,6.304821,6.38359,6.042257,5.7632823,5.2512827,5.5072823,6.547693,7.4141545,6.6461544,6.380308,6.442667,6.3474874,5.3103595,4.6867695,4.532513,4.201026,3.761231,3.9680004,3.9187696,4.3290257,4.6145644,4.4767184,3.892513,3.8071797,3.6562054,3.820308,4.210872,4.273231,3.892513,3.892513,3.6824617,3.2262566,3.006359,3.3608208,3.4756925,3.2065644,2.7273848,2.5337439,2.7766156,2.4352822,2.2022567,2.2121027,2.028308,1.9692309,1.9429746,2.048,2.2580514,2.4418464,2.1366155,1.6311796,1.2504616,1.1191796,1.1454359,8.024616,7.8047185,7.141744,6.5805135,6.304821,6.1538467,6.0717955,6.0750775,6.498462,7.3025646,8.073847,8.51036,7.8834877,7.066257,6.36718,5.5236926,5.4613338,6.4557953,7.3091288,7.581539,7.6012316,7.0137444,6.629744,6.0685134,5.435077,5.32677,4.713026,4.2994876,4.164923,4.414359,5.1889234,5.4153852,5.3727183,5.2414365,5.2315903,5.5991797,5.7796926,5.979898,6.741334,7.90318,8.608821,9.051898,9.521232,10.072617,10.6469755,11.067078,11.638155,12.905026,13.400617,12.343796,9.659078,9.554052,9.271795,9.501539,9.984001,9.501539,9.380103,9.747693,9.616411,9.002667,8.89436,8.018052,7.318975,6.764308,6.377026,6.2555904,5.970052,5.832206,5.428513,4.637539,3.6036925,2.9604106,2.2613335,1.6213335,1.1158975,0.81066674,0.60061544,0.41682056,0.27569234,0.19364104,0.15753847,0.101743594,0.06235898,0.032820515,0.013128206,0.009846155,0.0032820515,0.0032820515,0.0032820515,0.0032820515,0.0032820515,0.0,0.0,0.0032820515,0.013128206,0.01969231,0.118153855,0.72861546,1.9823592,3.3969233,3.882667,4.8377438,5.0609236,4.890257,4.6112823,4.4734364,4.2436924,2.3138463,0.69907695,0.118153855,0.013128206,0.013128206,0.006564103,0.0032820515,0.02297436,0.06235898,0.6432821,2.7076926,2.5993848,0.4397949,0.14441027,0.15753847,0.52512825,0.7122052,0.60389745,0.49230772,0.60061544,0.8730257,1.0272821,1.0305642,1.1060513,0.7581539,1.1290257,1.6968206,2.349949,3.373949,3.4625645,2.937436,2.5304618,2.3040001,1.6475899,2.8717952,2.5862565,2.4352822,2.7142565,2.3663592,3.31159,4.0467696,4.4964104,4.8672824,5.6418467,6.0783596,6.2490263,5.789539,5.0674877,5.1889234,6.1538467,6.747898,7.7325134,8.6580515,7.8506675,7.3452315,7.962257,9.094564,10.177642,10.696206,11.474052,11.818667,11.542975,11.405129,13.128206,12.924719,13.548308,14.043899,14.401642,15.553642,16.111591,15.77354,15.402668,15.596309,16.695797,17.444103,17.319386,16.964924,16.761436,16.853334,16.384,15.169642,14.5263605,14.7331295,15.028514,16.475899,16.42995,16.137848,16.088617,16.019693,15.8884115,16.190361,16.02954,15.067899,13.515489,14.221129,13.935591,13.206975,12.740924,13.407181,14.55918,15.776822,16.416822,16.679386,17.604925,18.786463,18.78318,19.026052,20.201027,22.239182,22.344208,20.94277,19.282053,17.96595,16.951796,17.91672,19.301744,19.67918,19.032618,18.747078,17.992207,18.139898,17.650873,16.088617,14.122667,14.39836,13.748514,12.721231,12.166565,13.22995,12.744206,12.1928215,11.69395,11.851488,13.748514,13.436719,12.179693,10.246565,8.536616,8.582564,8.6580515,8.598975,7.975385,7.056411,6.8004107,7.27959,6.744616,5.3924108,3.9909747,3.889231,3.8334363,3.7120004,3.8498464,4.2436924,4.525949,3.5971284,3.8301542,5.346462,7.529026,9.02236,7.53559,7.637334,8.300308,8.720411,8.329846,7.9425645,8.188719,8.441437,8.786052,10.013539,11.027693,10.738873,10.738873,11.730052,13.50236,10.660104,11.529847,13.279181,13.29559,9.189744,8.247795,8.4283085,8.211693,7.4469748,7.3714876,5.8453336,4.0369234,3.1081028,3.508513,4.9788723,3.314872,3.4100516,3.2000003,2.806154,4.5489235,3.6036925,2.7109745,1.9626669,1.6607181,2.3171284,3.7087183,4.9460516,5.674667,5.98318,6.426257,6.7872825,7.50277,7.2960005,6.235898,5.7632823,5.346462,4.0369234,3.8367183,4.9329233,5.674667,5.428513,5.4580517,5.280821,5.0084105,5.3234878,4.818052,4.594872,4.089436,3.0260515,1.404718,1.6410258,1.522872,1.3850257,1.6278975,2.7076926,2.2777438,2.5961027,2.917744,2.8947694,2.550154,2.9538465,2.609231,1.9528207,1.3653334,1.1618463,1.1684103,1.204513,1.1913847,1.0929232,0.9321026,0.9878975,1.3554872,1.6410258,1.6836925,1.5327181,1.7690258,1.9364104,1.975795,2.100513,2.7995899,3.4625645,4.0992823,4.716308,5.290667,5.7829747,6.5017443,6.616616,6.452513,6.0947695,5.398975,4.972308,4.2502565,3.4921029,2.92759,2.7437952,2.868513,2.2514873,1.7723079,1.7558975,2.0053334,2.0808206,2.3696413,2.7503593,3.0654361,3.1409233,3.058872,3.1048207,3.1474874,3.1277952,3.0785644,3.4297438,3.7940516,3.8038976,3.442872,3.0720003,2.6256413,2.231795,1.9692309,1.7920002,1.5163078,1.4408206,1.4605129,1.4080001,1.276718,1.204513,1.1355898,1.1979488,1.3357949,1.5622566,1.9561027,2.3040001,2.4648206,2.7634873,3.1245131,3.0654361,2.789744,2.2186668,1.6114873,1.214359,1.2668719,1.4112822,1.6082052,1.7624617,1.9823592,2.5895386,2.4943593,2.1530259,1.9364104,1.7526156,1.0601027,1.0338463,1.0272821,1.2471796,1.6410258,1.910154,2.0217438,2.3236926,2.553436,2.806154,3.5511796,3.9384618,4.0008206,4.086154,4.5062566,5.543385,6.2818465,6.422975,6.173539,5.8289237,5.7829747,5.425231,5.5696416,5.346462,4.535795,3.56759,3.6660516,3.5052311,3.629949,4.1780515,4.890257,4.1846156,3.8990772,3.9187696,4.312616,5.330052,5.605744,5.4186673,5.5138464,5.9602056,6.1374364,5.8978467,5.464616,5.2742567,5.3858466,5.4941545,5.0018463,4.919795,5.074052,5.3924108,5.8912826,5.3891287,4.9460516,4.713026,4.7589746,5.0642056,5.10359,5.32677,5.5302567,5.668103,5.8486156,5.402257,5.0642056,4.9788723,5.110154,5.218462,5.159385,5.2512827,5.4580517,5.543385,5.0871797,4.578462,4.4406157,4.5489235,4.824616,5.2315903,5.2447186,5.179077,5.3037953,5.7829747,6.692103,6.882462,7.3025646,7.830975,8.339693,8.713847,8.260923,8.267488,8.687591,8.868103,7.5421543,6.091488,5.431795,4.630975,4.818052,9.212719,11.257437,9.324308,9.084719,11.769437,14.194873,11.936821,13.541744,16.95836,18.710976,13.906053,19.456001,26.069336,26.63713,19.472412,8.346257,10.059488,11.69395,11.654565,13.08554,23.880207,17.742771,10.725744,9.728001,15.399385,22.117744,26.840618,35.55118,35.22954,26.22031,22.235899,44.5998,59.30667,53.84862,31.123695,9.458873,4.772103,4.709744,5.677949,6.23918,7.1187696,3.5446157,3.7152824,4.71959,4.706462,2.8849232,2.8192823,2.7602053,2.6387694,2.4516926,2.231795,2.1070771,2.2514873,2.3860514,2.284308,1.7558975,1.7723079,1.5655385,1.2406155,0.9517949,0.90256417,0.60389745,0.49230772,0.4135385,0.318359,0.29210258,0.24943592,0.33476925,0.47261542,0.58420515,0.58420515,0.508718,0.65969235,0.8730257,1.1388719,1.595077,1.3883078,1.3062565,1.4112822,1.6475899,1.847795,1.4080001,1.5064616,1.8313848,2.0545642,1.8313848,1.5064616,1.6869745,2.0086155,2.2383592,2.2744617,2.3433847,2.3827693,2.4155898,2.5829747,3.1343591,3.5478978,4.141949,4.273231,3.9122055,3.6562054,3.889231,4.6834874,5.3792825,5.8125134,6.301539,6.409847,7.0957956,7.7259493,8.100103,8.4512825,7.9261546,7.565129,7.765334,8.024616,6.941539,5.940513,5.431795,5.4613338,5.9602056,6.73477,6.8004107,6.1374364,5.937231,6.232616,5.87159,6.1374364,6.4032826,6.6428723,6.701949,6.2687182,5.792821,6.3606157,6.7938466,6.51159,5.543385,4.821334,4.9362054,4.57518,3.6036925,3.0391798,3.9286156,3.9286156,3.7710772,3.7973337,3.95159,3.387077,3.2886157,3.2032824,3.1015387,3.370667,3.3805132,3.2787695,3.0916924,2.934154,3.006359,3.1245131,3.0818465,2.9669745,2.8882053,2.9472823,2.9472823,2.5304618,2.2383592,2.169436,1.9692309,2.0841026,2.2711797,2.3269746,2.1956925,1.9889232,1.7132308,1.3095386,1.1126155,1.1979488,1.3883078,7.529026,7.5421543,7.017026,6.422975,6.0192823,5.8518977,5.684513,5.677949,5.832206,6.232616,7.062975,7.7718983,7.463385,6.8496413,6.3442054,6.0652313,6.3212314,6.889026,7.312411,7.4797955,7.643898,7.1122055,6.685539,6.245744,5.861744,5.7698464,5.7403083,5.097026,4.9296412,5.504,6.2490263,6.439385,6.262154,6.038975,5.979898,6.170257,5.98318,6.2063594,7.0334363,8.086975,8.43159,8.907488,9.065026,9.409642,10.164514,11.250873,12.327386,13.735386,13.968411,12.813129,11.369026,10.548513,9.810052,9.639385,9.829744,9.5146675,9.124104,9.120821,9.012513,8.818872,9.074872,8.01477,7.3452315,6.8233852,6.3277955,5.8256416,5.671385,5.4908724,4.9920006,4.1058464,2.9702566,2.162872,1.4736412,0.92225647,0.5349744,0.33805132,0.2231795,0.14441027,0.08861539,0.052512825,0.03938462,0.026256412,0.013128206,0.0032820515,0.0,0.0,0.0,0.026256412,0.026256412,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.016410258,0.06235898,0.6826667,1.910154,3.2820516,3.8301542,4.0500517,4.4274874,4.3716927,4.0434875,4.332308,2.9407182,1.4769232,0.512,0.15425642,0.052512825,0.02297436,0.013128206,0.009846155,0.009846155,0.01969231,0.47261542,2.1136413,2.0939488,0.4660513,0.17723078,0.10502565,0.25271797,0.3446154,0.3117949,0.30851284,0.6104616,0.9321026,1.0765129,1.1257436,1.4342566,1.3981539,1.6935385,1.8445129,1.972513,2.793026,2.9604106,2.7241027,2.6387694,2.6551797,2.1300514,2.9144619,2.9013336,2.8980515,3.1671798,3.4330258,4.972308,5.8256416,6.2162056,6.482052,7.066257,7.2270775,7.752206,7.9425645,7.7981544,7.9983597,8.553026,8.395488,8.864821,9.724719,9.160206,9.088,9.593436,10.112,10.6469755,11.762873,12.137027,11.992617,11.618463,11.61518,12.895181,13.098668,14.034052,14.546052,14.683899,15.701335,16.331488,15.793232,15.110565,14.992412,15.829334,15.419078,16.15754,16.469334,15.980309,15.514257,15.061335,14.516514,14.49354,14.903796,14.9398985,15.983591,15.954053,16.003283,16.426668,16.676104,16.482462,15.911386,15.163078,14.34913,13.459693,14.388514,14.408206,14.027489,13.728822,13.952001,14.076719,14.9628725,15.566771,15.904821,17.06995,18.51077,18.359797,18.392616,19.377232,21.06749,22.390156,22.144001,21.146257,19.790771,18.070976,18.294155,19.603693,20.082872,19.56431,19.61354,19.098257,19.928617,19.67918,17.801847,15.616001,15.793232,15.488001,14.28677,12.842668,12.842668,13.446565,13.348104,12.432411,11.736616,13.459693,13.482668,12.540719,10.998155,9.465437,8.802463,8.851693,8.87795,8.4512825,7.6274877,6.941539,7.4207187,7.0892315,5.914257,4.4406157,3.7842054,3.626667,3.5905645,3.5511796,3.5905645,3.9811285,3.570872,3.692308,4.890257,7.0793853,9.563898,8.379078,7.6209235,7.8539495,8.602257,8.349539,7.8014364,7.6603084,7.778462,8.362667,10.006975,11.001437,10.811078,11.224616,12.448821,13.082257,12.028719,12.455385,12.097642,10.466462,8.851693,8.487385,7.9917955,7.512616,6.8365135,5.4153852,4.2994876,2.8553848,3.239385,5.0215387,5.182359,3.8531284,3.495385,3.0851285,2.6847181,3.43959,4.020513,3.6824617,2.6945643,1.9889232,3.186872,3.7021542,4.2601027,4.6966157,5.0051284,5.3202057,6.514872,6.961231,6.6100516,5.986462,6.173539,5.861744,4.5587697,4.0500517,4.647385,5.218462,4.716308,4.706462,4.670359,4.525949,4.6244106,3.8071797,3.2886157,2.92759,2.4582565,1.4867693,1.5753847,1.3587693,1.1848207,1.3522053,2.1070771,2.4681027,2.6453335,2.9144619,3.2196925,3.1573336,3.4133337,2.681436,2.1202054,1.9954873,1.654154,1.273436,1.1684103,1.1520001,1.0962052,0.9156924,0.97805136,1.2865642,1.4966155,1.529436,1.5786668,1.7362052,1.9265642,2.0217438,2.0808206,2.3696413,3.1507695,4.1780515,5.218462,6.121026,6.8529234,7.076103,6.9349747,6.547693,6.0652313,5.6943593,4.95918,4.0500517,3.2886157,2.7798977,2.412308,2.0775387,1.6082052,1.4998976,1.8609232,2.4385643,2.4024618,2.546872,2.7569232,2.8882053,2.7766156,2.6617439,2.7273848,2.9144619,3.1507695,3.3509746,3.8334363,4.1222568,4.013949,3.5314875,2.92759,2.537026,2.297436,2.0808206,1.8182565,1.4998976,1.3489232,1.339077,1.2865642,1.1946667,1.2274873,1.211077,1.3095386,1.4244103,1.5885129,1.9790771,2.2055387,2.6486156,3.18359,3.5380516,3.2787695,3.0260515,2.3794873,1.8084104,1.4834872,1.2931283,1.404718,1.7493335,1.9692309,2.048,2.297436,2.353231,2.2646155,2.0512822,1.7657437,1.4998976,1.3357949,1.1979488,1.204513,1.3292309,1.404718,1.6311796,1.9823592,2.2646155,2.422154,2.546872,3.511795,3.8071797,3.9975388,4.388103,5.0215387,5.3825645,5.546667,5.421949,5.2545643,5.609026,5.7665644,5.5105643,5.1167183,4.673641,4.07959,3.757949,3.6102567,3.7809234,4.2863593,5.031385,4.4274874,3.8596926,3.698872,4.1846156,5.431795,5.0674877,4.2535386,3.9712822,4.4012313,4.9362054,4.8836927,4.663795,4.57518,4.630975,4.5522056,4.3585644,4.4964104,4.7917953,5.221744,5.937231,5.1265645,4.6276927,4.519385,4.6572313,4.670359,4.6769233,5.3005133,5.730462,5.8781543,6.373744,6.2129235,5.7042055,5.3070774,5.1232824,4.906667,5.037949,5.097026,5.2414365,5.3431797,4.9788723,4.4898467,4.46359,4.578462,4.7392826,5.080616,5.3858466,5.5991797,5.835488,6.235898,6.954667,7.066257,7.2927184,7.6110773,8.01477,8.5202055,8.408616,7.9819493,8.182155,8.65477,7.7456417,6.452513,5.1232824,4.1025643,4.493129,8.146052,9.67877,8.185436,7.683283,9.084719,10.223591,8.533334,10.469745,12.747488,13.410462,11.864616,16.282257,19.39036,18.865232,15.169642,11.565949,10.998155,10.528821,9.133949,8.805744,14.539488,13.239796,10.870154,14.631386,22.99077,25.688618,29.042873,38.334362,37.592617,25.938053,17.588514,25.380104,31.7079,32.768,25.951181,9.833026,6.0783596,8.661334,10.952206,9.826463,5.664821,4.384821,4.7261543,4.9854364,4.3651285,2.9768207,2.9571285,2.6945643,2.5009232,2.4516926,2.3827693,2.1464617,2.156308,2.1398976,1.9331284,1.4703591,1.4441026,1.3193847,1.1355898,0.9321026,0.74830776,0.65312827,0.5546667,0.4594872,0.380718,0.3446154,0.38400003,0.4004103,0.44964105,0.5218462,0.5415385,0.57764107,0.65312827,0.8336411,1.142154,1.5458462,1.2209232,1.1388719,1.1913847,1.3226668,1.529436,1.2373334,1.2373334,1.332513,1.4080001,1.4408206,1.3883078,1.5753847,1.8215386,2.0676925,2.3958976,2.4155898,2.4385643,2.477949,2.6354873,3.0982566,3.3641028,3.876103,3.9614363,3.6824617,3.820308,3.9876926,4.3684106,4.788513,5.1922054,5.6418467,5.9536414,6.616616,7.072821,7.282872,7.7357955,7.712821,7.450257,7.4371285,7.506052,6.810257,6.170257,6.0291286,6.2194877,6.4754877,6.413129,5.9995904,5.664821,5.668103,5.901129,5.85518,6.193231,6.5837955,6.803693,6.629744,5.835488,5.6943593,6.160411,6.5312824,6.373744,5.5072823,4.6605134,4.8147697,4.519385,3.508513,2.7076926,3.6036925,3.387077,2.9078977,2.7536411,3.2623591,2.9440002,2.9144619,2.6551797,2.2613335,2.4484105,3.1376412,3.170462,3.0752823,3.1015387,3.2262566,3.0096412,2.9144619,2.7864618,2.6486156,2.7142565,2.7109745,2.605949,2.3696413,2.044718,1.7788719,1.8215386,1.8740515,1.9035898,1.8412309,1.5556924,1.3620514,1.3620514,1.3620514,1.3193847,1.3751796,7.315693,7.3649235,7.003898,6.6133337,6.2687182,5.737026,5.47118,5.1889234,5.074052,5.3169236,6.12759,6.872616,6.885744,6.567385,6.311385,6.5083084,6.6625648,6.928411,7.1220517,7.2336416,7.4174366,7.1122055,6.7282057,6.547693,6.5772314,6.5706673,6.813539,6.2884107,6.1308722,6.6428723,7.2927184,7.4436927,7.1680007,7.026872,7.1844106,7.433847,7.3682055,7.64718,8.2215395,8.779488,8.736821,9.114257,9.088,9.222565,9.764103,10.660104,11.697231,12.71795,12.868924,12.27159,12.025436,10.79795,10.118565,9.701744,9.383386,9.137232,8.920616,8.982975,9.140513,9.330873,9.577026,8.789334,8.073847,7.3550773,6.6067696,5.83877,5.622154,5.0871797,4.240411,3.1967182,2.169436,1.4244103,0.86974365,0.49230772,0.26584616,0.13784617,0.09189744,0.06235898,0.04266667,0.029538464,0.02297436,0.016410258,0.006564103,0.0,0.0,0.0,0.0,0.026256412,0.026256412,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.02297436,0.46933338,1.5195899,2.7831798,3.318154,3.239385,3.826872,3.8367183,3.245949,3.2525132,1.8313848,0.9124103,0.39384618,0.15425642,0.059076928,0.029538464,0.032820515,0.032820515,0.03938462,0.10502565,0.3249231,1.014154,1.0043077,0.30851284,0.13456412,0.04594872,0.072205134,0.07548718,0.08205129,0.28882053,0.6170257,0.92225647,1.024,1.0568206,1.4703591,1.5819489,1.6246156,1.6016412,1.6377437,1.975795,2.1136413,2.550154,3.0884104,3.3969233,3.0260515,3.0490258,3.2262566,3.370667,3.6562054,4.6112823,6.0225644,6.741334,6.8463597,6.685539,6.889026,6.7938466,7.958975,8.950154,9.278359,9.383386,9.3078985,8.923898,8.920616,9.271795,9.229129,9.938052,10.518975,10.965334,11.523283,12.724514,12.304411,12.225642,12.304411,12.58995,13.37436,13.840411,14.319591,14.578873,14.838155,15.786668,16.075489,15.484719,14.759386,14.401642,14.680616,13.794462,14.739694,15.455181,15.163078,14.391796,13.840411,13.794462,14.368821,15.110565,14.998976,15.337027,15.110565,15.163078,15.67836,16.200207,16.118155,14.792206,13.515489,12.908309,12.898462,13.925745,14.506668,14.811898,14.985847,15.156514,15.074463,15.035078,15.320617,15.954053,16.679386,18.12677,18.323694,18.34995,18.740515,19.498669,20.62113,21.589334,21.910976,21.24472,19.40677,18.980104,19.856411,20.480001,20.36513,20.073027,19.843283,21.730463,22.216208,20.361847,17.818258,17.26031,16.692514,15.504412,13.883078,12.806565,14.070155,14.057027,13.206975,12.63918,14.155488,13.115078,12.521027,11.795693,10.7158985,9.435898,9.232411,9.051898,8.723693,8.178872,7.456821,7.460103,7.0498466,6.042257,4.7228723,3.826872,3.508513,3.4527183,3.4724104,3.5216413,3.7185643,3.6332312,3.882667,4.775385,6.4557953,8.917334,8.556309,7.5552826,7.4830775,8.2904625,8.293744,7.604513,7.1548724,7.13518,7.827693,9.6295395,10.515693,10.417232,11.001437,12.041847,11.434668,11.963078,12.324103,11.145847,9.084719,8.854975,8.635077,8.260923,7.5552826,6.1997952,3.7120004,3.0260515,2.1136413,3.259077,5.7009234,5.6451287,4.1452312,4.240411,4.46359,4.3290257,4.3290257,3.9778464,3.892513,3.2886157,2.553436,3.242667,3.1507695,3.4921029,3.9351797,4.3027697,4.57518,6.1407185,6.121026,5.8518977,5.940513,6.265436,5.9569235,4.7228723,4.010667,4.1911798,4.5522056,4.2305646,4.1911798,4.1058464,3.9384618,3.95159,3.117949,2.5961027,2.2580514,2.034872,1.9068719,1.7033848,1.5031796,1.3554872,1.3489232,1.6180514,2.2219489,2.3926156,2.7011285,3.1442053,3.1638978,3.0490258,2.5435898,2.425436,2.7175386,2.6912823,1.9922053,1.6246156,1.4080001,1.2209232,1.0010257,1.0633847,1.273436,1.4473847,1.5753847,1.8149745,1.9364104,2.0841026,2.2482052,2.3696413,2.353231,2.868513,4.007385,5.2315903,6.2818465,7.171283,7.2336416,6.9645133,6.49518,6.0291286,5.8223596,5.208616,4.3585644,3.5544617,2.8750772,2.2022567,1.6869745,1.394872,1.5031796,1.9659488,2.5173335,2.4713848,2.5993848,2.793026,2.9046156,2.7602053,2.605949,2.7011285,2.9538465,3.3050258,3.7120004,4.132103,4.269949,4.092718,3.56759,2.665026,2.3401027,2.1956925,2.0118976,1.723077,1.4375386,1.4145643,1.4342566,1.4145643,1.3620514,1.3850257,1.339077,1.4736412,1.5524104,1.6016412,1.910154,2.0873847,2.6880002,3.3017437,3.6004105,3.3444104,3.2164104,2.7470772,2.3040001,1.9856411,1.6246156,1.4900514,1.7296412,1.9200002,1.9561027,2.028308,2.0611284,2.2350771,2.1825643,1.913436,1.8018463,1.5655385,1.3817437,1.3128207,1.332513,1.3128207,1.6869745,1.9922053,2.2449234,2.3171284,1.9396925,2.6453335,3.2164104,3.6168208,3.9286156,4.3684106,4.57518,4.896821,4.9952826,4.9526157,5.2611284,5.6976414,5.5007186,5.0838976,4.716308,4.5128207,4.1878977,4.2141542,4.4045134,4.6572313,4.9788723,4.4242053,4.197744,4.2896414,4.7589746,5.737026,4.824616,3.626667,3.1343591,3.5183592,4.1091285,4.8016415,4.6178465,4.240411,3.948308,3.6332312,3.6758976,3.9975388,4.4077954,4.890257,5.586052,4.9099493,4.5423594,4.516103,4.6802053,4.6933336,4.7261543,5.3103595,5.691077,5.8486156,6.485334,6.413129,6.1046157,5.661539,5.169231,4.6769233,4.919795,5.0215387,5.159385,5.3103595,5.2611284,4.926359,4.8607183,4.824616,4.8377438,5.179077,5.5072823,5.8945646,6.1505647,6.3442054,6.7905645,6.954667,7.259898,7.5421543,7.79159,8.136206,8.339693,7.7718983,7.8112826,8.402052,8.080411,6.941539,4.965744,4.0402055,4.8016415,6.636308,7.6931286,6.8233852,6.1013336,6.3474874,7.1483083,6.1046157,7.197539,8.809027,9.557334,8.293744,9.93477,11.053949,11.437949,11.52,12.389745,11.37559,9.875693,6.8299494,4.1813335,6.87918,8.490667,10.289231,17.690258,26.77826,24.336412,21.051079,25.363695,25.002668,18.130053,13.338258,12.977232,14.053744,16.393847,16.456207,7.318975,6.189949,10.84718,13.13477,10.125129,4.132103,4.821334,4.9920006,4.585026,3.767795,2.937436,2.8717952,2.5271797,2.2711797,2.2350771,2.3269746,2.0053334,1.9856411,1.8510771,1.5163078,1.2406155,1.1684103,1.0601027,1.014154,0.98461545,0.79097444,0.8369231,0.7811283,0.65969235,0.52512825,0.42994875,0.41682056,0.380718,0.36758977,0.39056414,0.44964105,0.5349744,0.5907693,0.7581539,1.0305642,1.2537436,1.1093334,1.1388719,1.142154,1.1027694,1.1684103,1.0699488,1.086359,1.0305642,0.9878975,1.3128207,1.394872,1.522872,1.7001027,1.9561027,2.353231,2.3171284,2.4188719,2.540308,2.6945643,3.0293336,3.190154,3.3575387,3.4297438,3.5216413,3.9975388,4.056616,4.1911798,4.450462,4.785231,5.044513,5.4383593,6.0356927,6.436103,6.5969234,6.8266673,7.250052,7.3353853,7.243488,7.138462,7.197539,6.698667,6.2785645,6.173539,6.2555904,6.038975,5.681231,5.7107697,5.8420515,5.9536414,6.0685134,6.3442054,6.560821,6.554257,6.23918,5.61559,5.8847184,6.1472826,6.3967185,6.419693,5.789539,5.024821,4.9296412,4.571898,3.692308,2.7011285,3.2361028,3.0227695,2.3926156,1.913436,2.3893335,2.5206156,2.6256413,2.3926156,1.975795,1.9889232,2.7667694,3.0523078,3.1507695,3.2295387,3.2984617,3.0391798,2.8947694,2.7536411,2.6354873,2.6945643,2.7602053,2.6190772,2.2646155,1.8215386,1.5360001,1.5261539,1.5327181,1.5786668,1.5622566,1.2504616,1.270154,1.3850257,1.4441026,1.404718,1.339077,7.7292314,7.6176414,7.2631803,7.1122055,6.99077,6.091488,5.609026,4.890257,4.5390773,4.7622566,5.3727183,6.235898,6.6133337,6.619898,6.5017443,6.633026,6.442667,6.885744,7.197539,7.1515903,7.056411,7.0498466,6.921847,7.0465646,7.3780518,7.453539,7.4765134,7.430565,7.456821,7.6734366,8.165744,8.251078,8.096821,8.027898,8.195283,8.562873,9.035488,9.458873,9.6065645,9.527796,9.547488,9.69518,9.577026,9.517949,9.590155,9.603283,10.259693,10.660104,10.834052,10.870154,10.896411,10.056206,9.93477,9.668923,9.156924,9.061745,9.409642,9.865847,10.282667,10.463181,10.167795,9.819899,9.084719,8.109949,7.0400004,6.0225644,5.3792825,4.4012313,3.2754874,2.2088206,1.4276924,0.92553854,0.5546667,0.31507695,0.18707694,0.11158975,0.101743594,0.07548718,0.052512825,0.03938462,0.029538464,0.01969231,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.118153855,0.85005134,1.9429746,2.3138463,2.2580514,2.8160002,2.8422565,2.1530259,1.5163078,0.9321026,0.5349744,0.256,0.08205129,0.026256412,0.036102567,0.06564103,0.06235898,0.06564103,0.19692309,0.25928208,0.38400003,0.32164106,0.108307704,0.072205134,0.02297436,0.128,0.14769232,0.16738462,0.5874872,0.6826667,0.93866676,1.0338463,0.98133343,1.1290257,1.1848207,1.1815386,1.5130258,1.9823592,1.8051283,1.7723079,2.5337439,3.3050258,3.6693337,3.570872,3.2984617,3.56759,3.8564105,4.1911798,5.159385,5.937231,6.265436,5.9963083,5.4908724,5.6418467,5.658257,7.2861543,8.592411,8.854975,8.556309,8.316719,8.3823595,8.251078,8.060719,8.615385,9.849437,10.86359,12.114052,13.262771,13.197129,11.930258,12.796719,13.860104,14.227694,14.063591,14.588719,14.408206,14.181745,14.434463,15.55036,14.749539,14.053744,13.748514,13.827283,14.017642,13.574565,13.568001,13.745232,13.787898,13.29559,12.885334,12.86236,13.590976,14.634667,14.792206,14.729847,14.329437,14.001232,13.984821,14.34913,14.450873,13.15118,11.992617,11.749744,12.406155,13.269335,14.36554,15.281232,15.835898,16.09518,16.8599,15.770258,15.455181,16.23631,16.118155,17.67713,18.78318,19.088411,18.730669,18.304,18.185848,19.403488,20.657232,21.06749,20.171488,19.738258,20.20431,20.932924,21.192207,20.168207,20.164925,22.65272,23.899899,22.55754,19.643078,17.972515,16.659693,15.566771,14.50995,13.2562065,14.710155,14.7790785,14.444309,14.6182575,16.121437,12.964104,11.98277,11.782565,11.405129,10.33518,9.619693,9.081436,8.694155,8.402052,8.1066675,7.5946674,7.026872,5.930667,4.5489235,3.8432825,3.5774362,3.367385,3.5249233,3.889231,3.820308,3.511795,4.066462,4.8607183,5.802667,7.3386674,7.6635904,7.0793853,7.1220517,7.8769236,7.968821,7.1089234,6.8299494,6.9021544,7.4010262,8.700719,9.819899,10.003693,10.440206,10.94236,9.941334,10.397539,10.492719,9.668923,8.55959,8.996103,8.470975,8.119796,7.128616,5.2381544,2.7569232,2.284308,2.231795,3.6430771,5.684513,5.6320004,4.089436,4.9821544,6.340924,7.131898,7.276308,3.9056413,3.56759,3.511795,2.8816411,2.7076926,2.878359,3.4034874,3.9745643,4.33559,4.2962055,5.47118,5.1626673,5.3234878,6.160411,6.1374364,5.677949,4.5423594,3.9220517,4.013949,4.010667,4.073026,3.9614363,3.5872824,3.1770258,3.255795,2.986667,2.806154,2.425436,2.0020514,2.1103592,1.7001027,1.6475899,1.5589745,1.3817437,1.4309745,1.6705642,1.9856411,2.3991797,2.7175386,2.537026,2.1267693,2.4451284,2.865231,3.1967182,3.692308,3.0818465,2.487795,1.9429746,1.467077,1.0666667,1.0043077,1.1651284,1.4703591,1.8149745,2.0709746,2.2153847,2.2678976,2.3958976,2.5698464,2.5764105,2.8816411,3.9154875,5.031385,5.920821,6.6133337,6.7938466,6.7314878,6.514872,6.1472826,5.5302567,5.3103595,4.601436,3.692308,2.7798977,1.972513,1.7132308,1.5491283,1.6049232,1.847795,2.097231,2.2646155,2.5435898,2.8488207,3.0654361,3.0523078,2.9210258,3.0326157,3.2525132,3.5249233,3.892513,4.125539,4.076308,3.8432825,3.3509746,2.356513,2.1070771,1.972513,1.7723079,1.5064616,1.3423591,1.5524104,1.6902566,1.723077,1.6672822,1.5786668,1.4998976,1.6311796,1.657436,1.6049232,1.8313848,2.100513,2.6387694,3.1442053,3.4067695,3.314872,3.2295387,3.0490258,2.7273848,2.3433847,2.100513,1.6049232,1.4998976,1.6180514,1.8281027,2.0053334,1.7887181,1.9396925,2.100513,2.0611284,1.7526156,1.6114873,1.4408206,1.3784616,1.4178462,1.401436,1.6869745,1.9495386,2.2449234,2.425436,2.1300514,1.7526156,2.228513,2.7963078,3.2229745,3.8071797,4.1878977,4.5489235,4.7392826,4.7425647,4.6867695,5.0084105,5.3825645,5.179077,4.5489235,4.414359,4.6080003,4.7294364,4.97559,5.2315903,5.0609236,3.9712822,4.269949,4.9132314,5.4416413,5.976616,5.225026,3.9811285,3.4034874,3.751385,4.378257,5.858462,5.290667,4.3716927,3.7776413,3.1540515,3.0818465,3.3969233,4.007385,4.7294364,5.297231,5.0051284,4.821334,4.7491283,4.827898,5.113436,5.218462,5.333334,5.428513,5.6320004,6.265436,6.038975,6.048821,5.8256416,5.2676926,4.6605134,4.824616,5.028103,5.182359,5.330052,5.6320004,5.4941545,5.362872,5.169231,5.0543594,5.3792825,5.474462,5.83877,6.009436,5.9995904,6.301539,6.3934364,6.8594875,7.2960005,7.50277,7.4896417,7.893334,7.788308,7.9950776,8.425026,8.073847,7.3649235,5.4974365,4.59159,4.9329233,4.9821544,5.395693,5.546667,5.654975,5.8256416,6.048821,5.9569235,6.160411,7.7948723,8.717129,3.515077,3.6660516,6.2555904,9.196308,10.916103,10.371283,9.8363085,9.357129,6.226052,2.4910772,4.916513,6.0980515,9.019077,16.272411,23.32554,18.527182,8.444718,6.2687182,7.026872,8.461129,11.011283,10.259693,9.002667,8.625232,8.060719,3.7776413,4.1452312,8.441437,9.537642,6.1308722,2.7503593,4.240411,3.9811285,3.3969233,3.0818465,2.806154,2.5796926,2.2482052,1.9003079,1.7329233,2.041436,1.7165129,1.8084104,1.6804104,1.273436,1.1224617,1.083077,0.9288206,0.88287187,0.955077,0.98461545,0.96492314,0.9682052,0.86974365,0.67282057,0.49887183,0.29538465,0.24943592,0.26256412,0.30194873,0.380718,0.446359,0.52512825,0.6695385,0.83035904,0.892718,1.1093334,1.2668719,1.2307693,1.0404103,0.90256417,0.8992821,1.014154,1.0305642,1.0305642,1.3620514,1.3784616,1.4802053,1.6311796,1.8313848,2.1202054,2.172718,2.4582565,2.7011285,2.8225644,2.9243078,3.058872,2.8816411,2.9505644,3.3969233,3.9056413,3.9220517,4.1189747,4.3749747,4.601436,4.7261543,5.041231,5.464616,5.85518,6.173539,6.449231,7.017026,7.2237954,7.0957956,7.02359,7.778462,7.3058467,6.298257,5.6352825,5.5565133,5.664821,5.467898,5.8092313,6.173539,6.311385,6.2851286,6.6002054,6.6494365,6.380308,5.933949,5.6352825,6.3967185,6.921847,7.1154876,6.875898,6.11118,5.540103,5.0543594,4.5128207,3.8071797,2.8553848,2.92759,2.7306669,2.1497438,1.5491283,1.7591796,2.1989746,2.5140514,2.477949,2.1924105,2.0742567,2.300718,2.7437952,3.0752823,3.18359,3.1770258,3.05559,2.8717952,2.7963078,2.861949,2.986667,2.9210258,2.4516926,1.9593848,1.6246156,1.4211283,1.4473847,1.5392822,1.585231,1.4736412,1.1027694,1.3226668,1.211077,1.2176411,1.3981539,1.4112822,8.438154,8.267488,7.6931286,7.3583593,7.2992826,6.957949,6.262154,5.6943593,5.4186673,5.349744,5.142975,6.0324106,6.5870776,6.76759,6.6592827,6.439385,6.6592827,7.3353853,7.574975,7.128616,6.409847,6.810257,7.53559,8.109949,8.293744,8.086975,7.768616,8.057437,8.65477,9.094564,8.726975,8.618668,9.058462,9.153642,8.78277,8.576,9.905231,10.889847,11.047385,10.709334,11.001437,10.368001,9.760821,9.760821,10.092308,9.6295395,9.93477,9.058462,8.326565,8.27077,8.635077,8.845129,9.189744,9.324308,9.488411,10.512411,11.185231,11.516719,11.890873,11.936821,10.55836,9.938052,9.324308,8.408616,7.204103,6.058667,4.9460516,3.7349746,2.7470772,2.0512822,1.463795,0.90256417,0.52512825,0.2855385,0.17394873,0.19692309,0.23630771,0.20676924,0.14769232,0.07876924,0.029538464,0.01969231,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08205129,0.36430773,0.8369231,1.3718976,1.2865642,1.2307693,1.2668719,1.2964103,1.0535386,0.77128214,0.46276927,0.20020515,0.03938462,0.016410258,0.06564103,0.0951795,0.08205129,0.06564103,0.13784617,0.29538465,0.33476925,0.23958977,0.098461546,0.12143591,0.02297436,0.0,0.0,0.13456412,0.67282057,0.36758977,0.4266667,0.65969235,0.8598975,0.82379496,1.2504616,1.4506668,1.785436,2.1234872,1.8313848,1.9528207,2.359795,2.284308,1.9593848,2.5928206,3.2787695,4.1911798,4.8016415,5.024821,5.2348723,5.405539,5.100308,5.0149746,5.412103,6.117744,7.069539,8.03118,8.342975,7.958975,7.4469748,7.9458466,8.310155,8.303591,8.43159,9.93477,11.362462,12.514462,14.322873,15.599591,13.062565,10.925949,13.092104,15.40595,15.684924,13.732103,14.647796,14.464001,13.801026,13.50236,14.647796,13.610668,12.57354,12.921437,14.431181,15.274668,14.188309,13.403898,12.609642,11.746463,11.001437,11.96636,11.812103,12.294565,13.558155,14.145642,14.267078,13.764924,13.082257,12.458668,11.933539,12.153437,11.723488,11.556104,11.953232,12.58995,13.24636,14.191591,15.051488,15.632411,15.898257,17.38831,16.105026,15.212309,15.327181,14.496821,16.768002,19.265642,20.657232,20.292925,18.218668,17.375181,17.394873,17.785437,18.267899,18.770052,19.085129,20.36513,21.635284,22.084925,21.07077,21.060925,22.905437,24.041027,23.318975,21.011694,17.874052,16.019693,14.87754,14.01436,13.121642,14.769232,15.61272,16.052513,16.62359,17.988924,14.070155,11.756309,11.211488,11.506873,10.604308,9.701744,9.035488,8.503796,8.116513,7.9950776,7.2992826,7.2369237,6.0947695,4.1091285,3.4625645,3.6594875,3.387077,3.442872,3.9417439,4.332308,3.4297438,3.9745643,4.890257,5.58277,5.937231,6.045539,6.0356927,6.298257,6.8693337,7.430565,6.747898,6.87918,7.197539,7.5520005,8.28718,9.980719,10.203898,10.459898,10.94236,10.528821,9.577026,8.5891285,7.5913854,7.1647186,8.421744,8.677744,7.315693,5.796103,4.414359,2.3040001,2.487795,3.43959,5.47118,7.0990777,5.034667,3.948308,5.72718,8.467693,10.86359,12.20595,5.61559,4.5423594,3.82359,2.353231,3.0982566,2.878359,2.934154,3.511795,4.1124105,3.4789746,4.516103,4.70318,5.0149746,5.5762057,5.661539,5.2709746,4.9427695,4.969026,5.0609236,4.3651285,4.240411,4.082872,3.7054362,3.255795,3.2196925,2.7569232,2.612513,2.477949,2.2449234,2.0151796,2.0512822,1.847795,1.5688206,1.4441026,1.785436,2.1530259,1.9856411,2.1202054,2.537026,2.3663592,2.1202054,2.674872,3.186872,3.4724104,3.9975388,3.826872,3.4100516,2.8521028,2.228513,1.5556924,1.3357949,1.4276924,1.7591796,2.0841026,1.9987694,2.169436,2.156308,2.041436,1.9889232,2.2580514,2.9538465,3.9614363,4.9788723,5.7829747,6.2096415,6.2851286,6.7872825,6.9809237,6.49518,5.3103595,5.284103,4.5390773,3.4330258,2.3630772,1.7394873,1.5195899,1.5556924,1.5885129,1.5721027,1.6935385,2.1956925,2.4746668,2.6518977,2.8192823,3.0523078,3.1245131,3.3641028,3.626667,3.8334363,3.9680004,4.0041027,3.7382567,3.4198978,3.0654361,2.4418464,2.3204105,2.2153847,1.9035898,1.4900514,1.404718,1.719795,1.8543591,1.9035898,1.8838975,1.723077,1.723077,1.7427694,1.7132308,1.6738462,1.7690258,2.2449234,2.6584618,3.1048207,3.4724104,3.4494362,3.0687182,2.7011285,2.1956925,1.719795,1.7690258,1.5983591,1.6016412,1.7362052,1.9331284,2.0906668,1.785436,1.6344616,1.7887181,2.0578463,1.9232821,1.654154,1.4572309,1.3981539,1.4998976,1.7558975,1.7165129,1.5622566,1.654154,2.1070771,2.7766156,1.910154,1.6935385,1.9200002,2.3926156,2.930872,3.5511796,3.945026,3.945026,3.7218463,3.7842054,4.1747694,4.857436,5.32677,5.293949,4.6834874,4.525949,4.4045134,4.886975,5.6451287,5.4613338,3.9253337,3.9417439,4.3585644,4.71959,5.280821,5.8289237,4.785231,4.096,4.6112823,6.088206,6.2588725,4.4701543,3.0785644,2.7273848,2.349949,2.5698464,2.8980515,3.6496413,4.6145644,5.0674877,4.772103,4.9460516,5.110154,5.1626673,5.3694363,5.4941545,5.431795,5.333334,5.3005133,5.3858466,5.47118,5.464616,5.3924108,5.2348723,4.9296412,5.0642056,5.106872,5.106872,5.156103,5.402257,5.3398976,5.543385,5.668103,5.661539,5.7829747,5.661539,5.730462,5.7074876,5.72718,6.363898,6.2884107,6.2818465,6.5312824,6.87918,6.806975,7.072821,7.453539,8.050873,8.52677,8.086975,7.3682055,6.1440005,5.074052,4.128821,2.5796926,4.056616,5.3234878,6.4032826,6.9021544,6.012718,5.366154,4.8640003,5.2611284,5.211898,1.2832822,4.466872,6.9021544,8.277334,8.989539,10.161232,7.1122055,9.15036,8.39877,5.024821,7.24677,4.073026,6.009436,13.144616,19.639797,13.718975,5.3070774,3.3050258,4.4832826,7.213949,11.474052,9.974154,8.818872,8.421744,7.7456417,4.3027697,2.4713848,2.7470772,3.2000003,3.0785644,2.8225644,3.9811285,2.9801028,2.156308,2.2678976,2.487795,2.3401027,1.8740515,1.5327181,1.529436,1.847795,1.6377437,1.5425643,1.4080001,1.2570257,1.2832822,1.270154,0.9288206,0.7811283,0.9124103,0.9616411,0.75487185,0.8205129,0.9485129,0.9485129,0.65641034,0.37415388,0.24943592,0.256,0.3446154,0.44307697,0.56451285,0.6695385,0.764718,0.83035904,0.79425645,0.90256417,1.0765129,1.0699488,0.9288206,0.97805136,1.0010257,1.1093334,1.204513,1.2406155,1.1913847,1.1782565,1.3029745,1.4178462,1.4998976,1.6311796,2.231795,2.7569232,3.0982566,3.1671798,2.8980515,2.9472823,2.8488207,2.8324106,3.0030773,3.3575387,3.2951798,3.757949,4.086154,4.201026,4.59159,5.093744,5.172513,5.208616,5.5565133,6.5444107,6.557539,6.304821,6.242462,6.5345645,7.0334363,7.450257,6.774154,6.0980515,5.87159,5.920821,5.3694363,5.297231,5.737026,6.2588725,5.9667697,6.5772314,6.7183595,6.695385,6.626462,6.4557953,7.762052,9.330873,9.412924,7.6996927,5.356308,4.647385,3.9942567,3.3608208,2.930872,3.1113849,2.5862565,2.0086155,1.6738462,1.6246156,1.6475899,2.100513,2.678154,2.8192823,2.5271797,2.3794873,2.1956925,2.3893335,2.8225644,3.2131286,3.1277952,2.7142565,2.6190772,2.6486156,2.7306669,2.9144619,2.1464617,1.9167181,1.8248206,1.7263591,1.7394873,1.7165129,1.7001027,1.6082052,1.394872,1.0535386,1.0765129,0.90912825,0.94523084,1.2635899,1.6180514,8.146052,7.75877,7.4174366,7.174565,7.0104623,6.8365135,6.091488,5.481026,5.152821,5.07077,5.0215387,5.0116925,5.333334,5.76,6.2916927,7.1483083,7.709539,7.781744,7.433847,6.885744,6.5050263,7.3091288,7.8112826,8.316719,8.648206,8.149334,7.8703594,8.195283,8.582564,8.772923,8.789334,8.766359,8.979693,9.222565,9.40636,9.55077,9.875693,10.315488,10.43036,10.397539,11.0145645,10.555078,10.013539,9.842873,10.033232,10.115283,9.826463,8.815591,8.264206,8.464411,8.818872,9.7903595,10.748719,11.044104,11.001437,11.930258,11.858052,12.248616,12.35036,11.697231,10.082462,10.154668,9.252103,8.237949,7.253334,5.717334,4.6145644,3.7349746,2.8980515,2.0775387,1.404718,0.9682052,0.57764107,0.5349744,0.8730257,1.3587693,0.9747693,0.55794877,0.24287182,0.07876924,0.029538464,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.19364104,0.4397949,0.65641034,0.81066674,0.764718,0.77456415,0.88943595,0.9682052,0.67610264,0.5316923,0.38728207,0.20348719,0.036102567,0.03938462,0.13784617,0.1148718,0.068923086,0.052512825,0.07548718,0.32164106,0.3249231,0.21333335,0.11158975,0.14769232,0.068923086,0.20348719,0.20348719,0.0951795,0.28225642,0.25928208,0.4266667,0.6892308,0.90584624,0.90912825,0.7318975,0.9682052,1.4178462,1.785436,1.6968206,2.0841026,2.481231,2.9833848,3.446154,3.4855387,3.9351797,4.841026,5.3760004,5.2447186,4.673641,5.1659493,5.349744,6.0258465,7.138462,7.778462,8.2215395,8.457847,8.362667,8.103385,8.116513,8.28718,8.595693,8.769642,9.156924,10.725744,11.218052,11.631591,12.685129,13.7386675,12.780309,12.842668,13.801026,14.536206,14.713437,14.78236,14.066873,14.913642,15.07118,14.437745,15.038361,14.450873,13.108514,12.278154,12.540719,13.784616,13.059283,12.117334,11.703795,11.523283,10.233437,11.040821,10.5780525,10.35159,10.837335,11.47077,13.302155,14.10954,13.3940525,11.818667,11.175385,10.604308,10.768411,11.316514,11.969642,12.514462,13.476104,14.641232,15.074463,14.762668,14.631386,15.222155,15.212309,15.323898,15.442053,14.631386,16.508718,18.054565,19.295181,20.109129,20.22072,19.311592,18.645334,18.376207,18.057848,16.643284,16.580925,17.32595,18.632206,20.122257,21.267694,20.660515,21.72718,23.56513,24.467693,21.927387,18.271181,15.9573345,14.483693,13.702565,13.8075905,14.427898,16.20677,17.191385,17.289848,18.294155,15.576616,13.341539,12.1928215,11.913847,11.460924,9.764103,9.143796,8.700719,8.057437,7.3485136,6.564103,6.5312824,6.0324106,4.841026,3.69559,2.9144619,2.802872,3.0916924,3.4592824,3.5282054,3.2000003,3.764513,4.585026,5.2315903,5.4580517,5.737026,5.5926156,5.7632823,6.301539,6.5903597,6.2555904,6.8266673,7.515898,8.050873,8.677744,8.897642,9.330873,9.875693,10.295795,10.210463,9.668923,8.15918,7.273026,7.463385,8.057437,8.87795,6.5739493,5.077334,4.788513,2.5600002,2.5961027,2.8914874,3.9154875,5.100308,4.8147697,3.4756925,7.3649235,12.268309,16.23631,19.590565,11.067078,5.287385,2.4516926,2.03159,2.7667694,3.2131286,2.9144619,2.937436,3.43959,3.6758976,5.0051284,5.543385,5.658257,5.7403083,6.196513,5.9536414,5.546667,5.093744,4.7622566,4.778667,4.2469745,4.0500517,3.8301542,3.508513,3.318154,2.806154,2.487795,2.4943593,2.5796926,2.1103592,1.5819489,1.6114873,1.8116925,1.9626669,2.041436,2.4943593,2.28759,2.1136413,2.156308,2.0841026,1.9659488,2.1202054,2.4418464,2.858667,3.314872,3.3575387,3.2196925,3.0523078,2.7536411,1.9954873,1.6475899,1.782154,1.9200002,1.7460514,1.083077,1.020718,1.079795,1.3161026,1.7394873,2.3204105,3.1015387,3.9712822,4.6867695,5.0838976,5.0510774,5.172513,5.681231,6.229334,6.340924,5.4186673,4.818052,4.4242053,3.515077,2.2449234,1.6410258,1.5097437,1.6114873,1.6640002,1.6705642,1.9364104,2.3794873,2.5206156,2.605949,2.7667694,3.0260515,3.3345644,3.4494362,3.5938463,3.7710772,3.761231,3.4658465,3.131077,2.8816411,2.7175386,2.5140514,2.5796926,2.4615386,2.3072822,2.1858463,2.100513,2.172718,2.1366155,2.034872,1.8740515,1.6278975,1.4998976,1.463795,1.3981539,1.3456411,1.4998976,1.9954873,2.4648206,2.8849232,3.1376412,2.9965131,2.3827693,2.1169233,1.9528207,1.8084104,1.7690258,2.3105643,2.6617439,2.605949,2.2219489,1.8838975,2.048,1.9200002,1.6968206,1.5688206,1.7263591,1.7624617,1.6869745,1.6246156,1.6180514,1.6213335,1.7296412,1.5819489,1.5458462,1.7263591,1.9462565,1.8609232,1.8904617,2.0184617,2.2383592,2.550154,3.0260515,3.6102567,3.8071797,3.5774362,3.3444104,3.6758976,3.9122055,4.1682053,4.57518,5.284103,5.5532312,5.5236926,5.362872,5.097026,4.6211286,3.5807183,3.6562054,3.7448208,3.7054362,4.3651285,5.61559,5.4153852,5.0609236,4.785231,3.7316926,4.9985647,4.325744,3.7349746,3.7415388,3.3641028,3.495385,4.1025643,4.7655387,5.0084105,4.309334,4.269949,4.969026,5.674667,5.87159,5.2480006,5.077334,5.208616,5.100308,4.6867695,4.3716927,4.565334,4.529231,4.529231,4.640821,4.7458467,4.900103,5.211898,5.2414365,5.0609236,5.2545643,5.398975,5.5663595,5.6976414,5.7698464,5.796103,5.7009234,6.2194877,6.521436,6.557539,7.0465646,6.875898,6.665847,6.564103,6.6428723,6.892308,7.177847,7.709539,8.103385,8.208411,8.109949,7.939283,7.650462,6.5411286,4.5456414,2.225231,2.7241027,2.9046156,3.121231,3.82359,5.5597954,3.692308,3.3280003,4.266667,4.713026,1.2832822,7.9458466,8.694155,7.6668725,7.02359,6.9152827,7.778462,5.464616,3.255795,3.4002054,7.125334,4.460308,5.100308,9.741129,13.889642,7.8703594,3.7382567,5.6320004,7.1220517,6.7577443,8.070564,7.7292314,7.6209235,8.3823595,8.779488,5.7074876,3.876103,3.9384618,4.647385,4.972308,4.07959,3.4921029,2.9768207,2.3827693,1.8609232,1.8773335,2.0151796,1.6672822,1.4736412,1.5688206,1.6016412,1.6869745,1.5819489,1.332513,1.0732309,1.0502565,0.93866676,0.74830776,0.80738467,1.0043077,0.79097444,0.62030774,0.63343596,0.82379496,0.9878975,0.7056411,0.38400003,0.30194873,0.3511795,0.446359,0.5021539,0.5677949,0.5546667,0.6662565,0.8730257,0.90256417,1.0732309,1.0108719,0.88943595,0.88943595,1.2209232,1.0994873,1.079795,1.2471796,1.4408206,1.2635899,1.2504616,1.3751796,1.6147693,1.7985642,1.6213335,1.9364104,2.5271797,2.8225644,2.7011285,2.5206156,2.6683078,2.674872,2.7864618,2.9111798,2.5993848,3.623385,3.9876926,3.9811285,4.082872,4.972308,5.179077,5.3234878,5.297231,5.280821,5.7534366,5.832206,5.861744,6.058667,6.439385,6.813539,7.6012316,7.5979495,6.774154,5.786257,5.979898,5.6385646,5.366154,5.5991797,6.157129,6.235898,6.4754877,6.4656415,6.8955903,7.9524107,9.324308,10.259693,9.6065645,7.9852314,5.8190775,3.318154,3.6069746,2.8192823,2.3860514,2.8488207,3.882667,2.8488207,1.7624617,1.339077,1.5556924,1.6475899,2.0906668,2.5206156,2.8521028,2.9702566,2.733949,2.540308,2.4681027,2.409026,2.3794873,2.5304618,2.2613335,2.5698464,2.9768207,3.062154,2.4615386,1.9167181,1.7526156,1.8084104,1.9528207,2.0808206,1.8806155,1.6475899,1.404718,1.2438976,1.3226668,1.1126155,0.88615394,0.88615394,1.1323078,1.3981539,7.716103,7.1515903,6.7577443,6.426257,6.1768208,6.183385,5.917539,5.540103,5.3694363,5.405539,5.3202057,5.0215387,5.2578464,5.6418467,6.0160003,6.436103,6.547693,6.6395903,6.882462,7.131898,6.941539,7.75877,8.3134365,8.684308,8.621949,7.5487185,7.64718,7.6176414,7.5487185,7.6570263,8.300308,8.887795,9.012513,9.088,9.334154,9.787078,9.93477,10.082462,10.016821,9.882257,10.210463,10.279386,10.151385,10.013539,9.885539,9.6065645,9.380103,8.684308,8.346257,8.52677,8.720411,10.223591,11.428103,12.074668,12.258463,12.42913,12.143591,12.803283,12.685129,11.503591,10.394258,10.476309,9.330873,8.113232,7.0334363,5.346462,4.562052,3.8071797,2.986667,2.166154,1.5819489,1.0305642,1.0502565,1.7591796,2.553436,2.1070771,1.0666667,0.4594872,0.16082053,0.059076928,0.03938462,0.04594872,0.01969231,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.098461546,0.24615386,0.38728207,0.47917953,0.5316923,0.5513847,0.6071795,0.64000005,0.48902568,0.44307697,0.3708718,0.24287182,0.12471796,0.17394873,0.17394873,0.1148718,0.068923086,0.07876924,0.17066668,0.3511795,0.35774362,0.25928208,0.15097436,0.14441027,0.049230773,0.108307704,0.1148718,0.049230773,0.08205129,0.23302566,0.37743592,0.5349744,0.6465641,0.56451285,0.6301539,0.8402052,1.0633847,1.3850257,2.103795,2.2088206,2.428718,2.9472823,3.6430771,4.082872,3.698872,4.516103,5.2611284,5.602462,6.1440005,6.298257,6.196513,6.3934364,6.9054365,7.204103,6.9809237,7.253334,7.4896417,7.7456417,8.661334,9.110975,9.682052,9.780514,9.800206,11.116308,11.293539,11.595488,11.58236,11.257437,11.063796,12.632616,13.604104,14.004514,13.899488,13.397334,13.446565,14.106257,14.611693,14.788924,15.05477,14.716719,13.216822,11.69395,10.857026,10.978462,11.303386,11.211488,10.873437,10.354873,9.6295395,9.708308,9.353847,9.255385,9.5606165,9.869129,11.805539,13.124924,12.826258,11.460924,11.132719,11.008,10.925949,11.162257,11.651283,11.992617,13.574565,15.117129,15.599591,15.156514,15.07118,16.026258,16.410257,16.55795,16.531694,16.128002,17.302977,17.683693,17.929848,18.57313,20.007385,19.70872,20.38154,20.424206,19.265642,17.368616,17.624617,17.394873,18.021746,19.236105,19.14749,20.118977,20.473438,21.080618,21.185642,18.402462,16.229744,14.490257,13.482668,13.029744,12.475078,12.688411,15.780104,17.690258,17.529438,17.56554,15.55036,14.424617,13.945437,13.607386,12.632616,10.469745,9.747693,9.176616,8.208411,7.0400004,6.5280004,6.3868723,6.0947695,5.47118,4.670359,3.2131286,2.8422565,3.0851285,3.4724104,3.5544617,3.5413337,3.9154875,4.4734364,5.034667,5.4416413,5.172513,4.8705645,4.896821,5.2020516,5.32677,5.412103,6.2063594,7.059693,7.8080006,8.763078,9.094564,9.688616,10.174359,10.308924,9.947898,9.032206,7.6668725,6.7905645,6.957949,8.329846,7.6701546,5.2053337,3.5314875,3.1015387,2.2219489,2.5665643,2.6157951,4.332308,6.51159,4.788513,3.0851285,5.7140517,11.001437,16.01641,16.577642,10.177642,5.277539,2.7963078,2.4057438,2.5304618,2.7536411,3.0030773,3.117949,3.1474874,3.367385,4.46359,4.923077,5.366154,6.0980515,7.1023593,6.5936418,5.674667,4.926359,4.585026,4.516103,3.9844105,4.1091285,4.076308,3.748103,3.6627696,3.31159,2.6945643,2.4155898,2.5074873,2.428718,1.6640002,1.6935385,2.048,2.228513,1.719795,2.1891284,2.3466668,2.2055387,2.0053334,2.1956925,2.228513,2.284308,2.6486156,3.1803079,3.2984617,3.1113849,3.2131286,3.1442053,2.7076926,1.9790771,1.8346668,1.8281027,1.7624617,1.5130258,1.0272821,0.827077,0.82379496,1.0962052,1.6508719,2.425436,3.2754874,3.9712822,4.453744,4.7425647,4.926359,4.9952826,5.5302567,6.189949,6.452513,5.612308,4.9394875,4.3684106,3.5446157,2.540308,1.8543591,1.7001027,1.7263591,1.7263591,1.7099489,1.8904617,2.162872,2.3072822,2.412308,2.5206156,2.6289232,2.9505644,3.05559,3.1540515,3.2918978,3.3247182,3.1343591,2.8914874,2.7273848,2.7175386,2.8914874,2.8455386,2.6880002,2.5764105,2.5632823,2.5928206,2.802872,2.7733335,2.484513,2.0873847,1.913436,1.8412309,1.6935385,1.5622566,1.5392822,1.7165129,2.0512822,2.4582565,2.8225644,2.917744,2.4155898,1.7690258,1.6049232,1.6508719,1.7887181,2.0250258,2.4910772,2.6256413,2.5304618,2.231795,1.7033848,1.654154,1.6738462,1.5885129,1.4506668,1.5589745,1.7558975,1.8281027,1.8051283,1.7460514,1.7165129,1.5688206,1.4309745,1.3981539,1.4572309,1.4998976,1.595077,1.6902566,1.8313848,2.03159,2.2646155,2.6387694,3.0785644,3.2886157,3.2164104,3.0424619,3.1638978,3.3575387,3.7251284,4.33559,5.2480006,5.408821,5.2742567,5.179077,5.041231,4.3716927,4.073026,4.378257,4.2535386,3.69559,3.751385,4.709744,5.106872,5.2578464,5.0576415,4.0041027,3.9975388,3.4625645,3.4855387,4.1189747,4.3749747,4.457026,4.33559,4.4242053,4.604718,4.240411,4.4767184,4.8738465,5.113436,5.179077,5.3727183,4.7425647,4.4701543,4.352,4.2502565,4.092718,4.1222568,4.1222568,4.3585644,4.6802053,4.4996924,4.4800005,4.594872,4.7622566,4.9985647,5.4383593,5.4580517,5.5729237,5.8125134,6.121026,6.3474874,6.3277955,6.7249236,6.675693,6.2063594,6.2555904,6.3901544,6.2851286,6.173539,6.311385,6.9842057,7.4404106,8.2904625,8.556309,8.096821,7.5881033,7.243488,7.5552826,7.5421543,6.629744,4.663795,4.3618464,4.3290257,4.6900516,5.0609236,4.5587697,2.993231,2.8258464,4.125539,5.297231,3.058872,9.521232,11.83836,8.664616,3.2886157,3.6332312,4.962462,3.623385,2.1858463,2.6026669,6.1997952,4.7950773,4.965744,6.8529234,8.018052,3.4625645,3.3050258,6.2063594,7.5421543,6.695385,7.069539,5.9667697,6.5805135,8.556309,10.102155,7.9885135,5.7468724,6.774154,7.062975,5.5926156,4.3290257,3.6857438,3.2787695,2.605949,1.7558975,1.4145643,1.585231,1.5064616,1.4441026,1.4834872,1.5425643,1.4375386,1.4998976,1.4145643,1.148718,0.96492314,0.82379496,0.64000005,0.67610264,0.83035904,0.6301539,0.5218462,0.5513847,0.65312827,0.72861546,0.65312827,0.49887183,0.4201026,0.5152821,0.6859488,0.6465641,0.6826667,0.7122052,0.78769237,0.8763078,0.86646163,1.0568206,1.0436924,0.955077,0.94523084,1.2077949,1.086359,0.9485129,0.9747693,1.0994873,1.017436,1.0338463,1.1881026,1.4736412,1.8018463,1.9922053,2.2580514,2.7437952,3.1048207,3.2098465,3.131077,3.3444104,3.4067695,3.4166157,3.2951798,2.7667694,3.3805132,3.6332312,3.892513,4.342154,5.0116925,4.9329233,4.916513,4.854154,4.821334,5.0674877,5.3202057,5.7140517,6.1407185,6.514872,6.76759,6.928411,7.0465646,6.4754877,5.5958977,5.805949,5.730462,5.674667,5.7042055,5.8912826,6.311385,7.0859494,6.9021544,7.177847,8.579283,11.021129,9.796924,7.3091288,5.0510774,3.5741541,2.4681027,2.4352822,2.0742567,2.169436,2.878359,3.7349746,2.5698464,1.4933335,1.1224617,1.4408206,1.8215386,2.5632823,2.7733335,2.7700515,2.733949,2.7142565,2.6584618,2.5304618,2.5140514,2.6387694,2.7733335,2.5435898,2.6880002,2.865231,2.7733335,2.1497438,1.7558975,1.7165129,1.8543591,2.0545642,2.294154,2.2121027,1.8838975,1.5491283,1.3817437,1.4998976,1.2800001,1.0699488,0.96492314,1.0075898,1.1782565,7.1056414,6.452513,6.1341543,5.8289237,5.5171285,5.467898,5.4514875,5.3366156,5.4580517,5.789539,5.940513,5.5893335,5.5565133,5.602462,5.618872,5.6254363,5.5762057,5.7435904,6.2687182,6.8988724,6.9842057,7.8145647,8.661334,9.160206,8.986258,7.830975,7.512616,7.062975,6.747898,6.8299494,7.5618467,8.241231,8.480822,8.730257,9.176616,9.77395,9.924924,9.875693,9.642668,9.350565,9.235693,9.275078,9.179898,9.104411,9.015796,8.704,8.779488,8.346257,8.234667,8.602257,8.956718,10.548513,11.841642,12.790154,13.321847,13.321847,13.170873,13.6467705,13.239796,11.963078,11.332924,10.610872,9.242257,8.01477,6.9743595,5.4383593,4.854154,4.013949,3.1803079,2.4943593,1.9528207,1.6804104,2.0644104,3.0490258,3.6463592,1.9396925,0.7581539,0.3446154,0.21989745,0.13456412,0.068923086,0.059076928,0.03938462,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.07876924,0.22646156,0.45620516,0.56123084,0.5218462,0.44964105,0.40369233,0.37743592,0.36758977,0.30851284,0.23302566,0.18051283,0.18707694,0.13784617,0.09189744,0.07876924,0.12471796,0.256,0.36430773,0.33476925,0.30851284,0.2986667,0.20348719,0.068923086,0.08205129,0.09189744,0.052512825,0.016410258,0.23630771,0.32164106,0.39384618,0.45292312,0.4004103,0.7450257,0.8467693,0.90912825,1.2307693,2.2121027,2.1497438,2.353231,2.8488207,3.5380516,4.210872,3.6496413,4.1058464,4.70318,5.277539,6.373744,6.47877,6.1768208,6.183385,6.3967185,5.910975,5.622154,6.3343596,7.128616,7.8473854,9.101129,9.527796,10.043077,10.164514,10.148104,10.994873,11.126155,11.795693,11.88759,11.506873,11.972924,13.039591,13.643488,13.784616,13.456411,12.665437,12.694975,12.517745,12.87877,13.522053,13.193847,13.348104,12.609642,11.418258,10.249847,9.590155,9.95118,10.315488,10.049642,9.334154,9.199591,8.851693,8.769642,8.907488,9.101129,9.068309,10.594462,12.20595,12.714667,12.087796,11.444513,11.457642,11.277129,11.349334,11.769437,12.2847185,14.10954,15.356719,15.724309,15.563488,15.885129,16.784412,17.18154,17.316103,17.335796,17.319386,17.923283,17.847795,17.604925,17.824821,19.249231,19.728413,20.545643,20.854155,20.496412,19.99754,19.754667,18.550156,18.41559,18.95713,17.352207,18.313848,18.169437,17.94954,17.378464,14.874257,14.296617,13.426873,12.829539,12.475078,11.730052,11.684103,14.887385,17.32595,17.513027,16.479181,15.189335,14.985847,15.186052,15.153232,14.293334,11.556104,10.436924,9.662359,8.562873,7.076103,6.8266673,6.426257,6.1013336,5.874872,5.5729237,3.8859491,3.2656412,3.2820516,3.508513,3.5478978,3.7087183,4.092718,4.309334,4.5062566,5.3431797,4.768821,4.2896414,4.2174363,4.4045134,4.2502565,4.7360005,5.5105643,6.3376417,7.2336416,8.490667,9.409642,10.220308,10.663385,10.518975,9.6065645,8.67118,6.892308,5.602462,5.5958977,7.1220517,5.3431797,3.6857438,2.6617439,2.3893335,2.612513,2.7175386,2.7864618,4.7491283,7.0793853,4.7950773,2.8816411,3.31159,6.8463597,10.935796,9.724719,6.3606157,4.1156926,2.8816411,2.4320002,2.4188719,2.550154,3.0326157,3.3280003,3.3476925,3.4756925,4.2830772,4.8738465,5.504,6.2523084,7.02359,6.5083084,5.428513,4.6802053,4.4307694,4.082872,3.7349746,4.1583595,4.322462,4.0008206,3.7776413,3.623385,2.993231,2.4516926,2.3269746,2.6912823,2.1267693,1.9495386,2.1103592,2.2121027,1.5392822,1.8904617,2.1464617,2.1333334,2.034872,2.4057438,2.2416413,2.294154,2.809436,3.3903592,2.9997952,2.7470772,2.9801028,3.0194874,2.6453335,2.0873847,1.8215386,1.657436,1.4998976,1.3062565,1.0765129,1.0732309,1.1323078,1.3850257,1.9068719,2.681436,3.508513,4.2240005,4.709744,4.9887185,5.2315903,5.1200004,5.4153852,5.681231,5.5926156,4.9526157,4.8082056,4.332308,3.6758976,2.9505644,2.2088206,1.9298463,1.8609232,1.785436,1.6804104,1.719795,2.0151796,2.2121027,2.3368206,2.3958976,2.353231,2.5928206,2.7602053,2.8553848,2.917744,3.0358977,3.062154,2.9472823,2.8258464,2.8324106,3.0982566,3.1081028,3.0523078,3.0391798,3.117949,3.2656412,3.5971284,3.6168208,3.3280003,2.917744,2.7437952,2.5764105,2.2908719,2.044718,1.9331284,1.9790771,2.1956925,2.5173335,2.8324106,2.865231,2.1858463,1.5163078,1.3193847,1.3850257,1.5753847,1.8248206,2.0841026,2.1202054,2.0545642,1.9003079,1.5819489,1.2668719,1.2865642,1.3554872,1.3686155,1.3883078,1.4998976,1.6377437,1.7033848,1.6935385,1.6968206,1.4867693,1.4375386,1.4572309,1.4473847,1.3062565,1.4605129,1.5524104,1.7099489,1.9331284,2.100513,2.3860514,2.6190772,2.7569232,2.7963078,2.7798977,2.7175386,2.7766156,3.1343591,3.8400004,4.7917953,4.9296412,4.778667,4.778667,4.844308,4.3716927,4.5456414,4.95918,4.7622566,4.069744,3.9811285,4.263385,4.7228723,4.972308,4.8804107,4.5587697,4.210872,3.8301542,3.7973337,4.1517954,4.601436,4.916513,4.384821,4.0336413,4.1156926,4.1091285,4.59159,4.8147697,4.709744,4.6276927,5.349744,4.8049235,4.204308,4.0402055,4.2929235,4.414359,4.013949,4.096,4.6080003,5.1659493,5.034667,4.8607183,4.594872,4.7327185,5.2742567,5.6943593,5.8518977,6.311385,6.6002054,6.672411,6.9152827,6.813539,6.8660517,6.4689236,5.76,5.6287184,5.868308,5.7829747,5.8453336,6.311385,7.197539,7.525744,8.352821,8.677744,8.162462,7.141744,6.810257,7.3649235,8.001641,8.001641,6.744616,6.0061545,6.1472826,6.5936418,6.4295387,4.4077954,2.7241027,3.2886157,4.7261543,5.3431797,3.0949745,8.418462,11.52,8.018052,1.3357949,2.7044106,2.9604106,2.681436,2.0578463,2.0841026,4.5554876,3.5577438,3.692308,3.948308,3.3903592,1.1848207,3.7120004,5.618872,6.0750775,5.677949,6.449231,5.543385,5.61559,7.076103,8.976411,9.015796,7.384616,9.153642,9.117539,6.616616,5.549949,4.4340515,3.5282054,2.6387694,1.7887181,1.2242053,1.273436,1.3718976,1.404718,1.3981539,1.5031796,1.3128207,1.3718976,1.394872,1.2603078,1.020718,0.88615394,0.72861546,0.6629744,0.65969235,0.5677949,0.4955898,0.5316923,0.56123084,0.571077,0.65312827,0.6071795,0.48574364,0.5152821,0.65969235,0.6170257,0.65969235,0.77456415,0.84348726,0.82379496,0.7450257,0.8041026,0.8172308,0.8172308,0.8533334,0.9714873,0.8730257,0.7253334,0.7220513,0.8467693,0.8763078,0.98133343,1.2832822,1.6311796,1.975795,2.3401027,2.5731285,2.934154,3.3509746,3.7218463,3.9056413,4.141949,4.076308,3.8400004,3.5216413,3.1638978,3.2295387,3.4527183,3.817026,4.2502565,4.6276927,4.562052,4.417641,4.3716927,4.466872,4.59159,5.0543594,5.5663595,5.9536414,6.2227697,6.547693,6.0816417,5.920821,5.8256416,5.868308,6.419693,5.970052,5.7140517,5.6352825,5.7435904,6.0849237,7.1056414,7.0957956,7.1581545,7.8112826,8.982975,7.322257,5.858462,4.7458467,3.95159,3.249231,2.7175386,2.281026,2.2646155,2.612513,2.8947694,2.0906668,1.3029745,1.020718,1.3259488,1.9003079,2.9144619,3.0096412,2.6945643,2.3368206,2.169436,2.3827693,2.3171284,2.3433847,2.5304618,2.6715899,2.5961027,2.6289232,2.605949,2.4516926,2.172718,1.8838975,1.8346668,1.8412309,1.8970258,2.1530259,2.2121027,2.048,1.785436,1.5556924,1.4998976,1.3161026,1.214359,1.1224617,1.0568206,1.1355898,6.416411,5.8420515,5.717334,5.546667,5.2053337,4.9132314,4.768821,4.7392826,5.074052,5.6976414,6.23918,6.045539,5.7501545,5.464616,5.333334,5.540103,5.8453336,6.042257,6.23918,6.491898,6.813539,7.650462,8.667898,9.396514,9.511385,8.832001,7.5191803,6.770872,6.4656415,6.5017443,6.806975,7.072821,7.5487185,8.185436,8.838565,9.275078,9.330873,9.189744,8.963283,8.684308,8.320001,7.8703594,7.5454364,7.5585647,7.837539,8.03118,8.306872,8.044309,8.260923,9.094564,9.7903595,11.044104,12.084514,12.964104,13.650052,14.027489,14.263796,14.27036,13.696001,12.750771,12.199386,10.47959,9.173334,8.1755905,7.24677,6.0028725,5.3694363,4.33559,3.5183592,3.062154,2.6617439,3.1113849,3.7218463,4.2502565,3.8629746,1.1323078,0.33476925,0.28882053,0.33476925,0.21333335,0.08533334,0.03938462,0.04594872,0.03938462,0.013128206,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03938462,0.18707694,0.5481026,0.5973334,0.5021539,0.36102566,0.26912823,0.28882053,0.25928208,0.18707694,0.15097436,0.14112821,0.06564103,0.055794876,0.055794876,0.09189744,0.16082053,0.24287182,0.318359,0.26912823,0.3314872,0.47917953,0.4135385,0.23302566,0.27897438,0.23630771,0.07548718,0.04266667,0.24943592,0.29538465,0.32164106,0.39712822,0.4955898,0.90256417,0.8992821,0.94523084,1.2537436,1.7690258,1.8313848,2.2711797,2.8914874,3.498667,3.8990772,3.9122055,3.8400004,3.9844105,4.4242053,5.024821,5.395693,5.402257,5.7731285,6.166975,5.169231,5.4449234,6.2588725,7.0793853,7.827693,8.884514,9.055181,9.458873,9.7903595,10.029949,10.433641,10.594462,11.785847,12.970668,13.830565,14.759386,14.14236,14.063591,13.850258,13.354668,12.941129,12.064821,11.113027,10.998155,11.372309,10.617436,11.260718,11.497026,11.1064625,10.328616,9.878975,9.449026,9.622975,9.485129,8.973129,8.891078,8.625232,8.786052,8.966565,8.946873,8.687591,9.970873,11.802258,13.138052,13.331694,12.12718,11.59877,11.444513,11.602052,12.1238985,13.174155,14.815181,15.058052,14.976001,15.228719,16.032822,16.308514,16.790976,17.201233,17.414566,17.45395,17.732924,17.93313,18.031591,18.228514,18.94072,19.833437,19.314873,19.426462,20.755693,22.436104,21.090464,19.505232,18.983387,18.976822,17.10277,16.088617,15.504412,15.264822,14.838155,13.239796,13.53518,13.331694,12.908309,12.527591,12.409437,11.979488,14.03077,16.28554,17.073233,15.337027,14.946463,15.350155,15.940925,16.28554,16.121437,12.777026,11.047385,10.029949,9.02236,7.53559,7.3058467,6.432821,5.933949,6.0192823,6.114462,4.650667,3.8859491,3.5807183,3.4756925,3.2984617,3.5249233,4.082872,4.013949,3.6857438,4.8082056,4.6178465,4.0303593,3.9023592,4.141949,3.6857438,4.3027697,4.900103,5.618872,6.6133337,8.057437,9.235693,10.35159,10.886565,10.469745,8.871386,8.536616,5.943795,4.132103,4.027077,4.46359,2.9111798,2.4648206,2.9997952,3.9154875,4.1517954,3.1048207,3.4198978,4.7228723,5.796103,4.59159,2.917744,1.9987694,3.0687182,4.903385,3.82359,2.7864618,2.412308,2.1234872,1.8707694,2.1530259,2.5928206,2.8947694,3.2918978,3.7448208,3.9712822,4.7360005,5.5926156,6.0160003,6.0061545,6.088206,5.792821,5.037949,4.5062566,4.269949,3.7776413,3.56759,4.013949,4.309334,4.141949,3.6758976,3.5774362,3.2361028,2.7766156,2.5009232,2.917744,2.7273848,2.2744617,1.9954873,1.9462565,1.7985642,1.8707694,1.8182565,1.8904617,2.15959,2.5140514,2.0053334,2.048,2.6256413,3.1507695,2.4320002,2.4320002,2.6157951,2.7437952,2.678154,2.3794873,1.7001027,1.4473847,1.3259488,1.1979488,1.1027694,1.4375386,1.6377437,1.8806155,2.28759,2.9210258,3.7251284,4.529231,5.100308,5.3694363,5.435077,5.159385,5.142975,4.84759,4.2272825,3.7218463,4.07959,4.010667,3.6758976,3.1803079,2.5435898,2.1530259,2.0250258,1.9068719,1.7427694,1.7033848,2.097231,2.3236926,2.4549747,2.5074873,2.425436,2.5665643,2.7798977,2.878359,2.8849232,3.0654361,3.318154,3.3345644,3.245949,3.1737437,3.2361028,3.446154,3.5774362,3.69559,3.8498464,4.06318,4.3618464,4.394667,4.276513,4.07959,3.8498464,3.515077,3.1770258,2.8455386,2.553436,2.359795,2.5337439,2.7273848,2.930872,2.934154,2.3368206,1.654154,1.3095386,1.2209232,1.2471796,1.1946667,1.3357949,1.5556924,1.5721027,1.4112822,1.4211283,1.1290257,1.0043077,1.0371283,1.142154,1.1651284,1.1848207,1.3423591,1.4605129,1.4966155,1.5556924,1.5261539,1.5885129,1.6344616,1.591795,1.401436,1.5688206,1.591795,1.6968206,1.9003079,2.0151796,2.2088206,2.4352822,2.5698464,2.612513,2.674872,2.4549747,2.2153847,2.3466668,2.9801028,3.9581542,4.4865646,4.6900516,4.6802053,4.565334,4.4340515,4.781949,5.041231,4.785231,4.332308,4.7491283,4.493129,4.588308,4.532513,4.312616,4.414359,5.3103595,5.504,5.152821,4.6572313,4.6539493,4.854154,4.4077954,4.023795,3.9187696,3.8137438,4.194462,4.562052,4.6572313,4.650667,5.1331286,5.0018463,4.414359,4.2240005,4.5587697,4.8049235,4.1485133,4.3552823,4.955898,5.605744,6.0717955,5.87159,5.2709746,5.211898,5.7009234,5.8289237,6.4000006,7.4108725,7.6143594,7.056411,7.076103,6.770872,6.5083084,6.0356927,5.5204105,5.549949,5.536821,5.3070774,5.5630774,6.416411,7.387898,7.318975,7.79159,8.277334,8.224821,7.062975,7.062975,7.4830775,7.890052,7.939283,7.3616414,6.5083084,6.8693337,7.1056414,6.6034875,5.4974365,2.7864618,3.820308,4.854154,4.056616,1.5031796,5.4449234,7.2205133,5.172513,1.8609232,4.0434875,2.993231,2.2383592,1.6246156,1.4539489,2.477949,1.2504616,1.5130258,1.4408206,0.83035904,1.0896411,4.3749747,4.6867695,4.0041027,3.9909747,5.9995904,5.8157954,4.532513,4.1550775,5.366154,7.5388722,8.077128,10.541949,10.44677,7.8112826,7.141744,4.8607183,3.3247182,2.3663592,1.7624617,1.2209232,1.1585642,1.3193847,1.4211283,1.4145643,1.4867693,1.4145643,1.3095386,1.270154,1.2603078,1.079795,1.0043077,0.9156924,0.7778462,0.64000005,0.62030774,0.54482055,0.5349744,0.5874872,0.6695385,0.7417436,0.67938465,0.5152821,0.4201026,0.44307697,0.5152821,0.57764107,0.67938465,0.72861546,0.69251287,0.5940513,0.46276927,0.42338464,0.49230772,0.61374366,0.63343596,0.55794877,0.508718,0.6235898,0.8533334,0.9419488,1.1585642,1.6147693,2.0118976,2.2678976,2.5435898,2.7536411,3.0687182,3.4691284,3.9154875,4.3618464,4.5554876,4.276513,3.8071797,3.4133337,3.314872,3.3345644,3.56759,3.7054362,3.754667,4.0336413,4.1222568,3.9220517,3.9122055,4.141949,4.2535386,4.8705645,5.277539,5.405539,5.504,6.114462,5.654975,5.074052,5.346462,6.5050263,7.653744,6.449231,5.6287184,5.549949,5.930667,5.835488,6.245744,6.810257,7.145026,6.7774363,5.1232824,4.965744,6.3868723,7.076103,6.2555904,4.663795,4.1156926,3.1967182,2.4943593,2.1497438,1.847795,1.657436,1.273436,1.0732309,1.2406155,1.7788719,2.9472823,3.1770258,2.8717952,2.3105643,1.6475899,2.0118976,2.044718,1.9692309,1.9659488,2.1464617,2.28759,2.425436,2.425436,2.3171284,2.3269746,2.166154,2.0118976,1.8084104,1.6475899,1.7887181,1.8510771,2.0250258,1.9790771,1.6902566,1.4408206,1.3062565,1.3292309,1.3029745,1.2242053,1.3029745,5.8912826,5.671385,5.4416413,5.179077,4.8640003,4.4865646,4.3027697,4.0369234,4.1583595,4.650667,5.0051284,5.504,5.684513,5.6976414,5.832206,6.514872,7.066257,7.5881033,7.716103,7.522462,7.522462,7.9491286,8.3593855,8.749949,8.966565,8.697436,7.3550773,6.5050263,6.0717955,5.986462,6.196513,6.6100516,7.2172313,7.565129,7.529026,7.3091288,7.24677,7.3419495,7.453539,7.463385,7.2927184,7.000616,7.1187696,7.4240007,7.8014364,8.241231,8.349539,8.579283,9.4457445,10.656821,11.109744,11.864616,11.723488,11.749744,12.11077,12.084514,12.928001,13.210258,13.075693,12.58995,11.749744,10.223591,9.813334,9.107693,7.7718983,6.5772314,5.805949,4.6802053,3.876103,3.6857438,4.027077,5.10359,6.1046157,5.9930263,4.2207184,0.7187693,0.14441027,0.009846155,0.009846155,0.0,0.0,0.013128206,0.032820515,0.052512825,0.06564103,0.07548718,0.016410258,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02297436,0.108307704,0.3052308,0.15753847,0.15753847,0.17066668,0.16738462,0.2297436,0.16738462,0.098461546,0.04266667,0.016410258,0.016410258,0.026256412,0.03938462,0.08861539,0.14769232,0.12143591,0.15753847,0.25928208,0.3249231,0.4397949,0.8533334,0.63343596,0.6268718,0.39384618,0.029538464,0.15097436,0.3117949,0.31507695,0.25928208,0.24943592,0.39712822,0.9714873,1.020718,0.9682052,1.0010257,1.0994873,1.3062565,2.0545642,2.8160002,3.2886157,3.387077,3.6430771,3.2951798,3.4297438,4.1682053,4.670359,4.7655387,5.533539,5.832206,5.6320004,6.012718,6.7577443,6.23918,5.5532312,5.5630774,6.882462,7.637334,9.019077,9.580308,9.324308,9.688616,9.908514,11.283693,12.691693,13.561437,13.853539,13.367796,14.024206,14.204719,13.331694,11.85477,12.160001,11.35918,10.761847,10.824206,11.155693,11.336206,10.604308,9.82318,9.462154,9.596719,9.645949,9.895386,9.764103,9.170052,8.55959,8.461129,8.694155,8.841846,8.687591,8.224821,9.701744,11.434668,12.918155,13.7386675,13.581129,12.652308,11.605334,11.122872,11.562668,12.954257,14.565744,13.869949,13.351386,13.896206,14.8020525,15.251694,16.288822,17.046976,17.14872,16.708925,16.682669,17.007591,17.575386,18.356514,19.393642,19.797335,19.11795,18.753643,19.46913,21.421951,20.348719,19.751387,19.459284,19.114668,18.189129,16.246155,14.838155,13.860104,13.226667,12.849232,13.505642,13.515489,13.53518,13.689437,13.581129,12.553847,13.653335,15.179488,15.704617,14.070155,14.555899,16.200207,17.542566,17.893745,17.319386,13.925745,11.684103,10.299078,9.403078,8.55959,7.9983597,6.3474874,5.5302567,5.9569235,6.5312824,5.602462,4.59159,3.9384618,3.639795,3.249231,3.3476925,3.8038976,3.6496413,3.1245131,3.6627696,4.516103,4.0336413,3.7907696,4.027077,3.6627696,3.7120004,4.1911798,4.9526157,6.091488,7.936001,8.507077,9.980719,10.650257,9.714872,7.24677,7.529026,5.2381544,3.761231,3.6332312,2.546872,2.097231,1.9659488,4.125539,7.181129,6.363898,3.5052311,4.3684106,5.3136415,4.896821,3.8596926,3.2000003,2.917744,4.017231,5.0084105,1.9068719,2.3827693,1.7887181,1.3128207,1.273436,1.1126155,1.8084104,2.5435898,3.1967182,3.6660516,3.8596926,4.95918,5.435077,5.428513,5.356308,5.904411,5.3070774,4.8640003,4.5029745,4.1452312,3.692308,3.3280003,3.3805132,3.6430771,3.8859491,3.8596926,3.5052311,3.3805132,3.515077,3.6857438,3.4166157,3.1507695,2.5961027,1.8904617,1.529436,2.3958976,2.028308,1.654154,1.7526156,2.2350771,2.4418464,2.1956925,2.1989746,2.5107694,2.8488207,2.5796926,2.8225644,2.7470772,2.5829747,2.4549747,2.3794873,1.7099489,1.467077,1.394872,1.4080001,1.6016412,1.7723079,1.8707694,1.9626669,2.176,2.7011285,3.7382567,4.2371287,4.5029745,4.7524104,5.080616,4.972308,5.2381544,5.182359,4.529231,3.4166157,2.9046156,2.8225644,2.9210258,2.9604106,2.7175386,2.4582565,2.294154,2.2350771,2.2383592,2.228513,2.2514873,2.4516926,2.6453335,2.7569232,2.793026,2.8521028,2.9702566,3.062154,3.1540515,3.370667,3.9942567,4.2141542,4.2568207,4.197744,3.9680004,4.0402055,4.1583595,4.2207184,4.269949,4.4996924,4.7327185,4.7261543,4.667077,4.6211286,4.5456414,4.4734364,4.3552823,4.1156926,3.7743592,3.4330258,3.4691284,3.3608208,3.2065644,2.9735386,2.4713848,1.9331284,1.5261539,1.2274873,1.024,0.9156924,0.7811283,1.1224617,1.3259488,1.2012309,1.0075898,1.0568206,0.95835906,0.82379496,0.7515898,0.82379496,1.3620514,1.6410258,1.591795,1.4211283,1.6180514,1.5195899,1.5425643,1.5097437,1.5360001,1.9987694,1.8149745,1.5589745,1.4998976,1.6738462,1.8904617,1.9889232,2.6453335,3.0785644,3.0884104,3.0523078,2.5009232,2.1989746,2.1333334,2.284308,2.6387694,3.9581542,5.1954875,5.5007186,4.9460516,4.532513,5.2020516,5.0609236,4.4865646,4.125539,4.8836927,4.6867695,4.5095387,4.273231,4.023795,3.95159,5.6976414,6.7117953,7.0826674,6.961231,6.5444107,4.7622566,3.9253337,3.8334363,4.0467696,3.876103,3.2295387,3.515077,4.069744,4.571898,5.034667,4.4734364,4.1222568,4.07959,4.2436924,4.31918,4.4406157,4.8640003,5.0477953,5.182359,6.196513,6.121026,5.435077,5.228308,5.609026,5.7074876,6.416411,7.3780518,7.3682055,6.550975,6.514872,6.1505647,5.7632823,5.330052,5.0149746,5.172513,4.8049235,4.5029745,4.785231,5.7632823,7.1548724,6.8988724,7.240206,7.7456417,7.939283,7.2927184,7.3058467,7.197539,7.210667,7.3616414,7.4469748,6.554257,6.9743595,7.2664623,7.0957956,7.2172313,3.5314875,2.7109745,2.1924105,1.4572309,2.028308,2.9833848,2.6978464,2.2580514,2.7142565,5.080616,3.2000003,2.428718,1.5327181,0.47589746,0.4266667,0.39056414,0.81066674,0.702359,0.60061544,2.5796926,4.4110775,4.4832826,3.5807183,3.5577438,7.3550773,4.6211286,3.0293336,2.1202054,1.972513,3.2032824,7.1220517,11.98277,11.661129,7.020308,5.920821,3.3575387,2.2022567,1.7394873,1.463795,1.0994873,1.1716924,1.4998976,1.6672822,1.6082052,1.6311796,1.522872,1.4506668,1.2898463,1.0568206,0.88615394,0.94523084,0.8598975,0.78769237,0.764718,0.7187693,0.6301539,0.5546667,0.6892308,0.92553854,0.8402052,0.7778462,0.67282057,0.58092314,0.5874872,0.80738467,0.8205129,0.67610264,0.53825647,0.47261542,0.47261542,0.4004103,0.41682056,0.45620516,0.46276927,0.4266667,0.4266667,0.46276927,0.6104616,0.8336411,0.9911796,1.2373334,1.5622566,1.8313848,2.1267693,2.7602053,3.190154,3.5446157,3.8531284,4.128821,4.348718,4.44718,4.1780515,3.7185643,3.2525132,2.9604106,3.3641028,3.4625645,3.43959,3.4724104,3.754667,3.508513,3.1474874,3.0851285,3.4002054,3.8137438,4.414359,4.8640003,4.850872,4.772103,5.737026,6.2129235,5.4449234,5.4613338,6.7249236,8.116513,7.020308,6.2030773,6.186667,6.6034875,6.226052,5.2480006,6.5050263,8.14277,8.444718,5.8453336,6.0258465,7.7390776,7.9228725,6.0783596,4.273231,4.3716927,3.7710772,2.9243078,2.0939488,1.3718976,1.3850257,1.4703591,1.3686155,1.204513,1.5097437,2.8521028,3.5741541,3.6660516,3.2098465,2.3794873,2.294154,2.3827693,2.359795,2.2186668,2.2416413,2.3171284,2.4910772,2.477949,2.2416413,1.9823592,2.1169233,2.0611284,1.9364104,1.8116925,1.6771283,1.5556924,1.9823592,2.1431797,1.8674873,1.6475899,1.7099489,1.6771283,1.4473847,1.2307693,1.5721027,5.914257,5.4908724,5.0182567,4.7327185,4.6276927,4.4734364,4.4865646,4.466872,4.4964104,4.6834874,5.1626673,5.225026,5.5072823,5.720616,5.9536414,6.685539,7.2861543,7.752206,7.9491286,8.001641,8.303591,7.578257,7.456821,7.765334,8.224821,8.464411,7.259898,6.7085133,6.8332314,7.0826674,6.3540516,6.2916927,6.009436,5.8157954,5.98318,6.7610264,6.9710774,7.0990777,7.3452315,7.6603084,7.7325134,7.1483083,7.4404106,8.070564,8.621949,8.825437,8.92718,9.380103,9.888822,10.368001,10.939077,11.431385,11.467488,11.588924,11.766154,11.388719,11.956513,12.327386,12.465232,12.235488,11.382154,11.224616,11.083488,9.888822,8.096821,7.712821,6.3967185,5.1987696,4.650667,5.1167183,6.7872825,7.9097443,7.4207187,4.9394875,1.6475899,0.30194873,0.08861539,0.029538464,0.029538464,0.032820515,0.013128206,0.02297436,0.029538464,0.03938462,0.055794876,0.07548718,0.016410258,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.049230773,0.098461546,0.059076928,0.049230773,0.055794876,0.068923086,0.08205129,0.108307704,0.068923086,0.032820515,0.029538464,0.03938462,0.052512825,0.12143591,0.15097436,0.14441027,0.20676924,0.13784617,0.40697438,1.1060513,1.9068719,2.0873847,2.228513,1.6738462,1.0404103,0.8008206,1.2635899,0.8467693,0.39056414,0.39712822,0.7384616,0.64000005,0.7056411,0.6695385,0.63343596,0.6432821,0.6826667,0.97805136,1.5721027,2.1497438,2.6223593,3.117949,3.3280003,3.889231,4.194462,4.345436,5.169231,5.07077,5.172513,5.684513,6.3212314,6.3277955,6.242462,5.832206,6.2687182,7.456821,8.041026,8.132924,9.025641,9.163487,8.792616,9.970873,10.676514,11.30995,11.644719,11.861334,12.5374365,11.930258,12.681848,13.676309,14.181745,13.856822,12.104206,12.1468725,11.437949,10.020103,10.545232,11.126155,11.030975,10.249847,9.196308,8.707283,8.667898,9.278359,9.764103,9.754257,9.281642,9.025641,9.219283,9.117539,8.628513,8.323282,9.7214365,11.047385,12.114052,12.921437,13.640206,13.689437,13.275898,12.245335,11.300103,11.979488,12.475078,13.180719,13.384206,13.154463,13.3251295,14.25395,15.566771,16.183796,16.091898,16.305231,16.144411,16.640001,17.542566,18.31713,18.12349,18.399181,18.356514,18.185848,18.116924,18.422155,18.645334,18.533745,17.985641,17.293129,17.125746,16.66954,15.66195,14.496821,13.361232,12.199386,12.849232,13.74195,14.093129,13.866668,13.774771,12.87877,13.971693,15.169642,15.382976,14.326155,14.78236,16.866463,18.54359,18.65518,16.89272,14.933334,12.809847,10.866873,9.357129,8.438154,7.9458466,6.6395903,5.6287184,5.4941545,6.3245134,6.265436,5.5171285,4.6933336,4.0402055,3.446154,3.2295387,3.5774362,3.6069746,3.3641028,3.8334363,4.0533338,3.6594875,3.5774362,3.876103,3.7710772,3.761231,4.2502565,5.074052,6.23918,7.88677,8.303591,9.472001,9.626257,8.067283,5.159385,5.284103,4.6244106,6.0291286,7.6734366,3.0720003,1.9856411,1.975795,3.7349746,6.124308,6.1538467,3.4756925,2.8553848,4.240411,5.3694363,1.7723079,1.6508719,3.5807183,6.99077,8.470975,1.785436,1.5097437,1.3193847,1.1946667,1.3653334,2.3105643,2.546872,3.1803079,3.626667,3.5478978,2.8356924,4.8804107,5.2709746,5.074052,5.0149746,5.464616,5.159385,4.841026,4.565334,4.4045134,4.460308,3.889231,3.511795,3.2984617,3.2853336,3.5905645,3.3641028,3.2918978,3.626667,4.056616,3.7120004,3.4822567,3.2164104,2.6354873,2.0775387,2.5042052,2.4024618,1.9528207,1.7493335,1.913436,2.1103592,2.4155898,2.5895386,2.8816411,3.1540515,2.8947694,2.6617439,2.8160002,3.3542566,3.9318976,3.8695388,3.0523078,2.0709746,1.4276924,1.3062565,1.5885129,1.9364104,1.9987694,2.1333334,2.487795,2.993231,3.6004105,4.197744,4.6276927,4.8377438,4.8738465,4.7524104,4.9887185,5.024821,4.6211286,3.8334363,3.31159,2.989949,2.806154,2.6486156,2.3729234,2.4976413,2.546872,2.5961027,2.6715899,2.7273848,2.7733335,2.989949,3.1671798,3.239385,3.3050258,3.3969233,3.4527183,3.564308,3.7940516,4.1911798,4.9099493,5.152821,5.080616,4.850872,4.637539,4.585026,4.5554876,4.4832826,4.397949,4.414359,4.414359,4.4734364,4.598154,4.775385,4.97559,5.0871797,5.0149746,4.7261543,4.269949,3.761231,3.4198978,3.0818465,2.8717952,2.7241027,2.3991797,1.7263591,1.339077,1.1388719,0.99774367,0.7811283,0.7056411,0.86317956,1.0765129,1.1552821,0.92225647,0.98133343,1.017436,0.9419488,0.8205129,0.88615394,1.148718,1.3620514,1.4309745,1.3817437,1.3718976,1.5885129,1.5195899,1.4408206,1.5885129,2.169436,1.8609232,1.5195899,1.5655385,1.9528207,2.172718,1.8707694,2.0676925,2.4943593,2.878359,2.930872,2.3893335,2.0545642,1.9823592,2.225231,2.8225644,3.623385,4.6572313,5.395693,5.543385,5.031385,5.467898,5.362872,5.080616,4.893539,4.955898,4.565334,4.345436,3.826872,3.2328207,3.511795,5.0051284,5.6385646,7.6176414,10.066052,9.035488,5.5729237,3.751385,3.6562054,4.7556925,5.901129,4.2601027,3.564308,3.8071797,4.6769233,5.5597954,4.647385,4.0467696,3.8662567,3.9581542,3.9154875,4.007385,4.279795,4.6145644,5.0215387,5.6320004,5.7468724,5.428513,5.21518,5.3103595,5.586052,6.2523084,6.5280004,6.5739493,6.521436,6.4656415,5.622154,5.110154,4.7655387,4.5587697,4.6112823,4.8114877,4.585026,4.8114877,5.612308,6.3376417,5.8781543,6.2588725,6.7872825,7.030154,6.8430777,6.747898,7.1483083,7.637334,7.821129,7.312411,6.744616,7.328821,7.906462,7.958975,7.634052,6.8266673,6.550975,5.671385,3.9089234,1.847795,3.4330258,4.414359,4.4438977,3.9975388,4.3716927,4.31918,3.8367183,2.7963078,1.8740515,2.5271797,2.5206156,1.8937438,0.9878975,0.79097444,2.9440002,4.414359,4.20759,3.1540515,3.18359,7.3419495,3.3476925,1.9495386,1.6049232,2.1431797,4.7556925,9.084719,9.18318,7.062975,4.6145644,3.6135387,2.2514873,2.284308,2.297436,1.8116925,1.270154,1.3620514,1.4342566,1.5163078,1.5983591,1.6311796,1.3193847,1.2373334,1.1191796,0.8960001,0.7253334,0.9353847,0.88615394,0.7975385,0.7844103,0.85005134,0.6892308,0.636718,0.8960001,1.276718,1.1815386,1.014154,0.8795898,0.7778462,0.72861546,0.77128214,0.892718,0.8467693,0.67938465,0.49230772,0.47261542,0.3708718,0.3314872,0.35774362,0.446359,0.5874872,0.5677949,0.5546667,0.65312827,0.86646163,1.1126155,1.5327181,1.9331284,2.169436,2.2711797,2.4582565,2.8750772,3.2328207,3.6168208,3.9680004,4.07959,4.07959,4.210872,4.013949,3.436308,2.8488207,3.0194874,2.9735386,3.1376412,3.4002054,3.0949745,3.0949745,2.989949,2.7175386,2.4976413,2.8258464,3.6693337,4.4438977,4.5390773,4.1452312,4.2601027,5.7435904,5.730462,5.333334,5.3234878,6.1407185,5.8518977,5.7731285,6.0356927,6.3376417,5.970052,5.228308,5.3858466,5.943795,6.2916927,5.720616,5.543385,6.0816417,6.4065647,6.1407185,5.4580517,4.781949,3.7874875,2.7241027,1.8018463,1.1782565,1.3751796,1.7362052,1.8412309,1.7066668,1.7657437,2.8160002,3.2065644,3.2951798,3.2754874,3.186872,2.9735386,2.993231,2.9440002,2.7766156,2.6945643,2.5337439,2.553436,2.484513,2.2055387,1.7624617,2.1924105,2.3105643,2.1956925,2.0775387,2.3138463,1.9856411,1.9823592,2.0217438,2.0250258,2.100513,1.654154,1.5327181,1.3423591,1.1979488,1.7066668,5.5893335,5.1364107,4.962462,4.886975,4.8377438,4.8640003,4.8147697,4.6605134,4.585026,4.673641,4.893539,4.9296412,5.228308,5.661539,6.1374364,6.5837955,7.069539,7.680001,8.070564,8.139488,8.004924,7.50277,6.994052,7.066257,7.5454364,7.50277,7.427283,7.381334,7.387898,7.328821,6.941539,6.803693,6.1078978,5.805949,6.1768208,6.806975,7.2172313,7.0826674,7.2237954,7.6734366,7.6603084,7.719385,8.297027,8.736821,8.904206,9.18318,9.40636,9.842873,10.262975,10.706052,11.480617,11.828514,11.71036,11.782565,12.11077,12.166565,12.609642,12.4685135,12.511181,12.691693,12.153437,11.910565,11.378873,10.19077,8.874667,8.884514,6.770872,6.189949,6.2851286,7.2960005,10.541949,10.725744,7.7718983,3.7316926,0.56123084,0.108307704,0.04266667,0.029538464,0.032820515,0.029538464,0.006564103,0.009846155,0.013128206,0.01969231,0.029538464,0.029538464,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.02297436,0.026256412,0.016410258,0.013128206,0.016410258,0.02297436,0.036102567,0.06235898,0.055794876,0.06235898,0.09189744,0.118153855,0.18379489,0.18707694,0.128,0.101743594,0.32164106,0.27241027,0.63343596,1.0896411,1.4342566,1.5622566,1.6771283,1.9167181,1.785436,1.394872,1.4769232,1.017436,0.6826667,0.73517954,0.9517949,0.6104616,0.49887183,0.446359,0.38400003,0.42338464,0.86317956,0.7778462,1.2209232,1.6607181,2.0118976,2.6322052,2.7733335,3.2229745,3.7251284,4.056616,4.023795,4.709744,5.1298466,5.4613338,5.7468724,5.8880005,5.61559,5.737026,6.616616,7.9327188,8.687591,8.169026,9.088,9.609847,9.409642,9.682052,10.184206,10.338462,10.561642,10.778257,10.41395,11.434668,12.379898,13.200411,13.679591,13.453129,12.324103,12.202667,11.378873,10.059488,10.364718,10.459898,9.737847,8.914052,8.362667,8.116513,7.830975,8.39877,8.809027,8.887795,9.304616,9.298052,8.92718,8.52677,8.329846,8.464411,9.229129,9.80677,10.295795,10.7848215,11.323078,11.621744,11.890873,11.506873,10.955488,11.815386,11.487181,12.340514,13.069129,13.305437,13.61395,14.076719,14.966155,15.553642,15.734155,16.003283,15.8654375,16.265848,16.889437,17.335796,17.083078,17.224207,17.657436,18.090668,18.271181,17.972515,18.353231,18.002052,17.371899,16.86318,16.807386,17.19795,15.78995,14.490257,13.824001,12.944411,13.2562065,13.653335,13.745232,13.791181,14.693745,14.500104,14.91036,15.655386,16.229744,15.908104,15.760411,16.745028,18.23836,18.881643,16.594053,15.366566,13.548308,11.437949,9.527796,8.507077,8.1066675,7.076103,5.8157954,4.969026,5.4186673,6.436103,6.088206,5.106872,4.089436,3.495385,3.6102567,3.754667,3.6496413,3.3969233,3.4921029,3.4921029,3.2525132,3.3247182,3.7218463,3.9286156,4.0434875,4.522667,5.1200004,5.9634876,7.5618467,8.064001,8.635077,8.388924,6.99077,4.6572313,4.713026,4.381539,5.402257,6.813539,4.9329233,5.6287184,3.5249233,2.7241027,4.525949,7.4141545,4.33559,2.3926156,3.1015387,4.460308,0.95835906,0.9353847,2.7503593,5.2020516,6.048821,2.0217438,1.6082052,1.3357949,1.4178462,1.7755898,2.0217438,2.7536411,2.8488207,3.0293336,3.3312824,3.1081028,4.601436,4.916513,4.8738465,4.906667,5.0642056,4.919795,4.529231,4.1911798,4.1058464,4.3716927,3.8367183,3.5413337,3.1967182,2.8882053,3.1048207,3.0916924,2.9735386,3.2164104,3.7021542,3.7382567,3.3936412,3.2525132,3.0293336,2.7076926,2.5435898,2.609231,2.3105643,1.9528207,1.7132308,1.6443079,1.910154,2.3204105,2.7503593,3.0654361,3.131077,2.6584618,2.5928206,4.31918,6.695385,6.0192823,5.21518,2.8914874,1.394872,1.3357949,1.595077,2.1989746,2.5665643,3.05559,3.6036925,3.7448208,3.879385,4.073026,4.2272825,4.312616,4.3651285,4.345436,4.6112823,4.6933336,4.460308,4.1550775,3.4855387,3.0162053,2.8291285,2.7536411,2.3696413,2.4943593,2.5271797,2.550154,2.6223593,2.7995899,2.7963078,3.0654361,3.3444104,3.5807183,3.945026,3.9712822,3.8695388,3.9122055,4.204308,4.6966157,5.280821,5.8092313,6.009436,5.868308,5.6320004,5.3825645,4.962462,4.5456414,4.240411,4.092718,3.9942567,4.0500517,4.1485133,4.3716927,4.9985647,5.362872,5.287385,4.8705645,4.240411,3.5446157,3.308308,3.0752823,2.8882053,2.6912823,2.353231,1.6968206,1.3095386,1.0962052,0.9517949,0.77456415,0.69907695,0.7384616,0.892718,1.0502565,0.9747693,1.0404103,0.96492314,0.93866676,0.9911796,1.0010257,0.97805136,1.024,1.0666667,1.083077,1.1093334,1.4933335,1.5195899,1.5360001,1.7526156,2.2777438,1.9068719,1.7690258,1.8116925,1.9495386,2.0611284,1.8412309,1.7755898,2.0676925,2.5731285,2.806154,2.540308,2.2711797,2.1530259,2.228513,2.412308,2.7963078,3.6463592,4.5128207,5.100308,5.2676926,5.431795,5.228308,4.900103,4.630975,4.535795,4.381539,4.2568207,3.7054362,3.006359,3.1737437,4.4865646,4.8049235,6.180103,8.4283085,9.117539,8.165744,7.2303596,5.7074876,4.2141542,4.578462,5.4186673,4.3027697,3.7021542,4.3552823,5.2709746,4.8640003,4.201026,3.6857438,3.3805132,2.9997952,3.239385,3.7349746,4.342154,4.8804107,5.1364107,5.024821,5.0051284,5.041231,5.1954875,5.6352825,6.2063594,6.4689236,6.4754877,6.232616,5.6943593,4.781949,4.532513,4.338872,4.128821,4.352,4.890257,4.650667,4.7228723,5.35959,5.979898,5.435077,5.7731285,6.157129,6.3245134,6.5739493,6.744616,7.653744,8.146052,7.906462,7.453539,7.3747697,7.939283,8.267488,8.172308,8.165744,8.621949,8.490667,7.8539495,6.6133337,4.493129,5.3234878,5.7534366,5.8223596,5.72718,5.8157954,5.3858466,5.0149746,4.138667,3.1245131,3.2886157,2.9735386,2.2153847,2.03159,2.412308,2.3302567,3.18359,2.6486156,1.8970258,2.487795,6.370462,3.6135387,2.0184617,2.540308,4.785231,6.99077,12.373334,8.956718,5.4186673,4.647385,3.751385,2.4910772,2.172718,2.0086155,1.6968206,1.404718,1.404718,1.4375386,1.463795,1.4867693,1.5589745,1.2964103,1.2209232,1.0502565,0.8008206,0.8041026,0.97805136,0.9419488,0.88943595,0.8730257,0.8041026,0.83035904,0.8763078,1.014154,1.1881026,1.2209232,1.0929232,1.083077,0.9714873,0.827077,1.0108719,0.90912825,0.8598975,0.77456415,0.65641034,0.60061544,0.55794877,0.55794877,0.57764107,0.6104616,0.65312827,0.65641034,0.6235898,0.82379496,1.2340513,1.5392822,1.6935385,2.041436,2.3827693,2.5796926,2.5271797,3.0358977,3.2131286,3.2787695,3.3345644,3.3542566,3.5052311,3.7907696,3.8137438,3.495385,3.0687182,2.9538465,2.7963078,2.9144619,3.1113849,2.681436,2.3105643,2.5304618,2.6190772,2.4746668,2.6256413,3.2853336,3.876103,4.0992823,4.0369234,4.128821,5.408821,5.802667,5.5565133,5.1200004,5.1232824,5.2644105,5.2545643,5.287385,5.284103,4.890257,4.8344617,5.041231,5.0051284,4.601436,4.069744,3.8596926,4.4438977,5.106872,5.4941545,5.5958977,4.2469745,3.2065644,2.3171284,1.6049232,1.2931283,1.5097437,1.972513,2.300718,2.4451284,2.7011285,3.062154,3.2000003,3.117949,3.0293336,3.370667,3.0654361,2.9833848,2.9768207,2.9472823,2.8521028,2.612513,2.487795,2.5074873,2.4582565,1.9200002,2.156308,2.3958976,2.4484105,2.409026,2.6289232,2.4320002,2.4188719,2.2416413,1.9429746,1.9659488,2.15959,2.1169233,1.8937438,1.785436,2.297436,5.579488,5.0116925,4.8311796,4.8836927,5.034667,5.1889234,5.0576415,4.821334,4.775385,4.903385,4.8738465,5.031385,5.3234878,5.76,6.229334,6.5017443,6.9054365,7.3419495,7.6242056,7.719385,7.7292314,7.719385,7.2927184,7.13518,7.1647186,6.5444107,7.066257,7.450257,7.6242056,7.640616,7.650462,7.174565,6.51159,6.3310776,6.6100516,6.633026,7.174565,6.8955903,6.918565,7.430565,7.6767187,8.073847,8.539898,8.78277,8.884514,9.281642,9.521232,10.003693,10.499283,11.063796,12.048411,12.63918,12.491488,12.593232,13.069129,13.174155,13.312001,12.882052,12.832822,13.128206,12.724514,12.018872,11.355898,10.397539,9.416205,9.255385,7.27959,7.7259493,8.310155,9.120821,12.576821,12.534155,7.9163084,3.0949745,0.4201026,0.2100513,0.12143591,0.08861539,0.068923086,0.04594872,0.006564103,0.0,0.0,0.0032820515,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.016410258,0.016410258,0.0032820515,0.009846155,0.009846155,0.0032820515,0.01969231,0.055794876,0.07548718,0.09189744,0.12143591,0.18707694,0.21661541,0.16082053,0.072205134,0.04594872,0.2297436,0.2855385,0.6498462,0.90256417,0.9714873,1.142154,1.2996924,1.6082052,1.6738462,1.4211283,1.1093334,0.81394875,0.77456415,0.86974365,0.8763078,0.48246157,0.380718,0.44307697,0.4397949,0.47589746,1.0108719,0.75487185,0.97805136,1.1881026,1.3522053,1.9035898,2.3696413,2.865231,3.3280003,3.5938463,3.4166157,4.417641,4.890257,4.9493337,4.84759,4.95918,5.0149746,5.3858466,6.380308,7.7292314,8.595693,8.027898,8.940309,9.793642,9.915077,9.494975,9.613129,9.5606165,9.931488,10.354873,9.485129,10.509129,11.54954,12.084514,11.972924,11.457642,10.906258,10.712616,10.253129,9.718155,10.108719,9.892103,8.743385,7.8834877,7.755488,8.01477,7.643898,7.955693,8.004924,7.8802056,8.713847,9.012513,8.251078,7.5881033,7.568411,8.113232,8.5891285,9.055181,9.40636,9.580308,9.563898,9.531077,10.243283,10.5780525,10.535385,11.244308,10.679795,11.283693,12.3306675,13.275898,13.764924,13.850258,14.283488,14.966155,15.717745,16.28554,16.009848,16.278976,16.49231,16.548103,16.833643,17.05354,17.670565,18.330257,18.615797,18.051283,18.422155,17.96595,17.460514,17.293129,17.440823,16.882874,15.176207,14.099693,13.83713,12.964104,13.249642,13.472821,13.574565,13.984821,15.645539,16.521847,16.308514,16.315079,16.807386,17.03713,16.377438,16.44636,17.555695,18.507488,16.597334,15.074463,13.718975,12.032001,10.197334,9.094564,8.612103,7.765334,6.5017443,5.2676926,5.0116925,6.1440005,6.226052,5.4383593,4.2469745,3.4330258,3.8498464,3.9581542,3.7251284,3.3214362,3.1245131,2.930872,2.8849232,3.0949745,3.515077,3.9220517,4.3684106,4.9493337,5.287385,5.674667,7.0793853,7.8408213,8.008205,7.5618467,6.488616,4.7556925,4.634257,4.023795,4.394667,5.605744,5.904411,6.770872,4.345436,2.5600002,3.4592824,7.181129,4.709744,2.3040001,2.103795,3.062154,0.93866676,0.7975385,1.9922053,3.314872,3.5938463,1.6902566,1.5031796,1.3292309,1.5064616,1.7952822,1.3883078,2.3138463,2.2514873,2.4024618,2.9965131,3.2918978,4.309334,4.6572313,4.7228723,4.7261543,4.6900516,4.7228723,4.378257,3.9647183,3.767795,4.066462,3.8367183,3.5413337,3.1474874,2.806154,2.8422565,2.6912823,2.605949,2.806154,3.2131286,3.4756925,3.3772311,3.3214362,3.2853336,3.1343591,2.6289232,2.6880002,2.6354873,2.349949,1.913436,1.5885129,1.5458462,1.8543591,2.2908719,2.7208207,3.1113849,2.8127182,2.553436,4.7261543,8.192,8.277334,7.4765134,5.0018463,2.6289232,1.4408206,1.8412309,2.917744,3.308308,3.636513,4.0303593,4.128821,4.161641,4.1222568,3.9844105,3.7842054,3.626667,3.6693337,3.9745643,4.1911798,4.2338467,4.2896414,3.5938463,3.0720003,2.8225644,2.7076926,2.3269746,2.409026,2.4681027,2.484513,2.477949,2.5173335,2.5009232,2.7733335,3.170462,3.6036925,4.06318,4.1583595,4.1747694,4.3027697,4.571898,4.850872,5.2020516,5.933949,6.485334,6.6395903,6.5083084,6.1407185,5.5532312,4.9132314,4.397949,4.201026,4.0402055,4.066462,4.1583595,4.4373336,5.2742567,5.861744,5.789539,5.228308,4.4045134,3.6168208,3.3378465,3.1507695,2.993231,2.7700515,2.3466668,1.6508719,1.2438976,1.0108719,0.88287187,0.8172308,0.7811283,0.81066674,0.88943595,0.9682052,0.9616411,1.079795,1.0075898,0.9911796,1.0469744,0.9714873,0.96492314,0.92225647,0.8795898,0.88287187,0.9878975,1.3653334,1.4506668,1.5589745,1.8707694,2.4484105,2.2580514,2.2383592,2.1891284,2.103795,2.176,2.1267693,1.9954873,2.028308,2.2646155,2.5337439,2.550154,2.3991797,2.359795,2.4418464,2.412308,2.5928206,3.1606157,3.6857438,4.056616,4.4865646,4.5095387,4.381539,4.138667,3.95159,4.1124105,4.086154,3.876103,3.3608208,2.8356924,3.0030773,3.9778464,4.2338467,4.5489235,5.3234878,6.5870776,9.452309,9.271795,8.15918,6.5050263,2.9801028,4.9821544,4.6802053,4.0008206,4.017231,4.9460516,5.152821,4.6834874,4.020513,3.3969233,2.7602053,3.0162053,3.4789746,4.069744,4.594872,4.7392826,4.670359,4.6966157,4.7983594,5.0215387,5.47118,5.87159,6.170257,6.124308,5.7009234,5.07077,4.6178465,4.417641,4.07959,3.7448208,4.059898,4.585026,4.3618464,4.3290257,4.821334,5.5630774,5.579488,5.9930263,6.3277955,6.452513,6.5870776,6.8496413,7.906462,8.14277,7.5520005,7.7325134,7.9983597,8.001641,7.968821,8.1066675,8.592411,9.196308,8.904206,8.346257,7.6734366,6.5739493,7.5454364,7.318975,7.0531287,7.13518,7.197539,6.0619493,5.664821,5.097026,4.420923,4.6572313,3.9220517,2.8127182,2.5173335,3.4198978,5.1200004,2.9735386,2.044718,2.3204105,3.6791797,5.8880005,3.314872,2.1234872,3.2000003,5.940513,8.231385,11.559385,7.9294367,4.896821,4.637539,3.945026,2.7536411,2.0250258,1.657436,1.5425643,1.5688206,1.522872,1.5622566,1.522872,1.401436,1.3751796,1.2242053,1.2209232,1.086359,0.86317956,0.90256417,1.0043077,0.97805136,0.95835906,0.95835906,0.8566154,1.014154,1.0502565,1.0305642,1.0502565,1.2438976,1.1388719,1.2077949,1.1290257,0.96492314,1.1684103,0.94523084,0.86646163,0.9189744,0.9714873,0.7975385,0.7384616,0.764718,0.8041026,0.80738467,0.7384616,0.761436,0.8008206,1.017436,1.4145643,1.8182565,1.8970258,2.1300514,2.481231,2.809436,2.8488207,3.3017437,3.442872,3.31159,3.058872,2.9440002,3.1343591,3.31159,3.442872,3.4789746,3.3378465,2.8553848,2.553436,2.553436,2.681436,2.4582565,1.847795,2.041436,2.3926156,2.5961027,2.6847181,3.0752823,3.387077,3.6102567,3.8137438,4.1583595,4.8738465,5.333334,5.32677,4.844308,4.0992823,4.5423594,4.7458467,4.713026,4.4832826,4.138667,4.4996924,5.0182567,4.854154,3.9778464,3.1737437,3.2131286,3.8334363,4.348718,4.604718,4.9821544,3.6890259,2.7831798,2.0873847,1.5786668,1.3915899,1.6443079,2.162872,2.6256413,2.917744,3.1409233,3.0293336,3.2229745,3.1015387,2.8455386,3.4494362,3.1606157,2.868513,2.8455386,3.0227695,3.006359,3.0096412,2.7963078,2.6683078,2.5698464,2.0775387,1.9889232,2.2514873,2.5337439,2.737231,3.006359,2.8980515,2.7733335,2.3958976,1.9003079,1.7755898,2.2678976,2.3433847,2.2088206,2.1497438,2.537026,5.874872,5.218462,4.6834874,4.6112823,4.919795,5.113436,4.9887185,4.84759,4.919795,5.139693,5.1331286,5.3727183,5.681231,5.9634876,6.2523084,6.701949,6.928411,6.892308,6.8266673,6.9645133,7.565129,7.817847,7.8473854,7.64718,7.1680007,6.340924,6.6527185,7.171283,7.7259493,8.050873,7.7718983,6.921847,6.5969234,6.6461544,6.7249236,6.2818465,6.8332314,6.5870776,6.557539,7.0826674,7.8112826,7.860513,7.965539,8.274052,8.736821,9.120821,9.229129,9.800206,10.453334,11.16554,12.288001,13.259488,13.315283,13.574565,14.057027,13.673027,13.620514,13.35795,13.312001,13.321847,12.635899,11.851488,11.460924,10.624001,9.472001,9.147078,8.044309,9.478565,10.131693,9.990565,12.340514,12.176412,7.430565,2.8553848,0.6432821,0.4397949,0.26256412,0.19692309,0.14769232,0.07548718,0.01969231,0.009846155,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.013128206,0.0032820515,0.006564103,0.009846155,0.0032820515,0.0,0.059076928,0.098461546,0.098461546,0.101743594,0.20676924,0.14769232,0.07548718,0.02297436,0.0,0.0,0.16738462,0.4266667,0.7318975,1.0535386,1.3686155,1.7132308,1.1946667,0.8467693,0.84348726,0.5021539,0.40369233,0.5677949,0.72861546,0.7056411,0.4201026,0.4660513,0.71548724,0.83035904,0.79425645,0.9288206,0.86974365,0.86974365,0.80738467,0.8008206,1.2176411,2.097231,2.8553848,3.1081028,3.0752823,3.570872,4.0434875,4.141949,4.141949,4.1091285,3.9089234,4.325744,4.7228723,5.7534366,7.1614366,7.8014364,7.8014364,8.644924,9.488411,9.846154,9.613129,9.7214365,9.570462,9.938052,10.607591,10.361437,9.642668,10.299078,10.541949,9.921641,9.344001,8.694155,8.690872,8.749949,8.87795,9.659078,9.586872,8.704,7.9294367,7.702975,7.9917955,7.827693,7.817847,7.5946674,7.3452315,7.827693,8.231385,7.571693,6.8529234,6.698667,7.3386674,8.021334,9.068309,9.764103,9.82318,9.412924,8.845129,9.567181,10.125129,10.128411,10.233437,10.217027,10.594462,11.602052,12.829539,13.243078,13.472821,13.794462,14.624822,15.842463,16.764719,16.518566,16.833643,16.843489,16.62031,17.184822,17.56882,18.162872,18.658463,18.720821,17.975796,18.507488,18.179283,17.732924,17.641027,18.130053,15.868719,14.263796,13.63036,13.367796,11.9860525,12.416001,13.069129,13.673027,14.444309,16.09518,17.890463,17.572104,16.853334,16.626873,16.964924,16.39713,16.502155,17.214361,17.77559,16.73518,14.444309,13.446565,12.475078,11.113027,9.800206,9.212719,8.500513,7.4404106,6.2227697,5.4416413,5.674667,5.8978467,5.4974365,4.4734364,3.4527183,3.7316926,4.0008206,3.82359,3.2918978,3.0358977,2.5993848,2.7109745,3.045744,3.4100516,3.751385,4.565334,5.2447186,5.4482055,5.5269747,6.547693,7.5191803,7.702975,7.3485136,6.521436,5.0674877,4.594872,3.5478978,4.2141542,6.1768208,6.311385,5.549949,4.7983594,3.9844105,3.8006158,5.717334,4.4996924,2.300718,1.4769232,2.0184617,1.529436,1.723077,2.5140514,3.186872,2.9768207,1.0601027,1.0699488,1.2209232,1.4736412,1.6016412,1.1946667,1.6804104,1.9495386,2.2777438,2.7175386,3.0949745,4.059898,4.529231,4.5817437,4.4045134,4.279795,4.529231,4.2896414,3.8728209,3.6004105,3.8071797,3.9318976,3.515077,3.1343591,3.0096412,2.993231,2.3630772,2.284308,2.537026,2.878359,3.0654361,3.4494362,3.5314875,3.5314875,3.4034874,2.8455386,2.7602053,2.8947694,2.8356924,2.4943593,2.103795,1.723077,1.6607181,1.8871796,2.3236926,2.8389745,2.9078977,2.809436,4.841026,8.546462,10.729027,9.639385,8.385642,5.3234878,1.7952822,2.1497438,3.5216413,3.6496413,3.446154,3.4560003,3.8662567,4.096,4.1452312,3.9056413,3.4231799,2.8849232,2.9046156,3.1277952,3.442872,3.7448208,3.9581542,3.6102567,3.259077,2.92759,2.6223593,2.3072822,2.3236926,2.428718,2.4713848,2.4024618,2.2514873,2.3401027,2.550154,2.9636924,3.442872,3.6430771,3.895795,4.2305646,4.565334,4.788513,4.7622566,4.8738465,5.4941545,6.229334,6.7610264,6.8430777,6.4623594,5.9930263,5.3727183,4.785231,4.6244106,4.5062566,4.644103,4.886975,5.2348723,5.83877,6.308103,6.121026,5.4843082,4.6572313,3.9778464,3.446154,3.1048207,2.92759,2.740513,2.2449234,1.4933335,1.1060513,0.9124103,0.83035904,0.86317956,0.88615394,0.9747693,1.024,0.98133343,0.8467693,1.024,1.1093334,1.0962052,0.9944616,0.8467693,1.0535386,1.0338463,0.9353847,0.8960001,1.0436924,1.3259488,1.3686155,1.4966155,1.8838975,2.546872,2.7569232,2.7569232,2.6387694,2.5140514,2.5304618,2.5632823,2.5271797,2.3401027,2.1431797,2.3105643,2.4155898,2.294154,2.3794873,2.674872,2.7864618,2.8717952,3.0851285,3.0949745,2.9571285,3.1113849,3.1048207,3.2131286,3.242667,3.318154,3.889231,3.7021542,3.2754874,2.92759,2.8750772,3.239385,3.5905645,3.95159,3.895795,3.4231799,2.9604106,7.90318,8.149334,8.79918,9.4457445,4.1517954,3.495385,4.1189747,4.20759,3.7809234,4.699898,5.1232824,4.9788723,4.6211286,4.1878977,3.5971284,3.6857438,3.9122055,4.1878977,4.4340515,4.6080003,4.84759,4.7491283,4.71959,4.8705645,5.024821,5.2053337,5.3727183,5.297231,5.0149746,4.841026,4.972308,4.562052,3.9187696,3.4658465,3.7448208,4.0369234,3.889231,3.8596926,4.210872,4.896821,5.687795,6.3179493,6.8594875,7.1680007,6.8955903,6.8594875,7.6996927,7.748924,7.194257,8.077128,8.27077,7.512616,7.256616,7.817847,8.375795,8.73354,8.2904625,7.7325134,7.4043083,7.3058467,8.700719,8.493949,8.027898,7.8670774,7.8047185,6.5280004,5.970052,5.61559,5.546667,6.4754877,5.5269747,3.817026,2.3269746,3.006359,8.736821,3.9384618,3.0129232,4.135385,5.6418467,6.009436,2.425436,2.4188719,3.4756925,4.923077,7.9327188,7.0367184,5.5007186,4.33559,3.82359,3.501949,2.681436,1.9823592,1.5786668,1.5097437,1.6804104,1.6672822,1.6804104,1.591795,1.3883078,1.1684103,1.1191796,1.1881026,1.1815386,1.0732309,1.024,1.0568206,1.0404103,1.0305642,1.0502565,1.0633847,1.148718,1.0535386,0.9682052,1.0338463,1.332513,1.2077949,1.2668719,1.2373334,1.1158975,1.1585642,1.024,0.9878975,1.1388719,1.3029745,1.017436,0.90256417,0.9189744,0.98133343,1.0010257,0.90912825,0.9321026,1.0404103,1.1552821,1.3423591,1.8313848,2.1530259,2.3105643,2.5206156,2.8291285,3.1015387,3.370667,3.7087183,3.7152824,3.3641028,2.9997952,2.9669745,2.9078977,3.0293336,3.2722054,3.3247182,2.6354873,2.2416413,2.156308,2.2711797,2.353231,1.8609232,1.7165129,2.0151796,2.5435898,2.7667694,2.9440002,3.117949,3.2229745,3.318154,3.6135387,4.128821,4.4996924,4.5390773,4.066462,2.9243078,3.6069746,4.2502565,4.4438977,4.2207184,4.023795,4.1714873,4.7524104,4.709744,3.9647183,3.3969233,3.7743592,4.007385,3.9712822,3.8367183,4.076308,3.4330258,2.7634873,2.225231,1.8609232,1.5983591,1.8642052,2.3827693,2.8192823,2.986667,2.8389745,2.6978464,3.1671798,3.2065644,2.9078977,3.511795,3.4231799,2.878359,2.7306669,3.0358977,3.05559,3.383795,3.1343591,2.7634873,2.484513,2.2449234,1.9396925,2.048,2.4024618,2.8717952,3.383795,3.249231,2.8521028,2.3958976,2.028308,1.8346668,1.9626669,2.1169233,2.1792822,2.2153847,2.484513,5.8125134,5.5565133,5.07077,4.6080003,4.3585644,4.457026,4.4077954,4.322462,4.3749747,4.630975,5.034667,5.2545643,5.602462,5.943795,6.409847,7.384616,6.9087186,6.6625648,6.564103,6.550975,6.5772314,7.003898,7.322257,7.460103,7.50277,7.6603084,7.9524107,8.12636,8.146052,7.6996927,6.2096415,6.052103,6.11118,6.491898,6.892308,6.62318,6.987488,6.6592827,6.567385,6.9809237,7.506052,7.020308,7.328821,7.9852314,8.585847,8.743385,8.694155,9.068309,9.90195,11.057232,12.1928215,12.898462,13.157744,13.581129,13.988104,13.426873,14.198155,14.244103,14.083283,13.6467705,12.268309,12.25518,11.949949,10.679795,9.268514,10.023385,8.963283,10.71918,11.008,9.826463,11.474052,8.349539,4.713026,1.9462565,0.5973334,0.36758977,0.20676924,0.25928208,0.2231795,0.06564103,0.029538464,0.029538464,0.02297436,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.013128206,0.0,0.0,0.04594872,0.07548718,0.098461546,0.18379489,0.18379489,0.072205134,0.0,0.0,0.0,0.20676924,0.20348719,0.3446154,0.7811283,1.463795,1.8313848,1.3193847,0.5481026,0.0,0.0,0.14769232,0.29210258,0.574359,0.82379496,0.58092314,0.95835906,1.2898463,1.3883078,1.2077949,0.8533334,1.0010257,0.9747693,0.827077,0.764718,1.1454359,1.5360001,1.6869745,1.9790771,2.4352822,2.7175386,2.546872,2.7667694,3.2262566,3.5544617,3.190154,3.1638978,4.194462,5.333334,6.12759,6.5903597,7.3714876,8.612103,9.380103,9.55077,9.796924,10.834052,10.371283,10.473026,11.533129,12.251899,11.155693,10.41395,9.685334,9.101129,9.245539,9.321027,8.953437,8.569437,8.55959,9.291488,9.317744,8.920616,8.51036,8.054154,7.066257,7.3091288,7.059693,6.9842057,7.194257,7.2172313,7.328821,7.2172313,6.925129,6.669129,6.8496413,7.6209235,9.058462,10.082462,10.30236,10.010257,9.32759,9.511385,9.816616,9.9282055,9.964309,11.34277,11.523283,11.841642,12.560411,12.87877,13.633642,14.25395,15.1466675,16.07877,16.190361,17.115898,17.834667,18.048002,17.746052,17.19795,17.355488,17.98236,18.707693,19.049026,18.402462,18.963694,18.343386,17.293129,16.554668,16.8599,15.360002,14.01436,13.420309,13.121642,11.595488,11.388719,11.949949,13.164309,14.631386,15.655386,17.401438,17.673847,17.007591,16.134565,15.977027,16.46277,17.375181,17.70995,17.237335,16.479181,14.391796,13.138052,12.379898,11.483898,9.504821,9.26195,8.753231,7.752206,6.6002054,6.2096415,5.5762057,5.106872,4.6539493,4.20759,3.892513,3.4888208,3.8728209,3.95159,3.5380516,3.3411283,2.865231,2.9768207,3.4034874,3.7743592,3.6168208,4.4701543,4.903385,5.1298466,5.4153852,6.0717955,6.8299494,7.4043083,7.525744,7.02359,5.8125134,4.8607183,3.4166157,4.768821,8.214975,9.032206,8.507077,7.8736415,6.987488,6.232616,6.5017443,4.890257,2.4549747,1.4473847,2.1398976,2.8225644,4.9099493,5.156103,3.8695388,2.0841026,1.5721027,1.2406155,1.3522053,1.8281027,2.2547693,1.8773335,1.8773335,2.3433847,2.6912823,2.861949,3.3280003,3.764513,4.3060517,4.44718,4.1189747,3.692308,4.1189747,3.5938463,3.314872,3.511795,3.4625645,3.511795,3.4067695,3.308308,3.3247182,3.495385,2.4943593,2.0151796,2.166154,2.665026,2.8225644,3.1638978,3.4888208,3.8038976,3.882667,3.2361028,3.0162053,3.114667,3.2065644,3.1409233,2.9440002,2.3696413,2.1989746,2.1333334,2.1431797,2.4713848,2.5337439,3.0982566,5.9470773,10.55836,14.099693,12.022155,11.943385,8.539898,2.7831798,1.9528207,2.5271797,2.7241027,2.7011285,2.7306669,3.2196925,3.3903592,3.4592824,3.3214362,2.9702566,2.5173335,2.4681027,2.3105643,2.2678976,2.4188719,2.7011285,3.31159,3.5905645,3.5807183,3.308308,2.806154,2.4549747,2.3105643,2.2678976,2.3368206,2.6551797,3.045744,3.170462,3.3542566,3.5446157,3.3280003,3.4592824,3.7973337,4.1550775,4.457026,4.699898,4.578462,4.647385,5.228308,6.0356927,6.196513,5.865026,5.435077,4.9821544,4.6112823,4.4406157,4.7327185,5.4186673,6.0225644,6.2785645,6.117744,5.58277,4.850872,4.322462,4.0500517,3.767795,3.318154,2.7470772,2.4352822,2.294154,1.7690258,1.2340513,1.017436,0.9321026,0.88943595,0.8992821,0.86317956,0.94523084,1.0994873,1.1388719,0.74830776,0.90584624,1.0108719,1.0601027,1.0436924,0.94523084,0.9944616,1.017436,0.98461545,0.98133343,1.1913847,1.4703591,1.4769232,1.5622566,1.8412309,2.1825643,2.7798977,3.0490258,3.0851285,2.9210258,2.5173335,2.5895386,2.7569232,2.6880002,2.4943593,2.7011285,2.5435898,2.100513,2.0512822,2.3958976,2.4582565,2.2482052,2.1956925,2.2777438,2.4615386,2.7306669,2.609231,2.7634873,2.878359,3.045744,3.754667,3.314872,2.9571285,3.2131286,3.9351797,4.2863593,3.7021542,3.9680004,4.7917953,4.7917953,1.4966155,3.5478978,5.4875903,5.034667,4.568616,11.122872,3.7743592,2.5238976,3.0851285,3.4658465,3.9680004,3.9417439,3.9647183,4.4898467,5.221744,5.110154,5.0642056,5.5991797,5.6254363,5.097026,5.034667,5.156103,5.1331286,5.175795,5.146257,4.5456414,4.522667,4.588308,4.4734364,4.3027697,4.6080003,4.535795,4.1682053,3.6857438,3.4034874,3.767795,4.013949,3.9187696,3.948308,4.141949,4.1058464,4.5456414,5.349744,6.413129,7.3353853,7.4469748,6.8233852,7.4371285,7.8047185,7.762052,8.467693,7.968821,7.2861543,7.003898,7.0465646,6.669129,7.328821,7.282872,7.5979495,8.329846,8.513641,7.0859494,7.433847,7.88677,7.9786673,8.454565,7.4765134,6.636308,6.052103,5.914257,6.5017443,5.9634876,4.457026,2.556718,1.595077,3.6463592,4.1091285,4.5390773,4.2502565,3.9089234,5.5072823,2.9702566,4.3290257,4.8804107,4.3060517,6.698667,5.0642056,3.8662567,3.242667,3.1606157,3.4166157,2.868513,2.172718,1.6672822,1.4736412,1.5097437,1.5360001,1.4769232,1.4539489,1.4145643,1.1454359,1.2307693,1.2340513,1.2438976,1.3062565,1.404718,1.270154,1.2537436,1.2668719,1.2570257,1.2209232,1.1224617,0.90584624,0.86974365,1.0765129,1.3587693,1.273436,1.3686155,1.3226668,1.1355898,1.1585642,1.1224617,1.3062565,1.4112822,1.3456411,1.2373334,1.2471796,1.3062565,1.3193847,1.2635899,1.1913847,1.2012309,1.142154,1.1716924,1.3784616,1.7690258,2.3072822,2.5600002,2.6157951,2.612513,2.7470772,3.0260515,3.6102567,4.007385,3.879385,3.0358977,2.5731285,2.4648206,2.5074873,2.5796926,2.6387694,2.4188719,2.2547693,2.1464617,2.1333334,2.3040001,1.9987694,1.6935385,1.8215386,2.3762052,2.9144619,2.9144619,3.0982566,3.1474874,2.868513,2.1989746,3.501949,3.9844105,3.8071797,3.1671798,2.28759,3.0227695,3.6529233,3.9778464,4.010667,3.9975388,3.3280003,3.570872,3.508513,3.0424619,3.190154,3.6660516,3.4921029,3.3509746,3.4560003,3.5413337,3.1967182,2.8750772,2.7208207,2.6847181,2.5009232,2.4648206,2.806154,3.0129232,2.8750772,2.4713848,2.5928206,3.1376412,3.3805132,3.2328207,3.2196925,3.5971284,2.9505644,2.6026669,2.7634873,2.5173335,2.6026669,2.3138463,2.2514873,2.540308,2.806154,2.550154,2.2022567,2.1300514,2.4943593,3.249231,3.2131286,2.809436,2.4582565,2.297436,2.2121027,2.176,2.3302567,2.4910772,2.6683078,3.0818465,6.7282057,6.629744,6.0225644,5.356308,4.8344617,4.394667,4.345436,4.2830772,4.345436,4.604718,5.034667,5.5007186,5.8190775,6.235898,6.7938466,7.3616414,6.925129,6.5772314,6.36718,6.3901544,6.7840004,6.8299494,6.76759,6.6592827,6.7610264,7.525744,7.702975,7.5520005,7.1614366,6.5805135,5.832206,5.654975,5.973334,6.426257,6.7282057,6.6822567,6.8430777,6.2884107,6.163693,6.7314878,7.3714876,7.637334,8.43159,9.091283,9.567181,10.427077,11.0145645,10.696206,11.0145645,12.1238985,12.790154,12.803283,12.547283,12.698257,13.24636,13.476104,14.25395,14.230975,13.843694,13.302155,12.596514,12.35036,12.045129,11.392001,11.001437,12.393026,11.556104,12.445539,11.995898,10.338462,10.81436,6.7905645,3.3247182,1.1158975,0.26256412,0.24287182,0.14441027,0.13128206,0.108307704,0.06564103,0.07876924,0.059076928,0.14769232,0.26256412,0.27897438,0.02297436,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.036102567,0.03938462,0.0032820515,0.0,0.0,0.029538464,0.101743594,0.16738462,0.13456412,0.0951795,0.032820515,0.0,0.0,0.0,0.36430773,0.39384618,0.30194873,0.256,0.35446155,0.7384616,0.69251287,0.43323082,0.190359,0.21989745,0.25928208,0.318359,0.32820517,0.35446155,0.6301539,0.8795898,1.1946667,1.2931283,1.1126155,0.8172308,1.0535386,0.85005134,0.82379496,0.96492314,0.6301539,1.1290257,1.2931283,1.6311796,2.1267693,2.2514873,2.4910772,2.7798977,3.0949745,3.3345644,3.2984617,3.56759,4.630975,5.5696416,5.986462,6.0291286,6.8496413,7.637334,8.050873,8.493949,10.112,10.331899,9.800206,9.987283,11.152411,12.35036,11.9171295,10.755282,9.961026,9.724719,9.344001,9.672206,9.179898,8.628513,8.536616,9.170052,8.969847,8.832001,8.280616,7.3025646,6.3310776,6.058667,5.943795,6.3245134,7.1089234,7.778462,8.113232,8.257642,8.155898,7.9524107,7.9983597,8.592411,9.163487,9.590155,9.921641,10.400822,9.728001,9.6295395,9.6065645,9.577026,9.865847,11.352616,11.772718,11.992617,12.35036,12.658873,13.082257,14.10954,15.652103,17.004309,16.8599,17.611488,18.658463,19.410053,19.744822,20.017233,18.084105,17.631182,18.225233,18.901335,18.159592,17.539284,16.672821,15.868719,15.40595,15.553642,14.532925,13.525334,12.76718,12.3076935,12.012309,11.559385,11.234463,11.730052,13.062565,14.555899,15.82277,16.876308,16.997746,16.344616,15.95077,15.816206,17.060104,18.084105,18.087385,17.076513,14.959591,13.13477,12.104206,11.513436,10.14154,8.979693,8.349539,7.821129,7.3583593,7.3091288,6.058667,4.7327185,3.876103,3.6758976,3.9647183,3.9122055,4.1878977,4.4242053,4.325744,3.6726158,3.2229745,3.114667,3.4789746,3.9647183,3.7382567,4.210872,4.7622566,5.1987696,5.464616,5.6451287,6.3343596,7.197539,7.683283,7.394462,6.1078978,4.8607183,3.817026,4.7622566,8.621949,15.465027,14.775796,14.683899,12.475078,8.595693,6.6461544,6.73477,3.5216413,2.4615386,3.69559,2.0545642,4.240411,7.2336416,6.0980515,1.7952822,1.1946667,1.3522053,1.5556924,1.8116925,1.9495386,1.6213335,1.9823592,2.3204105,2.6617439,3.006359,3.314872,3.8301542,4.2535386,4.2863593,3.9187696,3.4231799,3.879385,3.442872,3.0654361,3.0720003,3.1573336,3.245949,3.2361028,3.0424619,2.9078977,3.4198978,3.1048207,2.3335385,2.097231,2.5140514,2.8488207,2.740513,3.2295387,3.5807183,3.570872,3.4789746,3.501949,3.5544617,3.6332312,3.6758976,3.5807183,3.1343591,3.0654361,2.8422565,2.425436,2.2777438,2.162872,2.7634873,6.180103,10.71918,10.8996935,14.119386,17.375181,15.747283,9.563898,4.4077954,2.2646155,1.7493335,1.847795,2.0086155,2.1464617,2.0611284,2.4057438,2.6617439,2.5895386,2.2383592,2.1891284,2.0742567,2.1431797,2.5271797,3.239385,3.8104618,3.8662567,3.7776413,3.6791797,3.4921029,3.1376412,2.8553848,2.5764105,2.3827693,2.484513,2.6223593,2.6683078,2.7864618,2.9833848,3.1081028,3.0949745,3.2918978,3.5774362,3.9089234,4.309334,4.381539,4.348718,4.634257,5.156103,5.3037953,5.3169236,5.228308,5.077334,4.919795,4.8049235,4.972308,5.1954875,5.4153852,5.549949,5.5072823,5.0510774,4.699898,4.466872,4.3027697,4.1091285,3.4625645,2.7273848,2.176,1.8248206,1.4276924,1.0962052,0.8566154,0.7318975,0.69907695,0.67938465,0.7811283,0.78769237,0.8172308,0.8369231,0.6629744,0.7811283,0.8763078,1.014154,1.1093334,0.9353847,0.9156924,0.9911796,1.0436924,1.0371283,1.020718,1.1618463,1.3620514,1.6475899,2.0217438,2.4516926,2.7569232,2.9669745,3.1277952,3.0654361,2.3696413,2.7273848,3.0523078,2.9407182,2.5107694,2.3958976,2.3729234,1.9790771,1.654154,1.5031796,1.3226668,1.4769232,1.5064616,1.522872,1.6246156,1.913436,2.0644104,2.5796926,2.8422565,2.9078977,3.508513,3.3542566,3.1409233,3.255795,3.7218463,4.201026,4.1911798,4.352,5.146257,5.861744,4.6080003,2.6157951,1.9429746,3.2525132,5.412103,5.47118,3.3280003,2.793026,2.7273848,2.9046156,3.9909747,4.6211286,4.4110775,4.6834874,5.6976414,6.6625648,6.2818465,6.311385,6.186667,5.661539,4.778667,4.775385,5.0838976,5.1889234,5.0051284,4.8640003,4.955898,4.8705645,4.2568207,3.4592824,3.508513,4.0041027,3.945026,3.876103,3.9089234,3.767795,4.20759,4.44718,4.453744,4.2240005,3.7874875,3.6791797,3.9811285,4.785231,5.8223596,6.4689236,6.3442054,7.0104623,7.2303596,6.941539,7.24677,7.3025646,7.177847,7.02359,6.688821,5.717334,4.7360005,3.3345644,3.3280003,5.1987696,8.086975,7.3616414,7.1089234,7.522462,8.585847,10.075898,9.636104,8.65477,7.7456417,7.4010262,7.9786673,7.197539,5.034667,3.5249233,3.2722054,3.43959,5.35959,5.7698464,6.0816417,6.163693,4.325744,4.2568207,4.8738465,4.6539493,4.128821,5.868308,4.9952826,3.2623591,2.6912823,3.4330258,3.7973337,3.0129232,2.353231,1.8182565,1.4933335,1.5589745,1.3981539,1.3817437,1.3784616,1.3062565,1.1454359,1.0732309,0.9878975,0.955077,1.020718,1.1946667,1.2471796,1.1749744,1.017436,0.86646163,0.8795898,0.9189744,0.88943595,1.024,1.2832822,1.3686155,1.4900514,1.6377437,1.6278975,1.5786668,1.9167181,1.6443079,1.404718,1.404718,1.5360001,1.3587693,1.2931283,1.3686155,1.4736412,1.5064616,1.3850257,1.3489232,1.1224617,1.1388719,1.5195899,2.0873847,2.097231,2.5632823,2.865231,2.9111798,3.1245131,3.3969233,3.5807183,3.639795,3.4789746,2.937436,2.4943593,2.356513,2.3696413,2.3893335,2.2744617,2.2482052,1.9561027,1.8510771,1.9823592,1.9856411,1.8182565,1.657436,1.8346668,2.3171284,2.7076926,2.7076926,2.9472823,3.0358977,2.8422565,2.5009232,2.7733335,3.186872,3.3903592,3.2196925,2.6912823,2.7503593,2.7798977,2.861949,2.9243078,2.7634873,2.3466668,2.6486156,2.7831798,2.6715899,3.0424619,3.498667,3.31159,3.0358977,2.9472823,3.0523078,2.6322052,2.6683078,2.8488207,2.9144619,2.674872,2.5304618,2.6157951,2.6322052,2.484513,2.2777438,2.4484105,2.930872,3.4166157,3.5774362,3.0358977,3.2787695,3.249231,3.1934361,3.1540515,2.9702566,3.0162053,2.5173335,2.1431797,2.2121027,2.6847181,2.028308,1.7263591,1.8543591,2.28759,2.7142565,2.8324106,2.7470772,2.8127182,3.0293336,3.0293336,2.3991797,2.3893335,2.5107694,2.5731285,2.7175386,7.131898,6.8233852,6.1538467,5.398975,4.772103,4.4242053,4.273231,4.276513,4.5029745,4.844308,5.034667,5.3103595,5.658257,6.1374364,6.705231,7.1909747,6.8430777,6.5837955,6.685539,6.99077,6.8988724,6.675693,6.7971287,6.9349747,6.9677954,6.997334,7.3714876,7.0793853,6.619898,6.186667,5.654975,5.3037953,5.47118,5.874872,6.2720003,6.452513,6.626462,6.482052,6.485334,6.7544622,7.0367184,7.269744,7.716103,8.224821,8.914052,10.161232,10.768411,11.329642,12.373334,13.5548725,13.673027,13.482668,12.918155,12.944411,13.505642,13.505642,13.636924,13.443283,13.065847,12.678565,12.47836,12.320822,12.297847,11.943385,11.58236,12.327386,12.219078,13.088821,12.934566,12.150155,13.53518,8.861539,4.3585644,1.3292309,0.1148718,0.08533334,0.052512825,0.03938462,0.032820515,0.026256412,0.036102567,0.026256412,0.072205134,0.16410258,0.21333335,0.059076928,0.5152821,0.26912823,0.01969231,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.013128206,0.016410258,0.009846155,0.016410258,0.036102567,0.029538464,0.0032820515,0.009846155,0.0032820515,0.02297436,0.08533334,0.13784617,0.049230773,0.029538464,0.009846155,0.0,0.0,0.0,0.16082053,0.33476925,0.27569234,0.049230773,0.029538464,0.18707694,0.21333335,0.28882053,0.4135385,0.4201026,0.64000005,0.49230772,0.380718,0.5284103,0.9878975,1.3029745,1.3259488,1.2012309,1.0272821,0.86317956,1.7132308,1.7132308,1.5885129,1.4605129,0.85005134,1.1848207,1.2635899,1.3981539,1.6475899,1.8051283,1.9593848,2.5796926,3.0096412,3.1540515,3.4822567,3.9548721,4.414359,5.1987696,6.042257,6.0816417,6.4065647,6.9809237,7.2303596,7.3682055,8.425026,9.032206,8.986258,9.642668,10.880001,11.083488,11.063796,10.492719,10.003693,10.066052,10.988309,10.8537445,10.095591,9.16677,8.464411,8.342975,7.8736415,7.9294367,7.6964107,7.0432825,6.5247183,6.304821,6.4065647,6.5706673,6.747898,7.0859494,7.8441033,8.169026,8.572719,9.091283,9.301334,9.728001,10.381129,10.781539,10.794667,10.65354,10.223591,9.895386,9.90195,10.098872,9.961026,11.099898,12.133744,12.649027,12.770463,13.161027,13.686155,14.28677,15.593027,17.217642,17.742771,18.041437,18.468103,19.14749,19.971283,20.594873,19.370668,18.15631,18.087385,18.743795,18.179283,17.066668,15.986873,15.38954,15.238565,15.018668,13.732103,12.721231,11.529847,10.473026,10.624001,10.673231,10.364718,10.788103,12.107488,13.558155,14.034052,15.382976,15.986873,15.596309,15.314053,14.670771,15.61272,17.083078,18.218668,18.353231,17.02072,14.168616,12.356924,12.015591,11.414975,9.754257,8.697436,7.955693,7.529026,7.719385,6.6527185,5.349744,4.3290257,3.8137438,3.7251284,4.457026,4.7261543,4.8607183,4.827898,4.210872,4.073026,3.5971284,3.6430771,4.073026,3.767795,3.7809234,4.3585644,4.890257,5.142975,5.2545643,5.83877,6.6067696,7.000616,6.7971287,6.1078978,4.8771286,3.570872,4.086154,7.3485136,13.302155,11.713642,11.644719,11.401847,10.115283,7.7357955,5.225026,2.6486156,1.7132308,2.1431797,1.6771283,2.5271797,3.945026,3.6135387,1.7033848,0.90584624,1.6344616,2.097231,2.2908719,2.2219489,1.913436,2.028308,2.2777438,2.6026669,3.058872,3.7874875,4.0303593,4.007385,3.882667,3.7152824,3.4560003,4.2436924,3.9581542,3.43959,3.1409233,3.1474874,3.2131286,3.387077,3.2656412,2.917744,2.861949,3.0326157,2.6026669,2.3860514,2.612513,2.917744,2.5009232,2.9965131,3.3969233,3.3312824,3.0720003,3.8104618,4.128821,4.1517954,3.9876926,3.748103,3.5511796,3.7087183,3.6496413,3.2754874,2.9768207,2.4549747,2.5173335,5.284103,9.258667,9.330873,13.932309,20.575182,22.764309,18.917746,12.370052,6.76759,3.767795,2.4320002,2.0118976,1.9593848,1.657436,1.8116925,2.3302567,2.8389745,2.678154,2.6683078,2.612513,2.733949,3.0785644,3.508513,3.9253337,4.1485133,4.266667,4.2272825,3.8531284,3.4494362,3.0523078,2.7700515,2.6387694,2.6518977,2.6945643,2.7831798,2.9735386,3.2065644,3.2886157,3.3444104,3.4100516,3.6168208,3.9056413,4.0369234,4.1747694,4.332308,4.6211286,5.034667,5.4383593,5.3891287,5.405539,5.609026,5.868308,5.7764106,5.7501545,5.4482055,5.2480006,5.225026,5.146257,4.9394875,4.397949,3.9089234,3.6430771,3.5380516,2.9669745,2.284308,1.7460514,1.4178462,1.1684103,1.0502565,0.8402052,0.6859488,0.65312827,0.7089231,0.69579494,0.8402052,0.8730257,0.7384616,0.5874872,0.7384616,0.86974365,1.0305642,1.148718,1.0043077,0.9517949,0.9419488,0.92553854,0.88943595,0.83035904,0.92553854,1.3226668,1.7624617,2.1070771,2.3630772,2.556718,2.6551797,2.7306669,2.6617439,2.1333334,2.2908719,2.8422565,3.1671798,3.05559,2.7208207,2.156308,1.7296412,1.3817437,1.1093334,0.94523084,1.2209232,1.3292309,1.339077,1.3357949,1.4244103,1.6377437,2.2350771,2.5895386,2.740513,3.4034874,3.3608208,3.4494362,3.639795,3.9253337,4.2994876,4.565334,4.5029745,4.8147697,5.4449234,5.579488,3.8629746,2.4516926,2.5042052,3.5249233,3.3542566,2.540308,3.3608208,4.2240005,4.204308,3.0358977,5.3760004,5.7665644,5.3858466,5.3825645,6.892308,6.7807183,6.6560006,6.452513,5.9995904,5.0084105,4.841026,5.0904617,5.3234878,5.402257,5.5007186,5.353026,5.21518,4.644103,3.761231,3.242667,3.2918978,3.4100516,3.6529233,3.889231,3.7973337,4.453744,5.159385,5.284103,4.818052,4.3749747,3.9056413,3.7710772,4.1517954,4.95918,5.8486156,6.121026,6.6527185,6.921847,6.885744,6.9710774,6.7249236,6.744616,6.8463597,6.521436,4.9362054,4.7261543,6.49518,5.668103,3.3608208,6.370462,7.204103,6.872616,6.7971287,7.571693,8.973129,9.216001,8.802463,8.753231,9.248821,9.609847,7.640616,5.297231,4.128821,4.269949,4.4406157,6.180103,6.242462,6.7577443,7.171283,4.2469745,3.8006158,3.945026,4.1747694,4.1124105,3.4921029,4.1714873,3.1737437,2.665026,3.1245131,3.3312824,2.8258464,2.349949,1.8609232,1.4375386,1.2603078,1.1848207,1.1388719,1.1323078,1.1191796,1.0075898,0.88943595,0.8336411,0.86974365,0.9517949,0.9353847,1.1126155,0.98133343,0.83035904,0.81394875,0.93866676,0.90912825,0.8763078,0.95835906,1.1651284,1.3915899,1.6049232,1.723077,1.7362052,1.7165129,1.8313848,1.5163078,1.4802053,1.5622566,1.6082052,1.4802053,1.467077,1.4112822,1.6180514,1.9495386,1.8379488,1.5983591,1.4408206,1.5261539,1.8642052,2.3138463,2.4385643,2.9210258,3.3411283,3.501949,3.43959,3.692308,3.6004105,3.2164104,2.7569232,2.5928206,2.4188719,2.2055387,2.1267693,2.1530259,2.044718,2.2678976,1.9889232,1.8445129,2.0053334,2.172718,1.8051283,1.6738462,1.8084104,2.1267693,2.4352822,2.3466668,2.5206156,2.8192823,2.9965131,2.6978464,2.2416413,2.3401027,2.678154,2.868513,2.4451284,2.3138463,2.2416413,2.281026,2.2711797,1.8707694,1.6278975,1.9626669,2.0217438,1.8149745,2.2186668,2.802872,2.9144619,2.9472823,2.9833848,2.802872,2.4352822,2.6683078,2.986667,3.0293336,2.5961027,2.4549747,2.5238976,2.556718,2.4385643,2.1530259,2.1464617,2.4910772,2.9997952,3.245949,2.550154,2.7306669,2.9833848,2.8882053,2.546872,2.5895386,2.793026,2.7864618,2.6026669,2.4582565,2.7634873,2.477949,2.2449234,2.2121027,2.3204105,2.294154,2.540308,2.6223593,2.7602053,2.9472823,2.9407182,2.550154,2.5206156,2.5961027,2.6486156,2.678154,7.069539,6.4590774,5.979898,5.366154,4.7425647,4.6145644,4.44718,4.5062566,4.7360005,4.9329233,4.7491283,5.0051284,5.5138464,6.042257,6.482052,6.8594875,6.6395903,6.6560006,6.944821,7.259898,7.0531287,6.7249236,7.000616,7.2172313,7.1023593,6.770872,7.145026,6.8660517,6.5936418,6.422975,5.8978467,5.405539,5.3891287,5.674667,6.1046157,6.554257,6.951385,7.197539,7.4240007,7.6964107,7.9885135,7.5421543,7.702975,8.260923,9.124104,10.295795,10.696206,11.71036,12.786873,13.4170265,13.128206,13.239796,12.891898,12.983796,13.410462,13.062565,12.931283,12.918155,12.744206,12.406155,12.166565,11.871181,12.130463,12.107488,11.933539,12.721231,12.826258,13.08554,12.412719,11.943385,15.028514,11.008,5.8453336,1.9331284,0.17723078,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.036102567,0.072205134,0.08861539,0.068923086,0.5874872,0.67610264,0.43651286,0.0951795,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016410258,0.12143591,0.25271797,0.21661541,0.108307704,0.049230773,0.01969231,0.006564103,0.009846155,0.006564103,0.055794876,0.08861539,0.06564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.18051283,0.18051283,0.0,0.0,0.0,0.0,0.128,0.35446155,0.48902568,0.73517954,0.6432821,0.6235898,0.81394875,1.0994873,1.6082052,1.4769232,1.1684103,0.9714873,1.020718,1.8806155,1.8773335,1.6836925,1.5327181,1.2242053,1.401436,1.3554872,1.3817437,1.5360001,1.6311796,1.6114873,2.1202054,2.6322052,3.0194874,3.5807183,3.9154875,4.076308,4.640821,5.4941545,5.8453336,5.9995904,6.3376417,6.692103,6.9349747,6.961231,7.8703594,8.385642,9.242257,10.223591,10.167795,10.266257,9.941334,9.93477,10.564924,11.753027,11.250873,10.072617,8.904206,8.064001,7.512616,7.197539,7.2927184,7.351795,7.141744,6.6592827,6.738052,7.1909747,7.328821,7.056411,6.885744,7.8080006,8.14277,8.690872,9.6065645,10.407386,10.758565,11.54954,12.005745,11.808822,11.080206,10.935796,10.505847,10.492719,10.725744,10.174359,11.050668,12.356924,13.190565,13.59754,14.552616,14.897232,14.6871805,15.0777445,16.259283,17.43754,17.286566,17.490053,18.202257,19.219694,19.96472,20.010668,18.458258,17.8839,18.550156,18.379488,17.72636,16.741745,15.924514,15.501129,15.402668,14.050463,12.458668,10.837335,9.622975,9.475283,9.682052,9.511385,10.026668,11.365745,12.740924,12.708103,13.869949,14.519796,14.208001,13.768207,13.594257,14.713437,15.91795,16.856617,18.031591,18.392616,15.973744,13.866668,13.167591,12.954257,10.706052,9.074872,7.9786673,7.4436927,7.5979495,7.240206,6.1505647,5.0674877,4.3290257,3.879385,4.850872,5.225026,5.182359,4.8804107,4.460308,4.57518,3.8531284,3.5314875,3.7940516,3.7743592,3.6496413,4.263385,4.857436,5.097026,5.0477953,5.691077,6.0947695,6.157129,6.0652313,6.308103,5.0477953,3.3017437,3.0260515,5.3366156,10.512411,7.6996927,7.6635904,11.047385,14.674052,11.539693,7.2205133,3.698872,1.6049232,0.9419488,1.0929232,1.0371283,1.0699488,1.273436,1.3915899,0.8336411,1.6147693,2.2482052,2.6486156,2.7011285,2.2744617,2.231795,2.3433847,2.422154,2.674872,3.6824617,4.007385,3.9318976,3.6758976,3.508513,3.757949,4.4898467,4.276513,3.7120004,3.2229745,3.0358977,2.9111798,3.1442053,3.255795,2.9702566,2.1956925,2.349949,2.4155898,2.4910772,2.6584618,3.0030773,2.605949,2.9768207,3.4198978,3.5314875,3.190154,4.082872,4.2896414,4.135385,3.8564105,3.6004105,3.5807183,3.876103,4.027077,3.9023592,3.692308,2.937436,2.6354873,4.5554876,8.011488,9.888822,12.416001,20.089437,25.800207,25.744411,19.403488,12.996924,8.228104,5.1856413,3.5478978,2.550154,2.665026,2.1825643,2.0841026,2.5632823,3.0523078,3.2918978,3.5314875,3.7316926,3.9318976,4.2535386,4.3552823,4.33559,4.345436,4.3552823,4.128821,3.6791797,3.2229745,2.9702566,2.9243078,2.8849232,2.9472823,2.986667,3.1671798,3.4855387,3.7842054,3.9023592,3.9023592,3.9975388,4.1583595,4.128821,4.315898,4.598154,4.9394875,5.284103,5.5663595,5.8190775,6.124308,6.5378466,6.9087186,6.8562055,6.51159,5.835488,5.1987696,4.8049235,4.6802053,4.824616,4.2962055,3.6890259,3.3542566,3.4198978,2.986667,2.3072822,1.7263591,1.3587693,1.0962052,1.0108719,0.82379496,0.6859488,0.6662565,0.7581539,0.58420515,0.6826667,0.73517954,0.6498462,0.56123084,0.63343596,0.7811283,0.96492314,1.1027694,1.0896411,0.97805136,0.88943595,0.827077,0.79097444,0.7581539,0.7581539,1.1027694,1.4703591,1.7132308,1.847795,2.0742567,2.162872,2.156308,2.103795,2.0545642,1.9265642,2.3893335,3.1081028,3.636513,3.4002054,2.349949,1.8674873,1.5655385,1.2898463,1.1093334,1.3653334,1.4408206,1.4244103,1.3850257,1.3522053,1.4375386,1.8970258,2.3433847,2.7273848,3.3411283,3.3050258,3.5249233,3.8071797,4.0533338,4.2436924,4.598154,4.594872,4.5554876,4.634257,4.7917953,4.571898,3.761231,3.1277952,3.0490258,3.495385,1.8576412,3.2754874,5.293949,5.7468724,2.7602053,4.135385,5.5663595,6.009436,5.8486156,6.8988724,6.8496413,6.5870776,6.3967185,6.163693,5.398975,5.2447186,5.366154,5.6287184,5.8978467,6.052103,5.5269747,5.152821,4.7491283,4.2863593,3.892513,3.498667,3.2787695,3.318154,3.5544617,3.7842054,4.279795,5.149539,5.5269747,5.2381544,4.821334,4.3618464,4.2994876,4.4832826,4.8640003,5.5138464,5.976616,6.6067696,7.1023593,7.2631803,6.9710774,6.4032826,7.1581545,7.13518,5.868308,4.516103,4.2371287,7.059693,6.2030773,2.6486156,5.142975,6.7085133,6.491898,6.173539,6.6461544,8.01477,8.448001,8.480822,9.127385,10.246565,10.545232,9.074872,8.136206,7.0892315,6.183385,6.5444107,7.6077952,6.567385,6.4065647,6.8004107,4.089436,2.8258464,2.8553848,3.6824617,4.0369234,1.8674873,3.9680004,3.8432825,3.245949,3.0227695,3.1113849,2.8914874,2.3926156,1.8871796,1.5360001,1.394872,1.2406155,1.014154,0.9616411,1.0371283,0.90912825,0.8008206,0.72861546,0.7811283,0.8763078,0.761436,0.86317956,0.78769237,0.7844103,0.90912825,1.0502565,1.0338463,0.90256417,0.86646163,1.0272821,1.3620514,1.6935385,1.7887181,1.8018463,1.7755898,1.6344616,1.4342566,1.6771283,1.7952822,1.6607181,1.585231,1.7165129,1.5983591,1.7657437,2.1792822,2.228513,2.048,2.103795,2.15959,2.225231,2.550154,2.7602053,3.373949,3.945026,4.1189747,3.6332312,3.7973337,3.5347695,2.9604106,2.3926156,2.349949,2.3105643,2.1267693,2.0053334,1.9889232,1.9298463,2.0742567,1.9528207,1.8346668,1.9232821,2.3794873,1.9003079,1.6738462,1.7033848,1.9495386,2.3368206,2.156308,2.172718,2.3958976,2.6322052,2.477949,2.0217438,1.8642052,2.041436,2.2678976,1.9200002,2.0020514,2.0742567,2.1202054,2.041436,1.657436,1.4211283,1.6114873,1.6344616,1.522872,1.9429746,2.4188719,2.5435898,2.6486156,2.7602053,2.5764105,2.359795,2.6551797,2.9997952,3.045744,2.5600002,2.3893335,2.2711797,2.28759,2.3630772,2.2449234,2.1202054,2.294154,2.7273848,3.058872,2.6256413,2.7831798,2.9046156,2.6978464,2.2514873,2.038154,2.228513,2.7798977,3.0129232,2.8521028,2.802872,2.9538465,2.7602053,2.553436,2.4320002,2.2646155,2.297436,2.225231,2.294154,2.4582565,2.412308,2.3893335,2.5107694,2.5928206,2.6026669,2.6683078,6.6822567,5.8814363,5.733744,5.4482055,4.9493337,4.8607183,4.8082056,4.821334,4.8344617,4.7392826,4.378257,4.71959,5.356308,5.910975,6.2588725,6.5345645,6.422975,6.672411,6.8660517,6.8988724,6.9645133,6.7216415,6.994052,7.0465646,6.8299494,6.987488,7.200821,7.017026,6.948103,6.994052,6.633026,6.163693,6.0750775,6.2687182,6.6395903,7.0957956,7.6570263,8.064001,8.5202055,9.120821,9.82318,8.874667,9.048616,9.737847,10.55836,11.365745,11.67754,12.245335,12.409437,12.104206,11.851488,12.3536415,12.314258,12.514462,12.87877,12.484924,12.704822,12.95754,12.941129,12.57354,12.022155,11.254155,11.785847,12.081232,12.47836,15.189335,13.725539,12.73436,11.195078,10.295795,13.446565,11.35918,6.770872,2.6387694,0.41025645,0.006564103,0.0,0.0,0.0,0.0,0.0,0.016410258,0.12143591,0.14112821,0.072205134,0.072205134,0.16410258,0.94523084,1.0010257,0.256,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.029538464,0.23302566,0.51856416,0.512,0.2231795,0.07876924,0.02297436,0.009846155,0.0,0.009846155,0.09189744,0.08861539,0.0,0.0,0.013128206,0.006564103,0.0,0.0,0.0,0.0,0.04266667,0.04266667,0.0,0.0,0.02297436,0.013128206,0.0,0.072205134,0.35446155,0.51856416,0.7122052,0.86646163,0.9682052,1.0535386,1.5786668,1.4933335,1.1913847,0.9911796,1.1224617,1.4736412,1.3193847,1.1585642,1.2176411,1.4572309,1.7099489,1.5589745,1.5195899,1.6738462,1.6836925,1.6311796,1.7001027,2.1103592,2.809436,3.4888208,3.5249233,3.8465643,4.2338467,4.667077,5.3169236,5.7468724,5.8125134,6.3245134,7.0104623,6.5050263,7.2172313,8.001641,8.667898,9.18318,9.645949,9.639385,9.229129,9.728001,10.925949,11.096616,10.614155,9.160206,8.083693,7.6635904,7.1187696,7.4371285,7.4207187,7.4207187,7.4174366,6.99077,7.4732313,8.15918,8.484103,8.260923,7.6767187,8.385642,8.648206,8.966565,9.67877,10.962052,11.211488,11.785847,12.091078,11.969642,11.69395,11.730052,11.401847,11.283693,11.273847,10.597744,11.21477,12.20595,13.167591,14.17518,15.793232,15.75713,14.976001,14.506668,14.867694,16.042667,15.681643,16.20677,17.050259,17.913437,18.763489,19.242668,17.85436,17.263592,18.005335,18.477951,18.517334,17.765745,16.482462,15.409232,15.766975,14.683899,12.727796,11.178667,10.315488,9.435898,9.202872,9.02236,9.468719,10.640411,12.163283,12.009027,12.678565,13.049437,12.714667,11.992617,13.039591,14.966155,15.465027,14.808617,15.868719,17.847795,17.490053,16.134565,14.795488,14.185027,11.290257,9.15036,7.821129,7.240206,7.200821,7.50277,6.6494365,5.6385646,4.9526157,4.5423594,5.080616,5.5236926,5.2512827,4.4340515,4.023795,4.269949,3.69559,3.2328207,3.2820516,3.7316926,4.0008206,4.673641,5.2578464,5.467898,5.2512827,5.8814363,5.970052,5.7074876,5.648411,6.7183595,5.4153852,3.3050258,2.038154,3.4297438,9.462154,6.488616,7.328821,13.948719,21.064207,16.141129,12.179693,6.6625648,2.7208207,1.1585642,0.446359,0.51856416,0.7187693,0.90912825,1.024,1.079795,1.3357949,1.9561027,2.674872,3.0096412,2.284308,2.4057438,2.4582565,2.28759,2.2186668,3.0326157,3.8104618,4.017231,3.7021542,3.4100516,4.197744,4.394667,4.0500517,3.5249233,3.0523078,2.7437952,2.3335385,2.4320002,2.7569232,2.7995899,1.8445129,1.5786668,1.8740515,2.2186668,2.4976413,2.9801028,2.92759,3.1573336,3.6069746,3.9876926,3.7809234,4.1911798,4.056616,3.69559,3.370667,3.2951798,3.3509746,3.6562054,3.9253337,4.0369234,4.0402055,3.3411283,2.9965131,4.1813335,7.177847,11.382154,10.712616,16.879591,23.880207,26.870155,22.180105,18.28431,14.25395,10.269539,6.75118,4.342154,4.663795,3.2853336,2.028308,1.8379488,2.8127182,3.4067695,4.1583595,4.6080003,4.8016415,5.287385,5.172513,4.571898,4.1156926,4.0434875,4.210872,3.7448208,3.3345644,3.1081028,3.0194874,2.865231,2.9636924,2.9505644,3.1113849,3.570872,4.276513,4.4701543,4.5522056,4.588308,4.6145644,4.630975,4.841026,5.07077,5.4186673,5.733744,5.605744,6.3934364,7.026872,7.456821,7.643898,7.5552826,6.8562055,6.0356927,5.074052,4.2502565,4.1550775,4.571898,4.3618464,3.9384618,3.6627696,3.8400004,3.629949,2.937436,2.2580514,1.7788719,1.3751796,1.1093334,0.8730257,0.73517954,0.7056411,0.7417436,0.49230772,0.3708718,0.39712822,0.512,0.5546667,0.46276927,0.5907693,0.7811283,0.9517949,1.0896411,0.9714873,0.88943595,0.8402052,0.81066674,0.7515898,0.65969235,0.761436,0.8992821,1.0272821,1.1881026,1.4572309,1.6344616,1.6607181,1.6935385,2.103795,1.8773335,2.0742567,2.865231,3.8334363,3.9614363,2.9735386,2.4549747,2.103795,1.7985642,1.5786668,1.7099489,1.6377437,1.5589745,1.5524104,1.5688206,1.5163078,1.8149745,2.294154,2.806154,3.2098465,3.1967182,3.370667,3.6562054,3.95159,4.135385,4.4045134,4.647385,4.57518,4.1485133,3.5774362,4.069744,4.1583595,4.2896414,4.525949,4.5390773,1.7723079,2.4713848,4.8607183,6.373744,3.6463592,2.0512822,3.820308,5.917539,6.9021544,6.918565,6.5247183,6.166975,6.058667,6.058667,5.661539,5.723898,5.8256416,5.98318,6.1472826,6.183385,5.4613338,4.785231,4.414359,4.4406157,4.8016415,4.4767184,3.8301542,3.387077,3.3903592,3.7743592,3.8334363,4.3552823,4.841026,4.9788723,4.6244106,4.4340515,4.673641,4.8771286,4.9526157,5.1626673,5.609026,6.6592827,7.4863596,7.643898,7.069539,6.3212314,7.653744,7.1483083,4.7589746,4.3027697,2.6847181,3.3641028,3.3936412,2.8553848,4.8607183,5.7042055,5.7731285,5.7764106,6.2851286,7.722667,8.018052,8.152616,9.035488,10.384411,10.752001,11.539693,12.977232,11.736616,8.4972315,7.939283,8.536616,6.419693,5.330052,5.4974365,3.623385,2.034872,2.2022567,3.3312824,4.0008206,2.156308,4.713026,4.8705645,4.1189747,3.4560003,3.387077,3.1638978,2.546872,2.0250258,1.8051283,1.8018463,1.3587693,1.0043077,0.92553854,1.020718,0.8992821,0.8763078,0.71548724,0.67282057,0.75487185,0.7056411,0.6629744,0.7187693,0.86974365,1.0469744,1.1290257,1.1946667,0.9747693,0.8598975,1.0043077,1.3259488,1.6804104,1.7427694,1.7624617,1.7788719,1.6246156,1.5885129,1.8707694,1.9167181,1.6869745,1.6738462,1.8838975,1.8051283,1.847795,2.103795,2.3466668,2.5928206,2.878359,2.8488207,2.6518977,2.92759,3.0227695,3.8006158,4.4832826,4.5587697,3.7809234,3.754667,3.4822567,3.062154,2.6190772,2.3269746,2.1792822,2.0775387,1.9922053,1.9396925,1.9823592,1.782154,1.8215386,1.7690258,1.7493335,2.3466668,1.9593848,1.6311796,1.5360001,1.7526156,2.2777438,2.103795,1.9856411,1.8838975,1.8281027,1.9068719,1.8937438,1.7066668,1.6508719,1.6902566,1.4276924,1.8149745,2.0676925,2.1267693,2.038154,1.9331284,1.657436,1.5983591,1.6705642,1.8674873,2.2580514,2.4451284,2.2908719,2.1792822,2.2482052,2.3729234,2.3204105,2.5698464,2.8849232,2.993231,2.605949,2.359795,1.9232821,1.8379488,2.1431797,2.3762052,2.3138463,2.3991797,2.7634873,3.2164104,3.249231,3.2853336,3.0916924,2.934154,2.7011285,1.9298463,1.7723079,2.481231,3.0391798,3.0424619,2.7306669,3.0982566,3.0326157,2.8389745,2.6683078,2.5238976,2.15959,1.7362052,1.7001027,1.9626669,1.9232821,2.0939488,2.3302567,2.4418464,2.4615386,2.6322052,6.196513,5.4514875,5.3825645,5.408821,5.2414365,4.896821,4.972308,4.7228723,4.4734364,4.414359,4.6244106,4.4274874,4.709744,5.284103,5.9602056,6.5444107,6.422975,6.4295387,6.47877,6.4032826,5.9503593,5.9634876,6.422975,6.557539,6.488616,7.2336416,7.709539,7.5520005,7.3583593,7.427283,7.781744,7.574975,7.4207187,7.702975,8.109949,7.643898,7.8145647,8.379078,8.966565,9.504821,10.240001,10.469745,10.538668,10.8307705,11.424822,12.084514,12.721231,13.016617,12.740924,12.340514,12.937847,13.098668,12.278154,12.27159,13.082257,12.924719,13.4859495,13.121642,12.786873,12.727796,12.498053,11.250873,12.324103,12.504617,13.124924,20.033642,13.748514,12.196103,12.20595,11.700514,9.6754875,9.734565,7.069539,3.5282054,0.7253334,0.029538464,0.006564103,0.0,0.0,0.0,0.0,0.036102567,0.24615386,0.32164106,0.20676924,0.12143591,0.08533334,0.65312827,0.82379496,0.40369233,0.0,0.0,0.0,0.0,0.0,0.0,0.036102567,0.036102567,0.08533334,0.23302566,0.48902568,0.20676924,0.072205134,0.01969231,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.072205134,0.036102567,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.12143591,0.06235898,0.0,0.0,0.0,0.47589746,0.7417436,0.8566154,1.0272821,1.6016412,1.4080001,1.2570257,1.214359,1.1585642,0.79425645,1.4276924,1.6968206,1.5491283,1.2832822,1.5425643,2.2744617,2.0808206,1.5885129,1.3062565,1.6475899,1.719795,1.9331284,2.0709746,2.3040001,3.1573336,3.3411283,3.626667,4.2240005,4.9854364,5.402257,5.9503593,5.940513,6.1078978,6.482052,6.409847,6.885744,7.3616414,7.896616,8.254359,7.890052,7.755488,8.280616,9.206155,10.108719,10.374565,10.059488,9.101129,8.477539,8.205129,7.3386674,8.438154,8.228104,7.653744,7.6274877,9.019077,10.056206,10.28595,10.20718,9.8363085,8.713847,9.042052,9.4457445,9.816616,10.167795,10.620719,10.400822,10.492719,10.338462,10.41395,12.20595,12.242052,12.288001,12.301129,12.1238985,11.490462,11.149129,11.483898,12.2847185,13.37436,14.634667,14.900514,14.585437,14.578873,14.992412,15.153232,15.00554,15.37313,15.707899,16.088617,17.211079,16.73518,16.09518,15.898257,16.502155,17.988924,17.257027,16.269129,15.00554,13.948719,14.083283,12.960821,12.678565,12.416001,11.657847,10.194052,9.521232,9.435898,9.4916935,9.96759,11.871181,11.579078,11.798975,11.963078,11.858052,11.628308,13.334975,15.904821,16.272411,14.477129,13.673027,15.113848,16.86318,17.424412,16.370872,14.342566,11.303386,8.979693,7.512616,6.885744,6.8955903,6.9349747,6.695385,6.114462,5.4449234,5.2480006,5.408821,5.5663595,4.890257,3.5249233,2.609231,3.0490258,3.3247182,3.2689233,3.121231,3.5249233,4.71959,5.4153852,5.737026,5.8978467,6.180103,6.058667,6.373744,6.0816417,5.609026,6.8660517,5.914257,3.5249233,1.7493335,2.3729234,6.9120007,7.2303596,10.906258,17.8839,22.98749,15.944206,12.150155,7.64718,3.8400004,1.4703591,0.64000005,1.2012309,1.332513,1.3029745,1.3620514,1.7394873,1.3620514,1.8510771,2.5796926,2.7831798,1.5885129,1.9528207,2.3729234,2.6322052,2.740513,2.9604106,3.9122055,3.892513,3.5840003,3.6135387,4.578462,4.2371287,3.4625645,2.865231,2.6223593,2.487795,1.9987694,1.8215386,1.975795,2.2580514,2.2580514,1.6738462,1.5622566,1.7526156,2.1234872,2.6256413,3.0523078,3.3509746,3.7185643,3.9778464,3.5872824,3.7316926,4.017231,3.6693337,2.917744,2.989949,3.1606157,3.5052311,3.7743592,3.9318976,4.1517954,3.5774362,3.0752823,3.259077,5.3037953,10.955488,10.138257,14.329437,18.83241,21.057642,20.50954,20.312616,20.657232,17.27672,11.1064625,8.283898,6.3212314,4.1550775,2.6387694,1.972513,1.6771283,2.300718,3.5282054,4.630975,5.277539,5.5072823,5.802667,5.2512827,4.457026,3.8465643,3.6627696,3.186872,3.0293336,2.9144619,2.6715899,2.2416413,2.2416413,2.5271797,3.045744,3.6758976,4.2272825,4.7622566,5.1626673,5.395693,5.4580517,5.3858466,5.4580517,5.5958977,5.976616,6.422975,6.422975,6.9382567,7.240206,7.5881033,7.824411,7.384616,6.518154,5.7534366,4.818052,3.9712822,3.9811285,4.3716927,4.1780515,3.892513,3.7185643,3.570872,3.948308,3.5872824,3.0654361,2.6453335,2.2416413,1.6935385,1.2537436,0.9485129,0.7778462,0.7187693,0.54482055,0.4201026,0.36758977,0.38400003,0.45620516,0.38400003,0.4660513,0.5874872,0.7122052,0.86974365,1.017436,1.0338463,0.9682052,0.82379496,0.58092314,0.6170257,0.65312827,0.71548724,0.8205129,0.9911796,1.1126155,1.3357949,1.4966155,1.6278975,1.9692309,1.9692309,2.4155898,2.9046156,3.3017437,3.754667,3.6069746,3.0752823,2.4713848,2.0644104,2.0906668,1.9692309,1.7362052,1.5885129,1.6049232,1.7394873,1.8740515,2.3204105,2.5928206,2.6486156,2.868513,3.0884104,3.3345644,3.5446157,3.8301542,4.4996924,4.4406157,4.525949,4.5029745,4.332308,4.210872,3.748103,3.495385,3.9811285,4.893539,5.0510774,2.8422565,1.7657437,3.0490258,5.3924108,4.9887185,3.511795,3.0227695,4.4340515,6.6002054,6.3310776,5.5893335,5.5663595,5.5663595,5.428513,5.540103,5.85518,6.0652313,6.0750775,5.901129,5.6451287,5.3169236,4.8049235,4.2305646,3.9581542,4.59159,4.824616,4.8738465,4.598154,4.141949,3.9220517,3.8728209,3.5314875,3.4527183,3.69559,3.8301542,3.767795,3.5249233,3.5741541,3.9548721,4.273231,4.588308,6.1538467,7.2861543,7.522462,7.584821,6.2785645,5.5302567,4.7425647,3.948308,3.8137438,1.972513,1.7755898,2.5829747,3.751385,4.6539493,3.7382567,4.5522056,5.3825645,5.720616,6.2720003,7.066257,7.3452315,8.766359,10.860309,11.030975,13.315283,15.770258,13.988104,8.562873,5.097026,5.730462,4.5522056,3.9975388,4.31918,3.5872824,1.6082052,1.8740515,3.1967182,4.414359,4.378257,5.684513,5.2053337,4.594872,4.3027697,3.570872,2.9965131,2.7076926,2.4451284,2.03159,1.3718976,0.77456415,0.827077,0.8992821,0.827077,0.8992821,1.1191796,0.90912825,0.7318975,0.7187693,0.65641034,0.8402052,0.88615394,1.0010257,1.214359,1.3718976,1.2635899,1.079795,0.9714873,1.0568206,1.4342566,1.3620514,1.2406155,1.3161026,1.5491283,1.6475899,1.6738462,1.6705642,1.6213335,1.6016412,1.785436,1.7001027,1.6246156,1.7165129,1.9429746,2.0906668,2.934154,3.308308,3.4067695,3.4264617,3.5872824,3.7185643,4.240411,4.647385,4.634257,4.073026,3.7940516,3.761231,3.6496413,3.242667,2.425436,2.0709746,1.8838975,1.847795,1.9823592,2.349949,2.03159,1.9167181,1.8182565,1.7723079,2.028308,1.7493335,1.5885129,1.404718,1.3259488,1.7394873,1.8018463,1.7690258,1.6344616,1.467077,1.4178462,1.3095386,1.3456411,1.4867693,1.5491283,1.2209232,1.4408206,1.7624617,1.9003079,1.8707694,1.9692309,1.9200002,1.8445129,1.8379488,1.9167181,2.0151796,2.2088206,2.103795,2.0676925,2.2153847,2.412308,2.3860514,2.5271797,2.7700515,2.8980515,2.5337439,2.2777438,1.8740515,1.7394873,1.913436,2.0611284,2.1825643,2.422154,2.8258464,3.2853336,3.5544617,3.0916924,2.9669745,3.2164104,3.442872,2.806154,2.0250258,2.2055387,2.5895386,2.7667694,2.6715899,3.1343591,3.5610259,3.639795,3.2820516,2.609231,2.3040001,1.7427694,1.5786668,1.847795,1.9823592,2.2514873,2.1169233,2.1924105,2.5600002,2.793026,6.2818465,5.907693,5.618872,5.58277,5.648411,5.32677,4.969026,4.709744,4.601436,4.588308,4.5029745,4.893539,4.7491283,4.9788723,5.756718,6.5083084,6.6592827,6.8463597,6.5706673,5.986462,5.8781543,6.445949,6.820103,7.197539,7.53559,7.5388722,7.604513,7.4863596,7.6603084,8.185436,8.684308,9.6295395,9.846154,9.442462,8.641642,7.765334,8.093539,8.969847,9.6525135,9.970873,10.325335,10.341744,10.581334,10.978462,11.746463,13.39077,13.929027,13.745232,13.679591,13.919181,14.001232,13.243078,12.73436,12.905026,13.252924,12.35036,12.599796,12.445539,12.314258,12.20595,11.690667,10.866873,11.772718,12.534155,13.804309,18.740515,14.290052,13.423591,14.043899,13.787898,10.003693,6.8430777,4.2994876,2.2482052,0.7581539,0.09189744,0.01969231,0.0,0.0,0.0,0.0,0.006564103,0.055794876,0.07548718,0.055794876,0.049230773,0.072205134,0.8369231,0.8960001,0.17723078,0.0,0.0,0.0,0.0,0.0,0.0,0.07548718,0.1148718,0.18707694,0.46276927,1.1946667,0.6432821,0.26256412,0.08533334,0.049230773,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.16738462,0.16082053,0.0,0.0,0.0,0.108307704,0.108307704,0.068923086,0.34133336,0.09189744,0.013128206,0.0,0.07548718,0.37743592,0.190359,0.44964105,0.7581539,0.90912825,0.90584624,0.86646163,1.086359,1.204513,1.1257436,1.014154,1.394872,1.3423591,1.4244103,1.719795,1.8084104,2.3663592,2.172718,1.9200002,1.9035898,2.0512822,2.2711797,2.5993848,3.0129232,3.3542566,3.3280003,3.3280003,3.5938463,3.9975388,4.46359,4.9854364,5.467898,6.304821,6.954667,7.030154,6.3245134,6.3901544,6.4754877,6.951385,7.4732313,7.0104623,7.2960005,8.385642,9.596719,10.620719,11.523283,10.210463,8.681026,7.634052,7.3550773,7.719385,8.2904625,7.506052,6.747898,7.273026,10.226872,10.660104,11.32636,12.015591,12.100924,10.518975,9.990565,9.987283,10.292514,10.679795,10.939077,10.59118,9.947898,9.26195,9.242257,11.047385,11.414975,11.897437,12.232206,12.2157955,11.697231,11.648001,11.546257,11.753027,12.422565,13.472821,13.869949,14.250668,15.337027,16.406975,15.287796,15.688207,15.048206,14.473847,14.611693,15.635694,15.346873,15.156514,15.409232,15.763694,15.182771,14.50995,14.903796,15.07118,14.585437,13.899488,12.875488,13.131488,13.338258,12.87877,11.851488,10.459898,9.665642,9.275078,9.416205,10.528821,10.929232,11.073642,11.126155,11.286975,11.785847,14.628103,16.564514,16.91241,15.970463,15.038361,14.70359,15.796514,17.076513,17.207796,14.769232,11.71036,9.301334,7.5979495,6.7314878,6.9087186,6.409847,6.2720003,6.2030773,6.0619493,5.8486156,5.106872,4.6605134,4.1156926,3.2886157,2.2055387,2.2153847,2.7503593,2.9571285,2.8324106,3.2065644,4.2568207,4.7360005,5.3924108,6.1013336,5.874872,5.832206,6.1078978,6.0160003,5.7534366,6.416411,5.87159,3.5872824,1.7427694,1.3489232,2.2383592,6.47877,11.08677,15.894976,17.54913,9.501539,8.65477,5.2348723,2.5238976,1.4769232,0.7253334,1.1913847,1.5819489,1.8642052,2.0775387,2.349949,2.3926156,2.3663592,2.5140514,2.6453335,2.1234872,2.2055387,2.4615386,2.7142565,2.9111798,3.131077,3.7907696,4.0500517,3.876103,3.6069746,3.9548721,3.5052311,2.7437952,2.1891284,2.0053334,1.9987694,1.8149745,1.6475899,1.7460514,2.0611284,2.2449234,1.9528207,1.5589745,1.4309745,1.7099489,2.3204105,2.8750772,3.5413337,3.9942567,4.0533338,3.6824617,3.43959,3.7349746,3.6036925,3.0523078,3.0752823,2.934154,3.186872,3.495385,3.7382567,4.017231,3.5511796,3.3772311,3.501949,4.8836927,9.442462,13.751796,11.825232,9.478565,11.23118,20.299488,21.861746,21.35959,18.41559,14.260514,11.716924,8.940309,6.7610264,4.4767184,2.4910772,2.3269746,1.913436,2.6551797,3.4034874,3.7448208,4.007385,4.788513,4.9920006,4.6900516,4.1780515,3.9548721,3.6069746,3.3575387,3.1245131,2.9472823,2.9997952,2.8816411,2.8225644,2.9604106,3.4166157,4.2863593,4.6966157,4.955898,5.031385,4.9427695,4.7524104,4.8049235,4.97559,5.2414365,5.4580517,5.349744,5.9995904,6.314667,6.616616,6.87918,6.7150774,5.98318,5.4514875,4.824616,4.1747694,3.9351797,4.0992823,3.8990772,3.6069746,3.3312824,3.0096412,3.2131286,3.1048207,2.92759,2.7766156,2.609231,2.3236926,1.9200002,1.4539489,1.014154,0.7187693,0.6629744,0.54482055,0.43323082,0.36758977,0.3708718,0.40697438,0.48574364,0.6170257,0.72861546,0.6629744,0.90584624,1.020718,0.9944616,0.8172308,0.4955898,0.5021539,0.6104616,0.7056411,0.7844103,0.955077,0.92225647,1.1782565,1.467077,1.6935385,1.9200002,2.0841026,2.3630772,2.6945643,2.9669745,3.0096412,2.9407182,2.92759,2.7470772,2.409026,2.1398976,1.9495386,1.7001027,1.5425643,1.6049232,1.9823592,2.176,2.300718,2.5206156,2.8553848,3.1737437,3.1409233,3.3017437,3.6168208,4.1222568,4.9394875,4.568616,4.46359,4.210872,3.945026,4.3716927,4.6966157,4.4077954,4.3618464,4.886975,5.76,4.709744,3.1967182,2.4910772,2.6420515,2.4746668,5.1200004,4.1452312,3.8990772,5.4153852,6.4065647,5.2611284,5.35959,5.602462,5.549949,5.4153852,5.431795,5.651693,5.8486156,5.9470773,6.0225644,5.7731285,5.7107697,5.3103595,4.630975,4.348718,4.6867695,5.1954875,5.3169236,5.1298466,5.349744,5.428513,4.2830772,3.6332312,3.8662567,4.0500517,3.5577438,3.3476925,3.4921029,3.876103,4.1747694,4.6867695,6.1440005,7.4469748,8.146052,8.4512825,5.835488,4.578462,3.9351797,3.7054362,4.204308,3.446154,3.170462,3.5807183,4.1485133,3.6168208,4.1452312,5.3727183,6.1538467,6.245744,6.294975,7.0400004,6.987488,8.044309,10.203898,11.556104,11.546257,11.516719,9.586872,6.0258465,3.242667,3.5544617,3.5971284,4.2207184,5.074052,4.6244106,2.9768207,4.2994876,5.218462,4.8607183,4.844308,5.024821,4.8082056,4.650667,4.5489235,4.023795,2.9997952,2.605949,2.28759,1.8313848,1.3489232,0.83035904,0.90912825,0.9419488,0.8205129,0.9616411,1.0929232,1.0436924,1.0272821,1.0535386,0.92553854,1.1093334,1.1454359,1.1257436,1.1158975,1.1651284,1.1158975,1.0568206,1.0535386,1.1355898,1.2865642,1.2832822,1.3554872,1.3423591,1.2931283,1.4900514,1.4834872,1.5327181,1.595077,1.6278975,1.5786668,1.7755898,2.0250258,2.0545642,1.9823592,2.3335385,2.9538465,3.387077,3.7349746,3.9187696,3.7087183,4.2436924,5.037949,5.3202057,4.9952826,4.647385,4.1517954,4.276513,4.010667,3.1737437,2.412308,2.2449234,1.9331284,1.7558975,1.8215386,2.0808206,1.8609232,1.7493335,1.7329233,1.7329233,1.5885129,1.4375386,1.2471796,1.1290257,1.1684103,1.4473847,1.2832822,1.3423591,1.3357949,1.211077,1.1618463,1.0929232,1.204513,1.2668719,1.1618463,0.892718,1.0929232,1.3423591,1.5589745,1.7329233,1.9200002,1.9987694,1.9823592,1.8838975,1.7952822,1.8904617,2.0775387,1.9889232,1.9429746,2.0578463,2.2646155,2.231795,2.3171284,2.546872,2.7241027,2.4352822,2.8422565,2.92759,2.6617439,2.1858463,1.8051283,2.1300514,2.3630772,2.7076926,3.117949,3.2984617,3.1967182,3.0162053,3.006359,3.05559,2.6847181,2.100513,1.9167181,1.9987694,2.2711797,2.7306669,2.7569232,2.993231,3.2098465,3.1573336,2.5862565,2.425436,1.8510771,1.5786668,1.7985642,2.166154,2.356513,2.2678976,2.2744617,2.3794873,2.231795,5.6320004,5.3891287,5.4383593,5.605744,5.674667,5.395693,5.3037953,5.3234878,5.3037953,5.1954875,5.037949,5.179077,5.041231,5.0543594,5.3202057,5.5926156,5.9470773,6.2523084,6.117744,5.681231,5.622154,6.2194877,6.5280004,6.8332314,7.1154876,7.020308,7.2664623,7.4830775,7.9458466,8.710565,9.596719,10.473026,10.371283,9.731283,8.966565,8.474257,8.6580515,9.6295395,10.394258,10.696206,11.040821,11.32636,11.657847,11.933539,12.458668,13.955283,14.086565,13.787898,13.90277,14.34913,14.139078,14.027489,13.791181,13.318565,12.731078,12.3536415,12.386462,12.081232,12.1238985,12.324103,11.634872,10.939077,11.572514,13.052719,15.29436,18.619078,16.699078,16.098463,16.075489,15.254975,11.631591,5.8125134,2.9965131,1.5130258,0.5349744,0.07876924,0.016410258,0.0,0.0,0.0,0.0,0.029538464,0.02297436,0.013128206,0.036102567,0.15753847,0.28225642,0.73517954,0.69251287,0.39712822,1.1520001,0.44307697,0.11158975,0.006564103,0.0,0.0,0.45292312,0.84348726,1.1946667,1.3128207,0.8041026,0.46933338,0.2986667,0.18379489,0.07548718,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.2231795,0.33476925,0.2986667,0.40369233,0.31507695,0.256,0.18379489,0.14112821,0.22646156,0.29538465,0.12471796,0.0,0.03938462,0.190359,0.33476925,0.4266667,0.5415385,0.7187693,0.9517949,0.9747693,1.1585642,1.3292309,1.3686155,1.2242053,1.5130258,1.5885129,1.4572309,1.3357949,1.657436,1.8904617,1.9429746,2.2153847,2.6256413,2.5993848,2.674872,2.930872,3.2787695,3.5478978,3.4625645,3.8531284,4.325744,4.6112823,4.821334,5.4580517,5.182359,5.917539,6.6560006,6.7872825,6.0717955,6.2785645,6.498462,6.925129,7.282872,6.8463597,7.4108725,8.385642,9.6754875,10.886565,11.32636,9.682052,8.011488,6.892308,6.5083084,6.669129,7.1876926,6.941539,6.9054365,7.762052,9.905231,9.777231,10.597744,11.739899,12.363488,11.418258,10.528821,10.299078,10.486155,10.962052,11.739899,11.661129,10.860309,9.787078,9.170052,10.016821,10.217027,10.387693,10.686359,11.004719,10.962052,11.132719,11.136001,11.316514,11.83836,12.708103,13.252924,13.771488,14.985847,16.216616,15.382976,15.642258,14.841437,14.217847,14.329437,15.051488,14.660924,14.5952835,14.50995,14.024206,12.704822,13.069129,13.804309,14.280207,14.427898,14.752822,13.787898,14.319591,14.519796,13.761642,12.632616,11.0145645,10.164514,9.734565,9.609847,9.908514,9.970873,10.203898,10.528821,11.1064625,12.337232,15.38954,16.091898,15.937642,15.622565,15.031796,14.516514,14.401642,14.930053,15.307488,13.715693,11.178667,9.222565,7.6734366,6.5837955,6.2523084,6.242462,6.180103,6.265436,6.4590774,6.482052,4.8377438,3.7940516,3.2000003,2.7667694,2.0611284,1.9856411,2.281026,2.4516926,2.5304618,3.0720003,3.757949,4.381539,5.0149746,5.651693,6.2194877,6.2916927,6.6592827,6.6822567,6.226052,5.671385,5.3694363,3.6594875,2.0906668,1.4211283,1.6082052,6.196513,10.601027,14.224411,14.14236,5.1232824,5.146257,3.6726158,2.1792822,1.3489232,1.086359,1.6213335,1.8543591,2.1169233,2.5271797,2.9965131,3.4494362,2.7733335,2.5009232,2.8455386,2.6880002,2.665026,2.5993848,2.6322052,2.7733335,2.8914874,3.4822567,4.0303593,3.95159,3.4002054,3.259077,2.9078977,2.28759,1.8346668,1.7099489,1.8313848,1.8543591,1.7001027,1.7526156,2.0808206,2.4451284,2.231795,1.6147693,1.4145643,1.8313848,2.4352822,2.993231,3.6463592,4.0434875,4.194462,4.450462,3.9384618,3.7349746,3.564308,3.370667,3.318154,2.8914874,2.9505644,3.2196925,3.5478978,3.8990772,3.570872,3.5774362,3.8564105,4.6933336,6.7282057,11.024411,10.9915905,9.068309,9.5835905,18.773335,24.234669,20.578463,15.849027,13.479385,12.288001,10.000411,8.710565,7.125334,5.100308,3.639795,2.103795,1.782154,2.1398976,2.7667694,3.4034874,4.59159,4.8672824,4.650667,4.4110775,4.670359,4.2929235,3.9778464,3.7743592,3.6857438,3.6660516,3.6562054,3.2820516,3.0391798,3.1934361,3.7710772,4.457026,4.923077,5.0543594,4.9526157,4.923077,4.699898,4.6834874,4.8738465,5.156103,5.3005133,5.802667,6.2096415,6.373744,6.2752824,6.0160003,5.720616,5.8256416,5.6352825,5.093744,4.781949,4.585026,4.1780515,3.6758976,3.1934361,2.8882053,3.1409233,2.9735386,2.878359,2.9669745,2.9669745,2.8258464,2.3926156,1.8116925,1.2274873,0.77128214,0.761436,0.6104616,0.44964105,0.36102566,0.3708718,0.3511795,0.39712822,0.51856416,0.6235898,0.53825647,0.6826667,0.81394875,0.8336411,0.7220513,0.5284103,0.46276927,0.60061544,0.6695385,0.6465641,0.7811283,0.8172308,0.9944616,1.2274873,1.4736412,1.7427694,1.7657437,1.8149745,2.1202054,2.5829747,2.740513,2.612513,2.6518977,2.6256413,2.3958976,1.9232821,1.6049232,1.5491283,1.5819489,1.6475899,1.8248206,2.1858463,2.4484105,2.809436,3.2262566,3.4067695,3.045744,3.2328207,3.692308,4.138667,4.2830772,4.086154,4.1452312,4.073026,3.9220517,4.161641,4.6933336,4.8705645,4.8836927,4.95918,5.349744,5.21518,4.640821,3.9844105,3.3936412,2.806154,3.5741541,3.751385,4.007385,4.8377438,6.560821,5.901129,5.8157954,5.737026,5.504,5.330052,5.293949,5.3825645,5.605744,5.924103,6.2752824,6.232616,6.058667,5.7009234,5.3136415,5.2480006,5.366154,5.7731285,6.0028725,5.9634876,5.927385,5.9995904,4.824616,4.1517954,4.342154,4.3716927,3.8071797,3.6135387,3.826872,4.263385,4.4996924,5.3366156,6.2785645,6.803693,6.747898,6.2884107,4.7589746,4.3027697,4.7983594,5.4908724,5.0084105,3.7874875,3.495385,4.1583595,5.0018463,4.44718,4.5095387,5.0510774,5.87159,6.2785645,5.0838976,5.1954875,5.3858466,6.2916927,7.781744,8.960001,9.304616,8.490667,6.685539,4.598154,3.4724104,3.4789746,3.767795,4.529231,5.2545643,4.7360005,3.892513,4.827898,5.5958977,5.6254363,5.737026,5.3234878,5.1265645,4.8672824,4.5029745,4.20759,3.2131286,2.7044106,2.0841026,1.3423591,1.086359,0.95835906,1.0436924,1.0108719,0.90256417,1.142154,1.0765129,1.0929232,1.204513,1.3620514,1.4506668,1.7066668,1.4900514,1.2406155,1.142154,1.1585642,1.3784616,1.6147693,1.7526156,1.7493335,1.6278975,1.6607181,1.6836925,1.6278975,1.5655385,1.6968206,1.522872,1.522872,1.6049232,1.6607181,1.5425643,1.9167181,2.03159,1.9790771,2.1103592,3.0654361,3.7776413,3.8465643,3.9712822,4.2272825,4.066462,4.4767184,5.074052,5.2611284,5.0149746,4.8836927,4.128821,3.9056413,3.7973337,3.4658465,2.6847181,2.5271797,2.048,1.7558975,1.7657437,1.8215386,1.6114873,1.4244103,1.332513,1.2996924,1.1881026,1.1093334,1.0962052,1.083077,1.0962052,1.2438976,1.0404103,1.148718,1.1552821,1.024,1.1093334,1.1848207,1.0994873,0.98133343,0.86974365,0.7187693,0.9124103,1.079795,1.3423591,1.7066668,2.0545642,1.9954873,2.048,2.100513,2.1234872,2.162872,2.3171284,2.228513,2.162872,2.2121027,2.2646155,2.1989746,2.3138463,2.4418464,2.4418464,2.2088206,2.7766156,3.0916924,3.1343591,2.8914874,2.3696413,2.5074873,2.4484105,2.5961027,2.9702566,3.2262566,2.993231,2.7437952,2.678154,2.7109745,2.4713848,2.0742567,1.7001027,1.6147693,1.8937438,2.425436,2.3466668,2.428718,2.5074873,2.4549747,2.176,2.1497438,1.6902566,1.5622566,1.8412309,1.9364104,2.0217438,1.972513,1.8543591,1.7657437,1.8445129,5.333334,5.031385,5.2480006,5.4908724,5.5269747,5.3825645,5.3070774,5.3136415,5.2742567,5.1922054,5.2020516,5.3005133,5.1626673,5.041231,4.962462,4.7327185,5.2545643,5.61559,5.6352825,5.4580517,5.5532312,5.986462,6.3179493,6.452513,6.419693,6.38359,6.8955903,7.4141545,8.1066675,9.042052,10.19077,10.453334,10.092308,9.741129,9.616411,9.488411,9.4916935,10.31877,11.122872,11.69395,12.4685135,12.754052,13.216822,13.574565,13.915898,14.720001,14.523078,14.490257,14.506668,14.437745,14.112822,15.067899,15.058052,14.293334,13.466257,13.7386675,12.944411,12.304411,12.2847185,12.672001,12.563693,11.74318,12.018872,14.093129,16.961643,17.91672,17.355488,16.886156,16.531694,15.442053,11.907283,6.701949,3.114667,1.0896411,0.2855385,0.06235898,0.04594872,0.04594872,0.029538464,0.0,0.0,0.029538464,0.036102567,0.09189744,0.18379489,0.21333335,0.45620516,0.58092314,0.6892308,0.9944616,1.8543591,0.61374366,0.128,0.006564103,0.009846155,0.02297436,0.5874872,1.0010257,1.5786668,1.8149745,0.37743592,0.21661541,0.20020515,0.19364104,0.13456412,0.01969231,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.14441027,0.25271797,0.3446154,0.6170257,0.4660513,0.4955898,0.42338464,0.2100513,0.055794876,0.36102566,0.28882053,0.25271797,0.3314872,0.26256412,0.41025645,0.4201026,0.48902568,0.6826667,0.93866676,1.2603078,1.3456411,1.3095386,1.2537436,1.2898463,1.4998976,1.6377437,1.4276924,1.1027694,1.3817437,1.3784616,1.9265642,2.5074873,2.8488207,2.934154,3.1638978,3.370667,3.6693337,3.9745643,3.9876926,4.4734364,4.9920006,5.093744,4.972308,5.47118,5.077334,5.609026,6.1997952,6.5017443,6.6822567,6.747898,7.4896417,8.260923,8.5202055,7.834257,8.369231,8.717129,9.636104,10.738873,10.469745,8.858257,8.100103,7.194257,6.1013336,5.7534366,6.0192823,6.422975,7.02359,7.975385,9.55077,9.114257,9.803488,10.650257,11.418258,12.609642,11.756309,11.030975,10.686359,10.935796,11.959796,12.557129,11.890873,10.660104,9.632821,9.626257,9.370257,9.393231,9.7673855,10.341744,10.755282,10.965334,11.136001,11.52,12.104206,12.629334,13.124924,13.371078,14.273643,15.537232,15.645539,15.123693,14.454155,14.260514,14.716719,15.53395,14.792206,14.04718,13.203693,12.22236,11.122872,12.051693,12.882052,13.53518,14.171899,15.209026,14.191591,14.237539,14.221129,13.590976,12.360206,11.585642,10.532104,9.984001,10.069334,10.256411,10.157949,10.174359,10.489437,11.244308,12.547283,15.202463,15.248411,14.759386,14.54277,14.148924,13.938873,13.446565,13.062565,12.750771,12.084514,10.509129,9.02236,7.77518,6.7610264,5.8190775,6.0356927,6.180103,6.2785645,6.370462,6.49518,4.5456414,3.314872,2.8553848,2.789744,2.297436,2.041436,1.9790771,1.975795,2.1202054,2.7076926,3.4822567,4.06318,4.568616,5.2020516,6.2490263,6.8332314,7.0498466,7.1680007,6.921847,5.5105643,5.182359,3.9712822,2.4976413,1.4441026,1.529436,5.0477953,8.874667,11.506873,10.65354,3.239385,3.4658465,2.674872,1.7001027,1.1158975,1.2504616,2.0151796,2.156308,2.2580514,2.609231,3.2164104,3.5577438,2.878359,2.6157951,3.058872,3.3345644,2.9604106,2.9078977,2.9472823,2.9440002,2.8914874,3.3017437,3.9089234,3.82359,3.0851285,2.6617439,2.484513,2.0841026,1.6968206,1.5327181,1.7690258,1.9626669,1.9593848,2.0611284,2.3893335,2.865231,2.7602053,1.9462565,1.6016412,2.0151796,2.5862565,3.0227695,3.5052311,3.7874875,4.017231,4.7360005,4.5522056,4.06318,3.8334363,3.9154875,3.8432825,3.3936412,3.2754874,3.31159,3.4625645,3.8137438,3.5577438,3.387077,3.570872,4.1124105,4.7524104,8.201847,10.912822,11.024411,10.692924,16.082052,22.212925,19.114668,15.596309,14.874257,14.585437,13.978257,12.005745,9.961026,8.1066675,5.677949,3.0391798,1.463795,1.1618463,1.8674873,2.8291285,3.9286156,4.2469745,4.309334,4.571898,5.402257,4.8607183,4.7327185,4.650667,4.4865646,4.348718,4.4832826,4.1124105,3.6496413,3.314872,3.1540515,3.754667,4.3749747,4.7327185,4.821334,4.923077,4.7294364,4.673641,4.788513,5.0543594,5.398975,5.72718,6.196513,6.2884107,5.9503593,5.5991797,5.5663595,5.989744,6.0816417,5.6976414,5.32677,4.9362054,4.4832826,3.9417439,3.4166157,3.1507695,3.31159,3.2361028,3.0916924,3.0391798,3.2295387,3.058872,2.5829747,1.9790771,1.401436,0.955077,0.8467693,0.74830776,0.6071795,0.44964105,0.380718,0.34789747,0.35774362,0.42994875,0.508718,0.47589746,0.53825647,0.63343596,0.702359,0.7089231,0.6432821,0.50543594,0.6301539,0.65969235,0.56123084,0.6301539,0.7778462,0.90912825,1.020718,1.142154,1.3226668,1.3226668,1.3554872,1.7558975,2.3696413,2.5632823,2.4484105,2.3893335,2.3827693,2.297436,1.8904617,1.4244103,1.3686155,1.4769232,1.595077,1.6771283,2.0578463,2.4352822,2.858667,3.2820516,3.570872,3.3641028,3.4921029,3.895795,4.2502565,3.9384618,3.7382567,3.8432825,3.948308,3.9811285,4.1124105,4.4373336,4.8344617,4.9460516,4.8049235,4.824616,5.07077,5.5138464,5.546667,5.0149746,4.2240005,3.3969233,3.5216413,3.7710772,4.2568207,6.0258465,5.9667697,5.9503593,6.0816417,6.170257,5.7468724,5.737026,5.986462,6.180103,6.3343596,6.7872825,6.5739493,6.2162056,5.933949,5.861744,6.048821,5.9667697,6.091488,6.23918,6.232616,5.901129,5.76,4.9821544,4.673641,4.893539,4.6572313,4.2305646,4.1124105,4.279795,4.522667,4.417641,5.5565133,6.23918,6.0783596,5.149539,3.9811285,3.4625645,4.4340515,6.0652313,6.9809237,5.2709746,3.0687182,2.665026,3.4560003,4.4077954,4.069744,5.7829747,5.3431797,5.284103,5.609026,3.8071797,3.748103,4.1747694,5.3202057,6.6822567,7.00718,7.3025646,6.803693,6.012718,5.3760004,5.2676926,4.906667,5.097026,5.717334,6.2227697,5.6451287,4.923077,4.969026,5.2545643,5.4908724,5.6352825,5.5007186,5.284103,4.7392826,4.076308,3.9647183,3.56759,2.7864618,1.9626669,1.3029745,0.88615394,0.9517949,1.0338463,1.0666667,1.1027694,1.2931283,1.1979488,1.2668719,1.401436,1.5491283,1.7001027,1.9068719,1.6443079,1.4244103,1.4178462,1.4408206,1.9331284,2.2121027,2.3401027,2.3433847,2.2121027,2.2482052,2.1300514,1.9790771,1.8674873,1.847795,1.7362052,1.723077,1.7952822,1.8806155,1.8543591,2.0939488,2.1891284,2.3433847,2.733949,3.515077,4.2863593,4.266667,4.315898,4.6112823,4.6539493,4.7917953,5.0477953,5.097026,4.893539,4.663795,4.082872,3.5577438,3.3509746,3.2689233,2.678154,2.5928206,2.1267693,1.7952822,1.7099489,1.5655385,1.3653334,1.1093334,0.9353847,0.86974365,0.8467693,0.9124103,0.9682052,0.9616411,0.94523084,1.0666667,0.9747693,1.020718,1.0043077,0.9419488,1.0535386,1.1126155,0.96492314,0.78769237,0.65969235,0.56451285,0.75487185,0.8763078,1.1552821,1.5655385,1.8412309,1.8149745,1.9167181,2.0709746,2.2055387,2.2547693,2.3302567,2.3433847,2.3926156,2.4352822,2.294154,2.3105643,2.3762052,2.3663592,2.3072822,2.349949,2.7437952,3.0227695,3.2853336,3.4133337,3.0490258,2.8521028,2.7142565,2.733949,2.9144619,3.1573336,2.7076926,2.3893335,2.2449234,2.2121027,2.1497438,1.8445129,1.6147693,1.6180514,1.8084104,1.9331284,1.8149745,2.028308,2.1300514,1.9856411,1.785436,1.9790771,1.6869745,1.6738462,1.9232821,1.6377437,1.6640002,1.6738462,1.5655385,1.401436,1.4145643,5.6320004,5.330052,5.405539,5.4941545,5.4908724,5.546667,5.1364107,4.7589746,4.5423594,4.5456414,4.7622566,5.182359,4.9329233,4.7458467,4.7392826,4.4406157,4.9296412,5.2480006,5.3234878,5.3169236,5.6320004,5.802667,6.2916927,6.445949,6.242462,6.2916927,6.5969234,7.200821,8.060719,9.114257,10.253129,9.993847,9.662359,9.764103,10.19077,10.236719,10.148104,10.79795,11.602052,12.498053,13.965129,14.168616,14.920206,15.563488,15.849027,15.894976,15.717745,16.032822,15.793232,14.998976,14.697027,16.019693,16.20349,15.852309,15.540514,15.832617,13.932309,13.285745,13.056001,13.049437,13.705847,12.819694,12.678565,14.989129,18.182566,17.43754,16.728617,16.059078,15.520822,14.280207,10.601027,7.7292314,3.5216413,0.77456415,0.12471796,0.049230773,0.07876924,0.4594872,0.42994875,0.013128206,0.009846155,0.006564103,0.04594872,0.21661541,0.38728207,0.19692309,0.48246157,0.60389745,1.0338463,1.6311796,1.6738462,0.40369233,0.03938462,0.013128206,0.02297436,0.049230773,0.4135385,0.48574364,1.0075898,1.529436,0.4135385,0.27569234,0.14769232,0.15425642,0.21333335,0.036102567,0.01969231,0.006564103,0.0,0.0,0.0032820515,0.006564103,0.068923086,0.0951795,0.14769232,0.4266667,0.30194873,0.5907693,0.63343596,0.30194873,0.0,0.26584616,0.36102566,0.5513847,0.7581539,0.5481026,0.34789747,0.36430773,0.52512825,0.7056411,0.761436,1.4178462,1.5031796,1.2471796,1.0043077,1.2406155,1.3193847,1.3128207,1.2537436,1.2242053,1.332513,1.3423591,2.281026,2.8816411,2.917744,3.2229745,3.5314875,3.6135387,3.9680004,4.522667,4.6572313,4.896821,5.2512827,5.1200004,4.713026,5.0477953,5.661539,6.340924,6.6592827,6.9120007,8.113232,7.6110773,8.65477,9.882257,10.371283,9.616411,9.764103,9.380103,9.5606165,10.04636,9.242257,7.9130263,8.461129,8.1066675,6.5772314,6.11118,5.8912826,6.4557953,7.072821,7.79159,9.45559,9.31118,9.938052,10.112,10.404103,13.144616,12.724514,11.664412,10.81436,10.689642,11.457642,12.750771,12.370052,11.227899,10.125129,9.731283,9.199591,9.42277,9.980719,10.607591,11.185231,11.398565,11.503591,11.884309,12.471796,12.740924,13.213539,13.157744,13.607386,14.631386,15.314053,14.293334,13.948719,14.316309,15.254975,16.459488,15.274668,13.705847,12.386462,11.493745,10.761847,11.30995,12.235488,13.193847,14.037334,14.785643,13.768207,12.911591,12.714667,12.747488,11.667693,11.963078,10.676514,10.052924,10.614155,11.16554,11.32636,11.152411,11.208206,11.644719,12.1928215,14.17518,14.358975,13.850258,13.239796,12.580104,12.678565,12.754052,12.0549755,10.889847,10.610872,9.911796,8.661334,7.778462,7.213949,5.976616,5.7764106,6.0061545,6.052103,5.83877,5.8256416,4.240411,3.242667,3.0424619,3.2032824,2.6289232,2.1858463,1.8970258,1.7099489,1.7263591,2.1792822,3.3378465,3.7120004,4.1911798,4.9952826,5.661539,6.941539,6.944821,7.128616,7.3583593,5.904411,5.2611284,4.2338467,2.6912823,1.1913847,0.97805136,3.121231,6.692103,8.454565,7.181129,3.6430771,3.6627696,2.1497438,1.1290257,1.1651284,1.3489232,2.2219489,2.537026,2.5238976,2.5173335,2.9538465,2.8356924,2.7044106,2.7142565,3.0030773,3.7054362,2.9965131,3.2623591,3.6135387,3.620103,3.3017437,3.3214362,3.754667,3.6168208,2.8389745,2.2646155,2.2022567,2.048,1.7493335,1.4966155,1.7460514,2.0906668,2.3729234,2.6256413,2.934154,3.436308,3.564308,2.665026,2.038154,2.162872,2.674872,2.9440002,3.249231,3.4592824,3.7021542,4.397949,4.8049235,4.46359,4.279795,4.457026,4.466872,4.1714873,4.013949,3.8334363,3.6627696,3.7349746,3.5938463,3.062154,2.858667,3.2623591,4.1058464,7.640616,11.096616,12.402873,12.160001,13.643488,15.753847,15.970463,17.024002,19.012924,19.40677,19.452719,15.392821,11.959796,10.41395,8.54318,5.9667697,3.0096412,1.4178462,1.5392822,2.3040001,3.1573336,3.7087183,4.0992823,4.6276927,5.7796926,5.2053337,5.3202057,5.32677,5.07077,5.041231,5.113436,4.9362054,4.4340515,3.6791797,2.9111798,2.9735386,3.4198978,3.945026,4.332308,4.466872,4.6178465,4.7228723,4.8114877,4.962462,5.3005133,5.5729237,5.973334,6.0717955,5.8125134,5.5138464,5.3825645,5.61559,5.7534366,5.579488,5.1200004,4.7917953,4.5029745,4.1780515,3.8400004,3.629949,3.5971284,3.6890259,3.4198978,2.989949,3.2754874,2.9801028,2.5435898,2.0545642,1.6016412,1.276718,0.9878975,0.9714873,0.8992821,0.6695385,0.41025645,0.41025645,0.39056414,0.39712822,0.42994875,0.44964105,0.5021539,0.5546667,0.64000005,0.7417436,0.77128214,0.5973334,0.65641034,0.6859488,0.6104616,0.5677949,0.71548724,0.86646163,0.9353847,0.9189744,0.8992821,1.0568206,1.270154,1.7296412,2.2482052,2.281026,2.231795,2.1234872,2.0939488,2.1234872,2.0217438,1.4933335,1.2635899,1.2931283,1.4802053,1.6640002,1.9298463,2.2711797,2.6354873,3.0523078,3.6332312,3.8334363,3.8498464,4.076308,4.378257,4.092718,3.6660516,3.620103,3.7021542,3.817026,4.023795,4.1091285,4.3716927,4.516103,4.529231,4.6867695,4.824616,5.668103,6.229334,6.1341543,5.6320004,5.4875903,4.269949,3.5971284,4.0500517,5.142975,5.412103,5.6976414,6.4656415,7.213949,6.49518,6.4000006,7.0531287,7.243488,6.9677954,7.4174366,6.872616,6.5083084,6.3179493,6.2490263,6.1997952,6.0980515,6.048821,6.088206,6.0980515,5.792821,5.395693,5.0838976,5.1626673,5.398975,5.0182567,4.788513,4.7491283,4.844308,4.818052,4.2207184,5.2578464,5.9667697,5.661539,4.44718,3.2032824,2.8291285,5.0149746,6.944821,7.076103,5.149539,2.2350771,1.9856411,2.4352822,2.5895386,2.4549747,6.747898,6.0652313,5.0018463,4.821334,3.4592824,3.7054362,4.066462,5.5269747,7.2205133,6.432821,6.235898,6.8266673,7.4207187,7.6570263,7.5881033,7.131898,7.1220517,7.509334,7.9163084,7.604513,6.2030773,5.5138464,5.113436,4.824616,4.709744,5.159385,4.9920006,4.3585644,3.6660516,3.5872824,3.8728209,2.7864618,1.9200002,1.6147693,0.955077,0.9419488,0.92553854,1.0535386,1.273436,1.3522053,1.4112822,1.595077,1.7033848,1.719795,1.8149745,1.723077,1.6410258,1.723077,1.9035898,1.8871796,2.4024618,2.553436,2.6420515,2.7503593,2.7536411,2.8258464,2.678154,2.4418464,2.2055387,2.0184617,2.0841026,2.0873847,2.0906668,2.1497438,2.3105643,2.4155898,2.793026,3.2886157,3.692308,3.761231,4.3060517,4.519385,4.6966157,4.962462,5.2742567,5.169231,5.110154,5.034667,4.785231,4.1091285,4.086154,3.7021542,3.2295387,2.8225644,2.4910772,2.5042052,2.1989746,1.8707694,1.6147693,1.3292309,1.148718,0.88287187,0.7187693,0.6826667,0.65641034,0.8205129,0.7844103,0.7122052,0.72861546,0.90584624,0.93866676,0.8402052,0.7811283,0.8041026,0.8533334,0.7975385,0.77128214,0.6662565,0.50543594,0.4266667,0.61374366,0.7220513,0.955077,1.2635899,1.3489232,1.5688206,1.719795,1.8740515,2.0545642,2.2219489,2.1858463,2.3040001,2.4549747,2.5074873,2.3204105,2.425436,2.3958976,2.3269746,2.3630772,2.7306669,2.806154,2.8324106,3.0096412,3.245949,3.1967182,2.9702566,2.9440002,2.8914874,2.8127182,2.9440002,2.4582565,2.0742567,1.8182565,1.7526156,1.9922053,1.6278975,1.6902566,1.8838975,1.9200002,1.4933335,1.2865642,1.7329233,2.041436,1.9331284,1.6377437,1.9889232,1.9035898,1.9200002,2.0053334,1.5688206,1.5261539,1.5327181,1.5163078,1.3784616,0.9878975,5.9503593,6.1472826,6.2129235,6.091488,5.937231,6.1341543,5.7796926,5.0609236,4.493129,4.276513,4.2863593,4.667077,4.384821,4.2272825,4.453744,4.8049235,4.6605134,4.8049235,5.0576415,5.277539,5.3858466,5.080616,5.874872,6.619898,6.9645133,7.3550773,6.3901544,6.8004107,7.7390776,8.740103,9.705027,9.570462,9.317744,9.212719,9.393231,9.856001,9.760821,10.650257,11.414975,12.1468725,14.158771,15.330462,16.62359,17.362053,17.371899,16.981335,17.312822,17.430975,17.23077,16.846771,16.662975,16.59077,16.97477,17.28,17.161848,16.479181,14.549335,15.104001,14.884104,13.472821,13.289026,12.960821,12.373334,14.345847,18.353231,20.539078,19.39036,17.51959,15.035078,12.297847,9.91836,5.2676926,1.9987694,0.37415388,0.036102567,0.0,0.0,1.8412309,1.8642052,0.059076928,0.04594872,0.032820515,0.07548718,0.2231795,0.380718,0.32164106,0.41682056,1.0371283,1.5622566,1.6738462,1.3587693,0.32164106,0.052512825,0.03938462,0.02297436,0.0,0.35446155,0.3249231,0.34133336,0.56123084,0.8533334,0.88943595,0.46933338,0.23302566,0.24287182,0.0,0.013128206,0.006564103,0.0,0.0032820515,0.016410258,0.03938462,0.33805132,0.47261542,0.3052308,0.0,0.0,0.0,0.24287182,0.48902568,0.0,0.3052308,0.15097436,0.22646156,0.47589746,0.12143591,0.47589746,0.36430773,0.2297436,0.38400003,1.0075898,1.2996924,1.4572309,1.6278975,1.6902566,1.2504616,1.1651284,1.0436924,0.97805136,1.1618463,1.9068719,2.284308,2.793026,3.495385,4.138667,4.1517954,3.1015387,2.6190772,2.9669745,3.876103,4.5456414,5.0116925,5.2447186,5.0084105,4.7425647,5.586052,7.9786673,9.179898,9.186462,8.723693,9.26195,8.310155,8.346257,9.196308,10.361437,11.030975,10.496001,9.957745,9.416205,8.704,7.506052,6.8233852,7.0925136,7.788308,8.408616,8.467693,8.139488,8.165744,8.123077,8.100103,8.697436,9.941334,11.280411,11.579078,10.788103,9.93477,10.420513,10.525539,10.433641,10.456616,11.017847,12.2617445,12.3076935,11.414975,10.184206,9.537642,9.659078,9.852718,10.233437,10.709334,11.001437,11.575796,11.286975,10.896411,10.9456415,11.766154,12.898462,13.11836,13.033027,12.908309,12.665437,13.226667,13.768207,14.477129,15.409232,16.49559,15.067899,14.326155,13.853539,13.164309,11.687386,11.457642,12.150155,13.069129,13.748514,13.932309,13.380924,12.402873,12.268309,12.727796,12.009027,11.336206,10.811078,10.866873,11.362462,11.58236,11.703795,12.484924,12.763899,12.265027,11.58236,12.960821,13.305437,12.773745,11.628308,10.223591,10.771693,11.195078,11.024411,10.354873,9.842873,8.976411,7.788308,7.397744,7.5388722,6.560821,5.805949,5.3694363,5.2348723,5.228308,5.0215387,3.9811285,3.2754874,2.986667,2.8717952,2.3335385,2.3236926,2.0808206,1.7887181,1.6771283,2.044718,2.861949,3.4888208,4.201026,4.844308,4.8082056,6.173539,6.6625648,6.803693,6.675693,5.904411,4.7327185,3.6627696,2.422154,1.3554872,1.404718,1.9298463,6.196513,7.834257,6.0258465,5.5236926,4.010667,2.1858463,1.654154,2.2646155,2.1070771,2.422154,3.0982566,3.2000003,2.7208207,2.5632823,2.5009232,2.4976413,2.422154,2.4484105,3.0227695,2.9472823,3.2787695,4.010667,4.571898,3.8137438,3.373949,3.6036925,3.5544617,2.934154,2.1070771,1.9364104,2.0578463,2.044718,1.8543591,1.8313848,2.294154,2.868513,3.2787695,3.5446157,3.9975388,4.4373336,3.7776413,2.9243078,2.5042052,2.8849232,3.0916924,3.2886157,3.5938463,3.9811285,4.2863593,4.420923,4.3552823,4.348718,4.493129,4.699898,4.345436,4.384821,4.525949,4.4077954,3.6004105,3.9187696,3.4198978,2.9210258,3.006359,4.0434875,7.8047185,11.47077,13.8765135,14.631386,14.145642,9.993847,8.352821,12.839386,20.896822,23.78831,19.088411,14.326155,11.687386,11.533129,12.373334,13.22995,8.490667,4.466872,3.255795,2.7306669,4.2568207,5.0609236,4.900103,4.4865646,5.4613338,5.5236926,5.3202057,5.179077,5.2742567,5.61559,5.139693,4.7917953,4.325744,3.7907696,3.508513,3.1803079,2.9505644,3.1770258,3.7218463,3.9680004,4.2240005,4.4438977,4.699898,4.9821544,5.2020516,5.546667,5.674667,5.723898,5.7107697,5.540103,5.074052,4.9329233,4.9854364,4.97559,4.4865646,4.3027697,4.1485133,4.056616,4.0303593,4.0434875,4.1780515,3.8629746,3.3805132,2.993231,2.9440002,2.6518977,2.477949,2.2777438,1.9954873,1.6771283,1.3128207,1.1749744,1.1323078,0.9944616,0.51856416,0.4201026,0.37743592,0.36102566,0.36430773,0.4135385,0.43651286,0.48902568,0.5316923,0.60061544,0.80738467,0.6629744,0.5973334,0.6892308,0.8008206,0.58092314,0.48246157,0.6301539,0.88287187,1.083077,1.083077,1.2800001,1.5458462,1.7362052,1.8149745,1.8773335,1.6804104,1.6705642,1.6508719,1.6311796,1.8018463,1.5064616,1.3423591,1.3686155,1.5163078,1.6016412,1.9068719,2.294154,2.678154,3.058872,3.508513,3.3378465,3.498667,3.8038976,3.9811285,3.6758976,3.3969233,3.308308,3.2361028,3.1081028,2.9604106,3.387077,3.6857438,4.1124105,4.637539,4.9427695,4.84759,5.398975,6.124308,6.633026,6.6067696,7.1187696,5.937231,5.297231,5.5926156,5.3858466,5.7042055,5.8945646,6.4557953,7.1056414,6.774154,6.2490263,7.0531287,7.3025646,6.892308,7.4929237,7.394462,7.1876926,6.948103,6.5903597,5.858462,5.8847184,5.943795,6.0980515,6.2916927,6.377026,6.0980515,5.9536414,5.8880005,5.8486156,5.799385,5.687795,5.5597954,5.8092313,6.088206,5.293949,5.2578464,5.661539,5.6320004,5.0215387,4.4242053,4.2174363,6.4000006,7.1089234,5.930667,5.904411,3.1081028,4.1517954,3.8695388,1.8937438,2.6256413,4.027077,5.0838976,5.504,5.3169236,4.850872,4.850872,4.850872,5.8847184,6.9349747,4.9427695,6.7872825,9.206155,9.885539,8.933744,8.89436,9.347282,8.874667,8.576,8.848411,9.399796,7.4207187,6.550975,6.088206,5.5630774,4.7458467,4.598154,4.562052,4.420923,4.138667,3.8465643,3.7973337,2.7963078,1.8116925,1.3456411,1.4178462,1.4080001,1.0469744,0.892718,1.083077,1.3259488,1.4736412,1.913436,2.1398976,2.1825643,2.609231,1.9003079,1.8346668,2.1267693,2.3991797,2.166154,2.1530259,2.5993848,3.0391798,3.1803079,2.8980515,3.2164104,3.3772311,3.318154,3.0654361,2.7602053,2.553436,2.4484105,2.2219489,2.0184617,2.3335385,3.1048207,3.882667,4.2305646,4.273231,4.699898,4.650667,4.7589746,4.7392826,4.785231,5.5532312,5.175795,4.844308,4.854154,4.8049235,3.570872,3.8990772,4.3585644,4.204308,3.4560003,2.868513,2.6978464,2.425436,1.9987694,1.4998976,1.1585642,0.9288206,0.7318975,0.71548724,0.81394875,0.7778462,0.62030774,0.52512825,0.53825647,0.6498462,0.80738467,0.7220513,0.54482055,0.36430773,0.28225642,0.4266667,0.574359,0.51856416,0.4201026,0.37743592,0.4266667,0.6235898,0.6892308,0.7581539,0.92225647,1.2504616,1.5688206,1.8313848,2.100513,2.4057438,2.7470772,2.612513,2.5238976,2.353231,2.1956925,2.3794873,2.2219489,2.3204105,2.3991797,2.425436,2.609231,2.3893335,2.097231,1.9429746,2.0151796,2.2580514,2.930872,2.6683078,2.349949,2.3335385,2.4582565,2.2744617,1.7985642,1.6016412,1.9068719,2.5796926,1.9692309,1.9265642,1.9790771,1.847795,1.4178462,1.1257436,1.273436,1.595077,1.847795,1.785436,1.8346668,2.0742567,2.172718,2.0676925,1.9823592,1.6771283,1.4178462,1.2898463,1.1979488,0.8533334,6.806975,6.2194877,5.789539,5.536821,5.5762057,6.1341543,5.671385,5.1364107,4.663795,4.3585644,4.312616,4.535795,4.4406157,4.466872,4.7327185,5.037949,5.330052,5.609026,5.805949,5.8256416,5.546667,5.5532312,6.0356927,6.5411286,6.957949,7.525744,7.643898,7.821129,8.448001,9.29477,9.498257,9.527796,9.6984625,9.7214365,9.603283,9.636104,9.590155,10.029949,10.909539,12.09436,13.367796,14.979283,16.400412,17.67713,18.487797,18.166155,18.231796,18.008617,17.952822,17.99549,17.529438,16.850052,16.584206,16.275694,15.799796,15.379693,13.50236,13.289026,12.727796,11.631591,11.641437,12.49477,13.659899,16.052513,18.83241,19.416616,17.769028,17.686975,17.608206,16.390566,13.285745,5.930667,2.1398976,0.8795898,2.6157951,9.324308,6.8463597,3.2820516,0.8566154,0.15425642,0.13128206,1.0371283,0.5481026,0.16738462,0.6826667,2.162872,3.0424619,3.249231,2.5238976,1.3620514,1.017436,0.58420515,0.26256412,0.09189744,0.13784617,0.46276927,0.16410258,0.0951795,0.2100513,0.35446155,0.256,0.34133336,0.45292312,0.5284103,0.48902568,0.24287182,0.128,0.068923086,0.029538464,0.009846155,0.052512825,0.016410258,0.45620516,0.48246157,0.07876924,0.08533334,0.016410258,0.21333335,0.38400003,0.34133336,0.0,0.06235898,0.30194873,0.7056411,1.0338463,0.8172308,0.9189744,0.8598975,0.8960001,1.0502565,1.1158975,1.4408206,1.6016412,1.4506668,1.1060513,0.95835906,1.2931283,1.3915899,1.2964103,1.2668719,1.7985642,2.156308,3.045744,3.7710772,4.0008206,3.761231,3.0424619,2.9735386,3.4067695,4.0402055,4.388103,5.398975,6.0783596,6.3573337,6.7117953,8.15918,9.878975,10.745437,10.381129,9.248821,8.664616,8.316719,8.858257,9.442462,9.718155,9.82318,9.6,9.544206,9.3078985,8.772923,8.057437,7.529026,8.188719,8.94359,9.278359,9.26195,8.795898,8.612103,8.858257,9.255385,9.101129,9.114257,9.8363085,10.617436,11.08677,11.1294365,10.709334,9.987283,9.685334,10.171078,11.444513,11.733335,11.480617,10.998155,10.253129,8.864821,9.642668,9.554052,9.586872,10.06277,10.660104,11.008,11.047385,11.0375395,11.211488,11.776001,12.002462,12.12718,12.281437,12.632616,13.384206,13.410462,13.643488,13.974976,14.562463,15.82277,15.645539,14.851283,14.329437,14.273643,14.155488,13.334975,13.282462,13.735386,14.198155,13.932309,13.761642,12.724514,12.635899,13.318565,12.6063595,11.057232,10.348309,10.374565,10.801231,11.07036,12.274873,13.305437,13.4400015,12.760616,12.156719,13.056001,13.318565,12.435693,10.866873,10.039796,10.541949,10.650257,10.489437,10.026668,9.07159,7.719385,6.9645133,6.701949,6.7577443,6.9152827,6.294975,5.4843082,4.8804107,4.598154,4.457026,4.125539,3.5183592,2.9965131,2.609231,2.0906668,2.1169233,2.0611284,1.9265642,1.8051283,1.8970258,2.737231,3.1015387,3.8104618,4.7425647,4.844308,5.3202057,5.579488,5.5565133,5.3727183,5.356308,4.2240005,3.045744,2.1169233,1.4900514,0.96492314,1.1782565,3.9318976,7.066257,10.59118,16.692514,8.51036,3.1277952,1.1946667,1.9364104,3.1540515,3.0720003,3.5741541,3.6857438,3.170462,2.5009232,2.5600002,2.6387694,2.678154,2.917744,3.9122055,3.9745643,3.7743592,3.9417439,4.322462,3.9844105,3.2820516,3.3641028,3.2196925,2.546872,1.7755898,1.6246156,1.972513,2.4418464,2.740513,2.6486156,2.5665643,3.1343591,4.1682053,5.1954875,5.4514875,5.0215387,4.1156926,3.2065644,2.740513,3.1277952,3.5807183,3.7809234,3.748103,3.8498464,4.788513,5.467898,5.07077,4.6966157,4.594872,4.138667,3.9318976,3.7940516,3.9975388,4.2830772,3.8564105,3.882667,3.4592824,3.4198978,3.7185643,3.4100516,6.045539,8.897642,11.506873,13.348104,13.814155,12.652308,8.690872,6.8529234,8.710565,12.471796,8.280616,7.0498466,7.5881033,9.813334,14.76595,14.976001,12.42913,10.108719,8.730257,6.7117953,5.805949,5.8814363,5.5138464,4.7360005,5.0477953,5.3136415,5.395693,5.353026,5.3431797,5.6287184,5.5696416,5.546667,5.146257,4.516103,4.352,4.0500517,3.6036925,3.3017437,3.2032824,3.1245131,3.3509746,3.6890259,4.056616,4.4274874,4.8114877,4.9887185,4.9526157,4.962462,5.113436,5.3431797,5.2414365,5.2545643,5.113436,4.8049235,4.571898,4.0467696,3.6890259,3.4592824,3.4231799,3.7382567,3.8038976,3.4494362,3.1507695,3.0260515,2.858667,2.546872,2.353231,2.166154,1.9922053,1.9462565,1.6968206,1.4506668,1.2668719,1.0699488,0.65312827,0.48574364,0.4135385,0.36430773,0.33805132,0.38728207,0.37415388,0.4135385,0.44964105,0.512,0.74830776,0.7778462,0.72861546,0.761436,0.81066674,0.5907693,0.4266667,0.46933338,0.6662565,0.9419488,1.204513,1.4998976,1.5130258,1.3751796,1.2340513,1.2668719,1.1585642,1.1323078,1.1520001,1.1749744,1.142154,1.0535386,1.1749744,1.3489232,1.463795,1.4309745,1.5885129,2.0644104,2.5337439,2.9472823,3.5446157,3.5511796,3.6594875,3.9647183,4.204308,3.761231,3.501949,3.3312824,3.121231,2.8980515,2.8389745,3.1474874,3.249231,3.4264617,3.8137438,4.381539,4.7622566,5.0838976,5.6943593,6.4032826,6.498462,7.460103,6.961231,5.4941545,4.263385,5.179077,3.9548721,4.5390773,4.886975,4.8377438,6.12759,5.4843082,5.8420515,6.1472826,6.170257,6.514872,6.6527185,6.5706673,6.7117953,6.951385,6.5805135,6.311385,6.3212314,6.449231,6.5345645,6.416411,6.2129235,5.861744,5.681231,5.8420515,6.3606157,6.485334,6.8397956,7.3485136,7.5979495,6.8463597,6.7314878,6.665847,6.2752824,5.789539,6.0619493,5.910975,6.166975,6.012718,5.225026,4.1846156,3.623385,3.0194874,2.7208207,2.7995899,3.0654361,4.535795,5.87159,6.436103,6.242462,5.9634876,6.665847,6.7544622,6.1440005,5.2020516,4.7360005,6.921847,7.968821,7.1909747,5.504,5.428513,7.0531287,7.282872,7.0859494,7.1647186,7.958975,6.498462,6.3310776,6.370462,6.301539,6.5772314,6.0783596,5.044513,4.210872,3.889231,3.9680004,3.6069746,3.1113849,2.281026,1.4145643,1.3226668,1.6607181,1.4473847,1.2570257,1.4408206,2.1333334,2.1333334,2.2350771,2.284308,2.3040001,2.487795,2.0906668,2.1169233,2.2547693,2.2383592,1.847795,2.1989746,2.6617439,2.8947694,2.878359,2.9111798,3.2984617,3.4231799,3.5249233,3.6069746,3.4560003,2.6354873,2.3729234,2.6223593,3.0654361,3.1409233,3.6463592,4.2830772,4.9460516,5.412103,5.3694363,4.9329233,4.7294364,4.827898,5.1200004,5.3234878,5.421949,5.5532312,5.477744,5.110154,4.522667,3.9253337,3.6594875,3.4625645,3.308308,3.4067695,2.7076926,2.0709746,1.6968206,1.5163078,1.1848207,0.9517949,0.82379496,0.7844103,0.7844103,0.72861546,0.60061544,0.49887183,0.45620516,0.45620516,0.42994875,0.3446154,0.32164106,0.27569234,0.21989745,0.26912823,0.34789747,0.3117949,0.28225642,0.32164106,0.4397949,0.51856416,0.702359,0.90584624,1.086359,1.2406155,1.5458462,1.7033848,1.913436,2.2416413,2.612513,2.8291285,2.609231,2.359795,2.28759,2.3926156,2.487795,2.5764105,2.678154,2.733949,2.5862565,2.3269746,2.169436,2.1136413,2.1431797,2.2219489,2.228513,1.9462565,1.7952822,1.8379488,1.7723079,1.657436,1.463795,1.4375386,1.6278975,1.8576412,1.9528207,1.9003079,1.7165129,1.4309745,1.1027694,1.0535386,1.2537436,1.585231,1.8609232,1.8084104,1.8379488,2.1202054,2.422154,2.5895386,2.5337439,2.0217438,1.6672822,1.276718,0.9517949,1.0994873,6.4590774,6.052103,5.8518977,5.658257,5.5269747,5.786257,5.658257,5.3202057,4.8705645,4.568616,4.8311796,5.080616,5.074052,5.172513,5.4482055,5.691077,5.9536414,6.3310776,6.678975,6.9152827,7.0137444,6.189949,6.038975,6.2752824,6.7117953,7.256616,8.283898,8.2904625,8.385642,8.766359,8.713847,8.868103,9.140513,9.416205,9.540924,9.3078985,9.475283,9.888822,10.489437,11.221334,12.051693,13.896206,15.570052,16.853334,17.608206,17.795284,18.294155,17.913437,17.536001,17.339079,16.794258,16.577642,15.927796,15.133539,14.614976,14.903796,13.292309,12.596514,12.015591,11.569232,12.100924,12.924719,15.0088215,16.754873,18.15631,20.801643,19.587284,17.024002,16.416822,17.063385,14.240822,5.402257,1.8116925,0.892718,1.6836925,4.84759,6.163693,3.56759,1.214359,0.6235898,0.6662565,3.2131286,2.1267693,0.8533334,1.142154,3.05559,4.8377438,4.2863593,2.8553848,1.5524104,0.9124103,0.55794877,0.24943592,0.07876924,0.16738462,0.6629744,0.13128206,0.013128206,0.18707694,0.35446155,0.04266667,0.08205129,0.2297436,0.43651286,0.56451285,0.37743592,0.318359,0.24615386,0.18379489,0.12143591,0.02297436,0.0032820515,0.19364104,0.2855385,0.20676924,0.12471796,0.026256412,0.10502565,0.29210258,0.4397949,0.34789747,0.18051283,0.190359,0.34789747,0.5874872,0.80738467,0.6629744,0.6301539,0.90584624,1.276718,1.1520001,1.401436,1.2668719,1.0601027,0.9189744,0.8041026,1.1913847,1.3981539,1.5031796,1.6475899,2.044718,2.612513,3.3805132,4.1485133,4.670359,4.650667,4.017231,4.2863593,4.325744,4.066462,4.5029745,5.799385,6.3934364,7.273026,8.480822,9.133949,9.892103,10.30236,10.023385,9.216001,8.523488,8.283898,9.38995,10.28595,10.210463,9.193027,9.032206,9.18318,9.222565,8.726975,7.2861543,7.7456417,8.999385,10.036513,10.528821,10.850462,10.696206,10.052924,10.134975,10.555078,9.31118,8.746667,9.196308,9.829744,10.581334,12.160001,11.779283,10.594462,9.826463,10.164514,11.779283,12.232206,11.395283,10.807796,10.515693,9.07159,9.317744,8.881231,8.582564,8.845129,9.685334,10.571488,11.063796,11.273847,11.346052,11.451077,11.451077,11.382154,11.628308,12.412719,13.804309,13.804309,13.650052,14.001232,15.113848,16.846771,17.001026,16.659693,16.164104,15.803078,15.796514,15.035078,14.647796,14.706873,14.729847,13.682873,13.610668,13.59754,13.90277,14.188309,13.525334,11.45436,10.505847,10.328616,10.541949,10.722463,11.884309,13.082257,13.673027,13.505642,12.947693,13.5318985,13.505642,12.248616,10.381129,9.747693,10.243283,10.039796,9.869129,9.6984625,8.717129,7.076103,6.2227697,5.9536414,6.11118,6.5739493,5.8486156,5.0182567,4.453744,4.3290257,4.601436,4.5456414,3.9154875,3.1606157,2.5173335,2.0118976,1.9954873,1.9462565,1.9659488,2.0841026,2.2449234,2.7602053,2.9997952,3.5314875,4.2535386,4.394667,4.4964104,5.0051284,4.9099493,4.3716927,4.7228723,4.0992823,3.2918978,2.5074873,1.7657437,0.9189744,0.8992821,2.359795,5.1298466,9.353847,15.494565,7.9786673,3.0818465,1.1355898,1.5163078,2.6322052,3.383795,4.066462,4.1485133,3.5872824,2.8160002,2.6912823,2.5600002,2.6617439,3.1409233,4.0336413,3.948308,3.6857438,3.8564105,4.3684106,4.420923,3.4625645,3.3936412,3.1081028,2.359795,1.785436,1.654154,1.8412309,2.409026,3.0949745,3.2918978,2.4418464,2.8324106,3.945026,5.041231,5.146257,4.529231,3.826872,3.1967182,2.9144619,3.3641028,4.263385,4.519385,4.338872,4.263385,5.142975,5.4908724,5.028103,5.044513,6.5837955,10.450052,5.1987696,3.5872824,3.4560003,3.636513,3.9680004,4.3651285,4.4734364,5.0149746,5.664821,5.0182567,5.408821,7.1909747,8.858257,9.974154,11.152411,10.427077,7.0925136,4.5817437,4.4307694,6.265436,4.076308,4.57518,5.979898,8.704,15.366566,13.334975,12.406155,11.490462,10.71918,11.431385,7.194257,5.8978467,5.602462,5.349744,5.182359,5.5007186,5.5204105,5.431795,5.4383593,5.76,6.0356927,6.11118,5.832206,5.333334,5.028103,4.647385,4.1780515,3.6791797,3.259077,3.0687182,3.3280003,3.4494362,3.7251284,4.201026,4.6769233,4.821334,4.59159,4.453744,4.535795,4.644103,4.850872,5.169231,5.1298466,4.7458467,4.5095387,4.493129,3.8531284,3.2656412,3.058872,3.2229745,3.3312824,3.2886157,3.1442053,2.9801028,2.937436,2.5928206,2.28759,2.0873847,2.0020514,1.9954873,1.7690258,1.591795,1.404718,1.1552821,0.7975385,0.61374366,0.48246157,0.39056414,0.34789747,0.39056414,0.33805132,0.37415388,0.4660513,0.5973334,0.761436,0.827077,0.8402052,0.8336411,0.7844103,0.5940513,0.508718,0.5874872,0.76800007,0.9714873,1.1257436,1.1881026,1.273436,1.1881026,0.9616411,0.8402052,0.7384616,0.74830776,0.77456415,0.7811283,0.77456415,0.77456415,1.014154,1.1848207,1.211077,1.2603078,1.4572309,1.8609232,2.2744617,2.609231,2.9144619,3.1671798,3.4888208,3.7021542,3.7021542,3.4560003,3.3214362,3.1277952,2.9111798,2.733949,2.6978464,2.9702566,3.2853336,3.5478978,3.8038976,4.240411,4.844308,5.1167183,5.540103,6.157129,6.5805135,7.3747697,7.433847,5.970052,3.7907696,3.2951798,5.037949,5.024821,4.5029745,4.381539,5.2414365,5.3694363,5.796103,6.055385,6.0816417,6.2063594,6.747898,6.675693,6.885744,7.384616,7.3091288,7.194257,7.026872,7.0137444,7.062975,6.7807183,6.4000006,6.0258465,5.858462,5.989744,6.409847,6.5247183,7.253334,7.768616,7.765334,7.453539,7.1056414,7.003898,6.7938466,6.6822567,7.450257,7.4896417,7.210667,6.560821,5.4974365,3.9909747,3.2754874,2.4188719,2.3105643,3.131077,4.3552823,4.8705645,6.0980515,7.1483083,7.568411,7.3583593,7.174565,7.1122055,6.114462,4.6605134,4.7655387,5.7468724,5.904411,5.0838976,4.1911798,5.2020516,5.3694363,6.2818465,6.9021544,6.987488,7.0957956,5.9470773,5.723898,5.684513,5.671385,6.117744,5.943795,5.1364107,4.4734364,4.138667,3.7316926,3.5872824,3.2262566,2.487795,1.6213335,1.2964103,1.5130258,1.6180514,1.7165129,1.9265642,2.3893335,2.2219489,2.5206156,2.7634873,2.7733335,2.7142565,2.1825643,2.100513,2.1497438,2.1169233,1.9167181,2.7208207,3.006359,3.0424619,3.0785644,3.3280003,3.7284105,3.754667,3.623385,3.4198978,3.0916924,2.934154,3.1540515,3.4789746,3.751385,3.9089234,4.5456414,5.1659493,5.5565133,5.7074876,5.805949,5.671385,5.034667,4.857436,5.228308,5.356308,5.3202057,5.4974365,5.4843082,5.175795,4.768821,3.8662567,3.5183592,3.18359,2.8225644,2.9078977,2.2547693,1.7788719,1.467077,1.2406155,0.9353847,0.8041026,0.78769237,0.8041026,0.76800007,0.5874872,0.48246157,0.40369233,0.34789747,0.30851284,0.27241027,0.23630771,0.24287182,0.21989745,0.17394873,0.19364104,0.25271797,0.27897438,0.28882053,0.3249231,0.45292312,0.63343596,0.82379496,0.9714873,1.0994873,1.3259488,1.5360001,1.7394873,1.9889232,2.2711797,2.4976413,2.858667,2.7437952,2.550154,2.5140514,2.678154,2.793026,2.737231,2.7503593,2.8127182,2.6322052,2.3958976,2.3138463,2.3040001,2.28759,2.1858463,1.8576412,1.6705642,1.6278975,1.6377437,1.529436,1.4539489,1.394872,1.3357949,1.3554872,1.6311796,2.0118976,1.8116925,1.4736412,1.2340513,1.1060513,1.0732309,1.1815386,1.3751796,1.5688206,1.6508719,1.6607181,1.8248206,1.9462565,2.034872,2.3302567,2.2383592,1.8116925,1.2438976,0.8336411,0.97805136,6.0225644,5.6320004,5.677949,5.664821,5.5007186,5.5007186,5.6418467,5.687795,5.4383593,5.07077,5.1364107,5.1954875,5.356308,5.6254363,5.8880005,5.8978467,6.1768208,6.7971287,7.1909747,7.381334,8.008205,6.5739493,6.055385,6.048821,6.314667,6.75118,7.939283,8.096821,8.136206,8.333129,8.310155,8.418462,8.795898,9.245539,9.5146675,9.265231,9.537642,9.82318,10.098872,10.377847,10.7158985,12.347078,14.322873,15.780104,16.554668,17.214361,17.736206,17.332514,16.764719,16.449642,16.44636,16.15754,15.271386,14.500104,14.345847,15.100719,13.558155,12.773745,12.130463,11.608616,11.769437,12.048411,15.258258,16.646564,16.810667,21.681232,20.20431,15.573335,13.3251295,13.587693,11.096616,3.8662567,1.148718,0.5021539,0.4004103,0.22646156,2.8947694,2.294154,1.2012309,0.83035904,0.8172308,2.9210258,2.0676925,0.955077,0.94523084,2.0611284,3.4100516,2.789744,1.7690258,1.1126155,0.764718,0.64000005,0.28882053,0.052512825,0.10502565,0.44964105,0.098461546,0.059076928,0.18379489,0.25928208,0.0,0.0,0.049230773,0.19692309,0.3446154,0.256,0.256,0.21333335,0.19364104,0.16738462,0.0,0.0,0.0,0.15097436,0.36758977,0.31507695,0.06235898,0.08205129,0.2100513,0.3314872,0.36102566,0.30851284,0.16082053,0.12471796,0.29210258,0.6432821,0.6432821,0.60061544,0.67938465,0.8402052,0.84348726,1.0436924,0.9124103,0.90912825,1.0272821,0.80738467,1.1815386,1.3522053,1.6213335,1.9331284,1.8543591,2.5698464,3.2951798,4.269949,5.1659493,5.077334,4.322462,4.6769233,4.716308,4.2994876,4.585026,6.308103,7.072821,8.228104,9.639385,9.701744,9.924924,9.869129,9.258667,8.3593855,7.9819493,7.896616,9.012513,9.846154,9.708308,8.717129,8.500513,8.507077,8.470975,8.086975,7.0137444,7.899898,9.275078,10.722463,11.772718,11.890873,11.670976,10.837335,10.617436,10.758565,9.5606165,9.383386,9.691898,9.842873,10.295795,12.619488,13.696001,12.2847185,10.850462,10.561642,11.286975,11.776001,11.155693,10.824206,10.840616,9.921641,9.619693,8.746667,8.073847,8.057437,8.861539,10.164514,10.998155,11.47077,11.618463,11.408411,11.503591,11.053949,11.08677,11.943385,13.285745,13.938873,13.935591,14.372104,15.589745,17.161848,17.782156,17.962667,17.48677,16.722052,16.636719,15.990155,15.350155,15.100719,14.841437,13.397334,13.856822,14.736411,15.31077,15.123693,13.978257,11.730052,10.981745,10.791386,10.738873,10.9226675,11.772718,12.704822,13.443283,13.791181,13.620514,13.915898,13.331694,11.825232,10.072617,9.485129,9.508103,8.986258,8.868103,9.088,8.576,6.747898,5.7468724,5.35959,5.4449234,5.927385,5.225026,4.5817437,4.2994876,4.381539,4.522667,4.97559,4.342154,3.387077,2.5698464,2.028308,1.8642052,1.7985642,1.9265642,2.2219489,2.5435898,2.8488207,3.058872,3.4166157,3.882667,4.125539,4.197744,4.562052,4.3716927,3.8038976,4.0467696,3.8564105,3.5938463,3.058872,2.297436,1.6016412,1.4802053,1.7526156,3.4330258,6.3376417,9.097847,6.1538467,3.2065644,1.4605129,1.211077,1.8445129,2.9013336,3.8038976,4.1025643,3.764513,3.1573336,2.7273848,2.4516926,2.5993848,3.1606157,3.8695388,3.6726158,3.623385,3.9614363,4.562052,4.9296412,3.6857438,3.5413337,3.2951798,2.5796926,1.8412309,1.7526156,1.7788719,2.2580514,2.993231,3.249231,2.3794873,2.8521028,3.7349746,4.352,4.266667,3.8990772,3.5807183,3.3542566,3.3805132,3.9417439,5.0149746,5.3398976,5.3070774,5.3169236,5.802667,5.349744,4.6539493,4.6900516,6.6527185,11.959796,6.1046157,3.8859491,3.3345644,3.5282054,4.6080003,6.12759,6.1078978,6.0356927,6.488616,7.1089234,5.8880005,6.422975,7.1122055,7.3550773,7.5552826,6.449231,4.778667,3.6168208,3.511795,4.46359,4.197744,4.768821,5.2611284,6.7774363,12.419283,9.938052,9.035488,8.113232,7.3419495,8.65477,5.677949,4.453744,4.5423594,5.1200004,4.97559,5.3070774,5.6943593,5.7632823,5.5007186,5.2578464,5.474462,5.3858466,5.280821,5.287385,5.3727183,4.965744,4.453744,3.95159,3.5544617,3.314872,3.3936412,3.3050258,3.43959,3.882667,4.414359,4.7327185,4.522667,4.269949,4.1682053,4.125539,4.352,4.7458467,4.8016415,4.450462,4.069744,4.322462,3.8465643,3.242667,2.8324106,2.6551797,2.6847181,2.8225644,2.9046156,2.9472823,3.1409233,2.9210258,2.537026,2.1792822,1.9364104,1.7952822,1.6246156,1.5524104,1.404718,1.1388719,0.8336411,0.67938465,0.5218462,0.40697438,0.36430773,0.39712822,0.3249231,0.36758977,0.5218462,0.7187693,0.8402052,0.86646163,0.86317956,0.82379496,0.74830776,0.6268718,0.6498462,0.80738467,0.9911796,1.0929232,1.0043077,0.85005134,0.9189744,0.88615394,0.702359,0.571077,0.5546667,0.6104616,0.61374366,0.571077,0.6104616,0.62030774,0.78769237,0.892718,0.9189744,1.0699488,1.4867693,1.7362052,1.9495386,2.1792822,2.3827693,2.6912823,2.92759,2.9833848,2.8816411,2.7634873,2.930872,2.9636924,2.9078977,2.8225644,2.7963078,2.9669745,3.3936412,3.8137438,4.135385,4.4373336,4.962462,5.172513,5.5138464,6.0619493,6.547693,7.128616,7.50277,6.738052,4.8705645,2.8882053,4.4438977,3.889231,4.197744,5.431795,4.713026,5.3169236,5.87159,6.3540516,6.6002054,6.3245134,6.8496413,6.6395903,6.616616,7.0432825,7.499488,8.04759,7.8408213,7.5520005,7.4240007,7.276308,6.7872825,6.5312824,6.4295387,6.482052,6.7577443,7.1614366,7.9195905,8.123077,7.7423596,7.6110773,7.2303596,7.003898,7.0104623,7.2336416,7.571693,8.3364105,8.198565,7.466667,6.3277955,4.84759,3.1409233,2.0578463,2.3794873,3.6562054,4.2207184,5.2644105,5.8814363,6.242462,6.7971287,8.260923,7.2336416,6.8430777,5.927385,4.8147697,5.333334,4.827898,4.522667,3.9253337,3.4034874,4.201026,4.348718,5.3103595,6.2687182,6.665847,6.2096415,5.034667,4.6802053,4.785231,5.1298466,5.6254363,5.7468724,5.287385,4.8607183,4.4964104,3.6332312,3.5216413,2.9472823,2.409026,2.0217438,1.5360001,1.6082052,1.8116925,2.1366155,2.477949,2.6518977,2.4976413,2.8980515,3.170462,3.1015387,2.9636924,2.356513,2.1825643,2.231795,2.349949,2.4484105,3.4198978,3.4231799,3.370667,3.5774362,3.761231,4.1025643,4.1091285,3.817026,3.4297438,3.2984617,3.4297438,3.6463592,3.9745643,4.466872,5.179077,5.4875903,5.8814363,6.012718,5.933949,6.0849237,6.1472826,5.5565133,5.280821,5.5958977,6.088206,5.674667,5.4383593,5.5138464,5.5630774,4.7622566,3.826872,3.6004105,3.1573336,2.4648206,2.3827693,2.03159,1.6475899,1.4178462,1.2832822,0.94523084,0.74830776,0.73517954,0.78769237,0.7515898,0.41682056,0.39384618,0.3446154,0.27897438,0.2231795,0.2100513,0.27241027,0.24943592,0.18707694,0.13784617,0.15425642,0.21661541,0.3446154,0.38728207,0.35774362,0.4266667,0.69251287,0.92553854,1.0305642,1.0765129,1.3095386,1.3981539,1.7001027,2.0020514,2.2153847,2.3794873,2.7306669,2.7503593,2.7437952,2.8389745,2.989949,2.8914874,2.7503593,2.7076926,2.740513,2.6518977,2.612513,2.3762052,2.2219489,2.15959,1.9167181,1.5753847,1.5491283,1.6049232,1.5983591,1.4802053,1.3883078,1.3915899,1.2964103,1.2307693,1.6705642,2.1202054,1.785436,1.4408206,1.3522053,1.2504616,1.1618463,1.1454359,1.1979488,1.276718,1.3161026,1.4703591,1.5786668,1.5753847,1.5721027,1.847795,1.8937438,1.5819489,1.1257436,0.79097444,0.892718,5.8190775,5.2512827,5.2742567,5.395693,5.408821,5.408821,5.579488,5.9667697,5.979898,5.5236926,4.9821544,4.667077,5.0116925,5.481026,5.7403083,5.6418467,6.1440005,6.961231,7.1515903,6.948103,7.7423596,6.5706673,6.163693,6.0324106,6.0356927,6.38359,7.076103,7.460103,7.821129,8.172308,8.274052,8.41518,8.937026,9.386667,9.6065645,9.744411,9.91836,9.813334,9.7673855,9.829744,9.737847,10.745437,12.665437,14.411489,15.642258,16.764719,16.78113,16.36431,15.839181,15.691488,16.564514,15.8884115,15.228719,14.969437,15.169642,15.570052,14.211283,13.59754,12.73436,11.618463,11.254155,11.195078,14.87754,16.20677,15.724309,20.601437,17.78872,12.875488,9.265231,7.525744,5.356308,1.9462565,0.4594872,0.029538464,0.036102567,0.08533334,0.30851284,0.36758977,0.45620516,0.5546667,0.4266667,0.44964105,0.41682056,0.33476925,0.2231795,0.1148718,0.108307704,0.068923086,0.06235898,0.18051283,0.5218462,0.8992821,0.51856416,0.128,0.036102567,0.108307704,0.06235898,0.15753847,0.16082053,0.08205129,0.13784617,0.20348719,0.08861539,0.059076928,0.118153855,0.0,0.0,0.0,0.049230773,0.098461546,0.0,0.0,0.0,0.13784617,0.3708718,0.46276927,0.12143591,0.23630771,0.26256412,0.08533334,0.02297436,0.25928208,0.21333335,0.25271797,0.43323082,0.50543594,0.8172308,0.79425645,0.5284103,0.25928208,0.39384618,0.574359,0.7811283,1.083077,1.273436,0.90584624,1.3095386,1.3981539,1.6607181,1.9265642,1.3620514,1.9922053,3.0293336,4.1780515,4.9854364,4.827898,4.125539,4.5062566,4.9099493,4.9427695,4.84759,6.921847,8.214975,9.324308,10.220308,10.226872,10.505847,10.121847,8.920616,7.50277,7.207385,7.1844106,7.8145647,8.1755905,8.077128,8.054154,7.8670774,7.4436927,7.1154876,7.141744,7.7390776,8.12636,9.094564,10.791386,12.386462,12.07795,11.588924,10.994873,10.463181,10.174359,10.315488,10.624001,10.794667,10.509129,10.364718,11.897437,15.028514,14.01436,12.150155,10.971898,10.253129,10.528821,10.663385,10.820924,10.935796,10.712616,10.633847,9.570462,8.549745,8.198565,8.769642,9.980719,10.896411,11.490462,11.713642,11.477334,11.67754,11.004719,10.742155,11.277129,12.09436,13.6237955,14.280207,14.838155,15.599591,16.374155,17.624617,18.166155,17.716515,16.79754,16.754873,15.977027,15.212309,14.998976,15.002257,13.99795,14.907078,15.803078,16.183796,15.638975,13.856822,11.779283,11.477334,11.401847,11.145847,11.444513,12.0549755,12.471796,12.872206,13.338258,13.846975,14.050463,12.921437,11.32636,9.941334,9.26195,8.65477,7.9163084,7.8112826,8.274052,8.41518,6.7117953,5.7632823,5.2545643,5.080616,5.353026,4.955898,4.4964104,4.3552823,4.417641,4.066462,5.0904617,4.673641,3.6726158,2.674872,2.0020514,1.723077,1.6705642,1.8084104,2.100513,2.4910772,3.1770258,3.3017437,3.367385,3.6529233,4.197744,4.3684106,4.194462,3.889231,3.6135387,3.511795,3.4264617,3.6135387,3.4822567,2.9801028,2.5731285,2.2711797,2.0611284,2.8160002,4.1189747,4.2436924,4.9099493,3.436308,1.785436,1.0404103,1.3981539,1.9922053,2.8980515,3.4789746,3.5478978,3.3903592,2.7864618,2.5238976,2.6847181,3.1671798,3.69559,3.5183592,3.7907696,4.2929235,4.8344617,5.2545643,3.8695388,3.6627696,3.6135387,3.117949,1.9823592,1.7920002,1.7657437,2.0808206,2.550154,2.6322052,2.6584618,3.4658465,4.0467696,4.027077,3.6758976,3.623385,3.6168208,3.7842054,4.135385,4.5390773,5.435077,5.8453336,6.1374364,6.416411,6.5312824,5.346462,4.2502565,3.6430771,4.2371287,7.069539,5.661539,4.164923,3.511795,3.95159,5.0609236,7.824411,7.637334,6.820103,6.954667,8.868103,7.003898,6.301539,6.422975,6.426257,4.768821,3.3772311,2.858667,2.7437952,3.1507695,4.772103,5.756718,6.0291286,5.349744,5.152821,8.546462,7.975385,5.858462,3.9122055,2.6322052,1.3029745,2.5271797,2.4516926,2.8914874,3.9942567,4.2305646,4.4767184,5.5302567,6.0258465,5.533539,4.571898,4.381539,4.07959,4.1452312,4.667077,5.3366156,4.9132314,4.378257,4.0041027,3.82359,3.639795,3.4100516,3.2656412,3.2886157,3.5052311,3.879385,4.3585644,4.348718,4.1222568,3.9056413,3.895795,3.9614363,4.20759,4.2601027,3.9778464,3.4625645,3.436308,3.373949,3.1048207,2.6518977,2.2416413,2.034872,2.0644104,2.3696413,2.8422565,3.2262566,3.2886157,2.934154,2.3794873,1.8543591,1.5885129,1.4572309,1.3817437,1.2438976,1.024,0.8172308,0.69251287,0.5415385,0.43323082,0.39384618,0.41682056,0.3708718,0.4135385,0.56451285,0.764718,0.88287187,0.892718,0.827077,0.7811283,0.77128214,0.7089231,0.7975385,1.0010257,1.1815386,1.2077949,0.955077,0.7187693,0.6235898,0.56123084,0.5021539,0.5021539,0.636718,0.69579494,0.6301539,0.512,0.5415385,0.5874872,0.57764107,0.60389745,0.7122052,0.90256417,1.4441026,1.5031796,1.5163078,1.723077,2.15959,2.3794873,2.3729234,2.3762052,2.4024618,2.228513,2.5895386,2.9505644,3.1343591,3.1409233,3.1540515,3.1442053,3.4658465,3.9220517,4.3684106,4.706462,5.074052,5.1987696,5.5007186,5.9995904,6.308103,6.9021544,7.328821,7.509334,6.9842057,4.9099493,3.0654361,2.0939488,3.629949,6.0028725,4.2502565,4.781949,5.58277,6.5444107,7.200821,6.738052,6.770872,6.4032826,6.163693,6.432821,7.4371285,8.530052,8.369231,7.7981544,7.397744,7.50277,7.0859494,7.026872,6.994052,7.000616,7.4174366,8.3593855,8.933744,8.805744,8.251078,8.178872,7.397744,6.816821,6.951385,7.3386674,6.554257,7.8473854,8.169026,7.53559,6.4065647,5.6976414,3.7054362,2.2777438,3.1540515,4.900103,2.9111798,5.2480006,4.919795,4.0992823,4.768821,8.694155,7.2992826,6.7872825,6.11118,5.477744,6.36718,5.0215387,4.338872,3.5741541,2.665026,2.2416413,4.2863593,4.6802053,5.333334,6.308103,5.8289237,4.312616,3.8432825,4.2896414,5.2020516,5.802667,5.927385,5.4449234,5.034667,4.670359,3.6430771,3.31159,2.4320002,2.1530259,2.409026,1.9396925,1.9495386,2.0578463,2.4516926,2.9997952,3.2295387,3.1474874,3.314872,3.2984617,3.0752823,3.0293336,2.5961027,2.4713848,2.5961027,2.8882053,3.2623591,4.013949,3.8629746,3.8629746,4.1682053,4.013949,4.3060517,4.381539,4.2141542,4.0467696,4.4045134,4.2469745,4.089436,4.46359,5.428513,6.6067696,6.232616,6.294975,6.380308,6.3343596,6.2523084,6.1374364,5.976616,5.904411,6.1505647,7.026872,6.3606157,5.586052,5.6254363,6.0028725,4.84759,3.9056413,3.6036925,3.0884104,2.3630772,2.284308,2.0775387,1.6672822,1.5360001,1.585231,1.1552821,0.8041026,0.6892308,0.71548724,0.6892308,0.28882053,0.3708718,0.3511795,0.27897438,0.20020515,0.18051283,0.32164106,0.256,0.15097436,0.10502565,0.14112821,0.20020515,0.4266667,0.5284103,0.4660513,0.45620516,0.67282057,0.95835906,1.083077,1.0633847,1.1520001,1.1815386,1.5458462,1.8609232,2.0217438,2.1989746,2.4582565,2.6453335,2.8947694,3.1409233,3.117949,2.7536411,2.6880002,2.6945643,2.674872,2.6617439,2.8356924,2.3893335,2.0118976,1.8642052,1.5425643,1.3653334,1.5589745,1.6771283,1.5622566,1.3587693,1.270154,1.339077,1.3062565,1.2800001,1.7165129,2.1464617,1.8215386,1.591795,1.6147693,1.3522053,1.273436,1.1454359,1.0994873,1.1454359,1.148718,1.4408206,1.5753847,1.6049232,1.5622566,1.4473847,1.2274873,1.142154,0.99774367,0.8566154,1.0043077,5.4153852,5.5007186,5.35959,5.3037953,5.3825645,5.3727183,5.4449234,5.5007186,5.402257,5.093744,4.59159,4.1911798,4.4012313,4.7491283,5.1167183,5.7534366,6.5083084,6.892308,6.672411,6.2030773,6.422975,6.3277955,6.3573337,6.3310776,6.3343596,6.7150774,6.994052,6.954667,7.0957956,7.456821,7.6143594,8.467693,8.956718,9.242257,9.682052,10.817642,10.817642,10.243283,9.6065645,9.26195,9.383386,9.67877,10.410667,11.769437,13.676309,15.763694,15.602873,15.031796,14.385232,14.221129,15.320617,15.990155,16.745028,17.079796,16.692514,15.471591,15.461744,14.897232,13.774771,13.049437,14.647796,15.235283,15.983591,16.210052,16.292105,17.683693,13.338258,7.958975,4.2535386,2.7306669,1.6935385,0.7187693,0.21661541,0.026256412,0.0,0.0,0.0,0.009846155,0.009846155,0.0,0.0,0.013128206,0.006564103,0.036102567,0.07876924,0.029538464,0.04266667,0.108307704,0.13456412,0.15425642,0.3511795,1.0699488,0.92225647,0.45620516,0.14441027,0.3511795,0.18051283,0.18379489,0.14112821,0.16082053,0.6859488,1.017436,0.4397949,0.29210258,0.5874872,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08533334,0.17066668,0.0,0.14769232,0.37415388,0.45620516,0.3052308,0.0,0.0,0.0,0.19692309,0.43323082,0.21333335,0.15425642,0.33805132,0.636718,0.80738467,0.5021539,0.57764107,0.8960001,1.2931283,1.4572309,0.9321026,1.332513,1.5524104,1.6278975,1.6180514,1.6180514,1.8970258,3.570872,4.315898,4.1091285,5.218462,5.474462,6.363898,6.5870776,6.0947695,6.058667,7.53559,9.140513,10.299078,10.689642,10.240001,10.801231,10.400822,9.55077,8.539898,7.4141545,6.51159,6.9087186,7.276308,7.1515903,6.941539,7.125334,6.2555904,5.9930263,6.944821,8.667898,8.264206,8.887795,10.161232,11.516719,12.176412,12.360206,12.212514,11.339488,10.633847,12.268309,11.132719,11.132719,10.889847,10.029949,9.202872,12.839386,13.764924,12.527591,10.522257,10.010257,10.791386,10.630565,10.374565,10.331899,10.28595,11.602052,11.264001,10.154668,9.284924,9.796924,10.528821,11.204924,11.204924,10.709334,10.696206,10.722463,10.771693,10.761847,10.837335,11.398565,12.937847,14.10954,15.104001,15.862155,16.082052,17.158566,17.874052,17.56882,16.584206,16.265848,15.117129,14.795488,15.465027,16.633438,17.135592,16.646564,16.387283,15.898257,14.992412,13.748514,12.186257,11.684103,11.385437,11.126155,11.444513,11.713642,12.11077,12.212514,12.294565,13.321847,14.102976,13.052719,11.464206,10.056206,8.956718,8.700719,8.050873,7.640616,7.683283,7.965539,7.243488,6.5444107,6.1046157,5.8157954,5.218462,5.3398976,4.8049235,4.1682053,3.7973337,3.8465643,4.529231,4.781949,4.073026,2.6847181,1.7099489,1.6836925,1.6147693,1.6278975,1.7690258,2.0151796,4.1878977,3.895795,3.1277952,3.1015387,4.273231,4.381539,4.1813335,3.8400004,3.5380516,3.4625645,3.18359,3.4888208,3.7185643,3.4756925,2.609231,1.585231,2.8914874,3.5511796,3.8301542,7.24677,4.269949,2.5074873,1.3850257,0.81066674,1.1913847,1.8609232,2.349949,2.605949,2.8521028,3.5872824,3.255795,2.9801028,3.0982566,3.4888208,3.5872824,3.4264617,3.9909747,4.7228723,5.1954875,5.097026,4.069744,3.639795,3.639795,3.570872,2.5928206,1.7755898,1.654154,1.7624617,1.910154,2.166154,3.387077,4.325744,4.7524104,4.588308,3.9056413,3.748103,3.7349746,4.240411,4.8049235,4.135385,4.854154,5.3825645,5.865026,6.2752824,6.409847,5.225026,4.0041027,2.6256413,2.038154,4.273231,3.9318976,3.249231,3.3247182,3.8629746,3.2032824,5.986462,7.975385,9.731283,10.94236,10.407386,7.817847,6.1472826,5.8945646,6.2096415,4.8672824,3.4133337,2.3466668,1.9495386,2.3072822,3.2951798,5.2381544,7.27959,7.6635904,7.499488,10.758565,12.186257,9.347282,7.259898,6.550975,3.4625645,3.0358977,2.3433847,2.3729234,3.0949745,3.4494362,3.2656412,4.263385,5.2447186,5.609026,5.3398976,4.778667,4.6834874,4.824616,4.9952826,5.0215387,4.312616,4.07959,3.9384618,3.8498464,4.1058464,3.8367183,3.767795,3.7152824,3.5380516,3.1573336,3.2689233,3.3411283,3.3476925,3.3476925,3.495385,3.6660516,3.9089234,4.0008206,3.817026,3.3411283,2.9636924,2.6683078,2.5074873,2.425436,2.2416413,1.7920002,1.6049232,1.8609232,2.409026,2.7634873,3.0785644,2.8750772,2.4057438,1.9659488,1.8904617,1.5392822,1.2406155,1.0305642,0.93866676,0.97805136,0.7811283,0.6235898,0.51856416,0.47917953,0.5021539,0.5513847,0.54482055,0.571077,0.636718,0.6859488,0.8467693,0.8566154,0.90584624,0.97805136,0.8533334,0.9156924,1.0962052,1.2176411,1.1979488,1.0535386,0.74830776,0.63343596,0.6662565,0.74830776,0.74830776,0.9321026,0.88615394,0.65312827,0.40697438,0.44307697,0.73517954,0.6268718,0.55794877,0.6826667,0.8533334,0.86646163,0.7515898,0.82379496,1.2209232,1.8937438,2.2580514,2.6978464,3.058872,3.1803079,2.8980515,2.7536411,3.045744,3.3280003,3.4494362,3.570872,3.4231799,3.6791797,3.9122055,4.096,4.6080003,5.2315903,5.395693,5.4186673,5.549949,5.9667697,6.7971287,7.1056414,7.6898465,8.402052,8.132924,7.2172313,5.0576415,3.2065644,2.4320002,2.7011285,3.249231,5.0182567,6.3343596,6.8365135,7.4469748,6.9809237,6.738052,6.87918,7.4240007,8.254359,8.4512825,8.050873,7.453539,6.9809237,6.882462,6.5903597,6.7183595,6.7216415,6.747898,7.6143594,8.700719,9.393231,9.55077,9.570462,10.374565,7.3485136,6.426257,6.8496413,7.250052,5.677949,5.4449234,6.521436,5.6418467,3.5380516,4.9296412,4.8311796,4.0467696,5.3760004,7.1483083,3.2032824,3.6562054,2.4976413,2.8750772,5.668103,9.475283,7.4240007,7.719385,7.6012316,6.7807183,7.4141545,6.51159,4.8771286,3.3641028,2.5961027,2.9768207,5.720616,5.5663595,6.1407185,7.7948723,7.5979495,5.6320004,4.57518,4.6834874,5.4974365,5.8125134,5.802667,5.074052,4.6769233,4.4865646,3.2032824,2.9604106,2.176,1.9692309,2.3302567,2.1366155,1.8806155,2.1267693,2.6715899,3.373949,4.1813335,3.7776413,3.511795,3.1409233,2.7634873,2.8225644,2.7011285,2.8160002,3.0194874,3.3247182,3.9220517,4.263385,4.4406157,4.598154,4.6112823,4.073026,4.5128207,4.630975,4.841026,5.1954875,5.4153852,5.661539,6.124308,6.4656415,6.6560006,6.9743595,6.619898,6.7872825,6.8496413,6.6067696,6.301539,5.924103,5.7829747,5.910975,6.2720003,6.7610264,6.294975,5.602462,5.284103,5.362872,5.2644105,4.2141542,3.245949,2.5764105,2.3236926,2.5173335,1.7723079,1.6968206,1.6902566,1.4375386,0.8992821,0.75487185,0.6071795,0.5284103,0.47261542,0.28882053,0.3511795,0.39384618,0.33805132,0.21661541,0.16738462,0.23958977,0.15753847,0.072205134,0.06564103,0.15097436,0.21333335,0.4397949,0.65312827,0.761436,0.74830776,0.80738467,0.9517949,1.0436924,1.0404103,0.9911796,1.1520001,1.4375386,1.719795,1.8838975,1.847795,2.0676925,2.6157951,3.0785644,3.2032824,2.8980515,2.5829747,2.7503593,2.9078977,2.8816411,2.806154,2.7602053,2.553436,2.2416413,1.8871796,1.5556924,1.4473847,1.9495386,1.975795,1.3587693,0.86974365,0.9682052,1.1848207,1.3489232,1.4211283,1.4966155,1.847795,1.782154,1.6836925,1.595077,1.204513,1.3522053,1.0962052,0.9485129,1.1848207,1.8313848,1.7329233,1.8281027,1.7920002,1.5688206,1.3718976,1.1520001,1.0896411,1.0896411,1.1257436,1.2373334,4.8672824,4.8738465,4.9526157,5.1659493,5.4383593,5.5532312,5.293949,5.0543594,4.8607183,4.6900516,4.4832826,4.0500517,3.9745643,4.2272825,4.6211286,4.824616,6.058667,6.994052,7.3091288,7.204103,7.3649235,7.1680007,6.8955903,6.3901544,5.8912826,6.055385,6.560821,6.892308,7.3649235,7.9228725,8.139488,9.383386,10.072617,10.423796,10.604308,10.732308,10.000411,9.124104,8.444718,8.077128,7.896616,8.549745,9.238976,10.400822,11.864616,12.868924,13.5318985,13.751796,13.974976,14.34913,14.7331295,16.459488,16.840206,16.410257,15.780104,15.642258,15.104001,14.519796,14.299898,14.677335,15.711181,14.148924,13.906053,14.549335,15.287796,14.998976,10.916103,6.409847,3.1934361,1.723077,1.1946667,0.636718,0.2855385,0.101743594,0.029538464,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0032820515,0.0,0.006564103,0.01969231,0.029538464,0.052512825,0.08533334,0.098461546,0.128,0.26584616,0.60389745,0.6662565,0.69251287,0.90584624,1.522872,0.8533334,0.33805132,0.06564103,0.032820515,0.13784617,0.20348719,0.08861539,0.3511795,0.702359,0.0,0.4201026,0.2100513,0.23302566,0.5152821,0.23302566,0.04594872,0.108307704,0.23958977,0.25928208,0.0,0.4004103,0.3052308,0.13456412,0.06235898,0.0,0.26256412,0.16738462,0.14441027,0.24943592,0.16410258,0.15097436,0.30851284,0.40697438,0.43651286,0.5874872,0.8566154,0.955077,0.9485129,0.95835906,1.1749744,1.1585642,1.1126155,1.2274873,1.4309745,1.3620514,2.6978464,3.8498464,4.4898467,4.97559,6.340924,5.681231,5.8486156,6.2851286,6.741334,7.2894363,9.110975,9.803488,10.04636,10.200616,10.33518,11.0145645,10.745437,9.980719,8.973129,7.781744,6.8988724,7.430565,7.6110773,7.017026,6.564103,6.0356927,5.5204105,5.799385,6.9349747,8.277334,8.52677,8.822155,9.636104,10.512411,10.089026,9.970873,11.096616,12.2617445,12.891898,13.026463,11.96636,12.389745,12.580104,11.67754,9.6754875,10.230155,11.667693,12.009027,10.9686165,9.947898,10.085744,10.33518,10.272821,9.737847,8.818872,9.494975,9.69518,9.45559,9.216001,9.856001,10.9226675,11.542975,11.464206,10.827488,10.171078,10.35159,10.617436,10.880001,11.053949,11.07036,12.547283,13.764924,14.880821,15.77354,16.032822,16.580925,17.201233,17.024002,16.065641,15.241847,14.004514,14.480412,15.675078,17.030565,18.428719,15.471591,15.07118,15.16636,14.746258,13.833847,12.35036,11.355898,10.866873,10.81436,11.053949,11.392001,11.424822,11.336206,11.395283,11.940104,12.908309,12.826258,11.651283,9.905231,8.700719,8.815591,8.792616,8.438154,7.9195905,7.781744,7.529026,6.9743595,6.7610264,6.7314878,5.937231,6.1472826,5.0051284,4.056616,3.9318976,4.322462,4.44718,4.4373336,3.7185643,2.4910772,1.7099489,1.595077,1.5688206,1.6705642,1.8051283,1.7591796,3.570872,3.446154,2.9801028,3.1376412,4.2601027,4.4964104,4.926359,4.6802053,3.8071797,3.3050258,3.0818465,3.3805132,3.6168208,3.5478978,3.2689233,3.7284105,3.9286156,3.2098465,2.6420515,5.0149746,2.8553848,2.048,1.3161026,0.62030774,1.1520001,1.5622566,1.8379488,2.0676925,2.3171284,2.609231,2.8258464,3.0260515,3.0523078,2.9243078,2.8160002,3.0982566,3.9548721,4.70318,4.9460516,4.594872,3.764513,3.2295387,3.1803079,3.367385,3.0949745,2.412308,2.1431797,2.2514873,2.7733335,3.7907696,4.325744,4.529231,4.562052,4.44718,4.066462,4.1878977,4.33559,4.709744,5.0543594,4.634257,5.2480006,5.7501545,6.196513,6.2851286,5.333334,9.668923,11.175385,10.601027,8.4283085,4.8836927,3.7021542,3.2196925,4.2305646,5.7009234,4.778667,5.901129,6.2129235,6.770872,7.6307697,7.8539495,7.2303596,6.377026,5.924103,5.8223596,5.3694363,4.529231,3.4560003,3.058872,3.5413337,4.394667,8.004924,9.4916935,10.249847,11.349334,13.515489,15.120412,13.643488,11.516719,10.118565,9.77395,6.76759,4.5390773,3.9089234,4.7261543,5.8420515,5.356308,3.8596926,3.0818465,3.2689233,3.2164104,3.767795,4.5390773,4.824616,4.6112823,4.5554876,4.522667,4.33559,4.1682053,4.069744,3.945026,3.7152824,3.4100516,3.2098465,3.1409233,3.0851285,3.1081028,3.3280003,3.5446157,3.639795,3.5905645,3.3542566,3.3772311,3.508513,3.5380516,3.2065644,2.7995899,2.4451284,2.2022567,2.0709746,1.9856411,1.8281027,1.6935385,1.6475899,1.7493335,2.0545642,2.537026,2.5206156,2.2613335,1.9692309,1.8051283,1.5688206,1.3522053,1.2012309,1.0929232,0.9156924,0.86646163,0.7581539,0.6465641,0.54482055,0.44307697,0.56123084,0.58420515,0.58420515,0.5973334,0.636718,0.827077,0.9682052,0.94523084,0.8041026,0.7811283,0.8992821,1.0962052,1.214359,1.1881026,1.0535386,0.8172308,0.7187693,0.82379496,1.0633847,1.2471796,1.1979488,1.1060513,0.8566154,0.5973334,0.77128214,0.7122052,0.6465641,0.64000005,0.69251287,0.7581539,0.96492314,0.9911796,1.0568206,1.2603078,1.5983591,2.2383592,3.0752823,3.4560003,3.3280003,3.2525132,3.1540515,3.1606157,3.1245131,3.058872,3.1442053,3.3280003,3.623385,3.826872,3.9614363,4.279795,4.647385,4.8377438,5.0182567,5.156103,5.0149746,5.658257,6.4557953,7.0400004,7.250052,7.1089234,6.633026,5.9503593,4.519385,2.7634873,2.0676925,2.0775387,3.95159,4.969026,5.024821,6.6395903,6.87918,6.8562055,7.0137444,7.637334,8.828718,8.546462,7.958975,7.529026,7.328821,7.066257,7.7390776,7.755488,7.5913854,7.571693,7.8834877,8.579283,9.078155,9.051898,8.14277,5.970052,4.601436,3.9778464,4.2929235,4.8082056,3.8695388,2.3696413,4.8771286,7.256616,6.885744,2.681436,4.420923,3.882667,3.626667,4.201026,4.1452312,4.5554876,2.3171284,1.5983591,4.023795,8.681026,7.830975,7.6570263,7.4141545,7.0925136,7.4141545,7.2237954,7.4010262,5.2512827,2.162872,3.5872824,6.038975,7.282872,8.320001,9.045334,8.2445135,6.698667,5.8190775,6.160411,7.141744,7.059693,6.813539,5.720616,4.466872,3.4560003,2.789744,2.4385643,1.9626669,1.8838975,2.2449234,2.6354873,2.1858463,2.0906668,2.3302567,2.8225644,3.4231799,3.4330258,3.7284105,3.7710772,3.370667,2.6880002,2.9078977,3.3017437,3.7415388,4.1156926,4.325744,4.2863593,4.4701543,4.709744,4.9362054,5.159385,5.3070774,5.169231,5.32677,5.835488,6.2227697,6.416411,6.49518,6.774154,7.145026,7.0826674,6.7577443,6.75118,6.6067696,6.2687182,6.0685134,5.917539,5.986462,6.2063594,6.3442054,6.0028725,6.0947695,6.038975,5.6976414,5.172513,4.8114877,3.9975388,3.255795,2.5107694,1.9692309,2.1136413,1.6049232,1.3292309,1.1913847,1.1257436,1.0962052,1.3587693,1.0436924,0.63343596,0.36102566,0.21661541,0.2100513,0.27897438,0.33476925,0.3446154,0.31507695,0.24943592,0.17066668,0.128,0.15753847,0.26256412,0.4594872,0.7187693,0.9419488,1.0699488,1.0765129,0.9911796,0.9156924,0.9616411,1.079795,1.0404103,1.2373334,1.3751796,1.5031796,1.6278975,1.6869745,2.0939488,2.5698464,2.8389745,2.8521028,2.802872,2.7175386,2.8947694,2.7700515,2.3171284,2.038154,2.1070771,2.0578463,1.9790771,1.8576412,1.5556924,1.6705642,1.8806155,1.8051283,1.3883078,0.88287187,0.9616411,1.1060513,1.2668719,1.401436,1.4966155,1.7132308,1.7657437,1.654154,1.4178462,1.1454359,1.3883078,1.2964103,1.2996924,1.5097437,1.7099489,1.7099489,1.8149745,1.7033848,1.401436,1.2635899,1.0633847,0.8730257,0.77456415,0.7844103,0.8467693,4.6211286,4.571898,4.6244106,4.8377438,5.1167183,5.2348723,5.0674877,4.716308,4.4340515,4.266667,4.0434875,3.895795,3.82359,4.1091285,4.6834874,5.1331286,5.917539,6.6034875,6.997334,7.213949,7.680001,7.79159,7.250052,6.685539,6.409847,6.439385,6.6067696,7.1122055,7.824411,8.454565,8.562873,9.649232,10.121847,10.292514,10.361437,10.400822,9.668923,9.101129,8.569437,8.1755905,8.254359,8.605539,9.058462,10.059488,11.346052,11.963078,12.347078,12.950975,13.771488,14.506668,14.569027,15.182771,14.7331295,14.27036,14.214565,14.375385,13.528616,13.479385,13.942155,14.631386,15.251694,14.12595,14.50995,14.660924,13.932309,12.763899,11.155693,7.456821,4.3618464,2.8160002,2.0118976,0.94523084,0.37743592,0.12143591,0.03938462,0.04594872,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.02297436,0.032820515,0.036102567,0.072205134,0.20676924,0.3708718,0.44964105,0.48574364,0.63343596,1.148718,0.88943595,0.36430773,0.036102567,0.0,0.0,0.0,0.0,0.14769232,0.29210258,0.0,0.2100513,0.10502565,0.21989745,0.54482055,0.5284103,0.10502565,0.23630771,0.33476925,0.24287182,0.21989745,0.53825647,0.36102566,0.20676924,0.19692309,0.072205134,0.20348719,0.17394873,0.15425642,0.19364104,0.22646156,0.42338464,0.52512825,0.52512825,0.49230772,0.5907693,0.8566154,0.73517954,0.78769237,1.1881026,1.6836925,1.3292309,1.2504616,1.3751796,1.8412309,2.9997952,3.367385,3.8859491,4.893539,6.180103,6.9710774,6.6133337,6.7282057,7.3058467,7.9917955,8.103385,9.449026,9.69518,10.115283,10.706052,10.197334,10.663385,10.502565,9.95118,9.153642,8.201847,7.5881033,7.4371285,7.1483083,6.678975,6.5247183,5.435077,5.2348723,6.042257,7.3682055,8.113232,8.858257,8.67118,8.697436,9.019077,8.651488,9.291488,10.761847,12.412719,13.604104,13.718975,12.35036,12.471796,12.599796,11.972924,10.555078,9.852718,10.738873,11.687386,11.618463,9.878975,10.000411,10.650257,10.610872,9.573745,8.15918,7.9261546,8.224821,8.474257,8.648206,9.304616,10.240001,10.689642,10.866873,10.824206,10.453334,10.834052,11.093334,11.638155,12.117334,11.45436,12.425847,13.558155,14.49354,14.989129,14.913642,15.665232,16.951796,17.109335,16.022976,15.120412,14.427898,15.126975,16.150976,16.416822,14.815181,12.045129,12.875488,14.267078,14.651078,13.938873,12.566976,11.634872,11.067078,10.807796,10.801231,10.971898,10.811078,10.706052,10.870154,11.339488,12.1698475,12.396309,11.795693,10.57477,9.386667,9.127385,9.147078,9.032206,8.585847,7.827693,7.716103,7.3058467,7.1844106,7.3091288,7.017026,6.7216415,5.356308,4.2568207,4.069744,4.788513,5.031385,4.381539,3.259077,2.156308,1.6344616,1.4998976,1.4802053,1.6246156,1.8313848,1.847795,3.1081028,3.259077,3.2328207,3.5380516,4.240411,4.5817437,4.9788723,4.670359,3.764513,3.255795,2.9243078,3.3444104,3.239385,2.6157951,2.737231,4.4406157,4.5095387,3.8400004,3.0293336,2.3860514,1.9856411,1.9035898,1.5327181,0.95835906,0.9517949,1.3161026,1.4998976,1.7493335,2.0775387,2.284308,2.5796926,2.8488207,2.7798977,2.4681027,2.4057438,2.8849232,3.7743592,4.5095387,4.7294364,4.3060517,3.6726158,3.1409233,3.1015387,3.4494362,3.5872824,2.9965131,3.045744,3.31159,3.692308,4.388103,4.7556925,5.0642056,4.9887185,4.57518,4.240411,4.276513,4.4865646,4.9132314,5.284103,5.0182567,5.654975,6.173539,6.4065647,6.055385,4.6802053,7.2172313,12.826258,16.850052,17.174976,14.263796,6.5083084,4.568616,4.778667,5.146257,5.366154,5.5663595,5.3891287,5.7435904,7.0498466,9.232411,7.7423596,6.7282057,6.232616,6.3474874,7.213949,7.4174366,6.521436,5.717334,5.677949,6.5903597,9.931488,10.985026,10.607591,10.827488,14.838155,16.01641,13.584412,11.605334,11.414975,11.618463,8.533334,5.6287184,5.106872,6.554257,6.961231,7.174565,5.805949,4.5128207,3.4888208,1.467077,1.7723079,2.8488207,3.442872,3.3575387,3.4527183,3.4166157,3.2984617,3.2328207,3.1934361,2.9801028,2.806154,2.605949,2.425436,2.3302567,2.3991797,2.6190772,2.9833848,3.1934361,3.1671798,3.0391798,2.8947694,2.9801028,3.1540515,3.245949,3.0654361,2.612513,2.3335385,2.2055387,2.1202054,1.8773335,1.8281027,1.8576412,1.7723079,1.6246156,1.719795,2.034872,2.2514873,2.2711797,2.100513,1.8674873,1.4539489,1.2668719,1.2307693,1.2373334,1.1388719,1.1191796,0.955077,0.7778462,0.63343596,0.49230772,0.54482055,0.6071795,0.6268718,0.636718,0.75487185,0.9124103,1.1290257,1.1158975,0.90912825,0.8730257,1.0502565,1.1355898,1.2537436,1.3489232,1.1716924,1.024,0.8795898,0.9419488,1.1782565,1.3357949,1.3062565,1.2471796,1.0469744,0.8172308,0.8992821,0.8336411,0.7778462,0.8041026,0.8992821,0.9419488,0.9878975,0.98133343,1.079795,1.270154,1.3883078,1.6804104,2.550154,3.18359,3.308308,3.1967182,3.1967182,3.4231799,3.5840003,3.5938463,3.5478978,3.692308,3.7710772,3.8006158,3.8432825,3.9942567,4.2338467,4.2371287,4.2994876,4.4734364,4.565334,5.113436,5.937231,6.4689236,6.629744,6.806975,6.665847,6.5280004,5.618872,3.895795,2.0250258,2.3958976,3.9778464,5.0149746,5.4580517,6.987488,6.957949,7.056411,7.0793853,7.177847,7.8736415,7.9097443,7.50277,7.2369237,7.276308,7.3583593,8.103385,8.109949,8.054154,8.086975,7.8112826,8.060719,8.323282,8.1066675,6.87918,4.07959,4.5554876,3.5446157,2.9571285,3.1474874,2.9243078,2.6354873,5.1954875,8.100103,8.349539,2.4320002,4.096,3.56759,3.7349746,4.5029745,2.7963078,5.182359,4.082872,3.1540515,4.315898,7.7423596,7.837539,7.755488,7.5618467,7.5454364,8.2215395,7.453539,8.185436,6.242462,2.8324106,4.5522056,7.1089234,8.569437,9.196308,9.284924,9.16677,7.830975,6.629744,6.189949,6.7085133,7.9458466,7.062975,5.8945646,4.5489235,3.2525132,2.3368206,2.172718,1.9922053,1.9298463,2.1202054,2.7175386,2.1858463,1.8674873,2.0053334,2.5435898,3.114667,3.0949745,3.5774362,3.9023592,3.7743592,3.259077,3.4264617,3.5446157,3.9089234,4.5029745,5.0018463,4.926359,4.9952826,4.9985647,5.034667,5.5236926,5.536821,5.756718,6.0750775,6.377026,6.5345645,6.7183595,6.951385,7.4010262,7.75877,7.256616,6.8955903,6.678975,6.3540516,5.930667,5.664821,6.114462,6.340924,6.4295387,6.363898,6.0324106,6.38359,6.235898,5.9569235,5.6352825,5.0838976,4.0500517,3.5544617,2.8192823,1.9068719,1.7033848,1.5819489,1.2832822,1.1520001,1.1913847,1.0994873,1.1290257,0.8402052,0.55794877,0.38728207,0.20676924,0.21333335,0.25271797,0.30194873,0.33476925,0.3249231,0.23302566,0.16082053,0.118153855,0.13128206,0.22646156,0.63343596,0.9353847,1.017436,0.9747693,1.0962052,1.1782565,1.017436,1.0272821,1.211077,1.1454359,1.3161026,1.4572309,1.5360001,1.5622566,1.6114873,1.8576412,2.4976413,2.8980515,2.8914874,2.7864618,2.7602053,2.8356924,2.612513,2.1398976,1.8904617,2.0250258,2.172718,2.1530259,1.9035898,1.4572309,1.6410258,1.7460514,1.6311796,1.3456411,1.142154,0.98133343,1.083077,1.3554872,1.654154,1.7887181,1.7427694,1.6607181,1.4211283,1.0962052,0.94523084,1.2504616,1.2898463,1.2800001,1.3522053,1.5688206,1.7033848,1.6771283,1.4572309,1.1355898,0.92553854,0.8763078,0.76800007,0.65969235,0.6268718,0.74830776,4.338872,4.384821,4.33559,4.4077954,4.6211286,4.8114877,4.6178465,4.2863593,4.059898,3.9811285,3.892513,4.023795,3.9286156,4.1780515,4.824616,5.395693,5.720616,5.907693,6.2030773,6.7774363,7.7292314,8.234667,7.778462,7.269744,7.030154,6.8004107,6.695385,7.197539,7.9524107,8.582564,8.677744,9.4916935,9.744411,9.849437,9.980719,10.082462,9.813334,9.69518,9.334154,8.864821,8.920616,9.009232,9.409642,10.148104,11.034257,11.634872,11.631591,12.153437,13.046155,13.824001,13.689437,13.574565,13.272616,13.105232,13.154463,13.252924,13.459693,14.490257,15.540514,16.154257,16.216616,15.468308,15.415796,14.884104,14.198155,15.195899,12.507898,7.8145647,4.210872,2.6354873,1.8904617,0.8795898,0.33476925,0.098461546,0.03938462,0.04594872,0.009846155,0.0,0.0,0.0032820515,0.01969231,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.029538464,0.1148718,0.20020515,0.24615386,0.22646156,0.2297436,0.45620516,0.512,0.23958977,0.029538464,0.013128206,0.072205134,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.108307704,0.30194873,0.4135385,0.09189744,0.256,0.33805132,0.2231795,0.23958977,0.65641034,0.45292312,0.256,0.23302566,0.10502565,0.14441027,0.256,0.42994875,0.58420515,0.5677949,1.1946667,1.014154,0.7417436,0.67282057,0.6662565,0.77128214,0.62030774,0.7844103,1.2964103,1.654154,1.5064616,1.6902566,1.9331284,2.3630772,3.511795,3.2623591,3.9318976,5.5204105,7.2927184,7.77518,7.9163084,7.9917955,8.352821,8.815591,8.6580515,9.547488,9.504821,9.757539,10.338462,10.098872,10.036513,9.82318,9.577026,9.209436,8.421744,7.8014364,7.27959,7.02359,6.9842057,6.885744,5.6943593,5.474462,6.2555904,7.5487185,8.3593855,8.835282,8.4053335,7.8769236,7.6242056,7.5585647,8.930462,10.857026,12.800001,14.070155,13.827283,11.776001,11.447796,11.910565,12.3306675,11.979488,10.633847,10.377847,11.122872,11.802258,10.384411,10.791386,11.434668,11.250873,10.033232,8.421744,7.4075904,7.4141545,7.827693,8.346257,8.969847,9.40636,9.757539,10.197334,10.725744,11.16554,11.625027,11.930258,12.35036,12.704822,12.3306675,12.875488,13.568001,14.158771,14.39836,14.034052,14.913642,16.433231,16.955078,16.226463,15.38954,14.985847,15.638975,16.219898,15.491283,12.117334,9.787078,11.37559,13.6008215,14.667488,14.260514,12.931283,11.989334,11.313231,10.86359,10.696206,10.755282,10.377847,10.223591,10.463181,10.771693,11.428103,11.723488,11.71036,11.303386,10.289231,9.268514,9.15036,9.350565,9.193027,7.9130263,7.7390776,7.5913854,7.5979495,7.6931286,7.6274877,7.2369237,6.0356927,4.821334,4.269949,4.9362054,5.1987696,4.325744,3.0654361,2.0118976,1.591795,1.3751796,1.3718976,1.6213335,2.0086155,2.2711797,3.0720003,3.4789746,3.8564105,4.20759,4.1714873,4.604718,4.8771286,4.578462,3.8038976,3.1474874,2.4582565,2.8816411,2.6912823,1.8248206,1.9068719,3.5938463,4.1878977,4.1550775,3.4067695,1.2996924,1.5392822,1.6049232,1.7033848,1.654154,0.8960001,1.1618463,1.3292309,1.7033848,2.166154,2.1858463,2.284308,2.425436,2.3991797,2.2482052,2.2514873,2.7273848,3.501949,4.2338467,4.5817437,4.2338467,3.7448208,3.4166157,3.5446157,4.0303593,4.3716927,3.9122055,4.0992823,4.2141542,4.1517954,4.4307694,4.781949,5.5729237,5.5565133,4.785231,4.601436,4.5029745,4.699898,4.9985647,5.1987696,5.10359,6.173539,6.452513,6.183385,5.356308,3.698872,3.4658465,11.050668,18.57313,22.183386,22.088207,10.131693,6.87918,5.720616,4.5029745,5.5302567,5.277539,4.7556925,5.4908724,7.7981544,10.801231,8.999385,7.6209235,6.695385,6.3540516,6.8365135,7.571693,8.746667,8.402052,6.672411,5.799385,7.965539,9.42277,9.38995,9.632821,14.441027,16.600616,12.937847,10.551796,11.168821,11.136001,10.292514,7.8014364,6.961231,7.75877,6.8988724,7.817847,6.944821,5.684513,4.394667,2.3762052,1.6213335,1.8346668,2.041436,2.041436,2.4155898,2.3204105,2.162872,2.2678976,2.553436,2.5304618,2.2744617,2.1464617,1.9593848,1.7296412,1.6738462,1.9298463,2.3335385,2.5304618,2.4484105,2.28759,2.300718,2.4320002,2.5928206,2.6978464,2.6617439,2.3893335,2.2547693,2.2383592,2.2186668,1.9692309,1.8838975,1.8642052,1.7887181,1.6705642,1.6475899,1.9068719,2.2153847,2.3991797,2.412308,2.3204105,1.7066668,1.332513,1.1946667,1.214359,1.2373334,1.2800001,1.1158975,0.9189744,0.75487185,0.5940513,0.60061544,0.6301539,0.6235898,0.6498462,0.8992821,1.0338463,1.2340513,1.2274873,1.0305642,0.94523084,1.1454359,1.2996924,1.522872,1.6968206,1.4834872,1.3522053,1.2603078,1.3062565,1.4276924,1.4112822,1.4309745,1.3653334,1.1913847,1.0108719,1.0338463,1.0994873,1.0633847,1.0469744,1.0896411,1.1126155,1.1323078,1.0699488,1.086359,1.214359,1.3653334,1.4834872,2.0053334,2.6026669,3.0030773,2.993231,2.9636924,3.43959,3.9351797,4.1452312,3.9581542,4.076308,4.069744,3.9122055,3.69559,3.6463592,3.8859491,3.8038976,3.879385,4.2272825,4.6145644,4.965744,5.5007186,5.865026,6.088206,6.5870776,6.8529234,6.7971287,6.121026,4.716308,2.6617439,3.0982566,4.201026,5.2447186,6.12759,7.39118,7.397744,7.5421543,7.456821,7.3058467,7.788308,8.1755905,8.064001,8.004924,8.224821,8.615385,8.73354,8.342975,8.077128,7.9458466,7.3353853,7.5881033,7.8637953,7.7357955,6.626462,3.8301542,4.7491283,3.6824617,2.7142565,2.6256413,2.8980515,3.1737437,5.602462,8.096821,8.178872,2.993231,3.4100516,2.9243078,3.6594875,4.6834874,1.9954873,5.356308,5.477744,5.1200004,5.5991797,6.820103,8.205129,8.201847,7.890052,7.8047185,7.958975,6.806975,7.5618467,6.232616,3.564308,5.041231,7.3583593,8.87795,9.613129,10.010257,10.94236,8.625232,7.381334,6.3474874,5.7796926,7.030154,5.8486156,5.093744,4.4734364,3.7251284,2.5993848,2.3762052,2.3729234,2.3171284,2.2744617,2.6486156,2.034872,1.8543591,1.9528207,2.2416413,2.681436,2.7733335,3.2525132,3.8400004,4.2469745,4.1517954,3.9844105,3.8629746,4.1583595,4.8344617,5.435077,5.4908724,5.346462,5.290667,5.435077,5.7140517,5.907693,6.4557953,6.813539,6.872616,6.954667,7.197539,7.6242056,8.01477,8.172308,7.958975,7.256616,6.6395903,6.0980515,5.691077,5.543385,6.11118,6.265436,6.265436,6.2194877,6.0685134,6.262154,5.7731285,5.4974365,5.549949,5.2676926,4.204308,3.7152824,3.05559,2.1464617,1.5688206,1.4867693,1.2504616,1.1552821,1.1716924,0.94523084,0.7220513,0.5677949,0.48246157,0.39712822,0.19692309,0.24287182,0.27569234,0.3117949,0.3511795,0.36758977,0.26256412,0.16738462,0.101743594,0.108307704,0.256,0.7122052,0.9682052,0.9616411,0.8402052,0.9747693,1.204513,1.1257436,1.1158975,1.2176411,1.1323078,1.2800001,1.4834872,1.5524104,1.5163078,1.6180514,1.7066668,2.300718,2.7142565,2.7569232,2.7306669,2.678154,2.678154,2.5074873,2.1924105,1.9954873,2.1300514,2.3729234,2.3204105,1.8806155,1.2964103,1.4539489,1.4966155,1.394872,1.2537436,1.3193847,1.1093334,1.2832822,1.595077,1.8510771,1.8937438,1.5589745,1.3620514,1.1290257,0.8730257,0.78769237,0.9616411,1.1716924,1.1913847,1.1257436,1.4145643,1.6640002,1.5556924,1.3193847,1.0535386,0.73517954,0.7450257,0.7056411,0.67282057,0.7122052,0.9189744,4.007385,4.201026,3.9975388,3.8564105,3.9909747,4.384821,4.201026,3.9778464,3.826872,3.82359,3.9778464,4.1878977,4.059898,4.266667,4.8344617,5.159385,5.4383593,5.3727183,5.612308,6.413129,7.634052,8.356103,8.326565,7.955693,7.529026,7.207385,7.1056414,7.4732313,8.093539,8.648206,8.73354,9.196308,9.344001,9.4457445,9.540924,9.435898,9.921641,10.161232,10.003693,9.577026,9.317744,9.517949,9.970873,10.400822,10.817642,11.529847,11.500309,11.644719,12.209231,12.839386,12.576821,12.921437,13.732103,13.925745,13.564719,13.850258,15.711181,17.903591,19.456001,19.954874,19.580719,17.742771,15.599591,14.792206,15.940925,18.642054,12.806565,6.439385,2.2646155,0.85005134,0.6301539,0.380718,0.17066668,0.059076928,0.04266667,0.059076928,0.049230773,0.01969231,0.0,0.006564103,0.036102567,0.006564103,0.0,0.0,0.0,0.0032820515,0.0,0.0,0.013128206,0.026256412,0.016410258,0.07548718,0.08861539,0.08205129,0.07548718,0.07876924,0.06564103,0.059076928,0.15097436,0.27241027,0.19692309,0.052512825,0.013128206,0.006564103,0.0032820515,0.01969231,0.0032820515,0.006564103,0.02297436,0.029538464,0.0,0.01969231,0.14769232,0.30851284,0.39712822,0.29538465,0.7187693,0.61374366,0.39712822,0.256,0.15097436,0.29210258,0.5677949,0.8467693,0.99774367,0.90256417,1.7755898,1.3193847,0.8566154,0.82379496,0.7778462,0.7581539,0.8533334,1.0469744,1.2832822,1.4572309,1.847795,2.3630772,2.733949,2.8160002,2.5862565,2.8717952,4.1058464,5.904411,7.6734366,8.602257,9.176616,9.16677,9.209436,9.334154,8.969847,9.488411,9.170052,8.861539,9.061745,9.91836,9.449026,8.946873,8.841846,8.881231,8.113232,7.2205133,6.957949,7.2664623,7.716103,7.506052,6.8660517,6.6428723,6.931693,7.709539,8.854975,8.759795,8.41518,7.6996927,6.957949,6.987488,8.963283,11.516719,13.689437,14.532925,13.10195,10.86359,10.522257,11.58236,13.013334,13.243078,11.434668,10.233437,10.496001,11.621744,11.565949,12.33395,12.527591,11.907283,10.55836,8.87795,7.7456417,7.4108725,7.781744,8.54318,9.163487,9.304616,9.659078,10.125129,10.758565,11.776001,12.1238985,12.501334,12.438975,12.235488,12.967385,13.607386,13.791181,14.129231,14.486976,13.99795,14.644514,15.763694,16.403694,16.193642,15.314053,14.795488,15.343591,15.566771,14.70359,12.596514,10.016821,11.211488,13.312001,14.611693,14.55918,13.318565,12.425847,11.762873,11.254155,10.866873,10.9456415,10.295795,9.931488,10.023385,9.898667,10.57477,11.10318,11.61518,11.82195,11.008,9.334154,8.986258,9.301334,9.370257,8.03118,7.6964107,7.821129,8.034462,8.070564,7.778462,7.643898,6.7544622,5.5762057,4.6867695,4.7622566,4.850872,4.201026,3.1409233,2.1103592,1.6475899,1.2931283,1.3029745,1.657436,2.2121027,2.6978464,3.3444104,4.076308,4.6933336,4.8738465,4.1813335,4.673641,4.8640003,4.6572313,4.010667,2.937436,1.9003079,2.0841026,2.0250258,1.4703591,1.3653334,1.8313848,3.1803079,4.2436924,4.345436,3.3017437,1.7329233,1.1651284,1.6443079,2.228513,0.9911796,1.0962052,1.2832822,1.7624617,2.2777438,2.0939488,2.0217438,2.0775387,2.1858463,2.2613335,2.2055387,2.6715899,3.3444104,4.0500517,4.5095387,4.33559,3.9647183,4.027077,4.4373336,4.969026,5.2447186,4.9099493,4.9296412,4.673641,4.20759,4.3060517,4.647385,5.7042055,5.7731285,4.919795,4.962462,4.637539,4.6572313,4.7392826,4.8344617,5.1298466,6.5936418,7.3452315,6.7872825,5.0215387,2.8488207,1.5556924,7.899898,15.737437,21.444925,23.945848,12.498053,9.019077,7.0465646,5.228308,7.3353853,5.973334,4.562052,5.5565133,8.694155,10.971898,10.210463,8.730257,7.716103,7.0137444,5.1200004,4.650667,8.375795,9.40636,6.2227697,2.6683078,3.3936412,5.408821,7.0925136,8.667898,12.196103,16.361027,13.019898,10.217027,10.282667,9.846154,11.687386,10.289231,9.202872,8.914052,6.8299494,7.276308,6.439385,5.5893335,5.3070774,5.467898,3.826872,2.4746668,1.5589745,1.270154,1.847795,1.8412309,1.5195899,1.657436,2.2547693,2.540308,2.1497438,1.9495386,1.7263591,1.4276924,1.1520001,1.2307693,1.529436,1.7591796,1.7887181,1.6508719,1.6935385,1.7624617,1.847795,1.9364104,1.9954873,2.034872,2.0709746,2.100513,2.1070771,2.0578463,1.9954873,1.7394873,1.6410258,1.7362052,1.7427694,2.1956925,2.4451284,2.605949,2.7634873,2.9702566,2.353231,1.6672822,1.2209232,1.0896411,1.1093334,1.2668719,1.1881026,1.0436924,0.8960001,0.69907695,0.67938465,0.63343596,0.58092314,0.6235898,0.9485129,1.1093334,1.2504616,1.2635899,1.1520001,1.0075898,1.1323078,1.522872,1.8806155,2.028308,1.9167181,1.7460514,1.8281027,1.9462565,1.9528207,1.7887181,1.7624617,1.6147693,1.404718,1.2274873,1.2077949,1.3161026,1.3554872,1.3587693,1.3522053,1.3686155,1.5524104,1.4309745,1.2438976,1.2012309,1.4834872,1.782154,1.847795,2.0873847,2.546872,2.92759,2.8258464,3.3378465,3.9811285,4.3684106,4.2174363,4.460308,4.4406157,4.135385,3.7316926,3.629949,3.95159,3.895795,4.0041027,4.414359,4.841026,4.9854364,5.139693,5.297231,5.5893335,6.2916927,6.997334,7.0498466,6.413129,5.2480006,3.9122055,3.754667,4.466872,5.412103,6.3245134,7.3353853,7.906462,8.073847,8.034462,8.146052,8.92718,9.527796,9.6525135,9.754257,10.026668,10.41395,9.636104,8.65477,7.88677,7.325539,6.521436,7.240206,7.9294367,8.218257,7.453539,4.699898,4.263385,3.623385,3.0293336,2.7963078,3.2820516,2.8422565,5.32677,7.6603084,7.8441033,4.955898,3.0096412,2.297436,2.8356924,3.6660516,2.8717952,5.3792825,5.914257,6.416411,7.0334363,6.117744,8.756514,8.690872,8.208411,7.817847,6.2588725,5.7042055,6.163693,5.435077,3.8990772,4.522667,6.3507695,8.116513,9.304616,10.112,11.464206,8.241231,7.4732313,6.692103,5.4514875,5.330052,4.013949,3.8859491,4.164923,4.194462,3.436308,3.0030773,3.0358977,2.9997952,2.7831798,2.681436,1.9626669,2.169436,2.2678976,2.0512822,2.1530259,2.612513,3.0391798,3.751385,4.565334,4.775385,4.4242053,4.378257,4.673641,5.156103,5.5007186,5.7468724,5.362872,5.428513,5.9634876,5.924103,6.5805135,7.243488,7.4436927,7.243488,7.240206,7.7718983,8.2904625,8.385642,8.283898,8.858257,7.7292314,6.7150774,5.9634876,5.586052,5.661539,5.8912826,5.927385,5.9930263,6.1078978,6.0619493,5.87159,5.0543594,4.706462,4.9788723,5.0642056,4.3290257,3.6594875,3.0358977,2.4188719,1.7788719,1.4375386,1.2307693,1.1093334,0.9944616,0.7581539,0.512,0.49230772,0.46933338,0.3511795,0.17394873,0.256,0.33476925,0.4135385,0.4660513,0.4397949,0.28882053,0.17066668,0.101743594,0.13784617,0.36430773,0.6892308,0.83035904,0.8467693,0.81394875,0.8467693,1.0929232,1.1782565,1.1651284,1.1191796,1.086359,1.2077949,1.4309745,1.4933335,1.4375386,1.6016412,1.7394873,2.0578463,2.3204105,2.484513,2.7044106,2.6354873,2.6289232,2.5895386,2.4582565,2.2022567,2.284308,2.4484105,2.284308,1.7558975,1.1979488,1.3128207,1.2438976,1.1913847,1.2471796,1.3817437,1.3128207,1.5458462,1.7690258,1.8281027,1.719795,1.2340513,1.083077,1.017436,0.9189744,0.8041026,0.7220513,1.0633847,1.1782565,1.0436924,1.2668719,1.5622566,1.5327181,1.3718976,1.1454359,0.80738467,0.79425645,0.76800007,0.8467693,1.0732309,1.3915899,3.9220517,4.007385,3.4691284,3.0293336,3.0916924,3.7382567,4.4832826,4.394667,3.9680004,3.5971284,3.5872824,3.623385,3.7874875,4.2502565,4.7950773,4.8049235,5.3694363,5.7468724,6.11118,6.5936418,7.27959,7.827693,8.2215395,8.3134365,8.329846,8.881231,8.805744,8.999385,9.458873,9.833026,9.429334,9.101129,9.07159,8.805744,8.178872,7.506052,8.960001,9.5146675,9.741129,9.878975,9.842873,10.453334,10.5780525,10.893129,11.588924,12.360206,12.603078,12.471796,12.832822,13.515489,13.321847,14.358975,15.826053,16.315079,16.219898,17.746052,19.173744,21.700924,23.568413,24.231386,24.352823,19.810463,15.37313,15.195899,16.896002,11.536411,9.265231,4.522667,1.1224617,0.18051283,0.108307704,0.068923086,0.06235898,0.04266667,0.068923086,0.28882053,0.23958977,0.09189744,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.0032820515,0.0,0.036102567,0.07548718,0.016410258,0.12471796,0.068923086,0.009846155,0.006564103,0.029538464,0.006564103,0.026256412,0.61374366,1.2242053,0.25928208,0.11158975,0.06564103,0.036102567,0.01969231,0.09189744,0.01969231,0.036102567,0.036102567,0.0,0.0,0.0,0.0,0.40369233,1.0633847,1.2964103,0.5284103,1.014154,1.2931283,0.92225647,0.45620516,0.761436,1.1684103,0.92553854,0.28225642,0.48902568,0.5481026,0.53825647,0.71548724,0.9485129,0.7187693,0.9616411,1.5163078,1.8281027,1.9692309,2.6387694,2.9801028,3.4067695,3.5840003,3.3280003,2.609231,3.8432825,4.4077954,5.1265645,6.4557953,8.467693,9.921641,10.322052,10.729027,10.824206,8.89436,8.467693,7.8670774,7.936001,8.648206,9.124104,9.222565,8.195283,7.578257,7.5421543,6.882462,5.979898,6.11118,6.7938466,7.581539,8.057437,8.704,9.478565,9.521232,9.002667,9.124104,9.6754875,9.517949,8.674462,7.683283,7.5979495,10.932513,13.37436,14.601848,14.17518,11.54954,11.355898,12.028719,12.786873,13.121642,12.816411,11.034257,10.197334,10.630565,11.943385,13.029744,14.14236,13.761642,12.1238985,9.852718,7.9491286,8.04759,7.972103,8.234667,8.920616,9.688616,10.788103,11.116308,11.1983595,11.32636,11.58236,11.654565,11.848206,11.414975,10.893129,12.100924,13.735386,14.162052,14.700309,15.330462,14.693745,14.998976,15.862155,16.022976,15.16636,13.945437,13.505642,13.991385,14.260514,14.244103,14.953027,11.963078,12.104206,13.282462,14.158771,14.145642,13.400617,13.489232,13.420309,12.747488,11.54954,11.648001,10.820924,10.023385,9.498257,8.789334,9.875693,11.162257,12.140308,12.363488,11.460924,9.885539,8.986258,8.779488,8.851693,8.362667,7.8506675,7.9228725,8.329846,8.6580515,8.316719,7.643898,6.7807183,6.121026,5.579488,4.578462,4.8836927,4.161641,3.1113849,2.2350771,1.8313848,1.4145643,1.3751796,1.6147693,2.0250258,2.5009232,3.442872,4.84759,5.464616,5.0838976,4.5456414,5.0116925,4.8705645,4.6145644,4.132103,2.7175386,1.9364104,1.6016412,1.2668719,0.99774367,1.3883078,0.54482055,2.359795,5.549949,8.562873,9.55077,3.131077,1.0765129,1.3226668,1.8937438,0.9321026,1.0666667,1.273436,1.522872,1.7755898,1.9823592,2.1530259,2.4615386,2.5665643,2.3762052,2.0611284,2.865231,3.6627696,4.2174363,4.4701543,4.532513,4.33559,4.8738465,5.4908724,5.76,5.477744,5.1232824,5.034667,4.84759,4.5128207,4.31918,4.709744,5.1167183,5.152821,4.8771286,4.7917953,3.7054362,3.2032824,3.5413337,4.568616,5.7534366,6.3868723,10.555078,11.0375395,6.9645133,3.8137438,2.1792822,5.4153852,11.090053,17.033848,21.333336,11.664412,9.127385,7.9425645,7.896616,14.342566,9.238976,6.042257,6.2129235,8.772923,10.299078,10.164514,8.986258,10.243283,12.104206,7.4141545,2.484513,4.70318,6.8266673,5.7665644,2.5928206,1.8379488,2.5009232,4.056616,6.055385,8.116513,12.5374365,12.678565,11.283693,9.846154,8.635077,10.039796,9.366975,10.312206,12.005745,9.002667,6.452513,5.786257,6.0849237,6.75118,7.506052,6.567385,4.519385,2.5304618,1.4572309,1.847795,1.8707694,1.3259488,1.017436,1.1979488,1.5885129,1.2931283,1.0469744,0.9616411,0.95835906,0.761436,0.761436,0.8730257,1.0666667,1.2603078,1.2964103,1.3226668,1.3095386,1.3029745,1.3128207,1.3128207,1.3620514,1.5753847,1.6738462,1.6311796,1.6771283,2.0578463,1.785436,1.6804104,1.9003079,1.9364104,2.6453335,2.868513,2.8455386,2.8488207,3.190154,2.934154,2.162872,1.4998976,1.1585642,0.97805136,1.1716924,1.1749744,1.1126155,1.0043077,0.74830776,0.60061544,0.574359,0.58092314,0.62030774,0.7778462,1.0469744,1.204513,1.3751796,1.4834872,1.2504616,1.142154,1.5622566,1.8609232,1.9396925,2.2580514,2.1366155,2.3696413,2.6157951,2.7175386,2.7175386,2.5337439,2.2580514,1.9462565,1.6246156,1.2832822,1.086359,1.3226668,1.723077,2.0742567,2.1956925,2.3433847,2.0611284,1.7066668,1.5064616,1.5556924,1.9232821,2.0151796,2.038154,2.3171284,3.2820516,3.4625645,3.7382567,4.092718,4.4865646,4.850872,5.2414365,4.7556925,4.345436,4.420923,4.8377438,5.228308,5.0149746,4.562052,4.279795,4.6080003,4.890257,4.8672824,5.0215387,5.5236926,6.2555904,7.1844106,7.8637953,7.6635904,6.6461544,5.586052,4.594872,5.3727183,6.2523084,6.616616,6.8955903,7.6898465,7.9819493,8.205129,8.681026,9.596719,10.696206,10.916103,10.909539,10.975181,11.047385,9.803488,8.851693,7.972103,6.948103,5.5696416,6.7183595,8.241231,9.124104,8.677744,6.5312824,3.7120004,3.2820516,2.9801028,2.4024618,2.9768207,2.4385643,4.6933336,7.722667,10.033232,10.679795,4.6145644,2.556718,2.166154,2.665026,4.8377438,6.045539,6.51159,7.312411,7.8506675,5.874872,8.36595,8.402052,8.283898,7.8080006,4.2568207,5.3924108,4.9362054,4.3684106,3.9614363,2.7766156,4.7917953,6.675693,6.8955903,5.858462,5.920821,5.395693,5.3366156,5.7698464,6.3442054,6.3310776,3.9384618,3.9187696,3.9253337,3.4494362,3.8137438,3.754667,3.7382567,3.6824617,3.4888208,3.0358977,2.2678976,2.6617439,2.8816411,2.5304618,2.1530259,2.8947694,3.31159,3.6594875,4.0303593,4.348718,4.6900516,5.0215387,5.175795,5.218462,5.4613338,5.914257,5.3760004,5.2480006,5.7632823,5.9963083,7.181129,7.9885135,8.01477,7.2861543,6.2851286,7.640616,8.36595,8.388924,8.198565,8.835282,7.8703594,7.017026,6.2096415,5.5893335,5.477744,5.8453336,6.265436,6.485334,6.5247183,6.6822567,6.377026,5.293949,4.9296412,5.2447186,4.6834874,4.3290257,3.6562054,2.8192823,2.156308,2.1825643,1.8904617,1.5327181,1.2274873,0.9878975,0.7318975,0.5874872,0.5677949,0.47589746,0.29538465,0.19692309,0.27241027,0.4266667,0.5973334,0.6465641,0.36758977,0.14769232,0.09189744,0.12143591,0.20348719,0.3511795,0.55794877,0.6662565,0.7384616,0.7975385,0.80738467,1.0765129,1.1716924,1.1585642,1.1585642,1.3423591,1.3686155,1.4834872,1.5064616,1.4178462,1.3587693,1.7985642,2.0184617,2.3040001,2.6912823,2.9604106,3.0096412,3.0030773,3.0752823,3.0818465,2.5928206,2.605949,2.481231,2.103795,1.6016412,1.3587693,1.5425643,1.276718,1.2635899,1.5655385,1.6016412,1.4572309,1.3817437,1.4506668,1.5885129,1.5885129,1.3062565,1.3456411,1.401436,1.3193847,1.0994873,0.9288206,1.1224617,1.2077949,1.1093334,1.1454359,1.401436,1.6475899,1.5195899,1.1126155,0.9911796,1.1126155,1.1716924,1.3292309,1.6836925,2.2580514,3.0293336,3.058872,3.1277952,3.1967182,3.3345644,3.7382567,4.4734364,4.588308,4.135385,3.5872824,3.817026,4.4307694,4.6966157,4.818052,4.97559,5.3202057,6.055385,6.377026,6.449231,6.482052,6.7183595,7.1581545,7.6570263,8.100103,8.484103,8.917334,8.825437,8.5661545,8.598975,8.930462,9.124104,9.03877,8.963283,8.982975,9.035488,8.910769,8.946873,8.694155,8.900924,9.596719,10.098872,10.492719,10.761847,10.857026,11.027693,11.848206,13.144616,13.988104,14.119386,13.919181,14.408206,16.498873,17.513027,17.801847,18.097233,19.515078,20.240412,22.885746,25.472002,25.875694,21.838772,19.124514,19.790771,21.097027,19.347694,9.888822,4.775385,1.782154,0.4201026,0.108307704,0.19364104,0.3117949,0.53825647,0.45620516,0.15097436,0.20348719,0.08861539,0.02297436,0.0,0.0032820515,0.013128206,0.0032820515,0.0,0.0,0.0,0.0032820515,0.0,0.0,0.016410258,0.036102567,0.016410258,0.20348719,0.21333335,0.15097436,0.10502565,0.128,0.06564103,0.098461546,0.27569234,0.40697438,0.08861539,0.07876924,0.03938462,0.006564103,0.0032820515,0.01969231,0.0032820515,0.006564103,0.006564103,0.0,0.0,0.0,0.013128206,0.13456412,0.3511795,0.56451285,0.7122052,1.0043077,1.142154,1.2832822,2.0217438,1.8182565,1.3718976,0.84348726,0.46276927,0.52512825,0.60389745,0.69251287,0.92553854,1.0994873,0.67938465,1.6082052,1.6377437,1.5556924,2.0086155,3.5314875,4.086154,4.647385,4.3585644,3.4166157,3.0490258,3.1376412,4.164923,5.4580517,7.026872,9.567181,11.116308,11.680821,11.96636,11.621744,9.212719,8.835282,8.297027,8.218257,8.421744,7.939283,6.944821,6.6395903,7.6077952,9.124104,9.140513,7.571693,6.7314878,6.76759,7.5552826,8.704,9.682052,9.091283,8.907488,9.360411,8.917334,9.494975,9.691898,9.586872,9.731283,11.152411,14.483693,16.833643,17.211079,15.648822,13.197129,12.291283,12.632616,12.822975,12.196103,10.81436,10.528821,11.168821,12.153437,13.115078,13.896206,14.040616,12.409437,10.9686165,10.253129,9.366975,8.87795,8.411898,8.592411,9.465437,10.505847,11.264001,11.667693,11.523283,11.096616,11.116308,10.535385,10.857026,11.23118,11.529847,12.356924,13.8765135,14.529642,15.113848,15.924514,16.745028,16.62031,16.534975,16.072206,15.192616,14.214565,13.794462,14.181745,14.457437,14.480412,14.903796,13.203693,13.4400015,14.641232,15.675078,15.241847,12.750771,12.235488,12.018872,11.529847,11.270565,11.963078,11.352616,10.308924,9.347282,8.631796,9.209436,9.770667,10.213744,10.564924,10.971898,10.528821,10.230155,9.593436,8.776206,8.582564,8.057437,8.260923,8.549745,8.621949,8.523488,7.5979495,6.8332314,6.3343596,5.924103,5.1265645,4.857436,4.2929235,3.4067695,2.4549747,1.9528207,1.6344616,1.585231,1.782154,2.1858463,2.7109745,3.3378465,4.0369234,4.8771286,5.5663595,5.4514875,5.474462,4.778667,4.4767184,4.384821,2.9965131,2.1464617,1.7394873,1.4375386,1.2504616,1.5360001,0.77128214,1.1093334,3.0851285,5.671385,6.2818465,4.3027697,3.629949,2.5665643,1.0929232,0.88287187,0.9878975,1.332513,1.6771283,1.9167181,2.0939488,2.1464617,2.477949,2.733949,2.678154,2.1956925,2.7864618,3.5577438,4.161641,4.5522056,4.9952826,5.32677,6.0685134,6.482052,6.193231,5.208616,5.0904617,5.21518,5.169231,4.854154,4.453744,4.6769233,5.1987696,5.402257,5.1298466,4.6933336,3.508513,3.3575387,4.0500517,5.0215387,5.32677,5.7534366,9.741129,11.556104,9.298052,4.890257,4.8147697,5.474462,8.464411,11.812103,9.96759,9.731283,6.770872,5.10359,6.3245134,9.6065645,10.246565,7.6635904,6.741334,8.854975,11.874462,12.383181,10.217027,10.532104,13.6697445,15.143386,8.989539,6.8463597,5.8453336,4.781949,4.1091285,4.2502565,5.654975,6.2884107,6.235898,7.702975,8.362667,8.717129,9.301334,9.760821,8.854975,9.557334,10.748719,11.418258,10.840616,8.598975,7.9130263,7.056411,7.017026,7.240206,5.602462,3.7448208,3.7382567,3.892513,3.387077,2.2744617,3.058872,2.4057438,1.4408206,0.8172308,0.7187693,0.63343596,0.5546667,0.46933338,0.39712822,0.39712822,0.4266667,0.4201026,0.512,0.7056411,0.86974365,1.0305642,0.9353847,0.8172308,0.79097444,0.8598975,0.9288206,1.0732309,1.2406155,1.3751796,1.4342566,1.6672822,1.7755898,1.7362052,1.7033848,2.0217438,3.4625645,4.1780515,4.332308,4.2436924,4.3618464,3.7710772,3.045744,2.3991797,1.9429746,1.6738462,1.6738462,1.5622566,1.3883078,1.1979488,1.0272821,0.84348726,0.761436,0.69907695,0.6629744,0.75487185,0.7975385,0.9747693,1.1946667,1.3653334,1.3981539,1.591795,1.7427694,1.7920002,1.8543591,2.2219489,2.4024618,2.809436,2.993231,2.9538465,3.117949,3.318154,3.1606157,2.733949,2.281026,2.172718,2.162872,2.4385643,2.8553848,3.2886157,3.626667,3.4100516,3.2918978,3.5380516,3.9614363,3.9122055,3.6627696,3.5774362,3.5971284,3.7251284,4.023795,3.9745643,4.07959,4.1911798,4.2535386,4.3290257,4.4832826,4.128821,3.9581542,4.348718,5.349744,6.042257,5.9503593,5.398975,4.900103,5.1331286,5.208616,4.9985647,5.037949,5.579488,6.5870776,6.9677954,7.4436927,7.0432825,5.612308,3.826872,4.4701543,5.3825645,6.009436,6.2752824,6.6034875,6.557539,7.450257,8.247795,8.628513,8.986258,9.176616,9.120821,9.238976,9.609847,9.938052,8.438154,7.4797955,6.885744,6.669129,7.0465646,7.4797955,8.267488,8.503796,7.506052,4.8082056,4.010667,3.9778464,3.0326157,1.9692309,4.0369234,2.7766156,4.3749747,6.554257,8.28718,9.813334,10.886565,7.765334,6.1046157,6.810257,6.045539,5.4580517,5.533539,6.1374364,6.482052,5.1298466,6.957949,6.921847,7.059693,7.13518,4.647385,4.493129,4.3290257,4.4242053,4.309334,2.7536411,5.3234878,6.820103,6.6560006,5.546667,5.5302567,4.896821,5.0904617,5.9634876,6.892308,6.7840004,5.435077,4.6867695,4.279795,4.027077,3.826872,3.6004105,3.4756925,3.1737437,2.793026,2.8291285,2.8914874,3.1474874,3.3509746,3.3345644,2.993231,2.878359,2.809436,3.1770258,3.945026,4.640821,5.32677,5.362872,5.47118,5.8978467,6.413129,5.9569235,4.9362054,4.6966157,5.5171285,6.6067696,7.7325134,8.342975,8.231385,7.702975,7.581539,7.64718,7.53559,7.496206,7.5388722,7.430565,7.9130263,7.4108725,6.675693,6.242462,6.4557953,6.088206,6.5017443,6.669129,6.485334,6.7807183,6.416411,5.3398976,5.1659493,5.6320004,4.6112823,4.588308,3.9680004,3.1015387,2.2416413,1.5360001,1.3784616,1.0568206,0.8041026,0.67610264,0.53825647,0.5481026,0.45620516,0.32164106,0.23630771,0.3314872,0.35774362,0.37743592,0.35774362,0.28225642,0.14769232,0.072205134,0.08533334,0.13784617,0.2231795,0.3511795,0.44964105,0.54482055,0.6465641,0.7220513,0.67282057,0.88287187,0.90584624,0.8730257,0.9189744,1.1716924,1.3718976,1.6114873,1.6377437,1.5392822,1.7624617,2.0545642,2.2514873,2.4910772,2.7175386,2.7044106,2.793026,3.0293336,3.249231,3.245949,2.7766156,2.612513,2.5764105,2.3236926,1.9889232,2.162872,1.8379488,1.6213335,1.5721027,1.5688206,1.332513,1.273436,1.522872,1.7099489,1.6935385,1.5885129,1.3062565,1.463795,1.5425643,1.4145643,1.3423591,1.4441026,1.5195899,1.6377437,1.7952822,1.9003079,2.041436,1.8838975,1.4867693,1.0896411,1.1126155,1.401436,1.7001027,1.9790771,2.1530259,2.0644104,2.9801028,3.045744,3.0982566,3.2098465,3.4067695,3.6824617,4.1222568,4.269949,4.1517954,3.9876926,4.1780515,4.6112823,4.965744,5.175795,5.395693,5.970052,6.294975,6.669129,6.816821,6.695385,6.5017443,6.6461544,7.384616,8.182155,8.763078,9.091283,9.015796,9.061745,9.363693,9.754257,9.744411,9.521232,8.858257,8.641642,8.94359,9.015796,8.530052,8.231385,8.375795,8.881231,9.31118,10.164514,10.361437,10.541949,11.096616,12.176412,12.947693,14.171899,15.025232,15.199181,14.907078,15.983591,16.692514,17.430975,18.38277,19.5479,21.398975,23.844105,24.280617,22.52472,20.808207,17.778873,19.987694,22.075079,20.552206,13.778052,4.388103,3.6890259,3.82359,1.9528207,0.25928208,0.6170257,0.8533334,0.86974365,0.6498462,0.26584616,0.13128206,0.04594872,0.009846155,0.013128206,0.032820515,0.029538464,0.016410258,0.009846155,0.009846155,0.01969231,0.03938462,0.04594872,0.036102567,0.02297436,0.02297436,0.16738462,0.17394873,0.14112821,0.12143591,0.1148718,0.108307704,0.36102566,0.39712822,0.16082053,0.01969231,0.18051283,0.08861539,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.128,0.3052308,0.3708718,0.5152821,1.1224617,1.4309745,1.5786668,2.5928206,1.9429746,1.4211283,1.0994873,0.9714873,0.98133343,0.9156924,1.1355898,1.3489232,1.3522053,1.0568206,1.6114873,1.5589745,1.7427694,2.5206156,3.7251284,4.601436,5.3169236,4.9854364,3.8038976,3.0752823,3.1442053,3.889231,5.031385,6.377026,7.827693,8.625232,9.301334,9.711591,9.869129,9.93477,9.7214365,9.330873,9.061745,8.897642,8.513641,8.109949,8.507077,9.754257,11.044104,10.71918,9.8592825,9.238976,9.005949,9.133949,9.432616,9.426052,8.746667,8.779488,9.53436,9.642668,10.30236,11.237744,11.71036,12.045129,13.604104,16.95836,18.993233,18.550156,16.144411,13.958565,12.4685135,12.678565,12.76718,12.097642,11.201642,11.559385,12.120616,12.928001,13.696001,13.810873,13.459693,11.963078,10.686359,10.043077,9.517949,9.462154,9.275078,9.829744,10.820924,10.765129,11.254155,11.385437,11.16554,10.84718,10.929232,10.778257,11.093334,11.533129,12.048411,12.859077,14.936617,15.392821,15.297642,15.42236,16.242872,16.449642,16.610462,16.164104,15.192616,14.401642,13.955283,14.034052,14.086565,14.060308,14.372104,14.464001,14.998976,15.990155,16.8599,16.433231,13.8765135,12.517745,11.670976,11.1064625,11.053949,11.98277,11.739899,10.633847,9.179898,8.086975,8.891078,9.570462,10.013539,10.220308,10.299078,10.71918,11.136001,10.57477,9.409642,9.360411,9.025641,8.933744,8.79918,8.556309,8.36595,7.3747697,6.5411286,6.173539,6.12759,5.7764106,5.421949,5.080616,4.3552823,3.2623591,2.231795,1.9528207,1.9823592,2.2153847,2.5895386,3.0916924,3.5544617,4.276513,5.211898,6.0061545,6.0160003,5.9503593,5.0116925,4.535795,4.4077954,3.058872,2.4385643,2.0053334,1.6902566,1.4572309,1.2964103,0.8598975,0.7581539,1.4145643,2.8422565,4.630975,4.926359,5.0674877,4.6572313,3.3378465,0.78769237,1.0765129,1.591795,2.028308,2.2416413,2.2580514,2.428718,2.4451284,2.537026,2.6847181,2.612513,3.0752823,3.879385,4.7589746,5.5958977,6.4032826,6.3606157,6.518154,6.3573337,5.8092313,5.2414365,5.284103,5.5958977,5.5565133,5.1659493,5.044513,5.2053337,5.2709746,5.146257,4.896821,4.7524104,3.9745643,3.8596926,4.201026,4.6211286,4.5587697,7.128616,8.457847,9.291488,9.580308,8.480822,9.728001,8.730257,9.170052,10.568206,8.27077,7.4863596,4.391385,2.9571285,3.9975388,5.156103,7.640616,7.6767187,7.8769236,9.344001,11.644719,15.399385,12.685129,9.993847,10.925949,16.20349,14.427898,10.180923,6.6494365,5.1856413,5.3202057,7.003898,8.172308,7.650462,6.4000006,7.5454364,8.464411,8.933744,9.45559,9.846154,9.258667,11.34277,11.542975,10.656821,9.360411,8.198565,8.182155,7.250052,6.055385,4.955898,4.010667,3.1442053,4.2240005,5.3005133,5.612308,5.5663595,4.9394875,2.8291285,1.2504616,0.7417436,0.37415388,0.24943592,0.21333335,0.18051283,0.14112821,0.16738462,0.19692309,0.19692309,0.24615386,0.3708718,0.54482055,0.702359,0.6695385,0.55794877,0.47589746,0.54482055,0.6859488,0.764718,0.8730257,1.0436924,1.2438976,1.4342566,1.7526156,1.8084104,1.6771283,1.8970258,3.4691284,4.2338467,4.5817437,4.706462,4.598154,4.1485133,3.7316926,3.2951798,2.7995899,2.2121027,2.103795,1.9626669,1.785436,1.6180514,1.5392822,1.3292309,1.1815386,1.017436,0.84348726,0.74830776,0.7056411,0.79097444,0.9616411,1.1979488,1.5163078,1.8576412,2.044718,2.1136413,2.1431797,2.2482052,2.5206156,2.9997952,3.2229745,3.1737437,3.2918978,3.7382567,3.9975388,3.8728209,3.5249233,3.4494362,3.5938463,3.5052311,3.5347695,3.761231,3.9909747,3.7874875,3.7710772,4.0467696,4.4996924,4.785231,4.6834874,4.601436,4.525949,4.4800005,4.5423594,4.5489235,4.6966157,4.84759,4.8771286,4.673641,4.601436,4.466872,4.2436924,4.1189747,4.4898467,5.221744,5.4547696,5.287385,5.0051284,5.080616,4.716308,4.5489235,4.781949,5.4153852,6.2096415,6.0225644,6.6002054,6.8332314,5.901129,3.2689233,4.31918,5.2676926,5.917539,6.1407185,5.8814363,5.8453336,6.8430777,7.6734366,7.9491286,8.103385,8.1755905,8.52677,9.074872,9.659078,10.033232,8.999385,8.001641,7.3714876,7.3091288,7.899898,7.4469748,7.6274877,7.755488,6.770872,3.242667,4.1091285,3.6758976,2.7536411,2.3893335,3.8728209,3.3903592,4.5423594,5.681231,6.3376417,7.2270775,10.663385,9.02236,7.525744,7.5913854,6.8496413,5.037949,4.7556925,5.1626673,5.4875903,5.0543594,6.47877,6.1505647,5.865026,5.6352825,3.6824617,4.4898467,4.6244106,4.4045134,3.9187696,3.0391798,4.972308,5.2611284,4.9952826,5.106872,6.373744,4.772103,4.850872,5.76,6.5378466,6.117744,5.933949,5.333334,4.7950773,4.4340515,4.0041027,3.6562054,3.436308,3.0982566,2.6880002,2.540308,3.0720003,3.3280003,3.3444104,3.1737437,2.865231,2.8717952,2.9801028,3.5905645,4.4832826,4.8147697,5.277539,5.2742567,5.5236926,6.052103,6.1768208,5.933949,5.4514875,5.2315903,5.58277,6.5936418,7.7718983,8.644924,9.130668,9.212719,8.966565,8.503796,7.2992826,6.6034875,6.669129,6.75118,7.174565,7.1089234,6.8463597,6.6592827,6.7905645,6.452513,6.7085133,6.954667,6.931693,6.741334,6.449231,5.8256416,5.7698464,5.8880005,4.5095387,3.9286156,3.5872824,3.3214362,2.7995899,1.529436,1.1355898,0.81394875,0.67610264,0.6498462,0.49887183,0.48902568,0.37743592,0.27897438,0.27897438,0.4397949,0.47261542,0.42994875,0.33476925,0.23958977,0.2297436,0.15425642,0.14112821,0.16410258,0.20348719,0.2231795,0.43651286,0.6826667,0.78769237,0.72861546,0.6301539,0.827077,0.9682052,0.98461545,0.9911796,1.276718,1.2406155,1.4211283,1.4506668,1.3784616,1.6771283,2.0512822,2.356513,2.6026669,2.806154,2.9702566,2.9702566,3.0260515,3.0654361,3.0227695,2.8488207,2.6880002,2.6617439,2.4910772,2.2383592,2.300718,1.9889232,1.8313848,1.7329233,1.6410258,1.5425643,1.6213335,1.7001027,1.7001027,1.5622566,1.2406155,1.2800001,1.5031796,1.6443079,1.657436,1.7165129,1.9659488,1.910154,1.9265642,2.1300514,2.356513,2.349949,2.1234872,1.7099489,1.3128207,1.2996924,1.4309745,1.7132308,1.913436,1.9462565,1.847795,3.6332312,3.6791797,3.6004105,3.495385,3.495385,3.757949,3.82359,3.9154875,4.20759,4.5522056,4.457026,4.70318,5.2020516,5.654975,6.0258465,6.5378466,6.488616,6.75118,7.076103,7.200821,6.875898,6.7314878,7.5520005,8.4283085,8.979693,9.347282,9.353847,9.672206,10.194052,10.522257,9.970873,9.426052,8.572719,8.303591,8.621949,8.65477,8.260923,8.320001,8.500513,8.700719,9.048616,10.148104,10.548513,11.053949,11.890873,12.694975,13.111795,14.336001,15.435489,15.747283,14.87754,15.018668,15.576616,16.692514,18.231796,19.797335,21.91754,22.806976,21.267694,19.206566,21.625437,17.864206,20.778667,21.691078,18.162872,13.99795,4.844308,4.9526157,6.189949,4.9920006,2.359795,1.0929232,0.73517954,0.71548724,0.6235898,0.21661541,0.12143591,0.04594872,0.013128206,0.026256412,0.068923086,0.118153855,0.10502565,0.06564103,0.026256412,0.02297436,0.052512825,0.055794876,0.049230773,0.06235898,0.13456412,0.72861546,0.6301539,0.41025645,0.31507695,0.28225642,0.24287182,0.43323082,0.380718,0.08533334,0.0,0.15425642,0.15097436,0.072205134,0.0,0.0,0.0,0.02297436,0.02297436,0.0,0.0,0.0,0.009846155,0.10502565,0.23302566,0.21989745,0.22646156,0.7318975,1.0075898,1.0896411,1.7887181,1.3259488,1.2406155,1.2603078,1.2438976,1.1585642,1.3292309,1.4375386,1.5130258,1.5458462,1.4900514,1.4309745,1.5195899,1.8543591,2.4582565,3.2623591,3.9712822,5.041231,4.926359,3.7021542,3.0752823,3.1409233,3.5183592,4.3552823,5.3398976,5.720616,6.485334,6.8430777,7.3583593,8.303591,9.6525135,9.895386,10.269539,10.361437,10.026668,9.393231,9.6065645,10.486155,11.707078,12.521027,11.759591,11.746463,11.34277,11.149129,11.093334,10.453334,9.508103,9.097847,9.225847,9.737847,10.345026,10.94236,11.933539,12.891898,13.8765135,15.42236,18.81272,20.555489,19.662771,16.843489,14.496821,12.918155,12.842668,12.583385,11.907283,12.022155,12.015591,12.517745,13.443283,13.958565,12.461949,12.2617445,11.812103,11.0145645,10.171078,9.957745,10.420513,10.532104,11.277129,12.3306675,12.048411,11.707078,11.316514,11.024411,10.857026,10.709334,11.188514,11.539693,11.782565,12.160001,13.13477,15.340309,15.75713,15.320617,14.795488,14.76595,15.445334,16.23631,16.17395,15.24513,14.375385,14.181745,13.99795,13.702565,13.53518,14.089848,16.019693,16.512001,16.748308,17.007591,16.708925,14.674052,13.331694,12.33395,11.631591,11.474052,12.268309,12.268309,11.16554,9.330873,7.817847,8.684308,9.662359,10.459898,10.801231,10.459898,10.696206,11.352616,10.994873,9.892103,10.020103,10.036513,9.668923,9.199591,8.868103,8.87795,7.709539,6.6067696,6.160411,6.242462,6.038975,5.9569235,5.9963083,5.543385,4.417641,2.858667,2.3893335,2.4188719,2.6847181,3.0391798,3.446154,3.7809234,4.7261543,5.6943593,6.2752824,6.235898,6.1407185,5.211898,4.6211286,4.352,3.186872,2.8455386,2.294154,1.8281027,1.522872,1.204513,1.0994873,0.81066674,0.71548724,1.3620514,3.4527183,3.892513,4.128821,4.2962055,4.325744,3.9614363,1.5721027,1.4998976,1.9987694,2.2416413,2.2777438,2.6486156,2.8521028,2.9440002,3.0358977,3.308308,3.748103,4.5817437,5.7698464,7.066257,8.021334,7.4863596,6.8430777,6.0356927,5.2676926,5.0182567,5.5762057,5.83877,5.612308,5.1987696,5.3924108,5.612308,5.3103595,4.965744,4.781949,4.70318,4.322462,4.240411,4.1846156,4.128821,4.3027697,6.8660517,6.4590774,6.8693337,9.015796,10.939077,12.57354,12.140308,11.605334,11.290257,9.862565,6.550975,3.3017437,1.8937438,2.2383592,2.359795,3.9844105,5.21518,6.557539,7.962257,8.845129,14.224411,12.786873,9.498257,8.500513,13.08554,15.553642,12.33395,8.835282,7.506052,7.8506675,9.107693,9.271795,8.169026,6.8233852,7.453539,10.033232,11.30995,11.487181,10.778257,9.40636,12.258463,12.27159,10.965334,9.6065645,9.202872,9.18318,8.704,6.2884107,3.4264617,4.571898,4.8738465,5.5204105,5.7632823,5.730462,6.419693,5.533539,3.249231,1.5524104,0.90584624,0.23958977,0.098461546,0.055794876,0.049230773,0.04594872,0.052512825,0.06564103,0.08861539,0.12143591,0.18051283,0.2986667,0.41025645,0.508718,0.49887183,0.4004103,0.33805132,0.48246157,0.54482055,0.65312827,0.8336411,1.0010257,1.2242053,1.5819489,1.7362052,1.6705642,1.6968206,3.131077,4.2371287,4.778667,4.785231,4.5554876,4.348718,4.0402055,3.6693337,3.255795,2.7864618,2.7142565,2.5042052,2.2219489,1.9561027,1.8313848,1.6246156,1.4802053,1.3292309,1.1355898,0.88943595,0.7253334,0.69579494,0.78769237,1.0404103,1.529436,1.913436,2.2646155,2.4155898,2.3794873,2.3696413,2.7011285,3.1245131,3.3378465,3.3542566,3.5052311,3.9712822,4.5423594,4.844308,4.8344617,4.785231,4.886975,4.5522056,4.194462,4.017231,3.9975388,3.9417439,4.1222568,4.31918,4.516103,4.890257,5.0018463,4.821334,4.5554876,4.3618464,4.345436,4.4373336,4.565334,4.7491283,4.9394875,5.024821,4.854154,4.841026,4.673641,4.2994876,3.9581542,4.1452312,4.5522056,4.906667,5.074052,5.0510774,4.457026,4.276513,4.5390773,5.097026,5.654975,5.182359,5.687795,6.311385,5.9602056,3.2689233,4.010667,4.886975,5.72718,6.2194877,5.910975,6.1078978,6.7314878,7.0990777,7.072821,7.069539,7.6274877,8.356103,9.110975,9.586872,9.3078985,8.874667,8.507077,8.201847,8.109949,8.536616,7.509334,7.2927184,7.3353853,6.416411,2.665026,3.7809234,3.114667,3.186872,4.013949,3.0851285,3.4166157,3.8432825,4.197744,4.535795,5.146257,7.3780518,8.139488,7.778462,7.128616,7.499488,5.3727183,5.1364107,5.549949,5.8453336,5.7435904,6.3343596,5.933949,5.2348723,4.414359,3.1573336,5.077334,5.159385,4.775385,4.5095387,4.1452312,4.5554876,4.2240005,3.8990772,4.2568207,5.8978467,4.8771286,5.1856413,5.920821,6.3606157,5.989744,6.2588725,5.914257,5.3103595,4.699898,4.2305646,3.7284105,3.3805132,3.0129232,2.6486156,2.4910772,3.0720003,3.3641028,3.3050258,3.0424619,2.9440002,3.314872,3.620103,3.9778464,4.352,4.571898,4.9887185,5.221744,5.605744,5.865026,5.146257,5.3169236,5.684513,6.0028725,6.308103,6.925129,7.906462,8.421744,8.881231,9.242257,8.996103,8.4972315,7.0990777,6.314667,6.442667,6.5870776,6.422975,6.5247183,6.675693,6.7544622,6.7117953,6.5837955,6.5378466,6.701949,6.8463597,6.363898,6.1308722,6.2030773,6.308103,5.9930263,4.6211286,4.1091285,3.5840003,3.308308,2.9702566,1.6640002,1.1191796,0.8336411,0.69907695,0.6170257,0.4660513,0.45620516,0.37743592,0.34133336,0.4004103,0.5316923,0.6104616,0.55794877,0.446359,0.3511795,0.3708718,0.21333335,0.18051283,0.20676924,0.24615386,0.27241027,0.5218462,0.7056411,0.76800007,0.7187693,0.62030774,0.7318975,1.0371283,1.1355898,1.0994873,1.4900514,1.3718976,1.4867693,1.5163078,1.4539489,1.6246156,1.9232821,2.231795,2.484513,2.740513,3.18359,2.9669745,2.9407182,2.917744,2.9078977,3.117949,2.9702566,2.806154,2.5764105,2.3072822,2.0939488,1.9528207,1.8773335,1.8313848,1.8445129,2.0217438,2.0742567,1.9429746,1.7099489,1.4080001,1.0436924,1.1815386,1.4309745,1.6508719,1.8051283,1.9396925,2.1497438,2.0808206,2.0578463,2.2449234,2.6322052,2.4910772,2.3138463,2.03159,1.7690258,1.8182565,1.6377437,1.7493335,1.8674873,1.8576412,1.7329233,4.565334,4.601436,4.4701543,4.141949,3.8334363,4.023795,3.7448208,3.8071797,4.3651285,4.9887185,4.663795,4.903385,5.3398976,5.910975,6.4754877,6.8233852,6.705231,6.810257,7.250052,7.755488,7.6931286,7.506052,8.14277,8.743385,9.032206,9.334154,9.577026,9.888822,10.368001,10.630565,9.793642,9.005949,8.628513,8.684308,8.920616,8.805744,8.720411,8.914052,9.028924,9.104411,9.563898,10.272821,11.0145645,11.979488,12.905026,13.065847,14.057027,14.92677,15.494565,15.593027,15.107284,15.130258,15.681643,17.001026,19.072002,21.605745,21.907694,21.192207,20.132105,20.09272,23.141745,19.328001,22.180105,20.532515,13.167591,8.812308,4.1485133,3.5282054,5.0084105,6.265436,4.59159,1.8379488,0.571077,0.15425642,0.0951795,0.055794876,0.01969231,0.0032820515,0.006564103,0.036102567,0.101743594,0.19692309,0.20676924,0.14112821,0.049230773,0.01969231,0.02297436,0.01969231,0.052512825,0.14441027,0.2986667,1.3981539,1.1913847,0.7450257,0.56451285,0.60389745,0.42338464,0.29210258,0.14441027,0.009846155,0.0032820515,0.006564103,0.15097436,0.14769232,0.0,0.0,0.026256412,0.055794876,0.04266667,0.0,0.0,0.0,0.016410258,0.01969231,0.009846155,0.01969231,0.06564103,0.04266667,0.101743594,0.27897438,0.47917953,0.5907693,0.90256417,1.1520001,1.1848207,0.95835906,1.6771283,1.5786668,1.5195899,1.6935385,1.6311796,1.3817437,1.7165129,1.910154,1.9003079,2.3040001,2.7733335,3.9253337,4.0369234,3.1606157,3.1245131,2.9768207,3.1474874,3.7120004,4.384821,4.5423594,5.8486156,5.7764106,6.3540516,7.8080006,8.52677,9.557334,10.9226675,11.835078,11.700514,10.112,10.361437,11.30995,12.557129,13.285745,12.274873,12.609642,12.032001,11.940104,12.288001,11.569232,10.125129,9.816616,10.000411,10.377847,10.978462,11.224616,11.713642,13.147899,15.432206,17.686975,21.00513,22.370462,20.955898,17.58195,14.720001,13.774771,13.354668,12.524308,11.602052,12.179693,11.529847,12.3536415,13.66318,13.833847,10.604308,10.633847,11.323078,11.277129,10.581334,10.774975,11.562668,11.802258,12.3306675,13.154463,13.459693,12.343796,11.621744,11.250873,10.994873,10.41395,11.319796,11.831796,11.946668,12.12718,13.302155,14.989129,15.717745,15.53395,14.7790785,14.066873,14.470565,15.494565,15.891693,15.307488,14.250668,14.342566,13.883078,13.328411,13.131488,13.748514,17.243898,17.26031,16.367592,15.875283,15.829334,14.529642,14.040616,13.512206,12.809847,12.504617,13.000206,12.895181,11.756309,9.90195,8.408616,8.776206,9.7673855,10.889847,11.631591,11.460924,10.837335,11.16554,10.912822,10.105436,10.354873,10.597744,10.174359,9.613129,9.3768215,9.865847,8.687591,7.2237954,6.422975,6.3277955,6.0652313,6.2194877,6.5936418,6.416411,5.395693,3.6890259,2.789744,2.6387694,2.9636924,3.4560003,3.7907696,4.1025643,5.1364107,6.0356927,6.416411,6.3507695,6.1046157,5.2742567,4.6769233,4.325744,3.4264617,3.2853336,2.5665643,1.8904617,1.5622566,1.5458462,1.5655385,0.9682052,0.69251287,1.1618463,2.281026,2.1267693,1.8937438,1.913436,3.43959,8.63836,2.4320002,1.1257436,1.4867693,1.8642052,2.1792822,2.7569232,3.56759,3.892513,3.8104618,4.1714873,4.7392826,5.684513,7.056411,8.546462,9.472001,8.651488,7.2927184,5.8978467,4.886975,4.6080003,5.8223596,5.8518977,5.408821,5.106872,5.4547696,5.8125134,5.395693,5.044513,4.9427695,4.6244106,4.4110775,4.338872,4.1222568,3.9417439,4.420923,4.906667,4.6276927,5.3202057,7.4436927,10.180923,12.002462,13.262771,13.252924,12.038565,10.456616,6.987488,4.125539,2.3072822,1.5622566,1.4933335,1.4703591,1.8707694,3.190154,4.7524104,4.7294364,8.41518,9.5606165,8.963283,7.955693,8.41518,11.552821,10.955488,9.908514,9.9282055,10.778257,9.501539,8.503796,7.827693,7.4699492,7.384616,10.57477,12.796719,13.249642,11.851488,9.219283,11.759591,12.534155,11.900719,11.090053,12.186257,11.513436,11.021129,7.955693,4.20759,6.294975,6.99077,7.3321033,6.2884107,4.4832826,4.201026,4.3716927,3.6496413,2.556718,1.3817437,0.17066668,0.0951795,0.04266667,0.016410258,0.013128206,0.013128206,0.013128206,0.029538464,0.049230773,0.08205129,0.14441027,0.21333335,0.380718,0.47589746,0.4266667,0.24287182,0.32164106,0.39056414,0.5481026,0.74830776,0.77456415,1.0436924,1.3161026,1.5360001,1.6344616,1.5360001,2.7503593,4.4077954,5.113436,4.7589746,4.529231,4.4373336,4.017231,3.5807183,3.3509746,3.4855387,3.436308,3.2032824,2.789744,2.3269746,2.0808206,1.8674873,1.7329233,1.657436,1.5589745,1.2668719,0.97805136,0.8172308,0.8205129,1.0108719,1.4145643,1.7657437,2.2383592,2.4385643,2.3794873,2.4910772,2.9702566,3.249231,3.3542566,3.4494362,3.8498464,4.273231,4.906667,5.5236926,5.930667,5.973334,5.8157954,5.3398976,4.70318,4.1222568,3.889231,3.9548721,4.338872,4.525949,4.460308,4.535795,4.6244106,4.3684106,4.027077,3.757949,3.620103,3.7415388,3.7874875,3.945026,4.3290257,5.0116925,4.8804107,4.916513,5.0543594,5.0871797,4.6834874,4.0336413,4.2207184,4.778667,5.2709746,5.293949,4.844308,4.562052,4.5554876,4.8114877,5.1922054,4.886975,5.1167183,5.504,5.333334,3.5282054,3.7907696,4.4701543,5.353026,6.170257,6.5936418,6.928411,7.1089234,6.921847,6.491898,6.2818465,7.1909747,7.778462,8.346257,8.572719,7.5454364,7.53559,8.306872,8.73354,8.67118,8.966565,8.034462,7.712821,7.5913854,6.5969234,3.006359,3.1343591,2.6518977,3.7316926,5.182359,2.4582565,2.993231,2.5632823,2.4582565,3.045744,3.764513,3.9548721,6.7905645,7.6767187,6.4656415,7.4436927,5.914257,6.048821,6.5017443,6.626462,6.445949,6.114462,6.0061545,5.1954875,3.9581542,3.7776413,5.61559,5.717334,5.618872,5.7009234,5.1954875,4.348718,4.342154,3.889231,3.2065644,4.0041027,5.2447186,6.0947695,6.4623594,6.49518,6.564103,6.6100516,6.308103,5.7140517,5.0116925,4.4996924,3.7743592,3.239385,2.7306669,2.3860514,2.6322052,2.9111798,3.1573336,3.2000003,3.1409233,3.3542566,3.9286156,4.263385,4.1058464,3.8038976,4.3027697,4.788513,5.169231,5.5729237,5.6320004,4.4734364,4.663795,5.467898,6.518154,7.3616414,7.4469748,8.001641,7.7981544,7.7423596,7.9852314,7.90318,7.5881033,6.875898,6.5805135,6.73477,6.62318,6.1341543,6.11118,6.265436,6.373744,6.2884107,6.304821,6.091488,5.979898,5.9634876,5.7140517,5.4941545,6.189949,6.482052,6.012718,5.398975,5.3136415,4.2994876,3.43959,2.8750772,1.8116925,1.3259488,1.0404103,0.78769237,0.54482055,0.43323082,0.48246157,0.43323082,0.4201026,0.49230772,0.5907693,0.65969235,0.6301539,0.56123084,0.49230772,0.4266667,0.18707694,0.18051283,0.25928208,0.35446155,0.47261542,0.6301539,0.56451285,0.5677949,0.67282057,0.65641034,0.61374366,0.98133343,1.1454359,1.142154,1.6672822,1.7263591,1.8281027,1.8149745,1.7165129,1.7394873,1.8313848,2.03159,2.2678976,2.5435898,2.9571285,2.6256413,2.7766156,2.8553848,2.8324106,3.2098465,3.170462,2.8816411,2.5665643,2.281026,1.9167181,1.9331284,1.913436,1.975795,2.169436,2.4648206,2.3860514,2.1858463,1.7887181,1.3128207,1.083077,1.0469744,1.2931283,1.5819489,1.8149745,2.034872,2.1267693,2.1103592,2.097231,2.225231,2.6518977,2.428718,2.3269746,2.3072822,2.3630772,2.4976413,2.0020514,1.9823592,2.0742567,2.0578463,1.847795,5.0674877,5.395693,5.175795,4.893539,4.706462,4.4242053,3.8137438,4.027077,4.5522056,4.9788723,5.0051284,5.077334,4.647385,4.9362054,5.979898,6.6527185,6.688821,7.0826674,7.522462,7.9261546,8.438154,8.720411,8.989539,9.081436,8.89436,8.408616,9.176616,9.488411,10.013539,10.6469755,10.512411,9.90195,10.236719,10.686359,10.817642,10.57477,10.502565,9.714872,9.147078,9.209436,9.796924,9.527796,9.974154,11.388719,13.052719,13.259488,15.530668,15.520822,15.589745,16.436514,17.11918,17.145437,17.818258,19.685745,22.593643,25.69518,22.327797,23.607798,26.994873,28.498053,22.688822,19.98113,19.393642,16.213335,9.875693,3.9680004,1.5885129,0.6071795,0.39384618,0.5874872,1.0994873,2.917744,1.394872,0.06564103,0.04266667,0.029538464,0.006564103,0.0,0.013128206,0.03938462,0.07548718,0.06564103,0.14441027,0.15425642,0.07876924,0.029538464,0.006564103,0.01969231,0.07876924,0.190359,0.33476925,0.45620516,0.38728207,0.30194873,0.3708718,0.761436,0.446359,0.26584616,0.118153855,0.0032820515,0.016410258,0.03938462,0.01969231,0.0,0.0,0.0,0.13456412,0.06564103,0.0,0.0,0.0,0.0,0.04594872,0.059076928,0.04266667,0.09189744,0.17723078,0.098461546,0.32820517,0.7844103,0.80738467,0.7844103,0.6498462,0.8467693,1.1913847,0.88615394,1.7394873,1.9626669,2.0611284,1.9823592,1.1290257,1.6410258,2.2908719,2.5009232,2.0611284,1.1454359,2.7076926,2.5665643,2.5600002,3.0654361,2.989949,3.0752823,3.0424619,3.170462,3.6135387,4.394667,4.9821544,5.356308,6.180103,7.4043083,8.27077,10.345026,11.605334,13.02318,13.761642,11.1983595,11.323078,11.756309,12.780309,13.568001,12.176412,12.297847,11.579078,11.244308,11.631591,12.1928215,10.105436,9.573745,10.518975,12.038565,12.406155,11.930258,12.672001,14.660924,17.847795,22.09477,25.012514,25.458874,22.216208,16.866463,13.778052,14.280207,14.011078,13.11836,12.032001,11.460924,11.483898,12.166565,13.02318,12.911591,10.056206,9.078155,9.8592825,10.374565,10.213744,10.604308,11.910565,12.373334,12.448821,12.2617445,11.628308,11.67754,11.588924,11.250873,10.729027,10.253129,11.474052,12.245335,12.504617,12.754052,14.083283,15.24513,16.439796,16.554668,15.872002,16.068924,14.28677,14.378668,15.0088215,15.202463,14.375385,13.994668,12.849232,12.4685135,12.760616,11.979488,16.617027,16.055796,14.352411,13.679591,14.329437,14.316309,14.375385,14.25395,13.909334,13.51877,13.98154,13.24636,11.946668,10.752001,10.361437,9.764103,10.226872,11.073642,11.851488,12.314258,11.641437,11.52,11.1983595,10.660104,10.633847,10.440206,10.125129,9.632821,9.304616,9.90195,9.7673855,8.067283,6.7314878,6.445949,6.6527185,6.3474874,6.5083084,6.2720003,5.3858466,4.2272825,2.7995899,2.3138463,2.8553848,3.9122055,4.3651285,4.9985647,5.861744,6.436103,6.6428723,6.8496413,6.2523084,5.3431797,4.7524104,4.414359,3.5872824,3.5610259,2.8422565,2.1333334,1.9003079,2.3663592,2.1202054,1.1257436,0.57764107,0.81394875,1.3259488,2.6223593,1.782154,1.6836925,3.757949,7.9819493,3.3050258,1.1651284,0.8533334,1.5327181,2.228513,3.0227695,3.8334363,4.2962055,4.4996924,4.9887185,5.917539,7.276308,8.598975,9.718155,10.742155,9.705027,7.716103,5.792821,4.6572313,4.7294364,5.865026,5.8092313,5.504,5.477744,5.8453336,6.3212314,5.7074876,5.169231,5.0642056,4.9296412,4.7458467,4.3060517,4.086154,4.07959,3.8006158,4.7622566,4.969026,4.059898,3.3214362,5.677949,9.655796,10.246565,10.66995,10.932513,7.8441033,7.3058467,6.7872825,4.585026,1.6738462,1.723077,1.9068719,1.6771283,1.6738462,2.0676925,2.5928206,2.0709746,4.713026,7.3353853,7.79159,4.95918,4.0434875,3.7316926,5.277539,8.264206,10.620719,7.066257,5.7501545,6.5444107,8.021334,7.4469748,7.9097443,9.32759,10.699488,10.965334,8.986258,11.930258,11.008,9.6525135,10.794667,16.8599,14.431181,11.0605135,8.434873,6.882462,5.356308,5.504,9.540924,9.911796,5.7632823,2.9440002,2.481231,3.370667,3.5971284,2.3794873,0.18379489,0.14769232,0.072205134,0.01969231,0.0,0.0,0.0,0.009846155,0.02297436,0.04594872,0.108307704,0.16738462,0.15425642,0.17394873,0.24287182,0.3052308,0.35446155,0.34789747,0.4135385,0.5907693,0.82379496,1.0436924,1.1716924,1.3915899,1.6213335,1.5097437,2.4615386,3.9745643,4.7622566,4.6276927,4.457026,4.2469745,3.9680004,3.6758976,3.629949,4.3027697,3.9122055,3.9614363,3.7710772,3.2886157,3.0818465,2.7536411,2.4320002,2.2613335,2.1825643,1.9364104,1.7657437,1.394872,1.2307693,1.2898463,1.204513,1.4605129,1.8379488,2.0742567,2.172718,2.3794873,3.1737437,3.318154,3.249231,3.4100516,4.2272825,4.9821544,5.540103,6.180103,6.803693,6.9120007,6.422975,5.3694363,4.348718,3.692308,3.4494362,3.5446157,3.7907696,3.9187696,3.8400004,3.6332312,3.5446157,3.7809234,3.879385,3.6562054,3.2032824,3.4231799,3.5971284,3.8596926,4.2535386,4.7294364,4.706462,4.9460516,5.533539,6.294975,6.820103,5.9667697,5.405539,5.2578464,5.4547696,5.720616,5.674667,5.3858466,5.0642056,4.850872,4.8377438,5.179077,5.356308,5.172513,4.663795,4.089436,4.2830772,4.6080003,4.8705645,5.3005133,6.5444107,6.889026,7.394462,7.3452315,6.7577443,6.377026,6.242462,5.927385,6.0685134,6.518154,6.3474874,6.5444107,7.9458466,8.904206,8.953437,8.818872,8.845129,8.786052,8.763078,7.6931286,3.31159,2.5796926,2.284308,2.1398976,2.2121027,2.9440002,3.2853336,2.6322052,2.0808206,1.847795,1.2373334,2.7864618,6.5247183,7.496206,5.549949,5.356308,4.9887185,5.2742567,5.2545643,4.9920006,5.5532312,5.602462,5.9634876,5.2545643,4.1091285,5.156103,5.1200004,6.547693,6.616616,5.0116925,3.9384618,4.1091285,4.6539493,4.0303593,2.6847181,3.0523078,6.0783596,7.0104623,6.678975,6.11118,6.514872,6.550975,6.196513,5.937231,5.720616,4.9296412,3.879385,3.0949745,2.3204105,1.8510771,2.546872,2.3663592,2.3269746,2.5238976,2.878359,3.1573336,3.7316926,4.1780515,4.4406157,4.644103,5.097026,4.890257,4.5522056,4.893539,5.7665644,6.0717955,5.609026,5.674667,6.6592827,7.7390776,6.8955903,7.1909747,7.5191803,8.050873,8.392206,7.5979495,7.427283,7.056411,6.688821,6.4623594,6.439385,6.488616,6.380308,5.8814363,5.287385,5.4482055,5.618872,5.937231,5.546667,4.772103,5.1265645,4.955898,5.7829747,6.11118,6.0947695,7.522462,6.117744,5.346462,4.630975,3.6332312,2.228513,1.8018463,1.273436,0.88287187,0.67610264,0.51856416,0.5677949,0.45292312,0.34789747,0.3708718,0.58092314,0.43323082,0.4135385,0.51856416,0.5973334,0.36758977,0.13456412,0.16738462,0.30194873,0.42338464,0.47261542,0.58420515,0.51856416,0.5316923,0.67938465,0.8402052,0.67938465,0.84348726,1.024,1.214359,1.6771283,1.8379488,1.9035898,1.7394873,1.5327181,1.8018463,1.972513,2.169436,2.3893335,2.4681027,2.0906668,2.2383592,2.6026669,2.553436,2.1366155,2.0742567,2.550154,2.5698464,2.484513,2.4057438,2.1956925,2.3794873,2.2613335,2.3040001,2.5140514,2.4418464,2.4910772,2.2547693,1.7723079,1.2406155,1.020718,0.98461545,1.2242053,1.522872,1.8412309,2.3040001,2.5107694,2.3696413,2.1891284,2.1136413,2.1530259,1.9068719,1.9462565,2.3991797,2.9243078,2.7175386,2.0578463,2.2219489,2.2711797,2.0808206,2.349949,4.893539,5.362872,5.2414365,5.044513,4.893539,4.535795,4.023795,3.69559,3.876103,4.529231,5.284103,5.3103595,4.8082056,4.9460516,5.865026,6.701949,7.781744,8.356103,8.5661545,8.759795,9.488411,9.465437,9.521232,9.468719,9.344001,9.432616,9.754257,9.577026,9.527796,9.793642,10.148104,10.19077,10.026668,10.036513,10.289231,10.561642,10.177642,10.138257,10.128411,10.259693,11.090053,11.172104,12.058257,13.016617,13.761642,14.467283,16.708925,17.798565,19.242668,20.896822,20.965746,21.293951,23.32554,26.725746,30.080002,30.897234,27.106464,29.22667,30.890669,27.690668,17.184822,12.530872,10.676514,8.769642,5.8190775,2.6847181,1.0272821,0.318359,0.118153855,0.16738462,0.36758977,0.7122052,0.52512825,0.56123084,0.85005134,0.702359,0.3052308,0.14112821,0.13784617,0.2100513,0.24615386,0.49887183,0.76800007,0.67282057,0.26912823,0.055794876,0.059076928,0.072205134,0.08861539,0.10502565,0.10502565,0.3052308,0.33476925,0.25928208,0.20348719,0.36102566,0.46276927,0.37415388,0.18707694,0.01969231,0.0032820515,0.006564103,0.0032820515,0.0,0.0,0.0,0.026256412,0.04266667,0.029538464,0.016410258,0.08533334,0.0951795,0.06235898,0.03938462,0.04594872,0.055794876,0.6662565,0.36102566,0.10502565,0.19692309,0.25928208,0.5677949,0.7220513,0.9353847,1.1618463,1.0929232,1.6640002,1.8970258,1.6771283,1.2898463,1.4211283,1.8871796,2.7864618,2.7569232,1.8642052,1.6311796,2.5698464,2.7273848,2.9571285,3.2886157,2.9407182,2.5600002,2.8980515,2.8750772,2.7208207,3.9811285,5.7764106,6.951385,7.3747697,7.702975,9.370257,10.807796,11.831796,12.6063595,13.036308,12.737642,13.095386,12.547283,12.370052,12.534155,11.687386,12.228924,12.048411,12.3766165,12.941129,11.959796,10.174359,8.759795,9.419488,11.703795,13.026463,13.410462,15.0777445,17.224207,19.764515,23.328823,24.809027,23.745644,20.217438,15.776822,13.459693,14.752822,15.488001,14.851283,13.003489,11.080206,10.676514,11.355898,12.068104,11.67754,8.969847,8.372514,8.677744,9.189744,9.521232,9.580308,10.555078,11.35918,11.730052,11.477334,10.492719,11.437949,11.611898,11.418258,11.040821,10.436924,10.633847,11.293539,11.569232,11.513436,12.081232,14.168616,15.202463,15.51754,15.514257,15.638975,15.264822,14.890668,14.854566,15.031796,14.8250265,14.447591,13.161027,12.898462,13.627078,13.331694,17.063385,19.094976,16.032822,10.758565,12.412719,12.242052,12.662155,13.24636,13.466257,12.665437,12.63918,12.645744,12.137027,11.352616,11.313231,10.755282,10.788103,11.191795,11.759591,12.301129,13.154463,13.367796,13.200411,12.612924,11.270565,11.063796,11.099898,10.489437,9.416205,9.147078,8.503796,7.781744,6.987488,6.380308,6.4689236,6.6822567,6.5345645,6.0947695,5.2742567,3.8104618,2.989949,2.6387694,3.0358977,3.9745643,4.7655387,5.910975,6.439385,6.5345645,6.442667,6.4722056,6.3934364,5.2447186,4.276513,3.8006158,3.1967182,3.2886157,2.428718,2.048,2.546872,3.2918978,2.806154,1.6968206,0.93866676,1.0338463,2.034872,4.197744,2.6387694,1.8182565,3.8990772,8.736821,8.54318,3.754667,0.7975385,1.270154,1.9462565,2.7798977,3.6824617,4.4734364,5.2053337,6.173539,7.0531287,8.083693,9.091283,9.846154,10.069334,8.992821,7.325539,5.723898,4.7917953,5.0609236,6.2063594,5.602462,5.1167183,5.464616,6.2227697,6.3376417,5.8092313,5.32677,5.034667,4.5489235,5.293949,4.7950773,4.3060517,5.028103,8.096821,7.000616,5.664821,4.5554876,4.082872,4.6145644,4.2863593,3.7940516,3.6069746,3.623385,3.1934361,5.3005133,8.198565,8.891078,6.436103,1.9429746,1.657436,2.6026669,3.9417439,5.2315903,6.4032826,2.6945643,2.8553848,3.8695388,4.46359,5.1167183,4.4964104,3.2032824,3.5413337,5.687795,7.6898465,9.393231,9.701744,8.021334,5.2447186,3.7710772,4.5489235,5.691077,7.259898,8.982975,10.256411,8.228104,8.94359,9.780514,11.080206,16.141129,14.296617,10.128411,7.7423596,7.9491286,8.247795,6.373744,6.872616,6.9677954,6.373744,7.315693,5.024821,3.7448208,2.7306669,1.7952822,1.3193847,0.40369233,0.08205129,0.009846155,0.0,0.0,0.0,0.009846155,0.02297436,0.032820515,0.04594872,0.16410258,0.19692309,0.18707694,0.17723078,0.20676924,0.3052308,0.318359,0.33805132,0.39384618,0.46933338,0.76800007,0.95835906,1.1257436,1.2340513,1.1454359,1.9790771,2.9636924,3.8038976,4.164923,3.6627696,3.639795,3.6758976,3.5446157,3.498667,4.266667,4.4406157,4.46359,4.141949,3.6463592,3.498667,3.2065644,2.7634873,2.409026,2.2219489,2.1333334,2.0217438,1.9200002,1.7985642,1.6475899,1.4736412,1.4178462,1.6475899,1.8970258,2.0151796,1.9790771,2.5862565,2.8225644,2.9407182,3.2000003,3.8728209,5.3037953,6.226052,6.7774363,7.0137444,6.889026,6.449231,5.477744,4.5423594,4.0533338,4.279795,4.2207184,3.9778464,3.754667,3.7349746,4.096,3.8137438,3.4527183,3.3936412,3.5741541,3.4855387,3.56759,3.757949,3.8859491,3.8990772,3.876103,4.125539,4.535795,5.221744,6.0685134,6.7610264,6.705231,6.416411,6.2063594,6.12759,5.9667697,5.858462,5.7534366,5.4416413,4.9821544,4.716308,4.969026,5.074052,5.0018463,4.7425647,4.2830772,4.578462,4.71959,5.3103595,6.413129,7.571693,7.5421543,7.171283,7.0400004,7.138462,6.87918,6.636308,6.62318,6.9087186,7.4207187,7.936001,8.5202055,9.202872,9.189744,8.51036,8.01477,8.369231,8.503796,9.383386,10.108719,7.9130263,4.5522056,2.7995899,1.7526156,1.1815386,1.5031796,1.4572309,1.273436,2.1989746,3.9844105,4.896821,5.9503593,7.2336416,7.2664623,6.196513,5.796103,5.536821,6.3376417,6.5345645,5.861744,5.4580517,6.73477,6.6625648,5.970052,5.110154,4.266667,6.5739493,7.6996927,8.329846,7.88677,4.5456414,3.2229745,3.2656412,4.6539493,5.8847184,3.9680004,5.579488,5.737026,5.5630774,5.8289237,6.954667,6.377026,5.9602056,5.681231,5.3398976,4.57518,3.817026,3.1507695,2.2908719,1.5458462,1.8051283,2.2646155,2.5862565,2.7667694,2.878359,3.062154,3.5282054,3.5807183,3.5544617,3.7776413,4.571898,5.146257,4.8147697,4.772103,5.169231,5.1331286,5.733744,5.861744,6.547693,7.3714876,6.482052,8.064001,8.480822,8.434873,8.27077,7.965539,7.207385,6.550975,6.180103,6.0816417,6.0356927,5.910975,5.9503593,5.609026,5.093744,5.349744,5.4908724,5.1626673,4.7360005,4.532513,4.857436,5.362872,5.924103,5.9963083,5.658257,5.6320004,5.546667,4.493129,3.761231,3.43959,2.4352822,2.1431797,1.6147693,1.0929232,0.7056411,0.46933338,0.4397949,0.47261542,0.41025645,0.27569234,0.2855385,0.2100513,0.21333335,0.23958977,0.25271797,0.24287182,0.18707694,0.16410258,0.25928208,0.43323082,0.5218462,0.56451285,0.57764107,0.61374366,0.7187693,0.9353847,1.0043077,1.2931283,1.3062565,1.1749744,1.6771283,2.1202054,2.2219489,1.9922053,1.6640002,1.6771283,1.8970258,2.1366155,2.5173335,2.793026,2.3466668,2.3368206,2.5337439,2.6289232,2.6354873,2.868513,2.7864618,2.9243078,2.993231,2.858667,2.5140514,2.6387694,2.6223593,2.5009232,2.359795,2.3433847,2.422154,2.2744617,2.028308,1.7362052,1.3883078,1.5556924,1.6771283,1.7952822,1.9593848,2.2186668,2.1825643,2.1792822,2.2777438,2.4484105,2.5435898,2.5042052,2.4188719,2.6486156,3.0030773,2.7273848,3.2229745,3.4691284,3.511795,3.2361028,2.3630772,3.8990772,4.2535386,4.519385,4.6276927,4.5817437,4.4438977,4.1878977,3.9581542,4.086154,4.601436,5.228308,5.533539,5.1954875,5.159385,5.677949,6.3376417,7.578257,8.621949,9.350565,9.819899,10.272821,10.381129,10.660104,10.561642,10.072617,9.724719,10.315488,10.443488,10.417232,10.364718,10.240001,10.79795,10.492719,10.226872,10.28595,10.368001,10.144821,10.666668,11.099898,11.382154,12.2387705,13.236514,14.201437,15.02195,15.776822,16.738462,17.91672,19.157335,21.051079,23.240208,24.408617,25.944618,29.397335,33.58195,36.93949,37.54339,35.127796,34.79303,33.17826,27.831797,17.191385,12.045129,9.577026,7.712821,5.4941545,3.0884104,1.6246156,0.78769237,0.41682056,0.4955898,1.1454359,1.4211283,0.92553854,0.56451285,0.636718,0.84348726,0.45620516,0.256,0.20348719,0.28225642,0.508718,0.90912825,0.90584624,0.67610264,0.36758977,0.098461546,0.06564103,0.07876924,0.10502565,0.12471796,0.108307704,0.41025645,0.43651286,0.37743592,0.32164106,0.24943592,0.34789747,0.30851284,0.17723078,0.03938462,0.0,0.0,0.0,0.0032820515,0.006564103,0.0,0.006564103,0.029538464,0.04266667,0.068923086,0.16082053,0.13128206,0.055794876,0.01969231,0.026256412,0.026256412,0.3314872,0.34789747,0.29538465,0.256,0.17723078,0.60389745,1.0929232,1.2898463,1.3029745,1.6935385,1.5556924,1.6114873,1.6410258,1.6114873,1.6607181,2.3958976,2.806154,2.6847181,2.1530259,1.6443079,2.1169233,2.1956925,2.484513,2.8816411,2.5895386,2.5009232,2.8389745,2.930872,3.0358977,4.332308,5.5532312,7.1876926,7.8441033,7.9917955,9.954462,11.565949,12.225642,12.914873,13.689437,13.673027,14.050463,13.869949,13.820719,13.856822,13.1872835,13.351386,12.389745,12.507898,13.410462,12.314258,10.824206,9.29477,9.708308,11.992617,14.017642,15.258258,17.427694,19.27877,20.568617,22.052105,21.907694,20.634258,17.811693,14.470565,13.078976,15.205745,16.374155,15.55036,13.069129,10.630565,9.685334,10.180923,10.880001,10.732308,8.907488,8.034462,8.119796,8.674462,9.238976,9.40636,9.760821,10.184206,10.663385,11.090053,11.260718,12.1238985,12.314258,12.245335,11.900719,10.811078,10.341744,10.86359,11.329642,11.533129,12.09436,13.298873,14.316309,14.916924,15.067899,14.930053,14.903796,14.473847,14.28677,14.441027,14.480412,14.073437,13.157744,13.318565,14.368821,14.322873,18.294155,20.17477,16.006565,9.281642,10.916103,11.529847,11.98277,12.675283,13.161027,12.150155,11.664412,11.552821,11.490462,11.349334,11.195078,11.011283,11.155693,11.441232,11.900719,12.78359,14.257232,14.79877,14.867694,14.404924,12.819694,12.435693,12.186257,11.487181,10.28595,9.068309,8.093539,7.680001,7.197539,6.5805135,6.340924,6.3901544,6.426257,6.196513,5.4580517,3.9548721,3.1606157,2.9997952,3.6693337,4.8836927,5.8912826,6.75118,6.9349747,6.7872825,6.416411,5.7107697,6.2851286,5.3398976,4.1846156,3.446154,3.0424619,3.114667,2.9538465,2.809436,3.1540515,4.706462,3.8990772,2.7831798,1.5753847,0.88615394,1.7099489,3.0654361,2.2613335,1.7723079,2.7076926,4.8082056,7.1187696,4.279795,1.5753847,1.1126155,1.8215386,2.5698464,3.6890259,4.781949,5.6943593,6.5247183,7.0826674,7.6209235,8.050873,8.300308,8.310155,7.9261546,7.138462,6.0356927,5.149539,5.4547696,6.3507695,5.6943593,5.2545643,5.737026,6.764308,6.196513,5.7009234,5.3891287,5.3070774,5.4449234,6.0849237,5.9602056,5.546667,5.7468724,7.9261546,5.684513,5.0674877,4.5095387,3.5347695,2.7733335,2.1398976,2.0086155,1.9035898,1.657436,1.3981539,3.0490258,5.7009234,7.4797955,7.174565,4.240411,2.2482052,2.3630772,4.1878977,7.000616,9.754257,5.474462,3.5413337,3.5183592,4.4832826,5.028103,4.647385,4.3716927,4.4734364,5.61559,8.845129,13.147899,11.753027,8.100103,4.926359,4.263385,4.076308,3.8531284,4.8738465,6.8332314,7.837539,7.4010262,8.769642,9.760821,10.512411,13.5089245,12.954257,8.861539,6.521436,7.243488,8.3593855,5.737026,5.428513,5.737026,6.242462,7.821129,6.2096415,5.2545643,4.4274874,3.9154875,4.604718,1.5885129,0.35446155,0.02297436,0.006564103,0.0,0.0,0.0032820515,0.009846155,0.013128206,0.02297436,0.08205129,0.15753847,0.190359,0.17066668,0.128,0.2231795,0.25928208,0.28225642,0.30194873,0.30851284,0.6826667,0.85005134,0.9616411,1.0371283,0.97805136,1.5360001,2.2153847,3.0752823,3.757949,3.508513,3.6004105,3.820308,3.9417439,4.007385,4.338872,4.450462,4.5095387,4.3651285,4.1058464,4.059898,3.8367183,3.3280003,2.9210258,2.737231,2.6223593,2.3466668,2.2547693,2.2186668,2.1333334,1.9068719,1.6836925,1.7690258,1.8773335,1.8871796,1.8412309,2.300718,2.6584618,2.930872,3.259077,3.9220517,5.182359,6.0750775,6.6461544,6.997334,7.276308,6.7610264,6.009436,5.211898,4.588308,4.394667,4.276513,3.8137438,3.4756925,3.5216413,4.0008206,3.9876926,3.8695388,3.9122055,4.1222568,4.269949,4.1485133,4.066462,3.9614363,3.82359,3.7087183,3.9089234,4.453744,5.1331286,5.733744,6.048821,6.173539,6.009436,5.914257,6.009436,6.173539,6.124308,6.173539,5.9503593,5.3727183,4.647385,4.6900516,4.9296412,4.854154,4.457026,4.2502565,4.4077954,4.8311796,5.7796926,6.921847,7.3616414,7.200821,7.4010262,7.5881033,7.5979495,7.460103,7.318975,7.315693,7.512616,7.8834877,8.329846,8.992821,9.373539,9.18318,8.6580515,8.562873,8.960001,9.222565,10.066052,10.692924,8.815591,3.8695388,2.1431797,1.3522053,0.8533334,1.6311796,2.3401027,2.7798977,3.7185643,5.0149746,5.612308,7.00718,7.4174366,7.138462,6.5903597,6.298257,6.747898,7.315693,7.072821,6.163693,5.8256416,5.976616,6.0685134,6.189949,6.1078978,5.287385,6.173539,6.6822567,7.4765134,7.64718,4.709744,2.7175386,2.7142565,3.9286156,4.9099493,3.508513,4.562052,4.768821,5.024821,5.6385646,6.314667,5.602462,5.1856413,5.0182567,4.8705645,4.3027697,3.3476925,2.665026,1.9331284,1.3784616,1.7723079,2.0742567,2.4549747,2.7437952,2.9636924,3.3214362,3.4527183,3.4560003,3.2623591,3.1277952,3.626667,4.269949,4.240411,4.3290257,4.6933336,4.844308,5.85518,5.9930263,6.3245134,6.925129,6.8627696,7.499488,7.584821,7.64718,7.8736415,8.093539,7.1548724,6.180103,5.4941545,5.2480006,5.395693,5.533539,5.61559,5.402257,5.07077,5.1987696,5.097026,5.0543594,4.886975,4.673641,4.7622566,5.142975,5.786257,5.756718,5.1922054,5.3136415,5.3366156,4.854154,4.1813335,3.515077,2.92759,2.3335385,1.7362052,1.2438976,0.90256417,0.6695385,0.51856416,0.4955898,0.43651286,0.36102566,0.47917953,0.46933338,0.42994875,0.3249231,0.19692309,0.15753847,0.20348719,0.29538465,0.3511795,0.3708718,0.43323082,0.5021539,0.57764107,0.7089231,0.88943595,1.0699488,1.0535386,1.204513,1.3915899,1.5360001,1.6311796,1.7952822,2.0151796,1.913436,1.5360001,1.3653334,1.8740515,2.1497438,2.425436,2.5961027,2.2186668,2.2711797,2.297436,2.2908719,2.3466668,2.6453335,2.5796926,2.7175386,2.6584618,2.3860514,2.2547693,2.4910772,2.5173335,2.3729234,2.1956925,2.2449234,2.4188719,2.4155898,2.2580514,1.9889232,1.654154,1.9035898,2.1267693,2.0775387,1.8838975,2.0676925,2.103795,2.2646155,2.4155898,2.5173335,2.6486156,2.7798977,2.7864618,2.8488207,2.9505644,2.878359,3.131077,3.1409233,3.3312824,3.6069746,3.3641028,3.3936412,3.5872824,3.8695388,4.086154,4.1747694,4.1682053,4.2174363,4.322462,4.6145644,5.0018463,5.149539,5.549949,5.5204105,5.4153852,5.5302567,6.11118,7.269744,8.516924,9.711591,10.614155,10.86359,11.073642,11.2672825,11.122872,10.774975,10.801231,11.208206,11.300103,11.392001,11.411694,10.893129,11.434668,11.030975,10.594462,10.55836,10.843898,10.883283,11.588924,12.133744,12.435693,13.154463,14.575591,15.711181,16.823795,17.742771,17.851078,19.18031,20.62113,22.432823,24.513643,26.397541,27.776003,31.399387,35.58072,38.915283,40.2839,38.485336,37.316925,34.310566,28.228926,19.06872,13.8075905,10.564924,8.152616,5.933949,3.820308,2.3302567,1.3259488,0.81394875,0.8992821,1.8051283,2.5731285,1.7296412,0.702359,0.3052308,0.7253334,0.4660513,0.28882053,0.20348719,0.23958977,0.43651286,0.77456415,0.7450257,0.6170257,0.46933338,0.16410258,0.108307704,0.0951795,0.108307704,0.118153855,0.108307704,0.33805132,0.41682056,0.48246157,0.53825647,0.47589746,0.39384618,0.27569234,0.14441027,0.03938462,0.0,0.0,0.0,0.0032820515,0.006564103,0.0,0.06564103,0.052512825,0.03938462,0.068923086,0.14441027,0.098461546,0.04594872,0.09189744,0.17066668,0.03938462,0.02297436,0.17723078,0.37415388,0.6071795,0.9944616,0.8598975,1.086359,1.2570257,1.3226668,1.6213335,1.8642052,1.7427694,1.7788719,1.9889232,1.8806155,2.4155898,2.3368206,2.2153847,2.1366155,1.6869745,1.8445129,1.9790771,2.231795,2.5206156,2.546872,2.5993848,2.7667694,3.2229745,4.023795,5.110154,5.4514875,7.5585647,8.661334,8.661334,10.131693,11.1294365,11.533129,12.018872,12.672001,13.013334,13.548308,13.6697445,14.116103,14.670771,14.152206,14.227694,12.809847,12.304411,12.911591,12.6063595,11.477334,10.427077,10.755282,12.524308,14.549335,16.577642,18.41231,19.272207,19.104822,18.586258,17.460514,16.406975,14.582155,12.514462,12.091078,14.516514,15.881847,15.369847,13.161027,10.427077,8.838565,9.238976,9.862565,9.875693,9.360411,8.027898,8.018052,8.704,9.442462,9.563898,9.705027,9.777231,10.066052,10.6469755,11.388719,12.018872,12.452104,12.678565,12.442257,11.241027,10.84718,11.178667,11.483898,11.766154,12.796719,13.197129,13.879796,14.483693,14.759386,14.555899,14.191591,13.725539,13.6008215,13.843694,14.060308,13.568001,12.950975,13.351386,14.434463,14.388514,17.112617,18.586258,14.933334,8.950154,10.105436,11.703795,12.153437,12.793437,13.466257,12.514462,11.844924,11.093334,10.8307705,10.975181,10.804514,10.699488,11.067078,11.339488,11.720206,13.203693,14.841437,15.629129,15.875283,15.501129,14.04718,13.492514,13.108514,12.484924,11.30995,9.347282,8.352821,7.890052,7.568411,7.145026,6.5017443,6.245744,6.363898,6.373744,5.8945646,4.650667,3.9286156,3.9253337,4.7392826,6.045539,7.1122055,7.351795,7.253334,7.076103,6.6527185,5.3694363,6.11118,5.431795,4.269949,3.3017437,2.937436,2.9801028,3.31159,3.3411283,3.5938463,5.7009234,5.579488,4.9952826,3.826872,2.425436,1.6246156,2.3401027,2.1792822,1.8412309,1.6344616,1.4933335,4.1124105,4.164923,2.609231,1.0469744,1.723077,2.359795,3.5544617,4.8049235,5.792821,6.38359,6.688821,6.7216415,6.5936418,6.567385,7.0400004,7.351795,7.1483083,6.5280004,5.927385,6.1308722,6.419693,5.8125134,5.5302567,6.0061545,6.8955903,6.0717955,5.5991797,5.3694363,5.395693,5.8420515,6.196513,6.3540516,6.633026,7.0892315,7.4863596,5.0477953,5.0543594,5.1167183,4.2174363,2.7175386,2.044718,2.0742567,2.1497438,2.1398976,2.422154,2.809436,3.4264617,4.2502565,5.139693,5.8420515,4.972308,3.9056413,4.7983594,7.962257,11.877745,9.429334,6.436103,5.5762057,6.442667,5.5105643,6.370462,7.939283,8.008205,7.2172313,9.065026,13.184001,11.602052,8.326565,6.052103,6.180103,5.76,4.7294364,4.965744,6.452513,7.276308,8.241231,8.641642,9.242257,10.240001,11.260718,10.35159,7.762052,6.3245134,6.7183595,7.466667,4.5029745,3.9220517,4.1156926,4.772103,6.8463597,8.533334,7.318975,5.1626673,4.0533338,6.0160003,2.546872,0.7778462,0.118153855,0.026256412,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.02297436,0.08205129,0.13784617,0.15097436,0.10502565,0.16410258,0.19364104,0.23630771,0.28225642,0.26584616,0.5481026,0.7089231,0.8402052,0.9485129,0.9353847,1.1749744,1.5688206,2.3105643,3.1507695,3.373949,3.5741541,3.9351797,4.273231,4.4340515,4.2962055,4.312616,4.5095387,4.5390773,4.3716927,4.2830772,4.164923,3.623385,3.2131286,3.0687182,2.9210258,2.412308,2.2646155,2.3335385,2.4320002,2.3335385,2.0676925,2.044718,1.9954873,1.8740515,1.8576412,2.294154,2.6945643,3.0260515,3.4067695,4.0992823,5.1889234,6.0291286,6.5706673,7.00718,7.762052,7.0925136,6.4065647,5.658257,4.890257,4.240411,3.9811285,3.498667,3.1277952,3.0916924,3.4756925,3.7842054,4.128821,4.352,4.453744,4.604718,4.338872,4.240411,4.2240005,4.2469745,4.2994876,4.6178465,5.1856413,5.5926156,5.733744,5.8092313,6.11118,6.055385,6.0356927,6.2129235,6.521436,6.4295387,6.49518,6.3245134,5.799385,5.093744,4.969026,4.95918,4.6572313,4.1485133,4.020513,4.086154,4.900103,6.242462,7.282872,6.5739493,6.7183595,7.6176414,8.116513,7.936001,7.686565,7.640616,7.702975,7.90318,8.146052,8.234667,8.641642,8.992821,9.127385,9.124104,9.32759,9.570462,9.567181,9.816616,9.412924,6.038975,2.3860514,1.591795,1.3981539,1.2373334,2.2022567,3.1934361,4.07959,4.841026,5.405539,5.674667,7.0104623,7.4075904,7.3485136,7.200821,7.177847,8.021334,7.9163084,7.020308,5.930667,5.684513,4.9526157,5.5072823,6.498462,7.138462,6.705231,6.925129,7.177847,7.1089234,6.294975,4.2207184,3.5446157,3.308308,3.5971284,3.9187696,3.1967182,3.9187696,4.2896414,4.7622566,5.3103595,5.4547696,5.034667,4.4701543,4.3060517,4.4077954,3.948308,2.9210258,2.2153847,1.6738462,1.3981539,1.7493335,2.1267693,2.4516926,2.737231,3.0424619,3.4494362,3.308308,3.4297438,3.242667,2.8225644,2.8750772,3.3050258,3.5577438,3.9844105,4.5489235,4.824616,5.6385646,5.6418467,5.9536414,6.7971287,7.522462,7.0990777,6.4689236,6.3606157,6.872616,7.460103,6.5870776,5.661539,4.9099493,4.5390773,4.7425647,5.0149746,5.024821,5.0018463,5.0904617,5.3431797,5.156103,5.284103,5.284103,5.100308,5.074052,5.2480006,5.618872,5.5072823,5.1331286,5.612308,5.3694363,5.2742567,4.7425647,3.826872,3.242667,2.4746668,1.8445129,1.4080001,1.1290257,0.86974365,0.67938465,0.56123084,0.4660513,0.43323082,0.5940513,0.60389745,0.5513847,0.40369233,0.2231795,0.14112821,0.256,0.37415388,0.40369233,0.36758977,0.40369233,0.49887183,0.6235898,0.8369231,1.083077,1.1618463,1.2274873,1.3193847,1.5983591,1.8642052,1.5524104,1.5031796,1.6607181,1.7132308,1.5589745,1.3029745,1.6968206,1.9856411,2.2022567,2.2711797,2.0217438,2.1858463,2.231795,2.1989746,2.166154,2.2744617,2.1989746,2.3040001,2.3368206,2.2514873,2.1989746,2.546872,2.556718,2.3860514,2.1825643,2.0939488,2.2186668,2.228513,2.1234872,1.9626669,1.8674873,2.0644104,2.2022567,2.0742567,1.8543591,2.100513,2.1825643,2.4681027,2.678154,2.740513,2.789744,2.937436,3.0490258,3.1671798,3.242667,3.1474874,3.3017437,3.3542566,3.6890259,4.1780515,4.194462,3.5840003,3.7152824,3.6496413,3.7382567,3.9417439,3.8104618,4.161641,4.5095387,4.9854364,5.3924108,5.211898,5.477744,5.7140517,5.5532312,5.3234878,6.042257,7.1909747,8.3134365,9.5606165,10.65354,10.886565,11.224616,11.057232,10.883283,11.172104,12.36677,12.225642,11.805539,11.828514,12.130463,11.67754,11.759591,11.234463,10.827488,10.994873,11.907283,12.228924,12.95754,13.377642,13.4859495,13.984821,15.186052,16.699078,18.182566,18.921026,17.811693,20.49313,22.419695,24.047592,25.632822,27.231182,27.789131,30.585438,33.920002,36.955902,39.69313,38.386875,39.03344,36.873848,30.536207,22.048822,16.144411,12.133744,9.26195,7.0400004,5.221744,3.3542566,2.048,1.3259488,1.2373334,1.8642052,3.0424619,2.284308,1.1158975,0.43323082,0.49887183,0.3446154,0.2231795,0.16410258,0.15753847,0.14769232,0.27897438,0.4594872,0.54482055,0.4594872,0.18707694,0.14769232,0.10502565,0.08205129,0.068923086,0.04594872,0.07876924,0.256,0.44964105,0.6104616,0.7450257,0.51856416,0.27897438,0.10502565,0.02297436,0.0,0.0,0.0,0.0,0.0,0.0,0.118153855,0.072205134,0.01969231,0.02297436,0.049230773,0.032820515,0.03938462,0.256,0.46933338,0.06235898,0.013128206,0.0032820515,0.24943592,0.84348726,1.7624617,0.97805136,0.7975385,1.1126155,1.4966155,1.1946667,2.425436,2.2055387,1.9823592,2.15959,2.0873847,1.9692309,1.8313848,1.7690258,1.7985642,1.8576412,1.9659488,2.297436,2.481231,2.5074873,2.7503593,2.8389745,2.8717952,3.5183592,4.7622566,5.910975,6.11118,8.3593855,9.642668,9.498257,10.020103,10.010257,10.394258,10.568206,10.748719,11.959796,12.452104,12.314258,12.859077,13.922462,13.853539,14.326155,13.39077,12.3995905,12.100924,12.635899,11.907283,11.618463,11.9860525,13.046155,14.677335,16.708925,17.460514,16.961643,15.55036,13.889642,12.875488,12.25518,11.372309,10.463181,10.65354,12.898462,14.424617,14.5952835,13.144616,10.161232,8.3593855,8.940309,9.383386,9.120821,9.547488,8.146052,8.27077,9.012513,9.642668,9.593436,9.875693,10.069334,10.171078,10.292514,10.676514,11.149129,11.730052,12.182976,12.166565,11.23118,11.37559,11.703795,11.798975,12.025436,13.50236,13.732103,13.748514,13.883078,14.129231,14.145642,13.4629755,12.937847,12.868924,13.1872835,13.4400015,12.911591,12.498053,12.980514,13.935591,13.748514,14.628103,16.134565,13.961847,9.842873,11.526565,12.452104,12.826258,13.51877,14.260514,13.633642,13.161027,11.785847,10.866873,10.729027,10.683078,10.233437,10.610872,10.840616,11.149129,12.983796,14.729847,15.786668,16.187078,15.908104,14.874257,14.132514,13.820719,13.361232,12.235488,10.003693,9.26195,8.569437,8.149334,7.821129,6.9842057,6.6592827,6.5312824,6.5969234,6.564103,5.8453336,5.3825645,5.5105643,6.2096415,7.213949,8.004924,7.650462,7.3025646,7.207385,7.0104623,5.7632823,6.0685134,5.467898,4.325744,3.1934361,2.789744,2.8324106,3.1967182,3.387077,3.8071797,5.7534366,6.885744,7.325539,6.688821,4.9788723,2.5600002,2.7241027,2.425436,1.8281027,1.1552821,0.67938465,2.038154,3.623385,3.0096412,0.98461545,1.5327181,2.162872,3.1737437,4.3716927,5.431795,5.8945646,6.193231,6.0619493,5.7764106,5.8486156,7.059693,7.7718983,7.5946674,7.1647186,6.928411,7.131898,6.744616,6.0258465,5.7731285,6.121026,6.5247183,6.091488,5.7435904,5.3694363,5.146257,5.549949,5.353026,5.612308,7.1187696,8.841846,7.9195905,6.2916927,6.294975,6.8397956,6.7577443,4.8114877,2.8750772,2.4385643,2.9111798,4.0402055,5.8912826,5.540103,3.945026,2.5009232,2.5665643,5.4416413,8.434873,7.0498466,6.4557953,8.546462,11.979488,12.327386,9.655796,8.385642,8.55959,5.861744,7.9097443,11.201642,11.789129,9.232411,6.5805135,9.275078,10.056206,9.019077,7.433847,7.7390776,8.237949,7.3780518,7.020308,7.7981544,9.097847,10.003693,8.87795,8.822155,10.075898,10.039796,7.8145647,6.9120007,6.6625648,6.6100516,6.51159,3.511795,2.8291285,3.3280003,4.7294364,7.6012316,12.07795,9.573745,4.785231,2.1366155,5.7764106,2.793026,0.99774367,0.19692309,0.03938462,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.026256412,0.059076928,0.098461546,0.1148718,0.15097436,0.14769232,0.20348719,0.28882053,0.256,0.33805132,0.512,0.7515898,0.95835906,0.9682052,0.92225647,1.0765129,1.6049232,2.3827693,2.9833848,3.3542566,3.698872,4.010667,4.1846156,3.9942567,4.076308,4.345436,4.3618464,4.096,3.9187696,4.0369234,3.5478978,3.1606157,3.0523078,2.8455386,2.1924105,2.041436,2.225231,2.5206156,2.6354873,2.4615386,2.3794873,2.228513,2.0512822,2.097231,2.6387694,3.0030773,3.2984617,3.6529233,4.2174363,5.2611284,6.2490263,6.885744,7.312411,8.1066675,7.2237954,6.409847,5.648411,4.900103,4.0992823,3.5577438,3.1081028,2.733949,2.5600002,2.8455386,3.2098465,3.817026,4.2338467,4.3552823,4.414359,4.125539,4.20759,4.4767184,4.844308,5.3431797,6.0028725,6.4754877,6.485334,6.2129235,6.2884107,6.892308,7.1581545,7.210667,7.174565,7.174565,6.892308,6.7840004,6.567385,6.245744,6.11118,5.8847184,5.2611284,4.6211286,4.161641,3.876103,3.9417439,4.850872,6.416411,7.4469748,5.7468724,6.262154,7.240206,7.781744,7.650462,7.2861543,7.450257,7.9491286,8.333129,8.388924,8.146052,8.320001,8.730257,9.216001,9.567181,9.524513,9.5146675,9.117539,8.612103,7.0465646,2.2416413,1.6410258,2.0578463,2.3204105,2.300718,2.9046156,3.3903592,4.2830772,5.0674877,5.5729237,5.9634876,6.626462,7.1647186,7.5454364,7.834257,8.155898,8.887795,7.906462,6.2588725,4.9526157,4.9329233,4.378257,5.3398976,6.8430777,7.893334,7.4863596,8.490667,8.851693,7.529026,5.1626673,4.076308,5.602462,4.7294364,4.056616,4.135385,3.4494362,3.9712822,4.2896414,4.578462,4.824616,4.8147697,4.8147697,4.069744,3.7940516,4.0041027,3.5216413,2.7503593,2.1070771,1.7001027,1.5589745,1.6344616,2.3794873,2.6978464,2.8914874,3.117949,3.3772311,3.1245131,3.3050258,3.2328207,2.8258464,2.609231,2.9013336,3.2918978,3.9122055,4.5817437,4.8049235,5.2480006,5.1167183,5.6287184,6.8365135,7.6012316,7.062975,6.058667,5.5696416,5.8157954,6.2687182,5.661539,5.179077,4.7228723,4.397949,4.5029745,4.6276927,4.4800005,4.6178465,5.1298466,5.664821,5.687795,5.661539,5.618872,5.609026,5.691077,5.8256416,5.622154,5.3858466,5.3924108,5.8912826,5.540103,5.3858466,5.044513,4.3651285,3.4133337,2.665026,1.9987694,1.5556924,1.2800001,0.94523084,0.7811283,0.62030774,0.50543594,0.4660513,0.54482055,0.5021539,0.44307697,0.3446154,0.23302566,0.18379489,0.3117949,0.36102566,0.39384618,0.4266667,0.4266667,0.51856416,0.6695385,0.9156924,1.1585642,1.1520001,1.4605129,1.6902566,1.9265642,2.0020514,1.4966155,1.4966155,1.4867693,1.6213335,1.7755898,1.5589745,1.463795,1.7132308,1.9495386,2.0217438,1.972513,2.172718,2.3762052,2.4549747,2.3630772,2.1530259,1.8576412,1.9889232,2.3630772,2.6880002,2.556718,2.9440002,2.9440002,2.7241027,2.3991797,2.041436,1.9528207,1.8445129,1.7657437,1.785436,1.9987694,2.100513,2.0118976,1.9331284,2.0184617,2.359795,2.3991797,2.7503593,3.0326157,3.0752823,2.9111798,3.0227695,3.1638978,3.4625645,3.7218463,3.4034874,4.056616,4.4012313,4.7491283,5.0018463,4.6276927,3.570872,3.8400004,3.7054362,3.7907696,4.007385,3.5544617,4.240411,4.46359,4.8114877,5.3103595,5.431795,5.737026,5.924103,5.412103,4.7491283,5.61559,6.810257,7.9261546,8.864821,9.468719,9.504821,10.568206,10.594462,10.528821,10.998155,12.3306675,12.596514,12.068104,11.766154,11.851488,11.641437,11.362462,10.906258,10.955488,11.638155,12.544001,13.371078,14.578873,15.041642,14.815181,15.120412,16.183796,18.087385,19.216412,19.193438,18.875078,21.828924,23.978668,25.790361,27.38872,28.550566,31.343592,34.113644,35.682465,37.22831,42.28267,45.174156,47.38954,45.59426,38.770874,28.212515,20.41436,16.81395,14.28677,11.58236,9.324308,6.186667,3.882667,2.4648206,1.8904617,1.9987694,3.062154,2.162872,1.4506668,1.2668719,0.16738462,0.0951795,0.0951795,0.14441027,0.21989745,0.3052308,0.28225642,0.2100513,0.108307704,0.016410258,0.016410258,0.016410258,0.006564103,0.02297436,0.059076928,0.04594872,0.068923086,0.17723078,0.22646156,0.24287182,0.4266667,0.26912823,0.128,0.04266667,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.013128206,0.0,0.02297436,0.03938462,0.38728207,0.7187693,0.0,0.013128206,0.02297436,0.26912823,0.5284103,0.13784617,0.28225642,1.079795,2.0676925,2.6617439,2.1366155,2.4648206,2.1825643,2.225231,2.5764105,2.2580514,1.8674873,2.2186668,2.2678976,1.8838975,1.847795,2.4320002,2.605949,2.7109745,2.7602053,2.4582565,3.4822567,3.620103,3.4560003,3.9220517,6.301539,7.6931286,8.700719,9.353847,9.688616,9.750975,10.725744,11.329642,11.792411,12.484924,13.899488,13.144616,12.58995,12.265027,12.386462,13.351386,14.011078,14.102976,13.37436,12.416001,12.635899,12.219078,12.5374365,12.87877,13.443283,15.333745,15.248411,14.762668,13.423591,11.421539,9.567181,9.82318,10.289231,10.295795,9.849437,9.6295395,11.923694,13.61395,13.643488,11.835078,8.881231,8.356103,9.55077,9.764103,8.690872,8.421744,8.021334,8.851693,9.170052,8.789334,9.094564,9.081436,9.993847,10.617436,10.765129,11.277129,11.286975,10.788103,10.758565,10.962052,9.947898,10.144821,11.126155,12.120616,12.980514,14.17518,14.089848,13.538463,12.694975,12.032001,12.314258,12.422565,12.09436,11.930258,11.963078,11.657847,11.352616,11.595488,12.566976,13.636924,13.380924,16.262566,17.11918,14.739694,12.42913,18.021746,13.61395,13.482668,14.434463,14.851283,14.693745,14.7790785,13.538463,12.20595,11.405129,11.122872,10.282667,10.226872,10.341744,10.59118,11.52,13.705847,15.304206,16.055796,16.180513,16.387283,15.2155905,14.519796,13.994668,13.164309,11.382154,10.94236,9.908514,8.815591,8.011488,7.643898,7.6701546,7.1154876,7.0367184,7.466667,7.430565,7.076103,7.4010262,8.018052,8.493949,8.346257,7.6996927,7.017026,6.9054365,7.1548724,6.7150774,6.3967185,5.5302567,4.1452312,2.802872,2.5928206,2.605949,3.1048207,3.501949,3.82359,4.716308,5.7403083,7.141744,6.8233852,5.1232824,4.8049235,2.5009232,1.5097437,1.0404103,0.764718,0.8402052,0.8402052,1.6443079,1.5885129,0.78769237,1.1290257,2.03159,2.6420515,3.5577438,4.634257,4.9887185,5.5630774,6.183385,6.5969234,7.069539,8.375795,9.353847,8.956718,8.077128,7.584821,8.316719,7.899898,6.7249236,6.0291286,6.0619493,6.0717955,6.3540516,6.3967185,5.5893335,4.71959,5.9667697,3.9023592,4.4865646,7.2631803,9.724719,7.3091288,7.578257,8.257642,9.412924,9.865847,7.2172313,3.5413337,2.8160002,4.7458467,8.1755905,11.093334,10.896411,8.247795,4.916513,2.6584618,3.2196925,8.5661545,8.51036,8.139488,9.025641,9.232411,10.683078,9.783795,9.330873,8.707283,3.8596926,3.895795,8.054154,11.191795,9.974154,2.868513,6.1407185,9.035488,9.298052,7.716103,8.116513,9.53436,8.989539,8.582564,8.851693,8.805744,12.406155,11.969642,10.023385,8.513641,8.818872,8.0377445,6.0028725,5.024821,5.4383593,5.586052,3.5216413,4.397949,7.899898,12.2387705,14.145642,14.500104,11.858052,6.5247183,2.674872,8.375795,2.4943593,0.41682056,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.032820515,0.04594872,0.055794876,0.09189744,0.16410258,0.16410258,0.19692309,0.24287182,0.18379489,0.256,0.37415388,0.7122052,1.1027694,1.0535386,0.7844103,1.020718,1.3915899,1.8018463,2.412308,3.0949745,2.937436,2.6978464,2.809436,3.370667,3.495385,3.370667,3.1113849,2.8947694,2.930872,3.626667,3.3969233,3.1277952,3.0030773,2.5009232,1.9790771,1.9003079,2.2186668,2.6617439,2.7470772,2.8455386,2.7503593,2.553436,2.4615386,2.793026,3.501949,3.8695388,4.076308,4.194462,4.1813335,4.71959,6.0980515,7.4469748,8.201847,8.116513,6.9809237,6.038975,5.405539,4.903385,4.073026,3.18359,2.5928206,2.284308,2.2711797,2.6256413,2.550154,3.0260515,3.692308,4.2535386,4.4865646,4.315898,4.0992823,4.164923,4.781949,6.1505647,7.003898,7.328821,7.259898,7.0104623,6.8496413,7.522462,8.625232,9.058462,8.674462,8.283898,7.8080006,7.3058467,6.951385,6.9152827,7.3550773,6.9645133,6.0061545,5.2545643,4.8640003,4.3651285,4.3027697,4.571898,5.756718,6.8562055,5.293949,5.330052,5.5597954,5.7731285,5.930667,6.1505647,7.076103,8.681026,9.281642,8.720411,8.375795,9.061745,9.3768215,9.609847,9.596719,8.743385,8.4512825,8.421744,7.384616,5.172513,2.7306669,2.8422565,4.096,4.5095387,3.9680004,4.210872,4.4438977,4.6834874,5.21518,5.8518977,5.9503593,6.1472826,6.2851286,6.7872825,7.634052,8.375795,8.999385,7.1056414,4.394667,2.7700515,4.332308,4.0533338,4.9887185,6.547693,7.719385,7.0957956,7.194257,7.3649235,6.2851286,4.906667,6.4689236,7.752206,6.038975,4.3684106,3.826872,3.570872,4.4734364,4.5456414,4.4045134,4.3651285,4.4242053,4.414359,3.889231,3.6332312,3.6562054,3.2032824,2.8127182,2.3696413,1.9462565,1.719795,1.9528207,2.3926156,2.9144619,3.2065644,3.2820516,3.4625645,3.170462,3.0687182,3.0260515,2.9505644,2.793026,3.3280003,3.764513,4.059898,4.2830772,4.6244106,5.3694363,5.435077,5.7829747,6.3212314,5.904411,6.186667,6.557539,6.5772314,6.1341543,5.4613338,5.366154,5.35959,5.2545643,5.1265645,5.3103595,5.2381544,4.926359,4.919795,5.2742567,5.5532312,6.0192823,6.1538467,6.012718,5.861744,6.180103,6.2162056,5.9503593,5.546667,5.3398976,5.8289237,5.792821,5.5893335,5.4514875,5.1364107,3.95159,2.986667,2.1136413,1.5721027,1.2865642,0.88615394,0.64000005,0.54482055,0.54482055,0.60389745,0.702359,0.54482055,0.32820517,0.23302566,0.256,0.24287182,0.256,0.37743592,0.46933338,0.45292312,0.3052308,0.36758977,0.54482055,0.761436,0.9353847,1.0075898,1.2274873,1.6738462,2.0545642,2.0939488,1.5556924,1.6049232,1.7624617,1.8740515,1.8773335,1.8149745,1.585231,1.6804104,1.7657437,1.8248206,2.166154,2.300718,2.4713848,2.612513,2.5895386,2.2121027,1.723077,2.03159,2.5337439,2.8750772,2.9604106,3.3378465,3.498667,3.2951798,2.8356924,2.4582565,2.162872,1.9889232,1.8379488,1.7558975,1.9364104,2.097231,2.1530259,2.2350771,2.409026,2.7011285,2.7995899,3.2164104,3.3378465,3.0227695,2.5928206,2.8980515,3.0293336,3.2918978,3.5872824,3.4034874,4.525949,4.7524104,4.893539,5.1987696,5.3694363,3.9122055,3.7907696,3.7185643,3.7316926,3.7152824,3.4198978,4.066462,4.4340515,4.8311796,5.2447186,5.346462,5.602462,5.930667,5.8978467,5.6976414,6.163693,7.312411,8.815591,9.298052,8.789334,8.749949,9.724719,10.131693,10.489437,11.001437,11.559385,12.36677,12.5374365,12.36677,12.196103,12.3995905,11.776001,11.946668,12.176412,12.084514,11.651283,13.095386,14.257232,15.366566,16.387283,17.014154,17.99877,19.75795,21.300514,22.626463,24.710566,27.605335,30.083284,32.7319,35.679184,38.606773,41.314465,42.10544,42.663387,45.9159,56.02462,57.951183,56.175594,50.799595,42.689644,33.4999,27.057232,22.436104,19.213129,16.377438,12.314258,8.825437,6.1472826,4.073026,2.5271797,1.5721027,1.8248206,1.2209232,0.69907695,0.574359,0.55794877,0.27897438,0.14769232,0.16410258,0.23958977,0.20676924,0.1148718,0.06564103,0.032820515,0.016410258,0.016410258,0.006564103,0.0,0.009846155,0.036102567,0.08205129,0.108307704,0.0951795,0.07548718,0.072205134,0.098461546,0.10502565,0.14441027,0.128,0.055794876,0.02297436,0.013128206,0.01969231,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0,0.0032820515,0.006564103,0.07876924,0.14441027,0.0,0.0032820515,0.032820515,0.36102566,0.8008206,0.7220513,1.0272821,1.467077,1.8642052,2.0611284,1.9167181,2.9604106,2.4418464,2.353231,2.8717952,2.3696413,2.484513,2.3762052,1.9462565,1.5688206,2.0775387,2.225231,2.1924105,2.3269746,2.6387694,2.809436,2.809436,3.1081028,3.511795,3.95159,4.4964104,5.0084105,5.2742567,7.24677,10.453334,12.009027,12.320822,12.389745,12.166565,12.491488,15.110565,15.182771,14.28677,14.342566,15.120412,14.217847,13.384206,12.757335,12.3766165,12.035283,11.2672825,12.297847,13.10195,13.75836,14.198155,14.188309,13.965129,13.39077,12.022155,9.96759,7.906462,8.848411,9.8363085,10.41395,10.276103,9.275078,11.139283,13.046155,13.459693,11.999181,9.40636,9.025641,9.416205,8.717129,7.259898,7.568411,7.8112826,8.3364105,8.6580515,8.766359,9.130668,9.498257,9.77395,9.905231,10.089026,10.788103,11.004719,10.643693,10.614155,10.929232,10.71918,11.07036,11.372309,11.963078,12.626052,12.599796,13.5318985,12.996924,12.196103,11.785847,11.910565,12.6063595,12.248616,11.116308,9.862565,9.498257,10.404103,11.339488,12.905026,14.647796,15.05477,18.71754,21.973335,18.944002,11.579078,9.672206,12.199386,13.302155,14.283488,15.366566,15.694771,16.072206,15.117129,13.558155,12.1468725,11.661129,11.237744,10.745437,10.587898,10.994873,12.022155,14.500104,15.337027,15.780104,16.315079,16.66954,15.983591,15.478155,15.327181,15.172924,14.093129,11.963078,10.325335,9.314463,8.710565,7.9130263,7.821129,7.581539,7.8834877,8.815591,9.872411,9.058462,8.621949,8.264206,8.123077,8.786052,8.441437,7.6931286,7.643898,8.257642,8.385642,7.4240007,6.0685134,4.3651285,2.8521028,2.556718,2.8422565,3.0129232,3.0523078,3.2951798,4.420923,4.345436,6.5903597,6.5837955,4.6572313,6.038975,3.8400004,1.910154,0.9288206,0.8992821,1.1684103,1.2570257,1.5491283,1.2603078,0.5677949,0.6170257,1.6475899,2.2580514,2.9111798,3.6562054,4.1485133,4.84759,5.72718,6.7610264,7.9294367,9.196308,9.488411,9.110975,8.247795,7.315693,6.9743595,7.5946674,6.8004107,6.11118,6.0750775,6.2916927,6.8660517,7.6209235,7.90318,7.7456417,7.857231,4.6244106,7.5487185,10.925949,11.365745,7.7981544,7.899898,8.516924,8.342975,6.7577443,3.8367183,5.277539,4.089436,2.681436,3.0293336,6.6494365,11.336206,15.386257,14.670771,9.741129,5.832206,5.933949,4.906667,4.5522056,5.097026,5.179077,8.644924,7.778462,5.7140517,4.46359,4.9099493,3.5807183,5.7042055,7.88677,7.955693,4.9329233,7.6077952,10.9686165,11.602052,9.544206,8.277334,9.291488,12.58995,12.301129,8.910769,9.232411,10.597744,11.122872,10.755282,9.869129,9.29477,6.4722056,5.2611284,5.6418467,6.5903597,6.0717955,4.342154,3.8006158,6.774154,11.575796,12.484924,13.863386,14.10954,9.557334,3.7349746,7.3649235,7.5946674,3.121231,0.059076928,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.036102567,0.059076928,0.06564103,0.09189744,0.1148718,0.12471796,0.15097436,0.19692309,0.23302566,0.20676924,0.24943592,0.47917953,0.8205129,1.017436,0.74830776,0.8960001,1.0994873,1.339077,1.910154,2.6715899,2.7602053,2.737231,2.868513,3.1277952,3.0358977,2.7241027,2.6551797,2.865231,2.9801028,3.4297438,3.373949,3.249231,3.1474874,2.8324106,2.3072822,2.3171284,2.3958976,2.4451284,2.733949,2.9111798,3.1048207,3.249231,3.3476925,3.501949,3.826872,3.9778464,4.2371287,4.71959,5.353026,5.8125134,6.636308,7.4929237,8.054154,8.008205,7.066257,6.2916927,5.7796926,5.32677,4.4274874,3.4002054,2.9604106,2.9407182,3.0916924,3.0654361,2.930872,3.2098465,3.757949,4.3552823,4.6933336,4.522667,4.673641,4.969026,5.395693,6.088206,6.7183595,7.322257,7.6668725,7.709539,7.6077952,7.8703594,8.369231,8.687591,8.776206,8.979693,8.651488,8.274052,8.034462,8.008205,8.136206,7.8145647,7.706257,7.50277,7.02359,6.2194877,5.796103,5.7468724,6.1997952,6.9021544,7.2369237,5.805949,6.262154,6.485334,6.0849237,6.3934364,7.00718,7.6931286,8.234667,8.723693,9.573745,9.271795,8.280616,7.4043083,6.889026,6.422975,6.452513,6.669129,6.3573337,5.3891287,4.194462,3.8662567,5.0838976,6.1538467,6.232616,5.333334,4.315898,4.378257,4.9329233,5.5236926,5.8157954,5.8847184,4.7425647,4.9493337,6.665847,7.643898,7.719385,5.609026,3.6004105,3.5314875,6.7610264,5.3694363,5.5663595,6.554257,7.128616,5.654975,4.2207184,3.8006158,4.2207184,4.962462,5.1889234,3.9023592,3.2032824,3.249231,3.5249233,2.8389745,4.5522056,4.466872,4.2371287,4.1813335,3.2656412,2.9801028,3.2722054,3.3772311,3.0785644,2.7044106,2.8324106,2.7109745,2.412308,2.1267693,2.172718,2.4549747,2.6683078,2.8389745,3.0916924,3.6332312,3.4592824,3.2787695,3.1409233,3.0884104,3.1343591,3.436308,4.164923,4.850872,5.3234878,5.733744,6.4295387,6.163693,5.7698464,5.5269747,5.159385,5.901129,6.564103,6.636308,6.0783596,5.32677,4.585026,4.493129,4.7950773,5.2381544,5.5663595,5.0149746,4.900103,4.9952826,5.333334,6.1997952,5.9995904,5.970052,5.920821,5.8420515,5.874872,5.8420515,5.83877,5.7009234,5.5105643,5.5958977,5.796103,5.1987696,4.7491283,4.535795,3.7809234,2.7766156,2.409026,2.0709746,1.5261539,0.90912825,0.79097444,0.6892308,0.6695385,0.69579494,0.6170257,0.5546667,0.446359,0.38728207,0.38400003,0.34133336,0.46276927,0.60389745,0.69907695,0.69579494,0.5481026,0.5218462,0.5940513,0.72861546,0.90584624,1.1060513,1.5097437,1.9396925,2.0151796,1.6705642,1.1520001,1.4867693,1.6640002,1.8084104,1.9922053,2.2416413,1.8445129,1.8281027,1.9561027,2.1431797,2.4484105,2.678154,2.5895386,2.6256413,2.7109745,2.225231,1.8346668,1.8445129,2.0020514,2.2350771,2.6420515,3.2853336,3.4297438,3.1967182,2.7142565,2.0906668,2.0906668,2.2547693,2.2121027,2.034872,2.2186668,2.425436,2.4451284,2.4024618,2.4155898,2.5895386,2.6978464,3.1113849,3.4100516,3.4264617,3.2525132,3.498667,3.1606157,2.989949,3.1671798,3.3050258,4.164923,5.6943593,5.917539,5.0084105,5.284103,4.273231,3.9942567,3.7809234,3.698872,3.7415388,3.8367183,4.1846156,4.5587697,4.8344617,5.0477953,5.3727183,5.474462,5.7731285,6.166975,6.744616,7.748924,8.15918,9.173334,9.472001,9.025641,9.07159,10.230155,10.696206,11.044104,11.487181,11.890873,12.507898,12.688411,12.291283,11.818667,12.432411,12.228924,12.42913,12.291283,11.894155,12.153437,13.200411,14.237539,15.465027,16.682669,17.257027,18.025026,19.209848,20.854155,23.194258,26.663387,28.649029,30.592003,33.3719,36.483284,38.029133,40.612106,40.70072,41.793644,45.712414,52.608006,50.05785,44.71467,38.272003,31.839182,25.93149,20.955898,16.843489,13.827283,11.411694,8.375795,6.058667,4.420923,3.0949745,1.9692309,1.1815386,1.1552821,0.90584624,0.63343596,0.4955898,0.6301539,0.33476925,0.256,0.23630771,0.190359,0.101743594,0.04266667,0.029538464,0.032820515,0.032820515,0.032820515,0.029538464,0.009846155,0.0032820515,0.016410258,0.055794876,0.072205134,0.059076928,0.06564103,0.08861539,0.068923086,0.08205129,0.18051283,0.18051283,0.072205134,0.013128206,0.006564103,0.009846155,0.006564103,0.0,0.0,0.04266667,0.026256412,0.006564103,0.0032820515,0.01969231,0.009846155,0.0032820515,0.0,0.0032820515,0.009846155,0.029538464,0.34133336,0.512,0.51856416,0.76800007,1.4539489,1.5885129,1.8412309,2.3138463,2.5665643,2.865231,2.7700515,2.7667694,2.7569232,2.038154,2.4155898,2.3302567,2.3040001,2.3794873,2.1267693,1.9593848,1.9954873,2.166154,2.540308,3.3378465,3.4330258,3.442872,3.7776413,4.1583595,3.623385,5.5696416,5.9667697,7.650462,10.765129,12.763899,12.488206,12.475078,12.4685135,12.905026,14.943181,15.671796,15.504412,15.264822,14.834873,13.144616,11.664412,11.303386,11.621744,12.20595,12.665437,13.22995,14.628103,15.314053,14.916924,14.230975,13.433437,12.074668,10.86359,9.875693,8.562873,8.339693,9.160206,9.957745,10.279386,10.28595,11.98277,13.088821,12.773745,11.16554,9.344001,8.818872,9.193027,8.444718,6.9054365,7.2631803,7.351795,7.643898,8.28718,9.048616,9.330873,9.494975,9.458873,9.53436,9.938052,10.794667,11.195078,10.834052,10.597744,10.692924,10.643693,10.742155,11.090053,11.690667,12.182976,11.82195,12.977232,13.13477,12.714667,12.097642,11.618463,11.487181,11.119591,10.312206,9.291488,8.700719,9.38995,10.541949,12.179693,13.984821,15.297642,17.076513,20.6999,20.312616,15.16636,9.626257,10.6469755,11.756309,13.472821,15.67836,17.631182,17.414566,16.423386,14.992412,13.676309,13.243078,12.73436,11.72677,11.227899,11.631591,12.740924,14.267078,15.048206,15.908104,16.800821,16.804104,15.560206,14.427898,14.762668,15.809642,14.716719,12.780309,11.208206,10.345026,10.069334,9.803488,9.7673855,9.462154,9.563898,10.331899,11.58236,10.20718,8.904206,8.01477,7.9491286,9.199591,9.40636,8.812308,8.539898,8.923898,9.501539,8.897642,7.2664623,5.2709746,3.5872824,2.8947694,5.681231,4.565334,3.4756925,3.764513,4.194462,3.7087183,5.175795,5.293949,4.132103,5.139693,3.5511796,2.0742567,1.0699488,0.6662565,0.7581539,3.5249233,5.333334,4.201026,1.1881026,0.38728207,1.083077,1.7985642,2.5600002,3.2787695,3.7448208,4.4701543,5.225026,6.163693,7.3386674,8.677744,8.953437,8.986258,8.5202055,7.5881033,6.5083084,6.8332314,6.370462,5.8880005,5.861744,6.4754877,7.1023593,7.0498466,9.577026,12.973949,10.555078,7.5913854,9.882257,12.412719,11.913847,6.885744,6.4032826,7.5520005,7.709539,6.5805135,6.1768208,5.5236926,3.9811285,3.5741541,4.6539493,5.924103,7.568411,10.157949,10.597744,8.930462,8.316719,9.787078,9.238976,7.328821,5.32677,5.1265645,7.197539,8.283898,7.8047185,7.020308,9.009232,7.7390776,5.723898,4.844308,5.3037953,5.6385646,6.0783596,9.321027,11.241027,10.512411,8.598975,9.662359,11.500309,11.339488,9.554052,9.6754875,9.025641,9.143796,10.709334,12.310975,10.450052,6.180103,6.196513,7.259898,7.4830775,6.3245134,5.943795,4.775385,5.2644105,7.003898,6.7314878,9.796924,11.418258,8.231385,2.989949,4.565334,4.6178465,1.9528207,0.13784617,0.072205134,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.026256412,0.055794876,0.08861539,0.118153855,0.12471796,0.15097436,0.19692309,0.24287182,0.25271797,0.20348719,0.2231795,0.3511795,0.6071795,0.9878975,0.73517954,0.86974365,0.9878975,1.0633847,1.4572309,1.9659488,2.4746668,2.7437952,2.7470772,2.681436,2.7569232,2.8258464,2.9046156,3.0326157,3.2918978,3.4855387,3.4231799,3.2164104,2.917744,2.546872,2.3466668,2.422154,2.3991797,2.3204105,2.6486156,3.114667,3.5216413,3.7316926,3.882667,4.417641,4.562052,4.8016415,4.9493337,5.156103,5.8847184,6.3967185,6.957949,7.2172313,7.0892315,6.744616,6.2194877,5.799385,5.5269747,5.2053337,4.4077954,3.5511796,3.2262566,3.1474874,3.0884104,2.861949,3.3542566,3.7842054,4.0500517,4.2207184,4.535795,4.699898,5.07077,5.6418467,6.2916927,6.7971287,7.3485136,8.14277,8.615385,8.690872,8.795898,8.953437,8.960001,9.035488,9.186462,9.18318,8.802463,8.73354,8.700719,8.635077,8.67118,8.562873,8.3823595,8.146052,7.8080006,7.2960005,6.820103,6.5083084,6.5247183,6.885744,7.456821,6.5017443,5.989744,5.2676926,4.6605134,5.474462,6.4295387,7.7292314,8.786052,9.120821,8.372514,8.018052,7.6176414,6.665847,5.467898,5.139693,5.5565133,5.5991797,5.5105643,5.4449234,5.4974365,4.8672824,5.297231,6.193231,7.1154876,7.77518,6.701949,5.907693,5.4186673,5.3694363,6.0028725,6.6395903,5.1987696,4.089436,4.279795,5.3103595,4.7655387,4.0434875,3.9909747,4.9132314,6.554257,6.3540516,6.7774363,6.557539,5.3070774,3.5282054,2.353231,2.6584618,3.7087183,4.7458467,4.9854364,3.6004105,3.4264617,3.6660516,3.7218463,3.2131286,3.8498464,3.8629746,3.82359,3.7743592,3.259077,3.1474874,3.4034874,3.2787695,2.7569232,2.5435898,2.5796926,2.3926156,2.2678976,2.3302567,2.556718,2.5665643,2.6715899,2.8488207,3.1015387,3.4658465,3.2853336,3.1606157,3.114667,3.186872,3.4297438,3.6529233,4.535795,5.0116925,4.926359,5.0609236,5.868308,6.091488,5.8190775,5.356308,5.2315903,5.586052,5.6943593,5.674667,5.5204105,5.074052,4.5817437,4.7655387,5.0838976,5.3005133,5.474462,4.919795,4.706462,4.854154,5.362872,6.2063594,5.907693,5.6418467,5.5138464,5.5597954,5.733744,5.684513,5.5696416,5.5729237,5.648411,5.5105643,5.182359,4.844308,4.312616,3.6890259,3.370667,2.9669745,2.6387694,2.2153847,1.7362052,1.4473847,0.9878975,0.88943595,0.88943595,0.8402052,0.69579494,0.51856416,0.4955898,0.5218462,0.54482055,0.57764107,0.5973334,0.65312827,0.69907695,0.69579494,0.60061544,0.5513847,0.57764107,0.6498462,0.77128214,0.9747693,1.2800001,1.4802053,1.5491283,1.5392822,1.5753847,1.6836925,1.6311796,1.6213335,1.7526156,2.0020514,1.7460514,1.8937438,2.166154,2.359795,2.3433847,2.7602053,2.7241027,2.6420515,2.5961027,2.3204105,2.0545642,1.8182565,1.7558975,1.9462565,2.3991797,2.740513,3.0326157,3.0194874,2.789744,2.7503593,2.2744617,2.15959,2.097231,2.0512822,2.2350771,2.4385643,2.5993848,2.6453335,2.6223593,2.674872,2.4976413,2.7667694,3.1343591,3.3608208,3.318154,3.3969233,3.3805132,3.56759,3.9187696,4.059898,4.493129,5.720616,6.298257,5.904411,5.346462,4.4734364,4.132103,3.820308,3.8859491,4.2568207,4.4340515,4.5062566,4.821334,5.0510774,5.156103,5.402257,5.549949,5.674667,6.166975,7.141744,8.418462,8.487385,9.025641,9.38995,9.573745,10.200616,11.490462,12.022155,12.12718,12.06154,12.035283,12.521027,12.859077,12.721231,12.448821,13.029744,12.73436,12.898462,12.809847,12.685129,13.659899,14.152206,14.657642,15.471591,16.305231,16.275694,16.928822,17.778873,19.134361,21.385847,24.98954,26.17436,28.146873,30.46072,32.68267,34.415592,37.14954,38.308105,40.595695,43.989338,45.745235,38.69539,31.753849,26.30236,22.229336,17.929848,13.37436,10.056206,7.7948723,6.163693,4.4996924,3.4789746,2.7503593,2.1924105,1.7001027,1.1749744,1.1323078,1.2603078,1.3062565,1.2077949,1.1093334,0.86317956,0.6465641,0.48246157,0.3314872,0.08861539,0.09189744,0.15097436,0.14769232,0.08205129,0.059076928,0.06235898,0.032820515,0.006564103,0.0032820515,0.02297436,0.032820515,0.04594872,0.07548718,0.101743594,0.08205129,0.068923086,0.15097436,0.15753847,0.06564103,0.006564103,0.0,0.0,0.0,0.0,0.0,0.04266667,0.026256412,0.009846155,0.01969231,0.049230773,0.016410258,0.0032820515,0.0,0.0032820515,0.009846155,0.055794876,0.3446154,0.4266667,0.42994875,1.0502565,2.0775387,2.1136413,2.231795,2.6715899,2.8356924,2.7766156,2.9571285,2.9210258,2.481231,1.7329233,2.4713848,2.3729234,2.3236926,2.4320002,2.034872,1.7263591,1.9823592,2.2646155,2.6683078,3.9351797,3.8564105,3.7743592,3.9581542,4.1583595,3.5905645,5.5893335,6.4295387,7.7456417,9.915077,12.087796,12.228924,12.4685135,12.665437,12.928001,13.61395,14.657642,15.40595,15.264822,14.135796,12.386462,10.65354,10.433641,11.057232,12.189539,13.824001,14.329437,15.973744,16.833643,16.305231,15.104001,13.279181,11.408411,10.256411,9.856001,9.5146675,8.516924,8.937026,9.465437,9.810052,10.692924,12.406155,12.882052,11.904001,10.069334,8.802463,8.789334,9.42277,8.963283,7.5552826,7.240206,7.4436927,7.571693,8.070564,8.73354,8.704,8.92718,9.110975,9.426052,9.970873,10.758565,11.280411,11.16554,10.909539,10.660104,10.230155,10.240001,10.962052,11.67754,11.910565,11.437949,12.763899,13.571283,13.499078,12.632616,11.497026,10.801231,10.33518,9.67877,8.933744,8.687591,8.838565,9.764103,11.204924,12.836103,14.273643,15.287796,19.062155,20.857437,18.323694,11.487181,10.492719,11.044104,12.796719,15.471591,18.84554,18.025026,17.237335,16.367592,15.501129,14.913642,14.283488,12.931283,12.117334,12.383181,13.564719,14.181745,14.959591,16.196924,17.411283,17.339079,15.478155,13.51877,13.495796,14.890668,14.605129,13.850258,12.337232,11.175385,10.827488,11.10318,11.733335,11.664412,11.493745,11.631591,12.327386,10.364718,8.828718,8.201847,8.598975,9.754257,10.102155,9.754257,9.396514,9.5606165,10.630565,10.568206,8.749949,6.3868723,4.345436,3.1770258,5.9470773,4.8607183,4.197744,4.716308,3.636513,3.5807183,4.1813335,4.3027697,3.892513,3.9975388,2.733949,2.1858463,1.4605129,0.60389745,0.5874872,3.8006158,5.681231,4.9362054,2.281026,0.43651286,0.8008206,1.529436,2.297436,2.9669745,3.5971284,4.532513,5.2053337,5.904411,6.8004107,7.939283,8.2904625,8.556309,8.54318,8.03118,6.7905645,6.9349747,6.7314878,6.3179493,6.0783596,6.6461544,7.24677,6.705231,9.120821,13.128206,11.910565,10.105436,10.9226675,11.989334,11.145847,6.4590774,4.322462,4.8607183,5.5269747,6.042257,8.379078,6.9645133,4.8114877,4.273231,5.142975,4.6539493,5.612308,7.6570263,8.992821,9.160206,9.028924,10.102155,10.643693,9.019077,6.058667,5.0674877,5.8420515,7.781744,8.625232,8.28718,8.887795,9.137232,6.951385,4.7950773,3.9811285,4.6572313,4.089436,6.409847,8.480822,8.805744,7.4896417,8.503796,8.349539,8.648206,9.268514,8.339693,7.4240007,6.8594875,8.861539,11.52,8.809027,5.474462,6.9152827,8.694155,8.500513,6.157129,6.5969234,5.684513,4.9460516,4.7360005,4.2371287,6.557539,8.43159,6.6461544,2.6026669,2.3302567,1.8609232,0.8566154,0.21333335,0.11158975,0.02297436,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.009846155,0.03938462,0.07876924,0.118153855,0.15753847,0.19692309,0.23958977,0.27241027,0.24615386,0.2231795,0.22646156,0.28225642,0.43651286,0.761436,0.7253334,0.82379496,0.8598975,0.8730257,1.1454359,1.522872,2.1956925,2.609231,2.5961027,2.3663592,2.5206156,2.7995899,2.9833848,3.114667,3.5052311,3.6857438,3.6594875,3.5577438,3.308308,2.6387694,2.353231,2.2186668,2.176,2.2777438,2.6683078,3.43959,4.1517954,4.315898,4.2371287,5.0182567,5.428513,5.7731285,5.940513,6.2096415,7.269744,7.568411,7.463385,7.062975,6.4590774,5.737026,5.661539,5.467898,5.2578464,4.9788723,4.417641,3.7284105,3.370667,3.0818465,2.7667694,2.5271797,3.114667,3.620103,4.07959,4.522667,4.955898,5.474462,5.8256416,6.3310776,7.026872,7.650462,8.04759,8.5891285,8.960001,9.133949,9.373539,9.688616,9.659078,9.573745,9.458873,9.078155,8.694155,8.805744,8.973129,9.015796,9.028924,8.828718,8.369231,8.0377445,7.9130263,7.7423596,7.397744,7.259898,7.2894363,7.2992826,6.941539,6.1407185,5.1298466,4.269949,4.1222568,5.431795,6.47877,7.893334,8.776206,8.39877,6.235898,7.026872,6.764308,5.4908724,3.9942567,3.826872,4.6145644,4.916513,5.172513,5.3169236,4.775385,4.594872,5.0018463,5.989744,7.3419495,8.625232,6.885744,5.3234878,4.5817437,4.821334,5.684513,6.47877,5.366154,3.9286156,3.1277952,3.3017437,3.006359,3.7120004,4.6834874,5.4875903,5.9930263,7.1515903,7.213949,5.5991797,3.1474874,2.1234872,1.7099489,2.8947694,4.1780515,4.965744,5.5597954,4.384821,4.1911798,3.8334363,3.1770258,3.1113849,3.1015387,3.4560003,3.7251284,3.6824617,3.3312824,3.4264617,3.4002054,3.121231,2.733949,2.6518977,2.356513,2.0644104,2.0611284,2.3433847,2.5993848,2.6584618,2.802872,2.937436,3.0391798,3.1737437,2.986667,2.8816411,2.9046156,3.1343591,3.6857438,4.1091285,4.818052,4.9788723,4.6244106,4.6572313,5.1331286,5.5204105,5.3924108,4.9821544,5.156103,5.395693,5.1922054,4.906667,4.6769233,4.420923,4.5062566,5.2611284,5.7796926,5.8190775,5.8092313,5.3694363,5.353026,5.5762057,5.914257,6.2818465,5.937231,5.5958977,5.431795,5.4843082,5.674667,5.6976414,5.402257,5.3234878,5.4580517,5.2742567,4.4767184,4.384821,4.0303593,3.3805132,3.3345644,3.18359,2.7011285,2.1956925,1.8970258,1.9462565,1.3259488,1.1323078,1.0929232,1.0075898,0.7515898,0.60389745,0.60389745,0.636718,0.67282057,0.74830776,0.67610264,0.6465641,0.6235898,0.5940513,0.55794877,0.5874872,0.65641034,0.67938465,0.6892308,0.827077,1.083077,1.1979488,1.339077,1.5589745,1.8018463,1.7394873,1.7165129,1.6738462,1.6344616,1.6771283,1.6508719,1.8609232,2.172718,2.3893335,2.2514873,2.5731285,2.4024618,2.1202054,1.9593848,2.0020514,2.0709746,1.8937438,1.8182565,1.9889232,2.3696413,2.4024618,2.6847181,2.7569232,2.6387694,2.8356924,2.4648206,2.359795,2.28759,2.2514873,2.484513,2.6847181,2.9111798,3.0096412,2.9965131,3.0818465,2.7798977,2.865231,3.1015387,3.2951798,3.31159,3.3542566,3.636513,3.8859491,4.017231,4.1025643,4.634257,5.7074876,6.4065647,6.311385,5.4875903,4.4800005,4.204308,3.9844105,4.332308,4.972308,4.84759,4.8705645,5.2020516,5.536821,5.7107697,5.7009234,5.901129,5.917539,6.304821,7.177847,8.198565,8.605539,8.887795,9.212719,9.878975,11.319796,12.599796,13.239796,13.11836,12.47836,11.920411,12.553847,13.223386,13.761642,14.063591,14.10954,13.115078,13.259488,13.702565,14.263796,15.409232,15.589745,15.432206,15.609437,15.921232,15.268104,15.770258,16.416822,17.289848,18.73395,21.35631,22.455797,25.4359,27.3559,28.534157,32.521847,35.154053,37.353027,39.880207,41.82318,40.592415,33.62462,27.43795,22.92513,19.259079,13.869949,9.494975,6.987488,5.467898,4.3651285,3.4067695,3.18359,2.8324106,2.4385643,2.0151796,1.5064616,1.6016412,2.0742567,2.409026,2.428718,2.3040001,1.9265642,1.2668719,0.90256417,0.79425645,0.2986667,0.27569234,0.33805132,0.28225642,0.118153855,0.072205134,0.072205134,0.049230773,0.01969231,0.009846155,0.01969231,0.01969231,0.04266667,0.059076928,0.059076928,0.04594872,0.03938462,0.07548718,0.08861539,0.059076928,0.02297436,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.009846155,0.032820515,0.06235898,0.01969231,0.0032820515,0.0,0.0,0.0,0.049230773,0.032820515,0.14441027,0.5415385,1.3292309,2.2711797,2.3663592,2.3335385,2.3827693,2.2088206,2.5731285,2.6518977,2.484513,2.1202054,1.6246156,2.477949,2.2711797,1.8510771,1.6935385,1.9232821,1.8313848,2.2613335,2.5895386,2.937436,4.1583595,3.4855387,3.7218463,3.9647183,3.9548721,4.076308,4.453744,5.5236926,7.2237954,9.229129,10.95877,12.005745,12.560411,12.744206,12.58995,12.025436,12.819694,14.086565,14.680616,14.148924,12.737642,11.021129,10.637129,11.034257,12.032001,13.820719,15.028514,16.420103,17.555695,17.782156,16.242872,13.423591,11.539693,10.361437,9.829744,10.052924,9.179898,9.222565,9.268514,9.301334,10.200616,12.09436,12.317539,11.050668,9.127385,8.03118,9.245539,10.174359,10.04636,8.923898,7.6996927,8.04759,8.093539,8.070564,8.008205,7.6964107,8.214975,8.940309,9.508103,9.888822,10.390975,10.919386,11.247591,11.218052,10.752001,9.819899,9.974154,10.925949,11.651283,11.697231,11.185231,12.616206,13.689437,13.856822,12.996924,11.431385,10.761847,10.213744,9.38995,8.667898,9.170052,8.982975,9.662359,10.9686165,12.3995905,13.190565,15.067899,19.137642,21.530258,19.606976,11.946668,11.392001,11.487181,12.47836,14.667488,18.402462,17.608206,17.35877,17.227488,16.866463,15.990155,15.540514,14.194873,13.223386,13.308719,14.536206,14.880821,15.589745,16.784412,18.031591,18.346668,16.466053,13.833847,12.616206,13.226667,14.332719,14.78236,13.200411,11.513436,10.781539,11.1983595,12.875488,13.266052,12.944411,12.458668,12.3306675,9.980719,8.874667,9.028924,9.954462,10.643693,10.505847,10.400822,10.259693,10.453334,11.812103,12.022155,10.016821,7.2303596,4.7655387,3.3936412,3.4855387,3.6135387,4.6834874,5.543385,2.9801028,3.3312824,3.8104618,4.1911798,4.2568207,3.7874875,2.359795,2.3335385,1.8707694,0.8763078,0.9878975,1.8182565,2.0808206,2.7306669,3.0720003,0.75487185,0.85005134,1.4834872,2.1070771,2.6584618,3.5610259,4.8147697,5.6451287,6.3442054,7.0432825,7.6996927,8.041026,8.15918,8.3134365,8.310155,7.522462,7.712821,7.7325134,7.430565,6.9776416,6.8562055,7.1876926,7.4240007,7.837539,8.776206,10.679795,10.896411,11.319796,11.145847,9.777231,6.8004107,3.6529233,2.6223593,3.1474874,4.9362054,7.972103,8.064001,5.504,3.318154,2.5271797,2.1398976,5.986462,10.33518,12.281437,11.008,7.8112826,5.58277,6.8660517,7.5191803,6.2916927,4.8049235,5.330052,6.1013336,6.6034875,6.38359,5.0576415,6.521436,7.509334,6.8430777,5.0871797,4.5587697,3.751385,4.2896414,5.0871797,5.536821,5.4843082,6.5772314,5.8781543,6.304821,7.496206,5.805949,5.835488,4.923077,5.7665644,7.427283,5.32677,4.1846156,6.2720003,8.356103,8.41518,5.6418467,6.0324106,5.681231,5.284103,5.2020516,5.47118,5.280821,6.8332314,6.1505647,3.2032824,1.9035898,1.9495386,1.0305642,0.28225642,0.08533334,0.052512825,0.009846155,0.0,0.0,0.0,0.006564103,0.01969231,0.032820515,0.06564103,0.12471796,0.19692309,0.27241027,0.29538465,0.29538465,0.28882053,0.25271797,0.25928208,0.2297436,0.23630771,0.30851284,0.42338464,0.69907695,0.764718,0.7417436,0.764718,0.98133343,1.3915899,1.8609232,2.231795,2.3827693,2.2514873,2.3269746,2.481231,2.7076926,3.0391798,3.564308,3.9253337,4.017231,4.194462,4.2174363,3.255795,2.5337439,1.9954873,1.9167181,2.2744617,2.7470772,3.761231,4.9493337,5.1265645,4.6276927,5.3103595,6.2523084,6.6625648,7.0498466,7.768616,9.028924,8.746667,7.906462,7.181129,6.62318,5.658257,5.8125134,5.674667,5.421949,5.1232824,4.7425647,3.9581542,3.4166157,2.934154,2.5140514,2.359795,2.3893335,2.8127182,3.820308,5.0674877,5.684513,6.3540516,6.6100516,6.8660517,7.3550773,8.113232,8.569437,8.700719,8.795898,8.963283,9.153642,9.593436,9.810052,9.682052,9.265231,8.769642,8.635077,8.746667,9.002667,9.265231,9.383386,8.861539,8.2904625,7.968821,7.9327188,7.9786673,7.893334,8.083693,8.267488,8.03118,6.813539,5.602462,4.972308,4.903385,5.4153852,6.5837955,7.2664623,7.857231,7.8441033,6.9842057,5.3136415,7.1614366,5.8157954,3.626667,2.1891284,2.349949,3.249231,4.2830772,5.1659493,5.149539,3.0194874,3.6758976,4.71959,6.0258465,7.0334363,6.7282057,4.161641,2.6190772,2.674872,3.9187696,4.9394875,5.1922054,4.6769233,4.023795,3.387077,2.4516926,3.4855387,4.8114877,5.3366156,5.1987696,5.7534366,7.387898,6.567385,4.069744,1.6475899,2.041436,1.8740515,3.4691284,4.781949,5.297231,6.0356927,4.6244106,4.2929235,3.4198978,2.1891284,2.6026669,2.9046156,3.5511796,3.9778464,3.9023592,3.3214362,3.3805132,3.114667,2.9013336,2.8553848,2.8258464,2.2219489,1.9298463,1.9692309,2.2022567,2.3368206,2.681436,2.8455386,2.865231,2.8488207,2.9833848,2.8258464,2.6322052,2.612513,2.9472823,3.8006158,4.5817437,4.926359,4.906667,4.7950773,5.034667,4.965744,5.0051284,4.818052,4.5554876,4.850872,5.346462,5.2381544,4.650667,3.9581542,3.8006158,4.309334,5.4908724,6.242462,6.3245134,6.370462,6.0192823,6.426257,6.75118,6.688821,6.4722056,6.0619493,5.858462,5.7435904,5.6287184,5.4580517,5.7107697,5.398975,5.093744,4.972308,4.818052,3.9286156,3.8662567,3.820308,3.6069746,3.6430771,3.2164104,2.6387694,2.1858463,2.0086155,2.1398976,1.8116925,1.4900514,1.3128207,1.1881026,0.79097444,0.86317956,0.80738467,0.73517954,0.7187693,0.764718,0.67938465,0.636718,0.58092314,0.5218462,0.5349744,0.69907695,0.8336411,0.8336411,0.764718,0.86646163,1.1520001,1.3489232,1.522872,1.6311796,1.5425643,1.4867693,1.7723079,1.8838975,1.7066668,1.5327181,1.6705642,1.7723079,1.9856411,2.2383592,2.225231,2.2153847,1.7624617,1.3292309,1.1979488,1.467077,1.8018463,1.9659488,2.0775387,2.2350771,2.5107694,2.3860514,2.4615386,2.4352822,2.2744617,2.2022567,2.4910772,2.7700515,2.8882053,2.917744,3.1442053,3.2787695,3.4067695,3.4297438,3.4166157,3.6036925,3.4724104,3.4133337,3.4264617,3.4658465,3.4494362,3.6036925,3.9712822,3.9154875,3.4691284,3.3509746,4.164923,5.477744,6.0685134,5.8190775,5.6943593,4.394667,4.529231,4.644103,4.919795,5.139693,4.699898,5.0674877,5.6418467,6.166975,6.554257,6.8955903,6.482052,6.8266673,7.456821,8.172308,9.065026,9.990565,9.764103,9.284924,9.426052,11.063796,12.3306675,12.868924,12.852514,12.616206,12.665437,13.397334,13.827283,14.431181,14.913642,14.204719,12.996924,12.786873,13.397334,14.628103,16.249437,16.324924,16.242872,16.210052,16.256,16.219898,16.000002,15.688207,16.341335,17.828104,18.82913,20.867283,25.186464,28.032001,29.640207,34.254772,35.160618,34.258053,33.73949,34.0119,33.70667,37.159386,33.28985,25.918362,17.690258,10.085744,8.425026,7.453539,5.8912826,3.9909747,3.5413337,3.748103,4.010667,3.3312824,2.03159,1.7394873,2.2022567,2.8947694,3.2754874,3.4264617,4.073026,3.0720003,1.7887181,1.3718976,1.6049232,0.88615394,0.58092314,0.39384618,0.2100513,0.049230773,0.06235898,0.013128206,0.01969231,0.029538464,0.029538464,0.029538464,0.029538464,0.03938462,0.052512825,0.059076928,0.04594872,0.059076928,0.068923086,0.08205129,0.08533334,0.06235898,0.049230773,0.01969231,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.036102567,0.01969231,0.0,0.0,0.0,0.0,0.0,0.029538464,0.13456412,0.36758977,0.28225642,0.3314872,0.49230772,0.7089231,0.9156924,1.4145643,1.3292309,1.3489232,1.5885129,1.5885129,1.270154,1.2537436,1.585231,2.0086155,1.9823592,2.789744,3.0654361,3.0260515,2.9636924,3.2196925,2.6322052,3.373949,3.9056413,3.9548721,4.516103,4.7360005,5.3234878,8.300308,12.045129,11.277129,11.72677,12.235488,12.691693,12.747488,11.795693,11.464206,12.583385,13.938873,14.519796,13.51877,12.310975,12.1928215,12.294565,12.576821,13.8075905,14.8709755,15.67836,16.659693,17.45395,16.89272,14.070155,12.150155,11.191795,10.932513,10.771693,9.7214365,9.452309,9.494975,9.685334,10.161232,12.4685135,12.038565,10.292514,8.434873,7.4469748,9.754257,11.034257,11.224616,10.505847,9.324308,8.283898,8.356103,8.39877,8.149334,8.208411,8.356103,9.32759,9.7214365,9.43918,9.659078,10.000411,10.47959,10.686359,10.407386,9.613129,9.6984625,10.14154,10.689642,11.063796,10.939077,11.648001,12.632616,13.144616,12.714667,11.139283,10.039796,9.757539,9.6295395,9.586872,10.148104,9.744411,11.008,12.662155,13.88636,14.313026,15.898257,19.30831,22.212925,21.00513,10.788103,11.142565,11.542975,12.153437,13.420309,16.082052,16.36431,16.607182,16.81395,16.771284,16.052513,16.295385,15.42236,14.6182575,14.644514,15.852309,16.452925,17.444103,18.195694,18.665028,19.410053,18.458258,15.425642,13.095386,12.649027,13.686155,14.322873,12.996924,11.497026,10.79795,11.076924,13.298873,13.499078,13.065847,12.675283,12.2847185,10.098872,9.40636,9.96759,11.18195,12.084514,11.047385,11.099898,11.411694,11.762873,12.557129,12.668719,10.433641,7.3452315,4.772103,3.9680004,3.1606157,3.1540515,4.4274874,5.533539,3.0654361,1.9331284,3.1671798,4.7622566,5.4974365,4.95918,3.2984617,2.5173335,1.8412309,1.2832822,1.6475899,0.9156924,0.82379496,1.5819489,2.3663592,1.3259488,0.8763078,1.4309745,2.156308,2.7667694,3.5249233,4.768821,5.970052,7.1220517,8.027898,8.283898,8.723693,8.487385,8.198565,8.146052,8.254359,7.450257,7.768616,8.362667,8.418462,7.1876926,6.491898,8.851693,9.842873,8.333129,6.514872,10.154668,12.931283,12.583385,9.472001,6.5903597,7.177847,5.6943593,5.2611284,6.163693,5.858462,3.0523078,1.591795,0.9189744,0.7844103,1.2373334,3.7251284,7.9917955,8.992821,6.678975,5.98318,3.6758976,4.279795,6.0849237,7.686565,7.9786673,7.6635904,6.3934364,5.5893335,5.618872,5.8125134,4.640821,4.824616,6.442667,8.881231,10.834052,6.744616,4.768821,4.325744,4.7392826,5.2644105,7.5585647,6.9349747,5.5007186,4.647385,5.0510774,4.6112823,3.8137438,3.5840003,4.2174363,5.402257,3.6430771,3.8531284,4.263385,4.397949,5.080616,5.412103,4.6867695,3.6004105,3.0293336,4.0434875,3.9712822,5.3169236,5.346462,3.9056413,3.4166157,1.8445129,0.9288206,0.36758977,0.03938462,0.016410258,0.0032820515,0.0,0.0,0.006564103,0.029538464,0.09189744,0.16082053,0.28225642,0.45620516,0.6268718,0.61374366,0.54482055,0.47917953,0.42338464,0.3511795,0.3249231,0.23958977,0.20020515,0.25271797,0.3511795,0.65641034,0.81394875,0.8467693,0.82379496,0.88615394,1.1158975,1.2668719,1.522872,1.8871796,2.166154,2.300718,2.425436,2.5961027,2.9538465,3.7218463,4.1124105,4.2469745,4.4242053,4.46359,3.7087183,3.0227695,2.3138463,2.038154,2.2580514,2.6256413,3.8334363,5.664821,6.091488,5.333334,5.858462,6.957949,7.5618467,8.2445135,8.89436,8.713847,7.686565,7.384616,7.4469748,7.3550773,6.439385,6.2818465,6.2785645,6.308103,6.157129,5.5236926,4.194462,3.4133337,2.9243078,2.6026669,2.4582565,2.225231,2.7076926,3.7087183,4.781949,5.2348723,5.7468724,6.242462,6.747898,7.256616,7.719385,9.271795,9.750975,9.43918,8.858257,8.772923,8.786052,8.79918,8.6580515,8.4053335,8.27077,8.809027,8.950154,9.07159,9.396514,9.993847,9.531077,9.084719,8.63836,8.3823595,8.713847,9.019077,8.746667,8.448001,8.339693,8.316719,7.9130263,7.7292314,7.8473854,7.9852314,7.522462,7.8637953,7.8506675,7.4404106,7.2303596,8.438154,8.4512825,5.605744,2.4943593,0.8369231,1.4966155,1.8379488,3.3312824,4.7983594,5.277539,4.0434875,4.604718,5.211898,5.8847184,5.677949,2.7011285,1.8346668,1.7558975,2.284308,3.3050258,4.7458467,4.2929235,4.2896414,3.754667,2.7667694,2.487795,5.4153852,6.422975,6.1505647,5.349744,4.896821,6.193231,5.6451287,3.698872,1.9331284,3.0654361,1.8937438,3.3312824,4.3716927,4.352,4.97559,3.5347695,3.8695388,3.5511796,2.5895386,3.4330258,3.7251284,4.0467696,4.076308,3.892513,3.9680004,3.626667,3.1277952,2.8225644,2.7634873,2.7175386,1.9954873,1.7624617,1.785436,1.972513,2.349949,2.605949,2.477949,2.4549747,2.7175386,3.1442053,2.9833848,2.6518977,2.5009232,2.7634873,3.5544617,4.4964104,4.7655387,4.6769233,4.630975,5.156103,5.402257,5.3694363,5.284103,5.218462,5.097026,5.32677,4.955898,4.352,3.9712822,4.348718,4.7524104,5.3924108,5.533539,5.35959,5.979898,5.786257,6.11118,6.4656415,6.5345645,6.180103,6.0324106,6.042257,5.9569235,5.5663595,4.699898,5.431795,5.421949,5.0215387,4.5489235,4.31918,3.5380516,3.5446157,3.639795,3.5938463,3.6332312,3.0096412,2.6518977,2.3663592,2.1136413,2.028308,2.3466668,2.097231,1.723077,1.401436,1.020718,1.2406155,1.0666667,0.81066674,0.65641034,0.65641034,0.55794877,0.6170257,0.63343596,0.5940513,0.65641034,0.8992821,0.9878975,1.0075898,1.0633847,1.2832822,1.3915899,1.5392822,1.6902566,1.6869745,1.2373334,1.0666667,1.4539489,1.7099489,1.6311796,1.4966155,1.654154,1.7296412,1.847795,1.9790771,1.9692309,1.8707694,1.5425643,1.3554872,1.4178462,1.6016412,1.4178462,1.8871796,2.300718,2.4516926,2.609231,2.2186668,2.1103592,2.1103592,2.1300514,2.166154,2.2416413,2.550154,3.3214362,4.1550775,4.059898,3.8990772,3.82359,3.7448208,3.6660516,3.6758976,3.8498464,3.7251284,3.7382567,3.8629746,3.629949,3.8137438,4.529231,4.7294364,4.132103,3.2032824,3.117949,3.8104618,4.5817437,5.218462,6.012718,4.2240005,4.4767184,4.519385,4.529231,4.6244106,4.857436,5.6352825,6.226052,6.6428723,6.9645133,7.3353853,6.550975,6.6034875,6.882462,7.1220517,7.4174366,8.704,8.973129,9.616411,10.962052,12.245335,12.481642,12.803283,12.947693,12.928001,13.056001,13.318565,13.574565,13.679591,13.673027,13.764924,13.6697445,14.12595,15.126975,16.282257,16.810667,16.259283,16.36431,15.983591,15.24513,15.560206,16.131283,15.819489,16.538258,18.15631,18.51077,20.374975,24.74995,28.235489,29.892925,31.264822,30.322874,31.494566,32.20349,32.692516,36.036926,45.32185,41.41621,30.365541,17.900309,9.426052,9.691898,8.854975,7.788308,6.8562055,5.8945646,4.578462,3.442872,2.356513,1.8018463,2.8750772,4.33559,4.315898,3.5807183,2.8914874,3.0129232,2.176,1.5064616,0.9616411,0.5940513,0.51856416,0.3511795,0.2855385,0.18707694,0.07548718,0.14769232,0.07876924,0.029538464,0.006564103,0.009846155,0.01969231,0.009846155,0.016410258,0.036102567,0.068923086,0.0951795,0.08861539,0.08861539,0.1148718,0.13128206,0.049230773,0.055794876,0.029538464,0.013128206,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.04594872,0.118153855,0.13456412,0.068923086,0.08861539,0.3052308,0.65312827,0.892718,1.6147693,1.4998976,1.4933335,1.7493335,1.6114873,1.3620514,2.097231,2.5435898,2.4024618,2.349949,2.678154,2.3991797,2.3236926,2.7667694,3.5478978,3.1770258,3.564308,3.6890259,3.511795,3.9548721,4.926359,5.970052,7.860513,9.924924,10.043077,11.119591,11.943385,13.37436,15.074463,15.51754,15.100719,14.759386,14.532925,14.155488,13.069129,13.499078,13.98154,14.50995,15.0777445,15.67836,16.66954,16.873028,17.027283,16.97477,15.671796,14.460719,13.321847,12.570257,12.212514,11.956513,11.024411,10.364718,10.089026,10.282667,10.9915905,12.448821,12.160001,10.217027,7.8736415,7.5191803,9.288206,10.985026,11.776001,11.434668,10.348309,9.409642,9.005949,8.917334,9.15036,9.954462,9.741129,10.459898,10.817642,10.243283,8.900924,8.960001,9.114257,9.432616,9.691898,9.357129,9.793642,9.754257,9.705027,9.980719,10.758565,11.339488,11.828514,11.9171295,11.828514,12.324103,12.317539,11.670976,11.172104,10.9915905,10.683078,10.328616,11.723488,14.122667,16.128002,15.668514,16.443079,17.401438,19.74154,20.073027,10.420513,9.944616,11.316514,12.504617,13.213539,14.897232,15.75713,15.983591,16.259283,16.551386,16.12472,16.75159,16.403694,15.51754,14.808617,15.304206,16.741745,18.103796,18.871796,18.914463,18.517334,16.443079,15.491283,15.018668,14.716719,14.601848,13.958565,12.813129,12.051693,12.137027,13.092104,14.444309,13.538463,12.3995905,11.861334,11.588924,10.525539,10.085744,10.617436,11.808822,12.681848,11.723488,12.2847185,12.826258,12.84595,12.888617,13.4170265,10.95877,7.2270775,4.132103,3.7842054,3.4756925,2.8816411,3.4822567,4.585026,3.31159,2.1464617,2.8980515,3.95159,4.630975,5.228308,5.920821,3.9909747,1.913436,1.0272821,1.5491283,1.2176411,1.5556924,1.7624617,1.4736412,0.7778462,0.7187693,1.1520001,2.0512822,3.1277952,3.817026,4.926359,5.7468724,6.7150774,7.53559,7.1876926,7.6274877,7.9819493,7.3714876,6.695385,8.621949,7.77518,6.7249236,6.951385,8.746667,11.21477,11.641437,11.641437,12.248616,13.078976,12.324103,7.965539,8.392206,7.453539,4.457026,4.1747694,5.3169236,5.2315903,5.3891287,5.549949,3.761231,1.9692309,1.4112822,1.8937438,2.9768207,3.9942567,3.4494362,4.0402055,4.391385,3.9712822,3.1015387,4.210872,5.940513,6.76759,6.301539,5.293949,4.352,5.402257,5.901129,5.2709746,4.9099493,4.1878977,3.8531284,4.5587697,6.4656415,9.258667,7.1515903,4.919795,3.4855387,3.7842054,6.741334,9.80677,10.121847,7.9261546,4.713026,3.2328207,4.0533338,4.010667,3.5971284,3.1442053,2.8258464,2.2678976,2.9472823,3.7251284,4.31918,5.32677,4.9329233,4.056616,2.8750772,1.9790771,2.3958976,3.7874875,3.9318976,3.3575387,2.858667,3.501949,1.9003079,0.88943595,0.47917953,0.41682056,0.19692309,0.16738462,0.108307704,0.04266667,0.02297436,0.1148718,0.36102566,0.5316923,0.5973334,0.60389745,0.636718,0.7811283,0.7975385,0.7318975,0.60389745,0.42338464,0.3314872,0.24943592,0.2100513,0.2297436,0.28882053,0.41025645,0.54482055,0.65641034,0.71548724,0.6892308,0.9321026,1.0896411,1.2800001,1.4802053,1.5556924,1.8970258,2.284308,2.546872,2.8356924,3.626667,3.5380516,3.6758976,3.879385,3.9089234,3.4756925,3.1638978,2.8455386,2.8291285,3.0982566,3.308308,3.82359,5.218462,6.0160003,6.0947695,6.688821,7.3485136,7.968821,8.372514,8.4283085,8.041026,7.522462,7.430565,7.171283,6.5870776,5.927385,5.58277,5.58277,5.5696416,5.330052,4.8049235,4.821334,4.135385,3.245949,2.5895386,2.5435898,2.553436,3.5380516,4.4898467,5.0543594,5.5269747,6.2555904,6.6395903,7.0892315,7.509334,7.328821,8.198565,9.084719,9.504821,9.275078,8.516924,8.684308,9.124104,8.956718,8.198565,7.768616,7.906462,8.146052,8.1755905,8.172308,8.809027,8.982975,9.156924,9.281642,9.337437,9.334154,9.268514,9.028924,8.667898,8.3364105,8.2904625,7.975385,7.9983597,8.392206,8.651488,7.7292314,7.574975,7.39118,6.7807183,6.3277955,7.584821,5.8092313,4.1583595,2.5993848,1.4112822,1.1913847,1.2668719,2.5140514,3.9154875,4.568616,3.6758976,3.2229745,4.017231,4.962462,5.113436,3.6758976,2.477949,2.294154,2.4943593,2.9472823,4.023795,3.9844105,4.4045134,4.565334,4.322462,4.1091285,5.9963083,5.651693,4.785231,4.457026,5.0674877,4.97559,4.640821,4.1911798,3.9581542,4.457026,3.6004105,2.9538465,2.3105643,1.782154,1.7887181,1.7920002,2.7241027,3.1606157,2.9702566,3.3345644,3.3444104,3.564308,3.7021542,3.6824617,3.636513,3.4330258,3.2196925,2.9997952,2.6617439,1.9593848,1.5425643,1.3817437,1.6377437,2.1464617,2.4484105,2.3827693,2.2744617,2.3138463,2.540308,2.8488207,3.2196925,2.865231,2.7011285,3.0523078,3.639795,4.1813335,4.6244106,4.6933336,4.4898467,4.4996924,4.9952826,5.5630774,5.756718,5.481026,4.9985647,4.585026,4.345436,4.381539,4.785231,5.6418467,6.0652313,6.2063594,5.8880005,5.6320004,6.665847,6.186667,6.560821,6.4590774,5.72718,5.3727183,5.7074876,5.4383593,5.3037953,5.3792825,5.077334,4.775385,4.903385,4.8016415,4.4110775,4.2568207,4.1485133,4.1714873,4.056616,3.8038976,3.6430771,2.9636924,2.553436,2.349949,2.1825643,1.785436,2.5895386,2.5796926,2.1530259,1.6705642,1.4506668,1.5031796,1.3259488,1.086359,0.86646163,0.6301539,0.6301539,0.82379496,0.88287187,0.8008206,0.8992821,0.9682052,0.88943595,0.83035904,0.86317956,0.96492314,1.083077,1.2340513,1.4539489,1.6344616,1.5031796,1.1782565,1.2931283,1.3686155,1.276718,1.2406155,1.6114873,1.8674873,1.9200002,1.8182565,1.7493335,1.7788719,1.8642052,1.8346668,1.6213335,1.2471796,1.142154,1.3817437,1.7329233,2.0578463,2.3040001,2.1103592,2.1956925,2.281026,2.297436,2.422154,2.6420515,3.05559,3.7284105,4.4242053,4.6080003,4.460308,4.31918,4.020513,3.7251284,3.9351797,4.1156926,4.0533338,3.9778464,3.8400004,3.3280003,3.5971284,4.06318,4.1025643,3.636513,3.117949,3.4034874,4.2338467,4.5456414,4.460308,5.3037953,4.44718,4.630975,4.7425647,4.8114877,4.8640003,4.906667,5.7042055,6.6002054,7.24677,7.381334,6.8233852,6.3474874,6.304821,6.557539,7.0137444,7.5979495,8.963283,9.898667,11.024411,12.27159,12.882052,12.635899,12.987078,13.220103,13.092104,12.842668,12.914873,13.51877,13.682873,13.430155,13.764924,14.10954,14.381949,15.028514,15.872002,16.118155,16.341335,16.787693,16.613745,16.049232,16.384,17.145437,17.509745,18.49436,20.09272,21.26113,24.756516,29.249643,31.72431,32.26913,34.06113,33.798565,36.296207,38.226055,39.1319,41.445747,52.355286,48.88944,35.99754,21.454771,15.852309,15.307488,13.312001,11.815386,10.850462,8.52677,5.8256416,4.266667,2.8389745,1.8412309,2.8488207,3.8006158,3.5183592,2.8324106,2.4320002,2.8291285,2.2482052,1.6114873,0.9616411,0.44307697,0.318359,0.23302566,0.19692309,0.14441027,0.09189744,0.15097436,0.11158975,0.052512825,0.009846155,0.0,0.006564103,0.0,0.01969231,0.059076928,0.0951795,0.08861539,0.09189744,0.1148718,0.11158975,0.07876924,0.04594872,0.06564103,0.04266667,0.01969231,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03938462,0.08205129,0.029538464,0.006564103,0.032820515,0.190359,0.65641034,1.7001027,1.8379488,1.6377437,1.4769232,1.4736412,1.5064616,1.3850257,2.028308,2.4188719,2.356513,2.4418464,2.225231,2.349949,2.878359,3.436308,3.245949,3.383795,3.4527183,3.6562054,4.06318,4.601436,5.402257,5.7435904,6.9710774,8.868103,9.642668,11.82195,12.950975,14.066873,15.363283,16.200207,16.449642,16.351181,15.904821,15.120412,14.017642,14.506668,15.468308,16.456207,17.19795,17.608206,17.575386,17.588514,17.319386,16.416822,14.496821,12.944411,12.274873,11.949949,11.546257,10.752001,10.397539,10.075898,10.128411,10.65354,11.510155,12.770463,11.963078,9.95118,7.9950776,7.748924,9.025641,9.787078,10.157949,10.167795,9.734565,9.632821,9.084719,8.950154,9.481847,10.31877,10.364718,10.6469755,10.81436,10.473026,9.179898,8.546462,8.054154,8.326565,9.130668,9.357129,9.478565,9.321027,9.019077,8.914052,9.540924,10.213744,10.912822,11.579078,12.2617445,13.111795,13.587693,13.29559,12.770463,12.091078,10.893129,11.047385,12.406155,14.148924,15.579899,16.12472,16.918976,17.24718,19.30831,19.636515,9.094564,9.613129,11.651283,12.918155,13.223386,14.50995,15.218873,15.566771,15.927796,16.154257,15.566771,16.141129,16.62031,16.370872,15.566771,15.202463,16.521847,17.939693,18.98995,19.255796,18.369642,15.596309,15.222155,15.730873,16.150976,16.049232,15.399385,13.718975,12.760616,13.269335,14.985847,16.01313,14.129231,12.645744,12.3995905,11.762873,11.126155,10.752001,11.424822,12.727796,13.052719,12.780309,13.541744,13.581129,12.885334,13.200411,13.797745,11.030975,7.2336416,4.276513,3.5840003,3.4297438,2.989949,3.2164104,3.8334363,3.3542566,2.3663592,3.367385,4.0303593,3.9745643,4.772103,5.658257,3.9056413,1.9561027,1.0371283,1.1520001,1.4736412,1.7591796,1.8740515,1.6640002,0.9419488,1.1027694,1.401436,2.0611284,3.0752823,4.194462,4.9952826,5.7468724,6.5345645,7.0859494,6.774154,6.875898,7.0400004,7.1154876,7.4797955,9.025641,9.5835905,7.650462,7.27959,9.094564,10.299078,10.217027,11.388719,12.678565,13.269335,12.672001,5.9963083,4.1747694,3.5610259,2.92759,3.4592824,3.4888208,3.7185643,4.519385,5.1200004,3.5741541,4.919795,4.457026,3.0818465,2.0184617,2.7995899,3.5807183,3.764513,3.6594875,3.1638978,1.7591796,4.6080003,5.481026,5.4875903,5.58277,6.5378466,5.7468724,6.0192823,5.7534366,4.6933336,3.9154875,3.6332312,3.570872,3.69559,4.1878977,5.4416413,4.8771286,4.7458467,4.1550775,3.6824617,5.3727183,7.860513,9.373539,9.875693,9.005949,6.0619493,6.0258465,4.7425647,3.6332312,3.1671798,2.858667,2.1858463,2.6847181,3.7185643,4.818052,5.7074876,4.325744,3.7021542,3.3214362,3.1474874,3.6135387,4.637539,4.6834874,4.332308,4.2305646,5.100308,3.6562054,2.284308,1.1191796,0.37743592,0.3708718,0.36430773,0.2231795,0.14441027,0.14441027,0.06564103,0.22646156,0.42338464,0.5481026,0.5907693,0.6498462,0.67282057,0.67282057,0.67610264,0.65641034,0.54482055,0.36102566,0.26584616,0.21333335,0.190359,0.20020515,0.25271797,0.38728207,0.57764107,0.7417436,0.71548724,0.8336411,1.024,1.211077,1.3554872,1.467077,1.7690258,2.1989746,2.537026,2.9013336,3.748103,3.5840003,3.5971284,3.7809234,4.020513,4.1058464,3.7251284,3.7152824,3.9154875,4.135385,4.164923,4.1846156,4.906667,5.789539,6.5444107,7.1154876,7.2992826,8.001641,8.500513,8.490667,8.067283,8.027898,7.77518,7.3025646,6.7249236,6.265436,5.904411,5.7501545,5.654975,5.4613338,4.9985647,4.781949,4.1846156,3.6430771,3.3280003,3.1573336,3.1015387,4.352,5.4941545,5.8880005,5.6451287,6.193231,6.5936418,7.000616,7.3616414,7.4075904,8.1755905,8.720411,9.176616,9.380103,8.89436,8.684308,8.887795,8.759795,8.362667,8.579283,8.021334,8.067283,8.044309,7.817847,7.79159,8.129642,8.612103,8.897642,8.848411,8.5661545,8.891078,9.120821,9.091283,8.704,7.939283,7.328821,7.4732313,8.001641,8.467693,8.323282,7.9327188,6.9087186,6.2129235,6.0980515,6.114462,4.3027697,3.006359,2.4648206,2.3466668,1.7460514,1.3620514,2.2646155,3.5478978,4.2962055,3.5872824,3.0752823,3.6890259,4.7360005,5.5729237,5.605744,4.273231,3.4133337,3.1474874,3.4198978,3.9909747,3.6726158,4.1714873,4.634257,4.6802053,4.388103,5.0018463,4.4832826,4.1517954,4.381539,4.6080003,4.0434875,3.892513,4.073026,4.322462,4.210872,4.2371287,3.7874875,3.2853336,2.937436,2.7306669,3.2886157,3.31159,3.2689233,3.4100516,3.7776413,3.5052311,3.4724104,3.370667,3.1671798,3.0785644,2.9538465,2.7700515,2.4681027,2.044718,1.5589745,1.6213335,1.9692309,2.3072822,2.4549747,2.3630772,2.2383592,2.3630772,2.553436,2.6978464,2.7602053,2.9669745,2.737231,2.7700515,3.242667,3.8071797,4.269949,4.781949,4.8344617,4.571898,4.8082056,5.3202057,5.654975,5.6943593,5.4416413,5.028103,4.850872,4.6145644,4.4964104,4.630975,5.1232824,5.6254363,5.602462,5.4843082,5.668103,6.5345645,5.9536414,6.1472826,6.183385,5.737026,5.044513,5.481026,5.1987696,4.955898,5.0116925,5.1167183,4.44718,4.4865646,4.571898,4.4996924,4.525949,4.2207184,4.1091285,3.9089234,3.5938463,3.4002054,3.0391798,2.7766156,2.605949,2.4648206,2.1989746,2.7536411,2.8980515,2.6551797,2.1989746,1.8412309,1.5360001,1.4441026,1.2898463,1.0010257,0.7089231,0.7384616,0.88943595,0.8992821,0.8041026,0.9517949,1.1224617,1.0765129,0.90256417,0.77128214,0.9321026,1.1552821,1.211077,1.2242053,1.2668719,1.3423591,1.2832822,1.2537436,1.1552821,1.0601027,1.2012309,1.4966155,1.7263591,1.8182565,1.7985642,1.7952822,1.7755898,1.8510771,1.7690258,1.4572309,1.0305642,1.1651284,1.3620514,1.6344616,1.9232821,2.0906668,2.28759,2.2383592,2.2121027,2.300718,2.3958976,2.4024618,2.8356924,3.4560003,4.010667,4.2141542,4.381539,4.338872,4.1517954,4.007385,4.1911798,4.161641,4.194462,4.1550775,3.9056413,3.3050258,3.8104618,4.266667,4.345436,4.0467696,3.6758976,4.2929235,4.6539493,4.7524104,4.8082056,5.2447186,4.59159,4.5390773,4.7622566,5.0477953,5.2447186,5.280821,5.7796926,6.774154,7.5552826,7.6077952,6.62318,6.2687182,6.2720003,6.675693,7.3386674,7.958975,9.278359,10.768411,12.084514,13.013334,13.466257,13.213539,13.666463,13.840411,13.5318985,13.334975,13.492514,14.221129,14.208001,13.656616,14.290052,14.34913,14.470565,14.746258,15.074463,15.16636,16.288822,16.613745,16.584206,16.65313,17.293129,17.51959,18.514053,19.958155,21.874874,24.612104,30.582157,36.368412,39.42072,39.968822,40.99939,41.652515,44.28472,47.13354,50.16944,55.12862,65.04698,58.673237,43.81867,29.443285,25.62954,23.46667,20.158361,17.660719,15.655386,11.536411,8.264206,6.052103,4.1025643,2.6387694,2.878359,2.9538465,2.4746668,1.9429746,1.785436,2.359795,2.1300514,1.4572309,0.8172308,0.4135385,0.16410258,0.13128206,0.15097436,0.15753847,0.13784617,0.13128206,0.12471796,0.08861539,0.03938462,0.0,0.0,0.009846155,0.06564103,0.14112821,0.18379489,0.108307704,0.07876924,0.08861539,0.068923086,0.029538464,0.052512825,0.06235898,0.059076928,0.03938462,0.01969231,0.036102567,0.02297436,0.006564103,0.0,0.0,0.006564103,0.0,0.0,0.0032820515,0.01969231,0.055794876,0.01969231,0.009846155,0.118153855,0.23630771,0.02297436,0.029538464,0.26256412,0.83035904,1.7165129,2.7798977,2.166154,1.7165129,1.5360001,1.6049232,1.7755898,1.7952822,2.169436,2.284308,2.1300514,2.294154,2.169436,2.5337439,3.117949,3.511795,3.1507695,3.5511796,3.5380516,4.017231,4.8705645,4.9493337,5.5991797,5.618872,6.5378466,8.260923,9.068309,11.316514,12.386462,13.505642,15.05477,16.548103,16.938667,17.06995,16.551386,15.638975,15.241847,15.320617,16.15754,17.404718,18.625643,19.324718,18.743795,18.054565,17.10277,15.803078,14.165335,12.087796,11.306667,10.906258,10.420513,9.842873,9.882257,10.026668,10.220308,10.564924,11.316514,12.800001,11.890873,9.911796,8.165744,7.9425645,8.845129,9.186462,9.248821,9.137232,8.789334,9.619693,9.330873,9.298052,9.947898,10.768411,11.149129,11.152411,11.050668,10.738873,9.728001,8.815591,7.752206,7.762052,8.763078,9.380103,9.399796,9.409642,9.216001,8.973129,9.209436,10.098872,10.620719,11.260718,12.100924,12.819694,12.967385,13.088821,13.046155,12.422565,10.532104,10.870154,12.032001,12.905026,13.456411,14.739694,16.308514,16.278976,17.191385,16.978052,8.966565,9.67877,11.286975,12.593232,13.489232,14.933334,15.645539,15.809642,15.688207,15.317334,14.506668,15.163078,16.150976,16.544823,16.17395,15.619284,16.659693,17.591797,18.54359,19.032618,17.972515,15.271386,15.041642,15.455181,15.812924,16.548103,16.265848,14.749539,13.568001,13.797745,16.006565,17.26031,14.54277,12.731078,12.908309,12.347078,11.224616,10.801231,11.680821,13.154463,13.203693,13.784616,14.775796,14.427898,13.121642,13.387488,13.804309,10.8307705,7.200821,4.588308,3.5840003,3.370667,3.242667,3.2525132,3.3050258,3.18359,2.8389745,4.516103,5.32677,4.9296412,5.546667,5.228308,3.7284105,2.5764105,2.0611284,1.2537436,1.5885129,1.5983591,1.8937438,2.1398976,1.0765129,1.2570257,1.5589745,2.162872,3.121231,4.345436,5.4843082,6.23918,6.744616,6.9087186,6.4032826,6.3376417,6.3540516,7.1581545,8.3823595,8.5661545,10.752001,9.8592825,8.723693,8.457847,8.474257,10.41395,11.523283,11.257437,10.052924,9.301334,5.287385,3.3542566,3.4067695,4.44718,4.578462,3.370667,3.1409233,3.95159,4.9821544,4.5062566,7.9195905,6.3474874,3.7120004,2.2383592,2.4320002,3.4921029,3.259077,2.802872,2.6584618,2.8127182,5.8518977,6.038975,6.0291286,6.770872,7.5191803,8.027898,7.1614366,6.0717955,5.1659493,4.1058464,3.249231,3.370667,3.5052311,3.3608208,3.3247182,3.8400004,4.7983594,5.077334,4.6211286,4.460308,5.398975,6.9349747,9.202872,10.738873,8.474257,7.256616,5.8518977,4.4274874,3.3936412,3.4264617,3.1737437,3.8137438,5.037949,6.160411,6.114462,4.312616,3.3969233,3.2032824,3.495385,3.9680004,4.571898,5.228308,5.609026,5.8157954,6.363898,4.2994876,3.0687182,1.8149745,0.6104616,0.45620516,0.48902568,0.3052308,0.19364104,0.20676924,0.15425642,0.13128206,0.23958977,0.36430773,0.47261542,0.5940513,0.5973334,0.5677949,0.5874872,0.63343596,0.58092314,0.3446154,0.24615386,0.19364104,0.15425642,0.15097436,0.20020515,0.2986667,0.4955898,0.7089231,0.7318975,0.7187693,0.86646163,1.1257436,1.3653334,1.3751796,1.5458462,2.03159,2.477949,2.9046156,3.7054362,3.8301542,3.8596926,4.0992823,4.4898467,4.630975,4.1813335,4.388103,4.7360005,4.9362054,4.9362054,4.706462,4.972308,5.861744,6.9710774,7.3780518,7.253334,7.860513,8.55959,8.809027,8.1755905,8.103385,7.680001,7.240206,6.9776416,6.9743595,6.629744,6.2063594,5.979898,5.858462,5.395693,5.041231,4.4964104,4.1714873,4.132103,4.066462,4.1124105,5.0051284,6.1013336,6.7249236,6.1538467,6.3540516,6.636308,7.030154,7.4141545,7.53559,8.2445135,8.530052,8.809027,8.982975,8.434873,8.123077,8.234667,8.234667,8.172308,8.681026,8.149334,8.083693,7.896616,7.4207187,6.931693,7.532308,8.247795,8.717129,8.861539,8.871386,9.317744,9.472001,9.40636,9.051898,8.205129,7.748924,7.565129,7.6143594,7.936001,8.644924,7.532308,6.183385,6.166975,6.921847,5.7665644,4.384821,3.7087183,4.33559,4.890257,2.0217438,2.1103592,2.6453335,3.7251284,4.647385,3.9089234,3.623385,4.0041027,4.7655387,5.658257,6.485334,5.5565133,4.493129,3.7940516,3.6791797,4.089436,3.7415388,4.1091285,4.59159,4.827898,4.716308,4.414359,3.8071797,3.6627696,3.892513,3.5511796,3.1540515,3.121231,3.5840003,4.1485133,3.9253337,4.338872,4.4865646,4.4406157,4.269949,4.0500517,4.46359,4.1452312,3.8137438,3.8071797,4.082872,3.7218463,3.4658465,3.1507695,2.802872,2.6223593,2.537026,2.300718,2.0020514,1.7690258,1.7657437,2.1300514,2.6322052,2.7766156,2.537026,2.356513,2.4549747,2.740513,2.9833848,3.0654361,2.9538465,2.8160002,2.7241027,2.937436,3.43959,3.9745643,4.4832826,4.844308,4.886975,4.7917953,5.07077,5.3366156,5.3727183,5.3366156,5.297231,5.211898,5.4186673,5.152821,4.70318,4.4406157,4.8114877,5.2644105,5.2348723,5.421949,5.937231,6.308103,5.76,5.5302567,5.605744,5.671385,5.1364107,5.2742567,5.10359,4.781949,4.525949,4.6178465,4.201026,4.1452312,4.279795,4.4077954,4.33559,3.9548721,3.8531284,3.636513,3.2787695,3.1245131,3.1967182,3.1277952,2.9243078,2.6978464,2.681436,2.9440002,3.131077,3.0129232,2.5764105,2.0118976,1.654154,1.6147693,1.4834872,1.1881026,0.96492314,0.90912825,0.9353847,0.9321026,0.8992821,0.96492314,1.0436924,0.99774367,0.8369231,0.7089231,0.8992821,1.0502565,1.0502565,0.99774367,0.9616411,0.9878975,1.1060513,1.0896411,1.0108719,1.0075898,1.276718,1.4441026,1.5983591,1.7329233,1.8346668,1.9035898,1.8806155,1.910154,1.7362052,1.3587693,1.024,1.1946667,1.3522053,1.5458462,1.7624617,1.913436,2.2219489,2.1169233,2.1103592,2.284308,2.284308,2.3335385,2.8980515,3.56759,3.9581542,3.7448208,4.1714873,4.391385,4.342154,4.1189747,3.9647183,3.9023592,4.135385,4.1485133,3.8137438,3.383795,3.7776413,4.2896414,4.6178465,4.594872,4.1813335,5.0149746,4.923077,4.7950773,4.8640003,4.6834874,4.6276927,4.3618464,4.644103,5.0609236,5.4153852,5.7074876,5.8912826,6.7117953,7.3747697,7.456821,6.8988724,6.439385,6.557539,7.0957956,7.722667,7.939283,9.160206,10.866873,12.251899,13.131488,13.935591,13.965129,14.5263605,14.624822,14.299898,14.624822,14.79877,15.195899,14.887385,14.27036,15.087591,14.539488,14.660924,14.8020525,14.716719,14.555899,15.91795,15.786668,15.763694,16.443079,17.417847,17.010874,18.44513,20.358566,22.774155,27.113028,34.727386,42.525543,47.91467,49.568825,47.4519,49.014156,51.78749,55.775185,62.0078,72.52349,77.79775,66.19898,50.353233,38.495182,34.45826,30.916925,27.103182,23.653746,20.148514,15.107284,11.831796,8.582564,5.986462,4.33559,3.6069746,2.937436,2.1792822,1.5589745,1.3193847,1.6968206,1.6344616,1.0601027,0.56123084,0.30851284,0.059076928,0.036102567,0.14441027,0.20676924,0.17394873,0.108307704,0.12143591,0.1148718,0.06564103,0.006564103,0.009846155,0.04594872,0.13784617,0.23302566,0.25928208,0.13784617,0.059076928,0.026256412,0.016410258,0.02297436,0.055794876,0.059076928,0.08205129,0.06235898,0.02297436,0.072205134,0.04266667,0.013128206,0.0,0.006564103,0.016410258,0.006564103,0.0032820515,0.013128206,0.04594872,0.12471796,0.055794876,0.02297436,0.25271797,0.54482055,0.28225642,0.35774362,0.8402052,2.0906668,3.442872,3.170462,2.4057438,1.8051283,1.7657437,2.156308,2.3040001,2.6518977,2.789744,2.5009232,2.0775387,2.3072822,2.7667694,2.9636924,3.0358977,3.1770258,3.6627696,3.8104618,4.1714873,4.827898,5.402257,5.034667,5.543385,5.927385,6.813539,8.096821,8.937026,10.489437,11.286975,12.632616,14.736411,16.712206,16.577642,16.361027,15.573335,14.887385,16.141129,16.160822,16.275694,17.174976,18.661745,19.682463,19.081848,17.51959,15.983591,14.890668,14.083283,12.340514,11.346052,10.5780525,9.984001,9.984001,10.036513,10.341744,10.269539,10.033232,10.683078,12.074668,11.595488,9.941334,8.241231,8.086975,8.562873,9.42277,9.7903595,9.350565,8.333129,9.547488,9.737847,9.941334,10.597744,11.565949,12.133744,11.999181,11.58236,10.985026,9.987283,9.317744,8.067283,7.765334,8.553026,9.193027,9.373539,9.737847,9.984001,10.036513,10.059488,11.175385,11.1064625,10.9686165,11.264001,11.877745,11.234463,11.414975,11.900719,11.795693,9.82318,9.980719,10.84718,11.211488,11.1983595,12.248616,14.562463,14.053744,13.699283,13.466257,10.295795,9.997129,10.57477,12.038565,14.076719,16.04595,16.787693,16.502155,15.635694,14.585437,13.718975,14.470565,15.478155,16.20677,16.41354,16.15754,17.043694,17.417847,17.91672,18.231796,17.09949,15.261539,15.264822,15.0088215,14.516514,15.940925,16.006565,15.484719,14.388514,13.866668,16.200207,17.897026,14.8480015,12.71795,12.918155,12.62277,11.227899,10.883283,11.72677,13.059283,13.351386,14.424617,15.770258,15.560206,14.083283,13.745232,13.633642,10.637129,7.204103,4.7950773,3.8400004,3.5971284,3.6069746,3.4822567,3.18359,3.0391798,3.3280003,5.733744,6.99077,6.6560006,7.076103,5.5893335,3.9909747,3.3772311,3.4789746,2.6978464,1.8248206,1.4145643,2.0742567,2.8455386,1.2274873,1.1520001,1.522872,2.3630772,3.4756925,4.44718,6.2884107,7.0400004,7.315693,7.181129,6.166975,6.265436,6.452513,7.181129,7.9852314,7.4797955,10.039796,11.283693,9.915077,7.4765134,8.333129,13.190565,12.27159,8.907488,5.7403083,4.716308,4.95918,4.768821,5.435077,6.5903597,6.1768208,4.7425647,4.1025643,4.1846156,4.6966157,5.10359,8.621949,5.973334,3.8137438,4.0533338,3.8531284,3.0949745,1.782154,1.1881026,2.0775387,4.70318,6.87918,7.3386674,7.6176414,7.8473854,6.747898,8.411898,7.1220517,6.2555904,6.4032826,5.3727183,3.314872,3.1409233,3.7054362,4.210872,4.2141542,5.2414365,5.5138464,5.7796926,6.0291286,5.4941545,4.7589746,4.969026,6.363898,8.057437,8.027898,6.413129,6.0619493,4.9329233,3.249231,3.4822567,4.2830772,5.61559,7.0334363,7.709539,6.422975,4.9427695,3.4100516,2.5665643,2.5928206,3.0982566,3.8104618,5.2578464,6.2884107,6.550975,6.491898,3.4724104,2.7109745,2.0808206,1.0108719,0.48246157,0.50543594,0.36102566,0.2231795,0.2100513,0.3708718,0.20676924,0.16082053,0.21333335,0.32820517,0.45620516,0.62030774,0.5940513,0.571077,0.5874872,0.5284103,0.30194873,0.21333335,0.16738462,0.13456412,0.15097436,0.2100513,0.26256412,0.39056414,0.574359,0.67282057,0.6170257,0.6826667,1.0108719,1.3817437,1.1946667,1.2635899,1.8642052,2.412308,2.8160002,3.4822567,3.9844105,4.161641,4.4701543,4.8377438,4.673641,4.315898,4.650667,5.110154,5.425231,5.6287184,5.674667,5.691077,6.2687182,7.210667,7.5552826,7.456821,7.830975,8.612103,9.147078,8.198565,7.5979495,7.1844106,6.9809237,7.0432825,7.4765134,7.351795,6.8004107,6.439385,6.298257,5.8289237,5.72718,5.333334,5.0149746,4.9329233,5.0510774,5.3202057,5.4843082,6.242462,7.2270775,6.997334,6.8332314,6.7971287,7.0925136,7.512616,7.4207187,7.890052,8.224821,8.421744,8.254359,7.269744,7.177847,7.3682055,7.397744,7.2894363,7.5421543,7.6931286,7.781744,7.4929237,6.9054365,6.5083084,7.3550773,8.201847,9.019077,9.780514,10.459898,10.65354,10.125129,9.537642,9.202872,9.081436,9.124104,8.470975,7.8539495,7.8145647,8.697436,6.3179493,5.208616,6.2227697,7.9524107,6.7216415,5.2480006,5.5072823,7.003898,7.3780518,2.4024618,3.1967182,3.1409233,3.9187696,5.156103,4.414359,4.279795,4.647385,4.890257,5.0674877,5.910975,5.717334,5.179077,4.3290257,3.692308,4.2830772,4.2305646,4.4110775,4.788513,5.1364107,5.024821,4.276513,3.620103,3.2918978,3.1048207,2.4549747,2.3860514,2.5435898,3.255795,4.1813335,4.2929235,4.6276927,4.903385,4.854154,4.5423594,4.3651285,4.33559,4.5489235,4.5062566,4.210872,4.1550775,3.9975388,3.5610259,3.1048207,2.740513,2.4385643,2.3433847,2.1103592,1.9823592,2.0775387,2.3762052,2.7241027,2.8750772,2.6880002,2.3729234,2.4943593,2.9144619,3.1015387,3.255795,3.370667,3.2196925,2.8816411,2.9801028,3.318154,3.7382567,4.135385,4.601436,4.670359,4.785231,5.0051284,4.9985647,4.9329233,4.8836927,4.955898,5.142975,5.333334,5.677949,5.398975,4.7983594,4.414359,5.0018463,5.405539,5.412103,5.6976414,6.242462,6.3343596,5.9995904,5.3037953,5.028103,5.2348723,5.2545643,5.1659493,5.1954875,4.903385,4.33559,4.0336413,4.066462,3.9548721,4.017231,4.138667,3.7743592,3.6332312,3.6660516,3.4658465,3.0884104,3.045744,3.3017437,3.3575387,3.1737437,2.92759,3.0096412,3.1245131,3.2032824,3.05559,2.6354873,2.0611284,1.9462565,1.8838975,1.7362052,1.5097437,1.3193847,1.083077,1.020718,1.0699488,1.1224617,1.0371283,0.82379496,0.7089231,0.65641034,0.6662565,0.81066674,0.8041026,0.827077,0.8598975,0.8533334,0.7187693,0.7778462,0.81394875,0.8730257,1.0043077,1.2668719,1.3259488,1.5163078,1.7263591,1.8904617,2.0020514,2.0742567,2.1464617,1.9462565,1.5031796,1.1355898,1.1224617,1.2077949,1.3915899,1.6278975,1.8215386,1.972513,2.0086155,2.172718,2.4155898,2.3696413,2.740513,3.43959,4.089436,4.269949,3.5446157,3.9680004,4.414359,4.4077954,3.9548721,3.5413337,3.7809234,4.2502565,4.2601027,3.751385,3.2754874,3.43959,3.9942567,4.578462,4.84759,4.4898467,5.2545643,5.1167183,4.7983594,4.535795,4.082872,4.9427695,4.893539,5.074052,5.2348723,5.2676926,5.218462,5.5958977,6.304821,6.744616,6.7774363,6.7282057,6.7183595,6.8955903,7.3682055,7.9294367,8.086975,9.101129,10.545232,11.861334,12.849232,13.640206,13.994668,14.6871805,15.028514,15.064616,15.563488,15.015386,14.933334,15.238565,15.625848,15.563488,14.966155,14.578873,14.578873,14.752822,14.496821,15.143386,15.074463,15.399385,16.170668,16.403694,16.672821,18.7799,20.795078,23.082668,28.320822,34.36308,42.866875,49.440823,51.003082,45.791183,50.087387,55.821133,62.53621,70.21621,79.30093,72.61211,59.375595,47.632416,40.756516,37.461338,32.99118,30.237541,26.73231,22.393438,19.50195,15.632411,11.851488,8.848411,6.744616,5.097026,3.7054362,2.6256413,2.0676925,2.0151796,2.1956925,1.5392822,1.1158975,0.79425645,0.47261542,0.108307704,0.04594872,0.15753847,0.18379489,0.08533334,0.06235898,0.12143591,0.08205129,0.03938462,0.032820515,0.04594872,0.13128206,0.20676924,0.21333335,0.15097436,0.07548718,0.026256412,0.016410258,0.016410258,0.01969231,0.029538464,0.10502565,0.12143591,0.072205134,0.0,0.0,0.0,0.0,0.006564103,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.026256412,0.07548718,0.06564103,0.032820515,0.25271797,0.7187693,1.1585642,1.4998976,1.8051283,3.0391798,4.0369234,1.5097437,2.0841026,2.0709746,2.103795,2.3171284,2.3663592,3.6102567,3.2984617,2.7175386,2.6256413,3.2361028,3.7710772,4.069744,4.1747694,4.2830772,4.7622566,4.138667,5.5565133,5.989744,5.3398976,6.439385,5.8518977,6.3277955,7.397744,8.996103,11.474052,13.633642,14.605129,14.592001,14.171899,14.283488,13.952001,13.3940525,12.675283,12.980514,16.617027,17.496616,16.771284,16.131283,16.226463,16.679386,15.238565,14.237539,13.636924,13.157744,12.251899,12.032001,11.933539,11.651283,11.024411,10.010257,9.924924,9.829744,9.468719,9.317744,10.57477,10.292514,9.947898,9.3078985,8.562873,8.329846,7.9294367,9.219283,10.404103,10.371283,8.713847,9.114257,9.527796,10.026668,10.722463,11.749744,12.49477,11.98277,11.191795,10.476309,9.596719,9.07159,8.264206,8.021334,8.372514,8.546462,8.372514,9.163487,10.121847,10.729027,10.742155,11.976206,11.936821,11.592206,11.510155,11.841642,10.827488,10.548513,10.509129,10.276103,9.4457445,9.800206,10.345026,10.509129,10.456616,11.076924,12.580104,12.242052,13.1872835,14.546052,11.444513,10.735591,11.510155,13.069129,15.081027,17.608206,17.266872,16.768002,16.091898,15.317334,14.634667,14.680616,15.507693,16.338053,16.610462,15.977027,16.597334,17.46708,17.890463,17.503181,16.282257,15.780104,16.111591,15.832617,15.038361,15.379693,15.894976,16.039387,15.081027,14.185027,16.416822,18.067694,15.914668,13.804309,12.87877,11.595488,12.632616,12.911591,12.954257,13.180719,13.899488,14.486976,16.170668,16.603899,15.563488,14.953027,13.673027,10.834052,7.5487185,4.962462,4.240411,4.352,4.2601027,4.066462,3.7973337,3.4166157,3.1015387,5.8223596,6.994052,6.052103,6.4557953,5.940513,4.276513,2.9505644,3.2722054,6.3474874,2.806154,1.7033848,2.9407182,4.460308,2.228513,1.5195899,1.7099489,2.678154,4.0434875,5.142975,6.692103,7.5454364,8.034462,8.024616,6.9120007,7.3025646,7.702975,6.806975,5.549949,7.125334,7.076103,8.474257,8.766359,8.444718,11.030975,12.265027,10.660104,7.322257,3.8104618,2.1530259,2.1989746,2.9997952,4.023795,4.906667,5.431795,5.4941545,5.8092313,4.9132314,3.259077,3.2361028,6.3343596,5.5072823,4.2338467,3.9778464,4.197744,2.8422565,1.7624617,1.5524104,2.2744617,3.4330258,4.59159,5.671385,4.9493337,3.5511796,5.4153852,5.1364107,3.5741541,4.201026,6.557539,6.23918,4.1517954,3.2853336,4.1025643,5.8978467,6.7905645,7.584821,7.2336416,6.5805135,6.5444107,8.116513,6.944821,5.536821,4.4077954,4.0467696,4.9132314,4.1189747,2.9702566,2.3335385,2.4681027,3.006359,3.8367183,5.901129,7.5979495,7.9261546,6.485334,5.618872,4.4964104,3.239385,2.609231,4.013949,4.7458467,6.521436,7.2303596,6.5017443,5.720616,3.2689233,2.1891284,1.4145643,0.6892308,0.58092314,0.45620516,0.43651286,0.380718,0.3117949,0.39712822,0.24943592,0.15097436,0.16738462,0.25928208,0.25928208,0.5513847,0.58092314,0.5546667,0.5513847,0.5021539,0.35774362,0.256,0.17066668,0.1148718,0.15097436,0.190359,0.28225642,0.34789747,0.41682056,0.6268718,0.6859488,0.79425645,1.024,1.2832822,1.2832822,1.3784616,1.9790771,2.4943593,2.8356924,3.4330258,3.895795,4.0500517,4.197744,4.391385,4.4406157,4.2207184,4.630975,5.2414365,5.858462,6.5312824,7.88677,7.381334,6.6428723,6.616616,7.568411,7.9458466,8.280616,8.864821,9.284924,8.408616,7.3091288,7.1089234,7.131898,7.0990777,7.1122055,7.8539495,7.785026,7.4141545,7.02359,6.6822567,6.121026,6.301539,6.4656415,6.294975,5.904411,5.930667,5.907693,6.409847,7.253334,7.522462,7.0465646,6.5805135,6.4754877,6.7150774,6.8955903,7.0432825,7.3649235,7.686565,7.7325134,7.1122055,6.8529234,6.5706673,6.124308,5.76,6.088206,6.4557953,6.957949,7.141744,7.02359,7.0957956,7.3747697,7.9786673,9.107693,10.469745,11.277129,11.667693,10.712616,9.649232,9.202872,9.5835905,9.449026,9.176616,9.048616,9.101129,9.124104,5.5729237,4.197744,5.1200004,7.1122055,7.6143594,4.8311796,5.32677,5.802667,5.221744,4.8049235,4.0008206,2.665026,3.0358977,4.6802053,4.4865646,4.414359,5.218462,5.2414365,4.5817437,5.080616,5.179077,5.35959,4.9920006,4.4438977,5.0674877,4.84759,4.9099493,5.287385,5.3398976,3.754667,2.7044106,3.0194874,3.5478978,3.4921029,2.3794873,2.1366155,2.8717952,3.9286156,4.7950773,5.110154,6.0028725,6.088206,5.543385,4.827898,4.670359,4.4865646,4.650667,4.827898,4.8049235,4.4865646,4.8147697,4.082872,3.2886157,2.8422565,2.546872,2.3171284,2.2678976,2.3893335,2.5961027,2.7306669,2.806154,2.5928206,2.3433847,2.284308,2.6387694,3.0916924,2.8291285,2.8488207,3.2065644,3.0358977,2.806154,3.3411283,3.9023592,4.197744,4.378257,4.46359,4.394667,4.601436,5.0116925,5.034667,4.900103,4.821334,4.8640003,4.969026,4.9427695,5.0904617,4.844308,4.3684106,4.0008206,4.2568207,5.0510774,5.110154,5.221744,5.737026,6.5903597,6.810257,5.970052,5.113436,4.71959,4.670359,5.402257,5.7665644,5.6943593,5.218462,4.4865646,4.352,4.089436,4.0336413,4.1058464,3.8006158,3.629949,3.6036925,3.4100516,3.1540515,3.387077,3.1540515,3.1245131,3.308308,3.508513,3.3280003,3.117949,2.8849232,2.6518977,2.4615386,2.3663592,2.2908719,2.162872,2.097231,1.9889232,1.5261539,1.1355898,1.1651284,1.2570257,1.2570257,1.2209232,0.97805136,0.8795898,0.77456415,0.6892308,0.82379496,1.0305642,1.0929232,0.9944616,0.8402052,0.8402052,0.85005134,0.69907695,0.67282057,0.81394875,0.8992821,0.75487185,1.2307693,1.7165129,1.9790771,2.1366155,2.294154,2.353231,2.2186668,1.8182565,1.0994873,1.0371283,1.1323078,1.4933335,1.9331284,1.9692309,2.1891284,2.3696413,2.6157951,2.8816411,2.989949,3.4297438,3.8334363,4.023795,3.895795,3.4330258,3.5544617,3.7776413,3.7973337,3.698872,3.9680004,4.785231,5.3103595,5.218462,4.325744,2.5796926,3.3476925,3.9614363,4.388103,4.6834874,4.9887185,5.159385,5.5236926,5.4186673,5.0609236,5.5236926,4.8082056,5.10359,5.2512827,5.2578464,5.284103,5.6451287,5.7501545,6.265436,6.8233852,7.2172313,7.4141545,6.9809237,7.515898,7.958975,8.083693,8.513641,9.409642,10.57477,11.595488,12.294565,12.724514,12.649027,13.236514,14.342566,15.474873,15.770258,14.752822,14.25395,14.39836,14.969437,15.40595,14.828309,14.562463,14.582155,14.772514,14.936617,15.543797,16.410257,17.106052,17.23077,16.426668,18.884924,20.54236,21.494156,23.194258,28.478361,34.589542,41.186466,45.2759,45.968414,44.48493,54.767593,60.944416,64.288826,65.01744,62.283493,51.06544,40.438156,32.16739,26.863592,23.998362,22.35077,20.946053,19.761232,18.730669,17.729643,15.629129,12.891898,10.525539,8.635077,6.439385,4.969026,3.7809234,2.8980515,2.3893335,2.3696413,1.463795,0.86646163,0.47917953,0.24287182,0.13128206,0.029538464,0.03938462,0.04266667,0.026256412,0.06235898,0.08205129,0.068923086,0.0951795,0.13128206,0.04594872,0.24943592,0.318359,0.24943592,0.12143591,0.07548718,0.055794876,0.036102567,0.02297436,0.016410258,0.01969231,0.08205129,0.08205129,0.049230773,0.009846155,0.0,0.0,0.0,0.009846155,0.02297436,0.0032820515,0.013128206,0.74830776,1.2635899,1.522872,2.3696413,2.172718,1.5327181,1.5425643,2.1792822,2.3072822,2.9210258,2.8488207,3.0162053,3.2229745,2.1333334,2.7175386,1.910154,2.0217438,3.0391798,2.609231,3.639795,3.6332312,4.2305646,5.349744,5.1987696,4.3716927,4.6867695,4.844308,4.6080003,4.821334,4.7458467,4.955898,5.5597954,6.2490263,6.2916927,5.8420515,7.204103,9.737847,12.530872,14.404924,15.051488,14.76595,14.454155,14.588719,15.186052,13.692719,12.685129,12.163283,12.790154,15.872002,16.75159,17.243898,16.79754,15.812924,15.638975,14.923489,14.716719,13.797745,12.3076935,11.766154,11.067078,11.073642,11.323078,11.434668,11.083488,10.089026,9.527796,9.019077,8.720411,9.304616,9.728001,9.813334,9.852718,9.8363085,9.478565,8.989539,9.321027,10.016821,10.663385,10.896411,10.978462,10.988309,11.126155,11.575796,12.49477,12.153437,11.864616,11.119591,10.105436,9.69518,9.120821,8.6580515,8.464411,8.507077,8.582564,8.214975,8.372514,9.373539,10.761847,11.290257,12.212514,12.363488,12.028719,11.500309,11.096616,10.364718,9.754257,9.337437,9.005949,8.467693,9.222565,9.475283,9.849437,10.604308,11.628308,12.484924,12.937847,15.1466675,16.489027,9.540924,9.055181,11.336206,14.27036,16.597334,17.913437,18.031591,17.408,16.810667,16.374155,15.573335,15.133539,16.101746,16.922258,16.768002,15.55036,16.01641,16.961643,17.27672,16.70236,15.852309,15.947489,15.983591,15.619284,14.976001,14.624822,16.170668,17.076513,16.292105,15.235283,17.762463,19.895796,18.884924,16.938667,14.949745,12.488206,14.336001,15.087591,15.251694,15.337027,15.842463,14.582155,15.635694,16.538258,16.33477,15.589745,12.763899,9.941334,7.778462,6.3212314,5.034667,5.106872,4.2436924,4.066462,4.3716927,3.1113849,6.4557953,6.8365135,5.9963083,5.110154,4.781949,5.421949,4.086154,3.0260515,4.381539,10.194052,5.832206,3.190154,3.5347695,5.47118,4.9362054,2.0512822,1.9167181,3.1638978,4.647385,5.435077,6.498462,7.4929237,7.6996927,7.020308,5.9963083,7.890052,8.192,7.709539,6.6461544,4.598154,4.647385,5.4186673,8.802463,12.586668,10.459898,7.8047185,6.803693,6.4032826,6.11118,5.98318,3.5905645,3.1277952,3.5774362,4.1714873,4.381539,7.499488,6.8299494,5.366154,5.5991797,9.521232,12.301129,8.900924,4.916513,3.4888208,5.3202057,4.06318,2.9407182,2.1333334,1.8379488,2.284308,4.7655387,4.069744,4.1485133,5.21518,3.7316926,5.5696416,6.12759,5.622154,4.9526157,5.677949,4.821334,3.2196925,3.255795,5.330052,7.8506675,7.141744,5.4482055,4.7425647,5.3858466,6.1407185,6.432821,7.4174366,6.488616,4.315898,4.841026,6.301539,4.962462,3.4921029,3.0851285,3.4560003,3.2918978,4.7360005,6.2916927,6.9349747,6.117744,5.907693,5.1298466,3.7448208,2.7503593,4.1846156,6.058667,7.5421543,7.8539495,6.928411,5.405539,3.9286156,2.5271797,1.3751796,0.69579494,0.761436,0.56123084,0.38400003,0.27569234,0.26584616,0.3708718,0.21661541,0.128,0.17066668,0.26584616,0.18707694,0.39056414,0.39712822,0.41025645,0.446359,0.30851284,0.30851284,0.3249231,0.25928208,0.14441027,0.15097436,0.20020515,0.2855385,0.31507695,0.30851284,0.41682056,0.55794877,0.69251287,0.8008206,0.8795898,0.9288206,1.2012309,1.8018463,2.294154,2.6945643,3.4560003,3.9614363,4.1682053,4.240411,4.378257,4.818052,4.6867695,5.179077,5.83877,6.554257,7.5552826,8.356103,7.719385,7.181129,7.24677,7.397744,7.6209235,8.008205,8.280616,8.303591,8.077128,6.987488,6.439385,6.2030773,6.2752824,6.8529234,7.7259493,7.762052,7.768616,7.817847,7.2336416,6.9842057,7.3649235,7.4075904,7.066257,7.2237954,7.512616,7.0367184,6.5411286,6.4689236,6.961231,6.9743595,6.5837955,6.436103,6.51159,6.12759,6.4000006,6.547693,6.6560006,6.8299494,7.1844106,7.0137444,6.636308,6.23918,5.976616,5.9536414,5.7435904,6.045539,6.3442054,6.432821,6.4000006,6.5936418,7.0925136,7.7357955,8.448001,9.225847,10.368001,10.151385,9.645949,9.481847,9.849437,9.219283,9.590155,10.029949,9.987283,9.3078985,6.5936418,4.5456414,4.824616,6.5017443,6.0750775,2.9210258,4.1583595,4.6112823,3.446154,4.1846156,3.1540515,2.1202054,2.176,3.0654361,3.1934361,4.2601027,4.8705645,4.972308,4.6834874,4.276513,4.138667,4.1058464,4.135385,4.322462,4.893539,4.529231,4.8705645,4.781949,4.2371287,4.338872,4.529231,4.06318,3.4034874,2.8750772,2.674872,2.2547693,2.865231,3.8662567,5.0543594,6.6625648,5.989744,5.933949,5.668103,5.0609236,4.670359,4.4865646,4.585026,4.713026,4.647385,4.194462,3.889231,3.3772311,2.917744,2.6518977,2.6322052,2.481231,2.356513,2.3860514,2.546872,2.681436,2.6387694,2.5895386,2.6617439,2.7733335,2.6387694,2.7011285,2.4516926,2.4549747,2.7733335,2.9636924,3.259077,3.7874875,3.9581542,3.882667,4.378257,4.7589746,4.857436,5.225026,5.7829747,5.8157954,5.35959,4.95918,4.7917953,4.84759,4.919795,4.772103,4.4077954,4.0402055,3.9351797,4.414359,5.159385,5.546667,5.622154,5.654975,6.12759,6.5345645,5.796103,4.8771286,4.3552823,4.4242053,5.0510774,5.35959,5.4613338,5.3398976,4.850872,4.1911798,4.007385,4.125539,4.2305646,3.895795,3.8038976,3.69559,3.3641028,3.0227695,3.314872,2.92759,2.865231,3.186872,3.564308,3.2525132,3.1638978,2.5993848,2.225231,2.28759,2.609231,2.3991797,2.1497438,2.0086155,1.8937438,1.4769232,1.1454359,1.3587693,1.3686155,1.0535386,0.9288206,0.90912825,0.8730257,0.8533334,0.8598975,0.8960001,1.0272821,1.1552821,1.1224617,1.020718,1.204513,0.98461545,0.764718,0.78769237,1.0010257,1.0469744,0.9485129,1.3718976,1.6804104,1.7690258,2.0644104,2.3302567,2.172718,1.7887181,1.3357949,0.9288206,0.7778462,1.0929232,1.595077,1.9626669,1.8346668,2.1792822,2.5698464,2.8488207,3.0720003,3.501949,4.020513,4.3716927,4.5554876,4.565334,4.384821,4.3618464,4.312616,4.125539,3.876103,3.8334363,3.8990772,4.066462,4.0500517,3.6562054,2.7995899,3.0391798,3.639795,4.384821,5.034667,5.330052,5.100308,5.028103,5.0904617,4.9854364,4.1189747,4.601436,4.893539,4.962462,5.225026,5.5630774,5.3234878,5.7403083,6.242462,6.8955903,7.634052,8.234667,7.6242056,7.581539,7.4863596,7.3616414,7.906462,8.92718,10.033232,10.8996935,11.487181,12.058257,12.694975,13.443283,14.431181,15.353437,15.465027,14.441027,14.204719,14.408206,14.746258,14.9628725,15.179488,14.818462,14.834873,15.537232,16.57436,16.761436,17.168411,16.984617,16.544823,17.322668,19.856411,21.38913,22.629745,24.848412,29.88308,36.785233,43.81867,47.458466,48.643288,52.772106,65.63775,68.73272,63.169647,53.454773,47.501133,39.624207,32.17067,25.504822,20.33231,17.683693,17.073233,15.43877,14.020925,13.105232,12.015591,10.794667,9.77395,8.484103,6.9677954,5.786257,4.955898,4.141949,3.3772311,2.737231,2.3663592,1.591795,0.94523084,0.512,0.27241027,0.101743594,0.049230773,0.036102567,0.036102567,0.036102567,0.032820515,0.068923086,0.12143591,0.17723078,0.19364104,0.118153855,0.2986667,0.39712822,0.33805132,0.17394873,0.0951795,0.098461546,0.068923086,0.04266667,0.032820515,0.02297436,0.055794876,0.068923086,0.04594872,0.0032820515,0.0,0.0,0.0,0.0032820515,0.013128206,0.009846155,1.595077,1.4966155,1.3357949,1.595077,1.6278975,1.1913847,1.3193847,2.1202054,3.0424619,2.8422565,2.5665643,2.993231,3.6758976,4.1550775,3.9745643,2.5074873,1.9823592,2.4320002,3.2000003,2.934154,3.370667,3.5347695,4.332308,5.7665644,6.9645133,5.477744,5.8223596,6.377026,6.6428723,7.2369237,6.314667,6.2129235,6.5706673,6.7314878,5.7435904,6.8955903,8.704,11.300103,14.099693,15.80636,15.179488,15.340309,15.589745,15.832617,16.548103,15.028514,14.112822,13.449847,13.279181,14.450873,15.730873,15.980309,14.976001,13.66318,14.145642,14.641232,13.860104,12.373334,11.172104,11.67754,12.274873,11.254155,10.640411,11.132719,12.120616,10.79795,10.010257,9.468719,9.193027,9.4916935,10.171078,10.482873,10.59118,10.482873,9.96759,9.432616,9.429334,9.819899,10.601027,11.910565,11.221334,10.512411,10.390975,10.988309,11.96636,11.949949,12.097642,11.500309,10.35159,9.947898,9.603283,8.812308,8.254359,8.201847,8.500513,8.214975,8.51036,9.403078,10.555078,11.273847,11.493745,11.779283,11.47077,10.79795,10.893129,10.482873,9.8363085,9.170052,8.6580515,8.444718,8.487385,8.641642,9.324308,10.499283,11.680821,12.225642,12.754052,13.275898,14.208001,16.367592,8.963283,10.200616,13.564719,15.842463,17.112617,18.002052,17.473642,17.06995,17.014154,16.193642,15.645539,16.25272,16.876308,16.748308,15.468308,15.9343605,16.981335,17.42113,16.889437,15.849027,16.324924,15.82277,14.959591,14.273643,14.224411,16.600616,18.17272,17.030565,15.074463,17.99549,20.246977,20.539078,18.871796,15.803078,12.471796,14.7790785,16.538258,17.243898,17.306257,18.021746,16.489027,16.649847,17.217642,17.09949,15.379693,11.306667,8.51036,6.892308,6.1013336,5.536821,5.0477953,4.634257,4.516103,4.650667,4.7491283,7.6668725,6.9842057,5.428513,4.391385,3.9154875,6.4754877,5.146257,3.2295387,3.876103,10.056206,7.6734366,5.7731285,7.1122055,9.16677,4.1517954,2.1792822,2.297436,3.3247182,4.345436,4.7294364,6.6067696,7.5487185,7.7292314,6.744616,3.626667,5.428513,5.87159,6.2063594,6.180103,4.0303593,3.7021542,4.1813335,6.157129,8.986258,10.709334,6.3212314,4.525949,3.9844105,4.397949,6.521436,4.4110775,3.9680004,4.637539,5.549949,5.5007186,4.70318,6.314667,6.0028725,4.141949,5.8125134,8.201847,6.0061545,3.4822567,2.6847181,3.4756925,2.7995899,2.225231,1.7362052,1.8051283,3.3903592,7.0990777,6.2030773,5.7074876,6.3967185,4.8311796,5.228308,6.0980515,6.2227697,5.5204105,5.044513,4.086154,2.7306669,3.0293336,5.1889234,7.578257,6.9809237,6.048821,5.474462,5.602462,6.422975,6.058667,7.076103,6.8627696,5.293949,4.7655387,6.3179493,6.0685134,4.8771286,3.7842054,4.020513,4.138667,4.9132314,5.979898,6.7282057,6.265436,5.609026,4.394667,2.9210258,2.15959,3.7218463,6.038975,7.171283,7.0465646,5.973334,4.667077,3.9384618,2.7044106,1.5097437,0.7253334,0.571077,0.47589746,0.2986667,0.16738462,0.14112821,0.19364104,0.1148718,0.13128206,0.15753847,0.20020515,0.3511795,0.37415388,0.39384618,0.4397949,0.44964105,0.27897438,0.23958977,0.21989745,0.21989745,0.21989745,0.15097436,0.18051283,0.23302566,0.25271797,0.25928208,0.33805132,0.4594872,0.58092314,0.6465641,0.67282057,0.74830776,1.1323078,1.8412309,2.5074873,3.0162053,3.5282054,3.8367183,4.06318,4.197744,4.3060517,4.565334,4.827898,5.7140517,6.6395903,7.5913854,9.130668,8.648206,8.024616,7.9228725,8.064001,7.207385,7.6242056,7.8408213,7.906462,7.9097443,7.958975,7.568411,7.0334363,6.6034875,6.38359,6.3507695,6.931693,7.4075904,7.702975,7.7456417,7.4436927,7.571693,7.755488,7.6734366,7.3649235,7.243488,7.2894363,6.951385,6.452513,6.0947695,6.2720003,6.616616,6.626462,6.557539,6.5017443,6.3573337,6.7216415,6.8004107,6.616616,6.436103,6.770872,6.633026,6.4689236,6.370462,6.2129235,5.664821,5.3169236,5.546667,5.914257,6.157129,6.196513,6.1341543,6.170257,6.449231,7.0826674,8.136206,9.334154,9.603283,9.645949,9.882257,10.43036,9.53436,10.358154,11.001437,10.121847,6.944821,6.370462,5.58277,5.622154,5.7698464,3.5577438,5.7534366,5.07077,3.170462,1.7493335,2.5271797,2.2383592,2.156308,2.162872,2.2153847,2.3269746,4.3060517,4.59159,4.4012313,4.210872,3.7448208,2.737231,3.0129232,3.4297438,3.5478978,3.626667,4.388103,5.156103,4.7360005,3.9844105,5.805949,5.3891287,4.450462,3.4231799,2.7109745,2.6551797,2.228513,2.8947694,4.0041027,5.172513,6.2818465,5.5105643,5.609026,5.5269747,5.156103,5.32677,5.5171285,5.546667,5.421949,5.093744,4.457026,3.8400004,3.4560003,2.9768207,2.4713848,2.4155898,2.3204105,2.3991797,2.5107694,2.5993848,2.6978464,2.8521028,2.7831798,2.9013336,3.1507695,3.0326157,2.8717952,2.737231,2.868513,3.255795,3.639795,3.751385,3.9548721,3.9778464,3.9220517,4.269949,4.706462,4.962462,5.32677,5.6451287,5.3431797,5.2020516,5.3202057,5.2644105,5.093744,5.3431797,5.2709746,5.172513,4.965744,4.7655387,4.886975,5.6418467,6.557539,6.8529234,6.436103,5.920821,5.4416413,5.3760004,5.149539,4.7524104,4.7392826,5.080616,5.182359,5.4580517,5.717334,5.1364107,4.4734364,3.9942567,3.9089234,3.9811285,3.5380516,3.7054362,3.7415388,3.3772311,2.8849232,3.1048207,3.114667,3.2820516,3.6430771,3.817026,3.0162053,2.8816411,2.5009232,2.2580514,2.2744617,2.4320002,2.8750772,2.6486156,2.1956925,1.7952822,1.5392822,1.2635899,1.3653334,1.3259488,1.0699488,0.9353847,1.083077,1.0929232,1.1093334,1.1684103,1.1815386,1.1946667,1.2471796,1.1684103,1.0305642,1.1224617,0.85005134,0.71548724,0.8172308,1.0272821,0.98133343,1.3161026,1.7296412,1.8051283,1.654154,1.9167181,2.0841026,1.6836925,1.3095386,1.1388719,0.9485129,0.8598975,1.2800001,1.8379488,2.1891284,2.048,2.353231,2.6715899,2.9078977,3.1803079,3.82359,4.2207184,4.4832826,4.640821,4.699898,4.630975,4.7622566,4.8311796,4.713026,4.3618464,3.8006158,3.7152824,3.6430771,3.9351797,4.1091285,2.8521028,2.868513,3.5314875,4.5587697,5.4843082,5.674667,5.1298466,5.3792825,5.5729237,5.2414365,4.273231,4.332308,4.493129,4.634257,5.031385,5.435077,5.077334,5.7534366,6.518154,7.273026,7.9917955,8.73354,8.060719,7.427283,7.1581545,7.3419495,7.8473854,8.753231,9.7903595,10.604308,11.158976,11.697231,12.724514,13.433437,14.070155,14.575591,14.592001,14.17518,14.572309,15.018668,15.0777445,14.63795,15.0088215,14.582155,14.720001,15.78995,17.178257,17.532719,17.312822,16.66954,16.564514,18.756924,20.420925,22.537848,25.232412,28.612925,32.768,40.795902,49.529438,54.564106,56.98298,63.379696,71.34196,67.36739,55.67016,42.768414,37.461338,32.512,27.024412,21.254566,16.262566,13.909334,12.337232,10.102155,8.237949,7.066257,6.1997952,5.914257,5.85518,5.435077,4.7360005,4.493129,4.266667,3.7710772,3.190154,2.6420515,2.176,1.6082052,1.0272821,0.5874872,0.3117949,0.101743594,0.098461546,0.07548718,0.055794876,0.049230773,0.04594872,0.068923086,0.15753847,0.23302566,0.27569234,0.31507695,0.36758977,0.45292312,0.4397949,0.3052308,0.13784617,0.12143591,0.098461546,0.08205129,0.072205134,0.049230773,0.108307704,0.12143591,0.072205134,0.0,0.006564103,0.009846155,0.009846155,0.006564103,0.006564103,0.009846155,1.6804104,1.204513,0.9682052,1.2964103,0.45620516,0.47917953,0.955077,1.8674873,2.8947694,3.4034874,2.2613335,2.6584618,3.2164104,3.3969233,3.4724104,2.041436,2.0020514,2.3729234,2.6256413,2.674872,2.737231,3.058872,3.4855387,4.1058464,5.2447186,4.8311796,5.6418467,6.99077,8.27077,8.986258,7.6996927,7.3485136,6.8988724,6.11118,5.5171285,7.427283,9.7673855,12.33395,14.742975,16.439796,15.107284,15.333745,16.039387,16.646564,17.096207,16.377438,15.327181,14.6642065,14.411489,13.899488,14.739694,14.693745,14.171899,13.873232,14.792206,15.14995,13.961847,12.47836,11.707078,12.406155,13.860104,12.672001,11.713642,11.923694,12.288001,11.109744,10.679795,10.423796,10.213744,10.374565,11.073642,11.405129,11.355898,10.939077,10.194052,9.488411,9.688616,10.387693,11.300103,12.27159,11.080206,10.075898,9.764103,10.223591,11.1294365,11.943385,11.858052,11.116308,10.308924,10.371283,10.28595,9.544206,8.763078,8.251078,8.011488,7.824411,8.392206,9.271795,10.036513,10.272821,10.325335,10.515693,10.315488,9.90195,10.148104,10.249847,9.875693,9.232411,8.576,8.198565,8.011488,8.218257,9.258667,10.758565,11.529847,11.930258,12.2157955,12.658873,13.709129,16.003283,8.402052,9.508103,12.553847,14.592001,16.505438,17.637745,16.964924,16.567797,16.807386,16.328207,16.213335,16.597334,16.81395,16.466053,15.425642,16.01313,17.174976,17.929848,17.769028,16.682669,17.122463,16.170668,15.126975,14.575591,14.401642,16.403694,17.670565,16.57436,14.788924,17.283283,18.73395,19.226257,18.070976,15.425642,12.301129,14.408206,16.905848,18.33354,18.789745,19.954874,19.301744,18.340103,17.723078,17.050259,14.844719,10.896411,8.3134365,6.692103,5.858462,5.8945646,5.211898,4.9329233,4.5489235,4.568616,6.5378466,7.6701546,6.705231,5.044513,3.6594875,3.0916924,6.774154,6.183385,4.6112823,4.5095387,7.463385,7.7357955,8.050873,8.900924,8.448001,2.556718,2.1858463,2.546872,3.3017437,4.197744,5.0543594,7.315693,8.198565,8.352821,7.069539,2.2580514,3.3017437,3.8400004,4.4832826,4.962462,4.1156926,3.495385,3.879385,4.273231,5.2053337,8.730257,5.208616,3.564308,2.92759,3.239385,5.2512827,4.2305646,4.4373336,5.284103,6.055385,5.874872,3.9384618,7.1844106,8.349539,6.2227697,5.6254363,5.543385,3.9154875,3.0358977,3.2853336,3.1343591,2.9768207,3.3345644,3.5610259,3.9909747,5.9470773,7.0826674,5.796103,5.0674877,5.3727183,4.6900516,4.6211286,4.9394875,5.5236926,5.737026,4.420923,3.6102567,2.809436,3.6036925,6.091488,8.89436,8.041026,7.6143594,6.8562055,6.1505647,7.017026,6.3376417,6.377026,6.373744,5.9667697,5.225026,5.208616,5.179077,4.4832826,3.4756925,3.5314875,4.397949,5.421949,6.301539,6.774154,6.6494365,5.3398976,3.383795,1.9561027,1.8904617,3.698872,5.5696416,6.1440005,5.730462,4.926359,4.6112823,3.761231,2.5140514,1.3883078,0.6662565,0.3708718,0.30194873,0.18379489,0.08861539,0.06235898,0.11158975,0.06564103,0.118153855,0.14112821,0.17066668,0.39384618,0.3314872,0.35774362,0.40369233,0.39384618,0.2297436,0.17394873,0.128,0.15425642,0.2100513,0.14112821,0.14769232,0.19692309,0.2231795,0.23958977,0.30851284,0.39712822,0.5218462,0.58092314,0.5874872,0.6629744,1.2603078,1.9396925,2.8455386,3.7185643,3.8990772,3.754667,3.9253337,4.1583595,4.312616,4.345436,4.9329233,6.439385,7.6242056,8.277334,9.216001,8.595693,8.218257,8.280616,8.39877,7.6242056,7.650462,7.5552826,7.525744,7.64718,7.893334,7.765334,7.256616,6.73477,6.3310776,5.937231,6.3507695,7.0925136,7.5552826,7.637334,7.7292314,7.7718983,7.709539,7.5388722,7.3025646,7.1122055,6.921847,6.8430777,6.7216415,6.426257,5.8486156,6.242462,6.416411,6.363898,6.226052,6.294975,6.567385,6.820103,6.73477,6.413129,6.413129,6.229334,6.265436,6.2523084,6.012718,5.4613338,5.1167183,5.172513,5.540103,6.0061545,6.245744,6.121026,5.989744,6.11118,6.616616,7.512616,8.487385,9.035488,9.344001,9.688616,10.436924,10.151385,10.8767185,11.221334,9.898667,5.7632823,6.7905645,6.416411,5.586052,5.549949,7.8736415,7.6767187,4.5587697,2.5042052,2.3827693,1.9528207,2.422154,2.8160002,2.4024618,1.719795,2.5731285,3.8038976,3.8498464,3.7743592,3.7973337,3.318154,1.9068719,2.412308,3.0129232,3.0851285,3.1606157,4.017231,4.857436,4.6112823,4.027077,5.651693,5.284103,3.9712822,2.802872,2.3335385,2.5928206,2.1234872,2.737231,3.817026,4.84759,5.4449234,4.9296412,5.156103,5.346462,5.431795,6.0356927,6.567385,6.5312824,6.189949,5.658257,4.896821,3.948308,3.5544617,3.121231,2.5698464,2.349949,2.3204105,2.4549747,2.5862565,2.6715899,2.7831798,2.930872,2.878359,3.0654361,3.4231799,3.370667,3.18359,3.2295387,3.4592824,3.8104618,4.1846156,4.1091285,4.1846156,4.269949,4.2929235,4.2338467,4.571898,4.926359,5.225026,5.353026,5.1298466,5.2676926,5.691077,5.717334,5.3825645,5.4547696,5.5565133,5.6320004,5.4547696,5.0215387,4.568616,5.146257,6.311385,6.9809237,6.813539,6.170257,5.4416413,5.4383593,5.3760004,5.110154,5.1232824,5.3202057,5.297231,5.6451287,6.0980515,5.549949,5.1856413,4.630975,4.33559,4.204308,3.5971284,3.6135387,3.623385,3.2984617,2.8488207,3.0358977,3.1606157,3.4822567,3.8104618,3.7776413,2.8389745,2.6322052,2.5074873,2.3958976,2.2908719,2.231795,3.006359,2.8356924,2.2482052,1.6935385,1.5195899,1.3915899,1.3161026,1.211077,1.0601027,0.9189744,1.1815386,1.2865642,1.3522053,1.4112822,1.4145643,1.4145643,1.3686155,1.2274873,1.0404103,0.9517949,0.7778462,0.7844103,0.94523084,1.1355898,1.1355898,1.6082052,1.9298463,1.9561027,1.8576412,2.1103592,2.041436,1.4834872,1.1060513,1.0568206,0.97805136,1.0732309,1.6049232,2.166154,2.4910772,2.4582565,2.5665643,2.5928206,2.737231,3.1540515,3.9351797,4.1517954,4.338872,4.453744,4.5062566,4.5456414,4.699898,4.7458467,4.7360005,4.5390773,3.8432825,3.8629746,3.6036925,3.639795,3.7218463,2.7667694,3.2032824,3.7809234,4.5817437,5.362872,5.5696416,4.7589746,5.0904617,5.293949,4.9952826,4.706462,4.1058464,4.082872,4.2962055,4.525949,4.7360005,5.0674877,5.805949,6.921847,7.8047185,8.326565,8.838565,8.188719,7.397744,7.3616414,8.04759,8.480822,9.107693,9.944616,10.755282,11.355898,11.605334,12.291283,12.770463,13.22995,13.607386,13.59754,14.217847,15.169642,15.793232,15.694771,14.76595,14.575591,14.244103,14.605129,15.711181,16.853334,17.499899,16.978052,16.761436,17.77559,20.404514,21.779694,24.871386,29.075695,33.57867,37.35631,48.01313,58.899696,65.92657,69.57949,74.922676,72.03118,59.17539,45.99795,37.4679,33.86749,28.393028,22.912003,17.43754,12.796719,10.6469755,7.604513,5.208616,3.5774362,2.7470772,2.674872,3.3542566,3.2787695,3.2262566,3.387077,3.3772311,3.314872,2.8553848,2.356513,1.9889232,1.7591796,1.3883078,0.9485129,0.5415385,0.24943592,0.12143591,0.15425642,0.128,0.07876924,0.052512825,0.108307704,0.128,0.18379489,0.27241027,0.38400003,0.508718,0.42338464,0.4397949,0.44964105,0.3708718,0.15753847,0.128,0.16410258,0.16738462,0.12471796,0.0951795,0.17394873,0.16738462,0.09189744,0.006564103,0.013128206,0.02297436,0.01969231,0.02297436,0.04594872,0.06235898,0.22646156,0.34789747,0.75487185,1.1257436,0.508718,1.4769232,1.6443079,1.7624617,2.409026,3.9942567,2.6453335,2.1464617,1.654154,1.1191796,1.2898463,1.6804104,1.782154,1.8281027,1.9364104,2.103795,2.0906668,2.4910772,2.556718,2.1792822,1.9035898,3.4034874,4.460308,6.166975,8.027898,7.958975,7.4896417,6.954667,5.927385,5.037949,5.9602056,7.3780518,10.262975,13.190565,15.369847,16.626873,15.442053,15.110565,15.760411,16.75159,16.699078,16.705643,15.409232,15.031796,15.399385,13.978257,14.083283,14.336001,15.031796,16.01641,16.682669,16.108309,15.481437,14.808617,14.25395,14.145642,15.061335,14.473847,13.840411,13.361232,11.98277,11.096616,11.316514,11.431385,11.149129,11.080206,11.713642,12.143591,12.228924,11.858052,10.962052,10.06277,10.571488,11.776001,12.852514,12.875488,11.611898,10.525539,9.7673855,9.508103,9.924924,11.349334,10.912822,10.075898,9.803488,10.5780525,10.939077,10.774975,10.082462,8.973129,7.6767187,7.3321033,7.781744,8.608821,9.18318,8.697436,8.989539,8.861539,8.828718,8.917334,8.677744,9.275078,9.373539,9.009232,8.320001,7.5454364,7.637334,7.9327188,9.219283,10.932513,11.158976,11.592206,11.602052,13.74195,15.346873,8.5202055,7.384616,9.462154,11.776001,13.5089245,16.009848,16.994463,16.09518,15.504412,15.750566,15.717745,16.33477,16.79754,16.626873,15.891693,15.209026,15.803078,17.11918,18.31713,18.730669,17.864206,18.01518,16.79754,15.812924,15.445334,14.838155,15.304206,15.638975,15.304206,14.9628725,16.46277,16.55795,15.993437,15.238565,14.244103,12.448821,13.735386,16.052513,17.939693,19.160616,20.722874,21.5959,19.784206,17.828104,16.44636,14.552616,11.569232,9.202872,7.318975,6.12759,6.166975,5.792821,5.044513,4.1156926,4.141949,7.210667,6.7774363,5.973334,4.785231,3.4330258,2.3696413,5.2676926,5.861744,5.901129,5.914257,5.228308,7.1122055,8.94359,7.939283,4.5390773,2.3926156,2.3302567,2.5009232,3.1442053,4.4110775,6.3442054,7.9327188,8.625232,8.776206,7.4896417,2.5993848,2.6912823,3.1113849,3.5741541,3.9056413,4.0303593,3.5413337,3.9581542,4.210872,4.204308,4.841026,3.626667,3.2196925,3.6726158,4.397949,4.1813335,3.9384618,4.2896414,4.6802053,4.827898,4.7228723,5.4613338,8.3134365,10.65354,11.277129,10.384411,7.0826674,4.7425647,4.266667,5.0871797,5.1331286,5.280821,6.0652313,6.5017443,6.803693,8.372514,4.6933336,2.6289232,2.3236926,3.0096412,2.9997952,3.9023592,3.8104618,4.2240005,4.9427695,4.076308,4.1517954,3.626667,4.381539,6.9645133,10.571488,9.619693,8.989539,7.778462,6.5345645,7.256616,7.4732313,6.564103,5.937231,5.920821,5.7665644,4.013949,3.1770258,2.7011285,2.3696413,2.297436,3.495385,5.405539,6.764308,7.128616,6.87918,4.972308,2.6912823,1.7526156,2.609231,4.453744,5.398975,5.2676926,4.7458467,4.417641,4.7491283,3.4494362,2.0151796,0.9911796,0.512,0.2855385,0.15097436,0.07876924,0.059076928,0.09189744,0.18707694,0.08533334,0.10502565,0.14441027,0.18051283,0.26256412,0.24615386,0.26584616,0.28882053,0.26912823,0.15753847,0.14112821,0.13128206,0.128,0.128,0.118153855,0.128,0.19692309,0.22646156,0.22646156,0.28225642,0.39056414,0.56123084,0.6268718,0.5907693,0.63343596,1.3981539,1.8313848,2.8849232,4.2502565,4.345436,3.8104618,3.8859491,4.2502565,4.57518,4.525949,5.3169236,7.325539,8.503796,8.372514,8.021334,8.211693,8.211693,8.136206,8.132924,8.39877,7.7259493,7.397744,7.3025646,7.381334,7.6307697,7.243488,6.7577443,6.2916927,5.976616,5.930667,6.3179493,6.944821,7.4240007,7.702975,8.060719,7.6603084,7.5388722,7.4207187,7.256616,7.213949,6.9120007,6.961231,7.240206,7.259898,6.183385,6.311385,6.170257,5.937231,5.72718,5.605744,5.7501545,6.2884107,6.5903597,6.5050263,6.38359,6.23918,6.3442054,6.173539,5.7534366,5.6385646,5.2315903,5.044513,5.330052,5.933949,6.308103,6.314667,6.445949,6.5969234,6.7905645,7.1909747,7.8112826,8.3823595,8.697436,8.920616,9.573745,10.262975,10.709334,10.617436,9.347282,5.920821,7.2631803,6.0816417,4.348718,5.3169236,13.51877,5.943795,2.3860514,2.6945643,4.3684106,2.5698464,3.4658465,3.5872824,2.5632823,1.5885129,3.4231799,3.006359,2.937436,3.318154,3.6135387,2.6551797,1.8149745,2.5173335,3.1048207,3.245949,3.9253337,3.6496413,4.1714873,4.312616,3.9745643,4.1189747,4.2338467,2.917744,1.7788719,1.6114873,2.3958976,2.0873847,2.540308,3.3575387,4.1550775,4.5554876,4.397949,4.6539493,5.139693,5.7403083,6.3934364,7.0367184,6.9743595,6.5345645,5.914257,5.1922054,4.0008206,3.501949,3.2000003,2.8717952,2.5665643,2.5600002,2.550154,2.5928206,2.7076926,2.8816411,2.8389745,2.9144619,3.255795,3.6496413,3.498667,3.442872,3.6890259,3.9417439,4.1058464,4.2863593,4.2502565,4.4274874,4.630975,4.637539,4.194462,4.453744,4.900103,5.225026,5.405539,5.681231,5.674667,5.914257,5.917539,5.579488,5.175795,5.2676926,5.362872,5.106872,4.4701543,3.7316926,4.073026,4.9296412,5.8092313,6.4000006,6.564103,6.2851286,5.858462,5.4613338,5.2578464,5.408821,5.61559,5.602462,5.861744,6.2555904,6.0258465,5.943795,5.6418467,5.297231,4.8804107,4.141949,3.6758976,3.4198978,3.1573336,2.9538465,3.1540515,2.9604106,3.2361028,3.4888208,3.3805132,2.7569232,2.5173335,2.5009232,2.4681027,2.359795,2.3072822,2.8553848,2.6551797,2.1366155,1.6311796,1.3784616,1.4211283,1.2931283,1.1257436,0.98133343,0.8533334,1.1782565,1.3784616,1.4605129,1.4506668,1.4309745,1.5163078,1.4441026,1.276718,1.0601027,0.82379496,0.8041026,0.9682052,1.1684103,1.3292309,1.4572309,1.7263591,1.8412309,1.9922053,2.2350771,2.5173335,2.2219489,1.6311796,1.1946667,1.0633847,1.079795,1.3686155,2.0086155,2.5435898,2.7634873,2.7241027,2.5993848,2.359795,2.4615386,3.0260515,3.8564105,3.9975388,4.2174363,4.345436,4.378257,4.4701543,4.3716927,4.1222568,4.1025643,4.201026,3.8104618,3.9876926,3.5840003,3.058872,2.7175386,2.7175386,3.698872,4.1124105,4.4012313,4.7655387,5.146257,4.3749747,4.338872,4.4406157,4.5489235,4.9821544,4.1058464,3.8006158,3.56759,3.495385,3.7874875,4.775385,5.72718,6.816821,7.9097443,8.726975,8.851693,8.385642,7.830975,7.653744,7.968821,8.530052,9.324308,9.842873,10.597744,11.460924,11.641437,11.897437,12.438975,13.069129,13.512206,13.426873,15.015386,15.842463,16.091898,15.95077,15.609437,15.43877,15.369847,15.868719,16.928822,18.051283,17.220924,16.456207,16.810667,18.707693,21.940514,25.504822,28.960823,32.68923,37.34318,43.838364,61.377647,74.32534,81.6476,85.64185,91.90401,79.3436,60.65888,46.070156,39.312412,37.62872,30.365541,23.194258,16.49231,11.122872,8.438154,6.5936418,4.926359,3.6562054,2.8488207,2.3958976,3.0424619,2.9768207,2.8356924,2.8291285,2.7306669,2.3171284,1.719795,1.2176411,0.97805136,1.0371283,1.0010257,0.7187693,0.3708718,0.108307704,0.06235898,0.17066668,0.20676924,0.15753847,0.098461546,0.18379489,0.318359,0.2855385,0.34133336,0.47261542,0.4135385,0.3249231,0.27897438,0.19692309,0.098461546,0.06235898,0.14769232,0.3511795,0.3511795,0.16738462,0.16738462,0.032820515,0.009846155,0.02297436,0.02297436,0.0,0.013128206,0.006564103,0.06235898,0.18379489,0.3052308,0.256,0.93866676,1.1093334,1.0338463,2.487795,3.7087183,4.2338467,3.889231,3.3247182,3.9811285,3.1409233,1.657436,0.8041026,1.0962052,2.3040001,1.5721027,1.2603078,1.7362052,2.553436,2.4582565,2.1989746,2.3663592,2.806154,3.3805132,3.9680004,5.408821,4.7524104,4.6900516,5.077334,2.930872,4.0041027,4.1911798,4.525949,5.4974365,7.0334363,8.218257,10.978462,14.316309,16.73518,16.23631,16.321642,16.387283,16.649847,16.869745,16.357744,15.504412,14.897232,14.87754,14.723283,12.635899,14.086565,15.110565,15.346873,15.120412,15.425642,16.06236,17.024002,17.618053,17.539284,16.89272,16.147694,14.769232,13.482668,12.76718,12.86236,11.851488,12.071385,11.992617,11.241027,10.604308,11.178667,12.393026,13.571283,14.10954,13.489232,12.757335,12.911591,13.558155,14.352411,14.998976,13.718975,11.592206,9.511385,8.008205,7.2631803,8.5202055,9.649232,9.833026,9.393231,9.796924,11.35918,11.510155,11.024411,10.203898,8.910769,7.860513,7.397744,7.5881033,8.01477,7.781744,7.5388722,7.056411,7.128616,7.565129,7.1876926,7.686565,8.251078,8.241231,7.680001,7.27959,6.6067696,6.8496413,8.011488,9.524513,10.269539,11.063796,10.948924,12.3536415,13.817437,10.010257,7.9950776,9.048616,10.70277,12.12718,14.129231,15.740719,15.284514,14.562463,14.276924,14.007796,14.995693,15.537232,15.488001,15.038361,14.710155,14.746258,16.30195,18.025026,18.842258,17.975796,18.146463,16.695797,15.126975,14.34913,14.677335,13.545027,13.873232,14.697027,15.668514,17.060104,16.508718,14.614976,13.308719,13.108514,13.108514,13.338258,14.04718,15.510976,17.43754,18.950565,21.418669,20.020514,17.992207,16.603899,15.153232,11.795693,9.088,7.269744,6.3868723,6.301539,6.1440005,5.280821,3.9745643,3.4756925,6.0258465,4.6834874,4.276513,4.7589746,4.972308,2.6387694,2.176,2.7733335,3.501949,4.59159,7.460103,8.585847,7.683283,7.0859494,6.9809237,5.431795,2.8192823,2.1497438,2.789744,4.3060517,6.4557953,6.7840004,6.7216415,7.1647186,7.1056414,3.6004105,2.540308,2.612513,3.370667,4.020513,3.4330258,3.6168208,4.201026,4.630975,4.325744,2.7175386,2.5074873,2.3827693,4.2272825,6.816821,5.8289237,5.7435904,4.1124105,3.062154,3.1606157,3.4166157,2.9538465,4.522667,7.8539495,10.811078,9.383386,6.8463597,5.61559,5.4449234,5.9634876,6.6822567,7.1844106,6.2752824,5.139693,5.2348723,8.283898,4.4045134,2.537026,2.231795,2.7667694,3.1573336,2.8914874,3.5741541,4.1714873,4.345436,4.457026,5.5663595,4.5062566,3.9712822,5.041231,7.200821,9.373539,9.284924,7.9425645,6.806975,7.781744,9.357129,8.267488,6.5411286,5.3398976,4.97559,3.764513,2.9407182,2.3269746,1.9561027,2.0906668,2.2613335,4.135385,6.7774363,8.41518,6.439385,3.6430771,2.3860514,2.9407182,4.585026,5.5991797,6.1374364,5.4482055,4.850872,4.417641,2.989949,2.6486156,1.5556924,0.6892308,0.36102566,0.21333335,0.1148718,0.04594872,0.0951795,0.2231795,0.25928208,0.101743594,0.17066668,0.20020515,0.15097436,0.21333335,0.22646156,0.28225642,0.29538465,0.256,0.24287182,0.20676924,0.20676924,0.17066668,0.108307704,0.108307704,0.15425642,0.19692309,0.20676924,0.2100513,0.25928208,0.5021539,0.7384616,0.79425645,0.69579494,0.67282057,1.0732309,1.1290257,2.03159,3.5774362,4.1517954,3.9680004,4.0500517,4.6244106,5.3202057,5.172513,6.3442054,8.119796,8.713847,8.093539,7.9950776,7.6767187,7.8834877,7.8408213,7.6767187,8.421744,8.228104,8.077128,7.7718983,7.2992826,6.8365135,6.616616,6.47877,6.2588725,6.1374364,6.636308,6.626462,6.8496413,7.174565,7.53559,7.9491286,7.509334,7.6307697,7.896616,7.88677,7.141744,6.6034875,6.626462,7.204103,7.90318,7.8441033,7.512616,6.5969234,5.914257,5.5565133,4.896821,5.32677,5.861744,6.193231,6.3474874,6.7150774,7.020308,7.131898,6.9677954,6.6527185,6.5312824,5.907693,5.6976414,5.802667,6.038975,6.1505647,6.1374364,6.564103,6.803693,6.8496413,7.325539,7.3616414,7.5454364,7.9458466,8.329846,8.132924,8.51036,9.567181,9.780514,8.116513,4.027077,4.6867695,3.5347695,3.117949,3.387077,1.6804104,0.71548724,1.5622566,2.8816411,3.508513,2.4713848,3.7284105,3.383795,2.5862565,2.2777438,3.2032824,3.1671798,2.9669745,3.259077,3.3641028,1.2504616,1.8379488,3.4297438,4.0041027,3.7054362,4.850872,4.1682053,4.417641,4.197744,3.5938463,4.1813335,2.2646155,2.0512822,1.654154,0.955077,1.6016412,2.359795,2.8127182,3.2656412,3.5314875,2.9440002,3.8596926,4.20759,4.6966157,5.4908724,6.2096415,6.73477,6.747898,6.229334,5.47118,5.080616,4.2994876,3.7284105,3.2722054,2.9440002,2.8849232,2.7011285,2.6912823,2.6847181,2.6847181,2.868513,3.0030773,3.2754874,3.6726158,3.9351797,3.570872,3.692308,4.1091285,4.3716927,4.348718,4.2272825,4.1911798,4.2371287,4.322462,4.279795,3.8137438,4.2896414,4.9854364,5.5958977,6.048821,6.5017443,5.8289237,5.87159,5.9634876,5.737026,5.1265645,4.713026,4.9920006,4.8147697,4.135385,4.013949,4.5489235,4.5095387,4.857436,5.6976414,6.2720003,5.5630774,5.687795,5.7731285,5.6287184,5.737026,5.8486156,5.8092313,5.835488,5.989744,6.2096415,5.989744,5.8814363,5.6320004,5.1298466,4.4110775,3.895795,3.3936412,3.1540515,3.1934361,3.2656412,2.8750772,2.9801028,3.1081028,2.9997952,2.609231,2.4024618,2.3401027,2.4615386,2.6978464,2.868513,3.259077,2.806154,2.1924105,1.6968206,1.2209232,1.2340513,1.3095386,1.204513,0.9878975,1.0371283,1.3292309,1.467077,1.401436,1.2242053,1.1749744,1.3095386,1.3062565,1.1782565,0.94523084,0.64000005,0.6892308,1.0305642,1.2931283,1.3718976,1.4342566,1.6902566,1.5721027,1.7558975,2.2613335,2.4582565,2.1989746,1.6311796,1.2603078,1.276718,1.5556924,1.8248206,2.4681027,2.937436,2.9210258,2.3335385,2.1398976,2.1267693,2.3893335,2.930872,3.6627696,4.027077,4.522667,4.84759,4.886975,4.716308,4.2272825,3.6660516,3.43959,3.5183592,3.4330258,3.7251284,3.2787695,3.2164104,3.5216413,3.0227695,3.2886157,3.8334363,4.2371287,4.5095387,5.097026,5.2414365,4.969026,4.97559,5.3366156,5.5072823,4.020513,3.820308,3.5938463,3.620103,4.0336413,4.8377438,5.868308,6.770872,7.8670774,8.848411,8.763078,8.172308,7.6603084,7.9130263,8.63836,8.553026,9.074872,9.662359,10.282667,10.857026,11.264001,10.758565,11.188514,11.98277,12.757335,13.305437,14.697027,15.064616,15.392821,15.924514,16.15754,15.675078,15.074463,15.37313,16.44636,17.014154,16.827078,16.502155,17.798565,20.98872,24.85826,29.059284,32.840206,37.248,43.776005,54.37375,70.04883,79.8556,86.39672,91.4478,95.93108,79.49457,62.020927,49.729645,43.234467,37.556515,28.816412,21.474463,15.461744,11.158976,9.403078,8.917334,7.4043083,5.612308,4.020513,2.8356924,2.7011285,2.789744,2.9243078,2.9571285,2.7798977,2.1398976,1.5819489,1.1388719,0.93866676,1.1946667,1.3259488,1.017436,0.60061544,0.2855385,0.15753847,0.17066668,0.190359,0.16738462,0.13456412,0.21989745,0.39384618,0.36430773,0.380718,0.45620516,0.37415388,0.2297436,0.12471796,0.059076928,0.072205134,0.21989745,0.81394875,0.93866676,1.0699488,1.2537436,1.1093334,0.32820517,0.06235898,0.016410258,0.016410258,0.013128206,0.06235898,0.36102566,0.892718,1.2570257,0.6465641,1.2832822,2.6715899,3.3345644,3.186872,3.5380516,3.3411283,3.3214362,3.370667,3.4756925,3.7251284,3.4494362,2.8258464,2.5764105,2.7142565,2.537026,2.231795,2.038154,2.156308,2.3663592,2.0053334,1.913436,2.412308,2.861949,3.0096412,2.989949,3.436308,4.1550775,4.338872,4.007385,4.017231,4.3585644,5.1889234,6.311385,7.4240007,8.132924,9.032206,10.453334,11.871181,13.065847,14.148924,15.218873,16.331488,17.427694,17.8839,16.49231,15.432206,14.011078,13.4629755,13.53518,12.511181,12.763899,13.236514,13.679591,14.01436,14.329437,15.254975,16.02954,15.698052,14.762668,15.169642,15.402668,14.247386,12.983796,12.448821,13.033027,12.947693,12.041847,11.264001,10.935796,10.752001,11.667693,13.105232,14.785643,15.694771,14.073437,12.416001,12.580104,13.699283,14.723283,14.41477,13.10195,11.329642,9.199591,7.325539,6.8233852,7.8769236,8.815591,9.481847,9.905231,10.308924,11.687386,12.435693,11.943385,10.630565,9.961026,9.03877,7.975385,7.2336416,6.921847,6.806975,7.000616,6.4689236,6.564103,7.3058467,7.3583593,7.253334,7.4240007,7.427283,7.1187696,6.669129,6.678975,6.698667,7.240206,8.4283085,10.013539,10.463181,10.955488,11.533129,12.678565,15.29436,9.4916935,9.268514,10.545232,11.395283,12.028719,14.03077,14.631386,14.437745,13.974976,13.666463,14.411489,14.844719,15.120412,15.199181,14.880821,14.145642,15.297642,17.168411,18.596104,18.41559,18.438566,16.62359,14.775796,13.863386,14.007796,13.302155,13.344822,13.801026,14.027489,13.056001,13.640206,13.131488,12.544001,12.435693,12.924719,12.901745,12.777026,13.29559,14.437745,15.42236,18.44513,18.198977,16.741745,15.182771,13.66318,11.08677,8.779488,7.171283,6.5411286,7.02359,6.550975,5.477744,4.7228723,5.156103,7.5881033,4.95918,3.5807183,5.4153852,8.349539,6.2030773,3.3772311,2.044718,1.9364104,3.5610259,8.205129,9.524513,9.074872,7.145026,5.7632823,8.704,5.691077,3.95159,2.993231,2.7306669,3.511795,5.297231,7.2369237,7.6734366,6.4557953,4.9427695,3.1409233,2.6026669,3.5216413,4.972308,4.923077,5.221744,5.802667,5.6976414,4.6572313,3.1442053,3.0523078,2.9046156,2.8980515,3.0884104,3.387077,4.2896414,4.322462,4.1025643,4.027077,4.2830772,3.058872,2.9210258,4.716308,6.957949,5.832206,4.5522056,3.826872,3.4166157,3.7218463,5.7796926,5.1659493,5.2676926,5.3398976,5.723898,7.857231,4.9132314,2.9965131,2.6518977,3.3312824,3.3903592,3.0227695,3.1474874,3.0096412,2.9505644,4.417641,4.201026,3.8859491,4.5029745,6.058667,7.5552826,8.664616,7.8112826,6.518154,5.868308,6.51159,7.197539,6.8693337,6.0980515,5.169231,4.069744,3.7120004,3.0490258,2.3630772,2.1792822,3.2623591,3.4822567,5.0904617,7.640616,9.340718,7.062975,3.6693337,3.2886157,4.44718,5.8814363,6.550975,6.99077,6.6428723,5.9536414,5.1364107,4.1878977,3.1606157,1.6705642,0.6629744,0.3446154,0.17723078,0.098461546,0.03938462,0.08533334,0.18379489,0.16082053,0.08205129,0.098461546,0.118153855,0.13128206,0.20020515,0.19364104,0.23302566,0.256,0.23302566,0.17066668,0.27241027,0.26912823,0.19364104,0.11158975,0.13128206,0.17066668,0.17723078,0.21333335,0.28225642,0.32164106,0.41682056,0.571077,0.73517954,0.84348726,0.83035904,0.86317956,1.1027694,1.8445129,2.8258464,3.2229745,3.7120004,4.073026,4.637539,5.179077,4.903385,7.0432825,8.306872,8.362667,7.6734366,7.506052,7.463385,7.397744,7.1647186,6.9677954,7.3616414,7.030154,6.8233852,6.567385,6.2523084,6.042257,6.0947695,5.9470773,5.654975,5.3694363,5.330052,6.491898,7.3747697,7.830975,7.9294367,7.975385,8.050873,8.28718,8.198565,7.716103,7.177847,6.875898,6.5903597,6.688821,7.0793853,7.1844106,6.9021544,6.738052,6.2851286,5.602462,5.21518,5.349744,5.5729237,5.730462,5.8945646,6.3474874,6.564103,6.816821,6.9054365,6.669129,5.979898,5.914257,6.196513,6.5772314,6.872616,6.941539,7.1154876,7.2237954,7.27959,7.381334,7.702975,7.955693,7.824411,8.188719,9.104411,9.816616,9.609847,9.209436,8.103385,6.23918,4.017231,3.511795,2.7273848,2.5238976,2.6223593,1.6049232,1.4112822,1.9396925,2.2088206,2.0709746,2.2153847,2.878359,2.989949,2.6715899,2.1858463,1.972513,2.4910772,2.5895386,2.3794873,2.1234872,2.228513,2.9013336,3.5052311,3.6693337,3.511795,3.6430771,2.5206156,3.9581542,4.417641,3.3280003,3.0949745,1.7066668,1.2865642,1.4506668,1.8707694,2.2744617,2.6880002,2.6551797,2.7634873,2.9538465,2.4943593,3.4691284,3.9680004,4.57518,5.3891287,6.052103,6.449231,6.4754877,6.121026,5.474462,4.70318,3.8728209,3.4002054,3.1081028,2.9243078,2.8717952,2.9702566,2.8488207,2.7963078,2.8980515,3.0523078,3.2262566,3.570872,3.82359,3.9187696,4.010667,4.023795,4.1780515,4.397949,4.5817437,4.6178465,4.640821,4.634257,4.466872,4.1550775,3.889231,3.9647183,4.2962055,5.041231,5.986462,6.5378466,5.933949,5.796103,5.661539,5.3792825,5.0904617,5.3694363,5.5958977,5.297231,4.70318,4.7589746,5.7140517,5.3858466,4.896821,5.0543594,6.3310776,5.664821,5.2709746,5.2644105,5.467898,5.4186673,5.4514875,5.901129,6.121026,6.0258465,6.088206,5.664821,5.618872,5.4580517,5.0116925,4.44718,4.2174363,4.135385,3.9647183,3.7316926,3.7185643,3.0129232,2.9078977,2.9243078,2.8160002,2.5731285,2.5009232,2.422154,2.605949,3.0194874,3.3575387,3.2295387,2.678154,2.0808206,1.595077,1.1585642,1.2012309,1.2570257,1.273436,1.273436,1.3292309,1.3686155,1.3784616,1.3292309,1.273436,1.3226668,1.467077,1.4506668,1.3226668,1.1257436,0.90912825,0.9189744,1.148718,1.2931283,1.2012309,0.8730257,1.401436,1.4900514,1.723077,2.1891284,2.4943593,1.8281027,1.332513,1.1716924,1.3292309,1.6311796,2.1431797,2.6715899,2.9111798,2.7963078,2.4943593,2.3762052,2.609231,2.9702566,3.3214362,3.626667,3.9122055,4.3585644,4.8771286,5.330052,5.5204105,4.5423594,4.0500517,3.95159,3.9975388,3.7743592,3.754667,3.6529233,3.4888208,3.3444104,3.3641028,3.7973337,4.397949,4.6966157,4.7589746,5.169231,5.5302567,6.0061545,6.701949,7.318975,7.1548724,3.255795,3.370667,3.6562054,3.882667,4.066462,4.450462,5.405539,6.380308,7.4797955,8.3823595,8.3593855,8.425026,8.274052,8.490667,8.887795,8.4972315,8.411898,8.874667,9.380103,9.833026,10.548513,10.203898,11.093334,12.018872,12.665437,13.61395,14.818462,15.002257,14.953027,14.995693,15.015386,15.442053,15.481437,15.796514,16.357744,16.423386,17.089642,17.923283,19.800617,23.056412,27.503592,31.133541,35.01949,40.320004,47.973747,58.70934,72.65149,84.4997,93.78462,97.79529,91.58237,70.12103,53.86503,42.93908,35.78749,29.161028,22.347488,16.04595,11.152411,8.152616,7.125334,6.8332314,5.789539,4.348718,2.9013336,1.8543591,1.5031796,1.5097437,1.9200002,2.5107694,2.793026,2.359795,1.9035898,1.529436,1.270154,1.1093334,1.1323078,0.95835906,0.6662565,0.37415388,0.2297436,0.18707694,0.24615386,0.23302566,0.16082053,0.20020515,0.28882053,0.26584616,0.27241027,0.3314872,0.34789747,0.190359,0.072205134,0.032820515,0.13456412,0.4594872,0.6826667,0.6104616,0.702359,0.9353847,0.8041026,0.45620516,0.2297436,0.108307704,0.07548718,0.08861539,0.16410258,0.86974365,1.2898463,1.142154,0.7975385,1.654154,2.8192823,3.190154,2.7241027,2.4549747,2.2547693,2.3926156,2.8849232,3.5216413,3.8367183,3.6496413,4.2174363,4.276513,3.6857438,3.4100516,3.1540515,2.7634873,2.5961027,2.5009232,1.8084104,2.038154,2.2482052,2.300718,2.169436,1.9396925,2.986667,3.7809234,4.201026,4.2830772,4.2338467,4.7589746,5.681231,7.0892315,8.67118,9.734565,11.047385,10.624001,10.331899,10.824206,11.539693,12.724514,14.191591,16.075489,17.375181,15.940925,15.291079,13.725539,12.35036,11.59877,11.244308,10.932513,11.670976,12.652308,13.302155,13.275898,15.097437,16.23631,15.812924,14.50995,14.565744,15.363283,14.998976,13.88636,12.872206,13.249642,13.830565,12.819694,12.114052,12.084514,11.565949,12.458668,13.869949,14.943181,15.051488,13.801026,13.138052,13.564719,14.358975,14.890668,14.605129,13.22995,11.546257,9.462154,7.6110773,7.3550773,8.214975,9.304616,10.098872,10.354873,10.098872,10.893129,12.1928215,12.143591,10.834052,10.305642,9.334154,8.602257,7.643898,6.698667,6.7085133,7.2237954,6.9809237,6.8988724,7.253334,7.64718,7.0465646,6.9087186,6.8397956,6.6560006,6.370462,6.38359,6.6067696,7.0892315,7.8408213,8.812308,9.281642,10.7848215,12.07795,13.4170265,16.544823,11.1983595,10.020103,10.512411,11.145847,11.35918,12.396309,13.718975,14.191591,13.768207,13.479385,13.656616,13.978257,14.5952835,15.136822,14.70359,13.51877,14.247386,16.196924,18.274464,18.97354,17.224207,15.537232,14.221129,13.413745,13.078976,12.803283,13.167591,14.050463,14.39836,12.219078,12.501334,13.013334,12.87877,12.491488,13.51877,13.814155,13.088821,12.507898,12.84595,14.467283,16.817232,16.603899,15.225437,13.538463,11.85477,9.993847,8.582564,7.2927184,6.498462,7.276308,7.003898,5.7009234,5.2578464,6.6822567,10.112,7.890052,4.604718,4.7327185,7.6898465,7.8473854,6.99077,4.46359,2.92759,3.2656412,4.594872,8.65477,8.503796,6.8627696,5.7632823,6.547693,7.387898,5.1364107,3.3312824,3.0818465,3.0523078,4.525949,6.810257,8.093539,7.6176414,5.681231,3.9647183,3.0785644,3.748103,5.218462,5.2676926,5.3858466,5.989744,6.121026,5.32677,3.6627696,3.6069746,3.820308,3.3017437,2.2383592,1.9889232,2.4648206,3.1245131,3.6758976,3.9220517,3.761231,2.7175386,2.2678976,3.1376412,5.0609236,6.7938466,9.212719,8.169026,5.4482055,3.9253337,7.578257,5.5302567,5.2414365,5.7534366,6.7840004,8.740103,4.923077,3.2229745,2.993231,3.387077,3.3476925,2.553436,2.7470772,2.7142565,2.5074873,3.4133337,3.5282054,4.1550775,4.9132314,6.488616,10.637129,10.44677,8.113232,5.720616,4.5423594,5.024821,5.648411,6.301539,7.131898,7.6603084,6.774154,5.2447186,3.7218463,3.498667,4.965744,7.6012316,7.650462,7.834257,8.188719,7.9228725,5.405539,2.8980515,3.2229745,4.5554876,5.540103,5.297231,5.83877,5.330052,4.6769233,4.2272825,3.8071797,3.2656412,1.7985642,0.7122052,0.35774362,0.15753847,0.08533334,0.036102567,0.06564103,0.16082053,0.24615386,0.14112821,0.101743594,0.0951795,0.118153855,0.19692309,0.20020515,0.18379489,0.18051283,0.18707694,0.13456412,0.21661541,0.2231795,0.18051283,0.14112821,0.16410258,0.16410258,0.16738462,0.19364104,0.23630771,0.24287182,0.3052308,0.5152821,0.77128214,0.9878975,1.1093334,0.892718,1.1520001,1.7033848,2.3630772,2.9440002,3.948308,4.397949,4.71959,5.028103,5.139693,8.523488,8.595693,7.6898465,7.020308,6.688821,7.315693,7.2237954,6.8496413,6.6395903,7.0400004,5.933949,5.7107697,5.684513,5.6385646,5.835488,6.0685134,6.052103,5.87159,5.5893335,5.2414365,6.445949,7.785026,8.474257,8.536616,8.805744,9.196308,8.960001,8.241231,7.39118,6.9776416,6.491898,5.98318,6.121026,6.8365135,7.3485136,7.5421543,7.529026,7.328821,6.925129,6.265436,6.0258465,5.648411,5.4974365,5.8289237,6.7872825,6.8955903,6.9710774,6.931693,6.619898,5.835488,5.7764106,5.976616,6.340924,6.8627696,7.634052,7.817847,7.8769236,7.975385,8.165744,8.36595,8.011488,7.6931286,8.274052,9.622975,10.614155,10.164514,9.248821,8.096821,6.921847,5.927385,4.9788723,3.9680004,3.6529233,3.9548721,3.9384618,3.3017437,2.5698464,2.1267693,2.2121027,2.930872,3.0162053,2.9440002,2.737231,2.4385643,2.0939488,2.4582565,2.1825643,1.8051283,1.9495386,3.3050258,3.0326157,3.1343591,3.1638978,2.917744,2.409026,1.9659488,3.2328207,3.495385,2.6322052,3.114667,3.0884104,2.2219489,1.7427694,1.910154,2.038154,2.1202054,2.9111798,3.2229745,2.740513,2.0512822,3.05559,3.3772311,4.0303593,5.0871797,5.691077,5.72718,5.9602056,5.868308,5.280821,4.3716927,3.570872,3.1934361,2.9735386,2.8488207,2.9702566,2.9702566,2.8225644,2.8192823,3.0818465,3.5741541,3.639795,3.882667,3.9942567,3.9811285,4.164923,4.2994876,4.4800005,4.775385,5.034667,4.8804107,4.70318,4.644103,4.568616,4.388103,4.0434875,3.9023592,4.1189747,4.9394875,6.0619493,6.629744,5.8814363,5.428513,5.0084105,4.6145644,4.4865646,5.346462,5.668103,5.0674877,4.1714873,4.6145644,5.874872,5.83877,4.95918,4.2896414,5.4875903,5.6254363,4.9296412,4.775385,5.2020516,4.9099493,5.0904617,6.4295387,6.8627696,6.114462,5.7009234,6.009436,5.8486156,5.395693,4.896821,4.667077,4.516103,4.338872,4.1550775,4.017231,4.0041027,3.6168208,3.6463592,3.4166157,2.8488207,2.4451284,2.6354873,2.6354873,2.861949,3.2754874,3.4067695,2.9440002,2.487795,1.9167181,1.3620514,1.1913847,1.1716924,1.2209232,1.2832822,1.3357949,1.4145643,1.3587693,1.3062565,1.2176411,1.1684103,1.3292309,1.6147693,1.5392822,1.4900514,1.4441026,0.9485129,1.014154,1.1946667,1.5163078,1.6902566,1.1093334,1.5819489,1.8281027,2.0676925,2.2711797,2.1464617,1.4998976,1.3686155,1.4244103,1.5622566,1.9035898,2.4713848,2.8882053,2.9735386,2.7995899,2.6715899,2.4188719,2.6978464,3.0982566,3.3903592,3.5347695,3.6562054,4.128821,4.7491283,5.421949,6.170257,5.1364107,4.4045134,4.0008206,3.8564105,3.8071797,3.5314875,3.3903592,3.2722054,3.2196925,3.43959,4.2371287,4.4307694,4.850872,5.5007186,5.58277,6.2884107,6.987488,7.128616,6.7807183,6.626462,3.370667,3.6660516,4.023795,4.197744,4.1911798,4.2469745,5.100308,6.0192823,6.944821,7.7423596,8.205129,9.147078,8.933744,8.615385,8.546462,8.379078,8.077128,8.4972315,8.940309,9.31118,10.112,10.102155,10.971898,11.634872,12.005745,13.033027,14.237539,14.644514,14.460719,14.050463,13.922462,14.900514,15.471591,15.730873,15.894976,16.265848,17.24718,18.944002,21.234873,24.362669,28.931284,32.469337,36.420925,42.243286,50.832413,62.529644,76.23221,89.104416,95.83263,92.28472,75.520004,54.57395,41.088,31.855593,24.82872,19.10154,14.381949,10.20718,7.259898,5.602462,4.673641,4.1452312,3.6791797,2.793026,1.6607181,1.1290257,0.77128214,0.6859488,1.0962052,1.8609232,2.487795,2.3663592,2.0118976,1.6246156,1.276718,0.9124103,0.81394875,0.8566154,0.69579494,0.35774362,0.23630771,0.20348719,0.26584616,0.2986667,0.27569234,0.26912823,0.20020515,0.17066668,0.18707694,0.22646156,0.23958977,0.118153855,0.03938462,0.029538464,0.13128206,0.4004103,0.40697438,0.32820517,0.36758977,0.48902568,0.43651286,0.65641034,0.5152821,0.30851284,0.19692309,0.2100513,0.26256412,0.84348726,1.0272821,0.7253334,0.7187693,1.7394873,2.0873847,1.9200002,1.6016412,1.6902566,1.9528207,2.3401027,3.0490258,3.9154875,4.4406157,4.5587697,5.10359,4.8804107,4.07959,4.3060517,3.6135387,2.9636924,3.006359,3.2754874,2.1989746,2.1070771,2.176,2.0742567,2.0217438,2.7831798,3.7743592,4.535795,5.225026,5.6451287,5.2578464,5.605744,6.2818465,7.387898,8.805744,10.194052,11.175385,10.220308,9.80677,10.630565,11.631591,11.936821,13.124924,14.992412,16.357744,15.061335,13.5318985,12.265027,11.283693,10.548513,9.977437,9.577026,10.236719,11.178667,11.881026,12.084514,14.165335,15.698052,16.118155,15.609437,15.140103,15.494565,15.186052,14.339283,13.4859495,13.590976,14.080001,13.46954,13.144616,13.164309,12.268309,12.422565,13.5089245,13.879796,13.282462,12.829539,13.13477,14.168616,14.907078,15.0777445,15.14995,14.162052,12.35036,10.148104,8.388924,8.283898,8.421744,9.366975,10.374565,10.834052,10.305642,10.466462,11.369026,11.588924,10.916103,10.361437,9.511385,9.137232,8.283898,7.0925136,6.7807183,7.39118,7.2237954,6.9842057,7.072821,7.574975,6.928411,6.7807183,6.76759,6.685539,6.4590774,6.5870776,6.8562055,7.1614366,7.4797955,7.8736415,8.375795,10.397539,12.442257,14.034052,15.744001,12.12718,10.637129,10.486155,10.929232,11.254155,11.687386,13.210258,14.053744,13.899488,13.869949,13.814155,13.584412,13.919181,14.644514,14.677335,14.188309,14.726565,16.183796,17.979078,19.052309,16.498873,14.624822,13.50236,13.010053,12.822975,13.049437,13.935591,15.126975,15.501129,13.147899,13.348104,13.794462,13.37436,12.626052,13.722258,14.480412,13.558155,12.773745,13.105232,14.700309,15.179488,14.65436,13.636924,12.3536415,10.761847,9.363693,8.51036,7.6143594,6.8365135,7.1056414,6.941539,5.85518,5.5138464,6.6625648,9.124104,8.4512825,5.0018463,3.511795,5.1364107,7.4797955,8.523488,6.491898,5.3366156,5.464616,3.7382567,6.058667,7.0400004,6.616616,5.4383593,4.84759,7.069539,6.0160003,5.041231,4.850872,3.5282054,4.2929235,6.2555904,8.018052,8.536616,7.1220517,5.540103,4.3552823,4.2962055,4.886975,4.460308,4.525949,5.7074876,6.38359,5.9602056,4.8771286,4.164923,4.276513,3.7973337,2.5731285,1.7033848,1.6968206,1.9659488,2.3696413,2.6420515,2.3991797,1.975795,1.8346668,2.878359,5.037949,7.2861543,11.063796,10.70277,7.6570263,4.857436,6.705231,5.9602056,5.5729237,5.3924108,5.9930263,8.690872,5.2644105,3.5183592,3.0982566,3.43959,3.751385,3.0949745,3.4888208,3.4724104,2.9538465,3.2032824,4.092718,5.221744,6.183385,7.578257,11.027693,10.696206,8.63836,6.052103,4.309334,4.962462,6.944821,8.03118,8.539898,8.487385,7.581539,6.23918,5.6418467,6.36718,8.27077,10.482873,10.164514,9.452309,8.28718,6.5837955,4.20759,2.8914874,3.5249233,4.325744,4.525949,4.381539,4.2272825,3.623385,3.190154,3.2262566,3.6758976,2.9702566,1.6771283,0.69907695,0.3117949,0.14112821,0.06564103,0.029538464,0.036102567,0.1148718,0.28882053,0.17066668,0.10502565,0.08205129,0.108307704,0.19692309,0.190359,0.15097436,0.13784617,0.14769232,0.13456412,0.17394873,0.17066668,0.17066668,0.17723078,0.18379489,0.18707694,0.190359,0.29538465,0.4004103,0.21333335,0.26912823,0.47589746,0.7187693,0.9682052,1.273436,1.0962052,1.273436,1.6836925,2.2580514,2.9997952,4.2962055,4.9985647,5.297231,5.4383593,5.737026,8.448001,7.6734366,6.73477,6.616616,5.9930263,6.7249236,6.6133337,6.3277955,6.301539,6.747898,6.0324106,5.8453336,5.8157954,5.868308,6.2129235,6.2785645,6.2851286,6.340924,6.4754877,6.62318,7.512616,8.283898,8.641642,8.677744,8.858257,9.304616,8.822155,7.8637953,6.997334,6.9087186,6.2490263,5.7501545,6.012718,6.889026,7.463385,8.39877,8.628513,8.375795,7.7948723,6.997334,6.3967185,5.8453336,5.664821,5.9963083,6.8004107,7.171283,7.1056414,6.931693,6.636308,5.865026,5.405539,5.5729237,6.124308,6.944821,8.044309,8.060719,8.149334,8.333129,8.5202055,8.51036,8.034462,7.6996927,8.139488,9.189744,9.856001,9.895386,9.544206,8.953437,8.3134365,7.8736415,6.370462,6.042257,5.76,5.3169236,5.4482055,3.9253337,2.9407182,2.5796926,2.7142565,2.9801028,2.7602053,2.477949,2.2219489,2.0578463,2.038154,1.9200002,1.5458462,1.4211283,2.1333334,4.312616,3.5610259,3.7218463,3.5741541,2.8914874,2.425436,2.6683078,3.1245131,2.7864618,2.2088206,3.495385,4.0533338,3.2918978,2.3794873,1.9331284,2.0151796,1.7788719,2.6387694,3.5577438,3.5840003,1.847795,3.1540515,3.255795,3.5183592,4.2994876,4.923077,4.7392826,5.1298466,5.0477953,4.312616,3.626667,3.2065644,3.0752823,3.0326157,3.0129232,3.1048207,2.9833848,2.8356924,2.92759,3.3247182,3.879385,4.017231,4.1714873,4.135385,3.9975388,4.1091285,4.2240005,4.5522056,4.896821,5.106872,5.044513,4.7228723,4.6145644,4.6276927,4.601436,4.3060517,4.1583595,4.3618464,4.969026,5.6976414,5.933949,5.5236926,5.1987696,4.8377438,4.4767184,4.322462,5.3825645,5.802667,5.1659493,4.1747694,4.644103,5.943795,6.0717955,5.225026,4.2174363,4.4800005,5.362872,5.0674877,4.8049235,4.896821,4.788513,5.0576415,6.51159,7.0367184,6.311385,5.805949,6.432821,6.23918,5.8092313,5.4383593,5.152821,4.706462,4.4438977,4.3716927,4.3585644,4.138667,3.9286156,4.132103,3.751385,2.802872,2.3105643,2.609231,2.7700515,2.9997952,3.2295387,3.1015387,2.8192823,2.412308,1.7952822,1.204513,1.1651284,1.1585642,1.3226668,1.4933335,1.5524104,1.4441026,1.404718,1.3915899,1.3653334,1.3292309,1.3259488,1.6016412,1.4966155,1.5885129,1.7591796,1.1815386,1.0666667,1.3259488,1.7263591,1.9265642,1.4736412,1.8543591,2.0906668,2.2580514,2.2514873,1.7788719,1.4211283,1.4933335,1.5819489,1.6836925,2.2153847,2.7437952,3.045744,3.0654361,2.8947694,2.809436,2.5600002,2.789744,3.1934361,3.4822567,3.4067695,3.5314875,4.135385,4.8147697,5.3891287,5.920821,5.152821,4.4110775,3.9417439,3.7842054,3.757949,3.2131286,3.0424619,3.0851285,3.2787695,3.6332312,4.969026,5.211898,5.7435904,6.7085133,7.003898,7.2237954,7.2960005,7.056411,6.626462,6.4065647,4.1846156,4.384821,4.3749747,4.345436,4.348718,4.312616,5.10359,5.8453336,6.5772314,7.3550773,8.264206,9.645949,9.088,8.188719,7.827693,8.15918,8.149334,8.592411,8.996103,9.317744,9.954462,10.161232,10.476309,10.640411,10.843898,11.707078,12.944411,13.653335,13.722258,13.50236,13.794462,14.316309,14.634667,14.788924,15.110565,16.20349,17.09949,19.058874,21.392412,24.264208,28.694977,32.95508,37.38585,43.392002,52.430775,66.04472,80.36431,89.92493,87.72267,73.22913,52.397953,37.851902,28.015593,20.667078,14.815181,10.686359,7.50277,5.796103,4.965744,4.381539,3.3575387,2.7963078,2.7273848,2.172718,1.2438976,1.142154,0.79425645,0.761436,0.9747693,1.3784616,1.9298463,1.9593848,1.6672822,1.2438976,0.8566154,0.6859488,0.571077,0.76800007,0.65969235,0.26256412,0.2100513,0.21989745,0.2231795,0.2855385,0.3708718,0.34133336,0.17066668,0.13128206,0.15097436,0.16082053,0.07548718,0.026256412,0.0032820515,0.01969231,0.068923086,0.15097436,0.2855385,0.5218462,0.64000005,0.5940513,0.512,0.8369231,0.6859488,0.42338464,0.26912823,0.2986667,0.30194873,0.36102566,0.4594872,0.62030774,0.9321026,1.7263591,1.276718,0.9124103,1.2668719,2.2908719,2.8225644,3.1048207,3.5347695,4.1222568,4.4964104,4.886975,4.650667,4.128821,3.8006158,4.276513,3.1015387,2.5337439,3.0720003,3.8662567,2.7208207,1.9331284,2.5140514,2.789744,2.9702566,5.146257,5.218462,6.045539,6.820103,7.1023593,6.806975,6.491898,6.6395903,7.1089234,7.8637953,8.979693,9.199591,9.081436,9.665642,11.168821,12.973949,12.593232,13.466257,14.693745,15.225437,13.843694,11.221334,10.535385,10.66995,10.620719,9.494975,9.222565,9.275078,9.662359,10.331899,11.162257,12.796719,14.460719,15.852309,16.515284,15.832617,15.343591,14.457437,14.112822,14.381949,14.473847,14.152206,13.561437,13.272616,13.108514,12.150155,11.588924,12.242052,12.301129,11.641437,11.831796,12.360206,13.88636,14.920206,15.120412,15.330462,14.923489,13.2562065,11.096616,9.3768215,9.173334,8.237949,8.507077,9.813334,11.257437,11.224616,10.909539,10.811078,10.896411,10.896411,10.295795,9.80677,9.442462,8.743385,7.706257,6.764308,7.145026,6.918565,6.6822567,6.744616,7.1515903,6.951385,6.8529234,6.9152827,7.020308,6.8660517,7.207385,7.2927184,7.2927184,7.387898,7.77518,8.155898,9.993847,12.104206,13.7386675,14.605129,12.3076935,10.9456415,10.456616,10.70277,11.480617,12.120616,13.308719,14.204719,14.611693,14.979283,14.844719,13.912617,13.538463,14.083283,14.930053,15.570052,16.275694,17.10277,17.956104,18.592821,16.633438,14.427898,13.213539,13.259488,13.883078,13.994668,15.117129,16.265848,16.354464,14.201437,14.992412,14.752822,13.751796,12.790154,13.200411,14.145642,13.459693,13.3940525,14.404924,15.179488,13.233232,12.481642,12.038565,11.355898,10.230155,9.238976,8.500513,8.0377445,7.653744,6.9349747,6.5837955,5.8814363,5.4908724,5.543385,5.6320004,6.0291286,4.082872,2.3762052,2.5600002,5.35959,6.948103,6.432821,6.882462,8.041026,6.3212314,3.1409233,4.8640003,5.533539,4.210872,4.972308,5.4580517,7.0367184,7.936001,7.076103,4.066462,4.5029745,5.7435904,7.131898,8.2215395,8.753231,7.3321033,5.9995904,5.110154,4.46359,3.3247182,3.4494362,5.113436,6.1407185,6.114462,6.3967185,4.8147697,4.3618464,3.8564105,2.9111798,1.9232821,1.7591796,1.3489232,1.1093334,1.1355898,1.2274873,1.6410258,1.7788719,3.2656412,5.6254363,6.2720003,8.293744,9.133949,8.011488,5.4908724,3.4724104,5.2512827,5.504,4.453744,3.8662567,7.059693,6.193231,4.420923,3.3312824,3.3936412,3.945026,3.8531284,4.345436,4.2830772,3.748103,4.0303593,5.1987696,6.554257,8.136206,9.403078,9.248821,9.176616,8.362667,6.5936418,5.044513,6.2851286,9.993847,11.388719,10.47959,8.247795,6.6494365,6.6133337,7.830975,9.176616,10.085744,10.568206,9.77395,9.032206,7.8145647,6.0750775,4.2207184,3.8662567,4.4438977,4.332308,3.6529233,4.2601027,3.170462,2.5862565,2.353231,2.5928206,3.692308,2.5796926,1.4145643,0.58092314,0.19692309,0.11158975,0.049230773,0.026256412,0.01969231,0.059076928,0.21989745,0.14769232,0.08533334,0.068923086,0.118153855,0.21661541,0.18379489,0.16410258,0.14441027,0.13128206,0.15097436,0.17066668,0.16410258,0.190359,0.23958977,0.21989745,0.24287182,0.23958977,0.4266667,0.62030774,0.25928208,0.2986667,0.42338464,0.57764107,0.79425645,1.2176411,1.2898463,1.4178462,1.7460514,2.3138463,3.0720003,4.460308,5.467898,5.98318,6.114462,6.2129235,7.0367184,6.1472826,5.8518977,6.294975,5.467898,5.874872,5.8289237,5.8125134,6.0324106,6.4032826,7.02359,6.994052,6.882462,6.944821,7.125334,6.931693,6.8365135,7.076103,7.702975,8.576,8.930462,8.516924,8.237949,8.241231,7.939283,8.136206,7.77518,7.062975,6.5247183,7.000616,6.377026,6.0980515,6.442667,7.1515903,7.4240007,8.809027,9.337437,8.907488,7.939283,7.3550773,6.5772314,6.265436,6.2916927,6.449231,6.4689236,7.171283,7.1909747,7.066257,6.820103,5.986462,5.2020516,5.3858466,6.1341543,7.0892315,7.939283,7.939283,8.116513,8.333129,8.441437,8.283898,8.113232,7.7981544,7.680001,7.8408213,8.103385,8.828718,9.540924,9.665642,9.298052,9.219283,7.8703594,8.684308,8.057437,5.7796926,5.041231,3.511795,3.3050258,3.4133337,3.2656412,2.7437952,2.1858463,1.9692309,1.6410258,1.3029745,1.6147693,1.1257436,1.017436,1.4736412,2.7076926,4.9526157,4.903385,5.47118,4.896821,3.501949,3.692308,3.9286156,3.6594875,2.809436,2.15959,3.3575387,3.6660516,3.3542566,2.6453335,2.0250258,2.2350771,1.9593848,1.9364104,3.1934361,4.4274874,2.0020514,3.501949,3.4921029,3.1967182,3.308308,3.9614363,3.7776413,4.0336413,3.7218463,2.9111798,2.7700515,2.9505644,3.058872,3.18359,3.2722054,3.1113849,3.0424619,2.9801028,3.2065644,3.6562054,3.9286156,4.269949,4.352,4.1911798,3.9417439,3.895795,3.8564105,4.2994876,4.6112823,4.6834874,4.9329233,4.7458467,4.670359,4.6802053,4.70318,4.6178465,4.519385,4.644103,4.890257,5.0609236,4.890257,5.1200004,5.156103,5.0838976,4.9362054,4.6802053,5.586052,5.9995904,5.648411,5.0051284,5.293949,6.2752824,6.180103,5.681231,5.0674877,4.2469745,5.093744,5.651693,5.3891287,4.6900516,4.850872,5.2348723,6.0356927,6.482052,6.370462,6.0750775,6.550975,6.5280004,6.38359,6.189949,5.691077,4.8016415,4.598154,4.6933336,4.6966157,4.2207184,3.8859491,4.010667,3.5872824,2.6551797,2.2744617,2.412308,2.7602053,3.0162053,3.0227695,2.7602053,2.8389745,2.3630772,1.7066668,1.204513,1.1224617,1.1979488,1.5360001,1.8609232,1.9364104,1.5786668,1.5983591,1.6311796,1.6902566,1.6804104,1.3981539,1.4998976,1.4145643,1.6246156,1.9626669,1.6278975,1.214359,1.591795,1.8412309,1.7066668,1.591795,1.9823592,2.0873847,2.1431797,2.0906668,1.5885129,1.5392822,1.522872,1.522872,1.7165129,2.4746668,2.8947694,3.0884104,3.0654361,2.917744,2.806154,2.8389745,3.0720003,3.442872,3.7021542,3.4067695,3.5741541,4.312616,5.0051284,5.277539,5.0018463,4.663795,4.240411,4.0303593,3.9811285,3.6890259,2.9505644,2.8356924,3.0523078,3.4527183,4.023795,5.7468724,6.5312824,7.0859494,7.765334,8.579283,7.8473854,7.194257,7.1515903,7.456821,7.066257,3.767795,3.6463592,3.8006158,3.9876926,4.1058464,4.164923,4.9460516,5.8190775,6.806975,7.6668725,7.8736415,8.533334,8.395488,7.8080006,7.328821,7.719385,8.050873,8.280616,8.572719,8.979693,9.429334,9.91836,10.075898,10.200616,10.522257,11.23118,12.048411,12.379898,12.662155,13.305437,14.710155,14.050463,13.282462,13.59754,14.86113,15.593027,16.997746,19.026052,20.41108,22.019283,26.840618,31.625849,37.69108,44.17313,52.017235,63.980312,77.138054,78.61826,67.79734,49.67385,34.868515,26.59118,18.395899,11.592206,6.7807183,3.876103,3.436308,3.1606157,2.9243078,2.733949,2.7470772,2.8816411,2.6387694,2.034872,1.3620514,1.1913847,0.82379496,1.079795,1.3620514,1.4539489,1.5261539,1.3292309,1.079795,0.7811283,0.5152821,0.44307697,0.39384618,0.45620516,0.36430773,0.17394873,0.25928208,0.25928208,0.15753847,0.10502565,0.12143591,0.12143591,0.098461546,0.06564103,0.04594872,0.03938462,0.016410258,0.0032820515,0.0,0.02297436,0.1148718,0.33476925,0.27569234,1.083077,1.5524104,1.3193847,0.8533334,0.574359,0.256,0.06564103,0.06564103,0.21333335,0.22646156,0.27569234,0.512,1.1651284,2.5337439,1.6049232,1.2996924,1.6968206,2.6715899,3.889231,4.1583595,3.6496413,3.0818465,2.6026669,1.785436,1.2603078,1.8970258,2.540308,2.5895386,2.028308,1.332513,1.7362052,2.2055387,2.294154,2.1366155,1.6114873,3.5774362,4.6867695,4.670359,6.3179493,6.439385,6.626462,6.8463597,6.941539,6.636308,6.173539,5.435077,5.5072823,6.3310776,6.6822567,7.781744,8.149334,8.562873,9.163487,9.4457445,11.07036,12.711386,13.797745,13.732103,11.900719,12.025436,12.12718,11.608616,10.65354,10.240001,9.957745,9.649232,9.997129,10.906258,11.503591,13.078976,14.546052,15.350155,15.284514,14.464001,14.562463,13.945437,14.588719,16.282257,16.646564,15.376411,13.164309,11.74318,11.319796,10.57477,11.136001,11.697231,11.769437,11.562668,11.979488,12.514462,13.410462,14.171899,14.473847,14.145642,13.4859495,13.174155,12.1238985,10.502565,9.734565,8.283898,7.4699492,8.746667,11.346052,12.297847,11.749744,11.631591,11.32636,10.686359,10.039796,9.941334,9.396514,8.736821,7.9852314,6.8496413,6.5936418,6.87918,6.8594875,6.564103,6.882462,7.3452315,6.675693,6.4065647,6.9021544,7.3550773,7.197539,7.312411,7.5552826,7.9097443,8.484103,8.582564,9.997129,11.579078,12.95754,14.555899,12.786873,11.254155,10.492719,10.834052,12.419283,13.275898,13.764924,14.775796,16.150976,16.662975,15.599591,14.805334,14.339283,14.378668,15.199181,15.172924,16.403694,17.831387,18.60595,18.080822,16.384,14.851283,14.486976,15.360002,16.617027,14.54277,15.067899,16.246155,16.275694,13.505642,14.772514,14.890668,14.381949,13.5548725,12.481642,12.895181,12.763899,13.354668,14.667488,15.412514,11.736616,10.919386,10.358154,9.314463,8.910769,8.838565,8.379078,8.385642,8.582564,7.568411,6.944821,5.756718,5.2414365,5.6320004,6.1341543,4.450462,2.809436,1.7723079,1.5622566,2.0742567,4.699898,4.450462,4.161641,5.028103,6.5772314,2.6453335,1.2800001,1.4802053,2.481231,3.7382567,4.8607183,8.759795,10.417232,8.326565,4.457026,5.1265645,4.8016415,5.2348723,6.75118,8.241231,7.7259493,6.820103,5.832206,4.8016415,3.495385,3.3345644,3.5971284,4.2338467,5.2742567,6.8365135,5.76,5.0904617,4.059898,2.605949,1.3718976,0.7515898,0.84348726,1.1716924,1.4834872,1.7394873,3.2787695,3.131077,3.1967182,4.391385,6.636308,7.026872,6.8233852,6.3245134,5.474462,3.876103,3.2886157,4.1222568,4.31918,3.8596926,4.775385,7.387898,6.695385,4.571898,2.5665643,1.9068719,1.6377437,2.1300514,2.9735386,3.8596926,4.59159,4.9099493,7.1581545,9.42277,10.873437,11.762873,9.4457445,6.7971287,5.024821,5.0051284,7.2631803,10.374565,13.561437,14.355694,12.471796,9.810052,8.310155,7.634052,7.686565,8.418462,9.810052,8.579283,7.6668725,6.665847,5.4547696,4.197744,4.673641,5.149539,4.6900516,3.5774362,3.2951798,3.1113849,2.2416413,1.7001027,1.7394873,1.8609232,2.6912823,1.4998976,0.38728207,0.11158975,0.07548718,0.052512825,0.04594872,0.03938462,0.049230773,0.12143591,0.15753847,0.08533334,0.07876924,0.18051283,0.28882053,0.27897438,0.24615386,0.19364104,0.13784617,0.13784617,0.15097436,0.19692309,0.28225642,0.36758977,0.36758977,0.29210258,0.26584616,0.25928208,0.25928208,0.25928208,0.25928208,0.39712822,0.52512825,0.65641034,0.9616411,1.1815386,1.4933335,1.7558975,2.0841026,2.8521028,4.2207184,5.0215387,5.5565133,5.87159,5.737026,7.069539,6.5411286,5.720616,5.2381544,4.7622566,5.6287184,6.117744,6.308103,6.36718,6.560821,7.2205133,7.5946674,8.018052,8.444718,8.467693,8.674462,8.5891285,8.67118,8.953437,9.065026,8.149334,7.571693,7.5421543,7.719385,7.2172313,6.8397956,6.452513,5.9930263,5.865026,6.928411,6.5378466,6.5312824,7.0367184,7.7423596,7.890052,8.461129,8.55959,8.5661545,8.549745,8.27077,7.75877,7.3714876,7.325539,7.4469748,7.200821,7.2861543,7.6767187,7.748924,7.243488,6.2555904,6.0356927,5.687795,5.7435904,6.304821,7.0498466,7.830975,8.283898,8.484103,8.576,8.759795,7.9163084,7.3682055,6.75118,6.3573337,7.125334,7.2861543,8.267488,9.028924,9.501539,10.57477,12.563693,12.566976,9.747693,5.5663595,3.7842054,4.969026,4.6867695,4.345436,4.453744,4.6244106,2.865231,2.9210258,2.5961027,1.6869745,1.9692309,1.723077,1.4802053,2.5665643,4.46359,4.8049235,6.564103,7.3682055,6.0324106,3.9122055,4.9132314,4.194462,4.023795,3.2361028,1.9790771,1.7099489,2.428718,1.719795,1.2504616,1.4769232,1.6475899,2.1366155,1.9659488,2.044718,2.4648206,2.5009232,3.0162053,3.0523078,2.930872,2.9604106,3.4494362,3.2656412,2.8258464,2.428718,2.356513,2.868513,3.3312824,3.2000003,3.0720003,3.0490258,2.7306669,2.92759,3.2328207,3.6529233,4.06318,4.197744,4.4406157,4.2994876,4.07959,3.8728209,3.5544617,3.6036925,4.010667,4.2174363,4.138667,4.1517954,4.5423594,4.713026,4.8082056,4.8738465,4.8377438,4.4964104,4.31918,4.562052,5.0609236,5.218462,5.3398976,4.9394875,4.7589746,4.8771286,4.7294364,5.4383593,5.677949,5.612308,5.6352825,6.3934364,6.6625648,6.160411,6.124308,6.49518,5.920821,5.3694363,6.232616,6.1078978,4.7655387,4.1189747,5.110154,5.658257,5.8781543,5.7468724,5.110154,6.173539,6.485334,6.1374364,5.605744,5.7534366,4.9099493,4.663795,4.650667,4.6244106,4.4406157,4.135385,3.629949,3.0851285,2.6518977,2.4582565,2.225231,2.7076926,3.1343591,3.1770258,2.9440002,2.553436,1.9790771,1.5163078,1.2931283,1.2832822,1.3686155,1.7001027,2.0217438,2.1530259,1.9692309,2.0184617,1.8740515,1.7329233,1.6672822,1.6180514,1.6410258,1.5753847,1.7099489,1.9692309,1.9068719,1.6508719,1.9364104,1.9167181,1.5064616,1.3718976,1.8609232,1.9462565,1.972513,1.9561027,1.6016412,1.5425643,1.3259488,1.4539489,2.0118976,2.6715899,2.865231,2.9505644,2.8225644,2.5731285,2.487795,3.0490258,3.508513,3.8038976,3.9056413,3.8465643,3.564308,4.2272825,4.8311796,4.9296412,4.6244106,4.6966157,4.5489235,4.397949,4.164923,3.495385,2.8717952,2.6617439,2.8750772,3.4724104,4.3651285,5.720616,6.7183595,7.2369237,7.466667,7.9195905,7.4929237,7.8145647,7.9327188,7.5881033,7.24677,3.4034874,3.748103,4.1813335,4.338872,4.266667,4.384821,5.4416413,6.052103,6.8693337,7.781744,7.9097443,7.955693,8.050873,7.9327188,7.53559,6.987488,7.532308,8.41518,9.222565,9.7214365,9.882257,9.764103,9.793642,10.112,10.679795,11.280411,12.038565,12.314258,12.281437,12.356924,13.184001,13.042872,12.438975,12.461949,13.410462,14.788924,16.026258,17.51959,19.429745,22.386873,27.510157,31.64226,37.75672,44.875492,53.983185,68.043495,76.22237,69.6878,54.803696,38.21949,26.86031,20.007385,13.10195,7.8769236,4.8311796,3.2032824,2.8225644,2.3893335,2.0512822,1.8740515,1.8051283,1.9987694,1.9987694,1.8051283,1.4966155,1.2406155,0.75487185,0.7187693,0.9353847,1.2635899,1.6114873,1.394872,1.0108719,0.7056411,0.57764107,0.56451285,0.4955898,0.43651286,0.3446154,0.256,0.28225642,0.23630771,0.13784617,0.07548718,0.072205134,0.072205134,0.029538464,0.013128206,0.009846155,0.006564103,0.0032820515,0.009846155,0.049230773,0.118153855,0.20348719,0.2855385,0.3052308,0.6268718,0.9878975,1.1848207,1.0633847,1.1126155,0.60061544,0.23630771,0.2297436,0.2855385,0.26912823,0.71548724,1.7591796,2.6880002,1.9462565,2.7864618,3.1507695,3.3509746,3.387077,2.92759,3.5971284,2.7306669,2.2088206,2.3827693,2.103795,1.9790771,2.5337439,2.5600002,2.0512822,2.2121027,2.0742567,1.9200002,2.1300514,2.793026,3.698872,3.751385,4.5423594,4.857436,4.906667,6.3277955,5.3760004,5.1265645,5.5072823,6.1374364,6.3212314,5.1922054,4.457026,4.6112823,5.671385,7.1581545,7.3485136,6.626462,7.0367184,8.39877,8.297027,9.882257,11.405129,12.560411,12.596514,10.315488,10.837335,10.9456415,10.305642,8.982975,7.456821,8.598975,9.6525135,10.512411,10.9915905,10.79795,11.963078,13.574565,14.12595,13.328411,12.11077,13.124924,13.564719,14.181745,15.1466675,16.049232,15.717745,13.013334,10.601027,9.337437,8.280616,9.3768215,11.011283,11.959796,12.163283,12.73436,13.252924,13.423591,13.59754,13.584412,12.668719,12.301129,12.232206,11.910565,10.988309,9.321027,8.375795,8.3364105,8.917334,10.144821,12.347078,12.763899,12.947693,12.356924,11.2672825,10.735591,9.711591,9.035488,8.3134365,7.5388722,7.0957956,6.554257,6.6822567,6.892308,7.017026,7.2960005,7.762052,6.928411,6.439385,6.7840004,7.2927184,7.427283,7.719385,8.057437,8.339693,8.484103,8.697436,9.442462,10.568206,12.11077,14.276924,13.755078,12.163283,10.988309,11.2672825,13.5548725,14.995693,14.677335,15.38954,17.362053,18.287592,17.51631,16.662975,15.665232,15.113848,16.22318,16.042667,16.948515,18.028309,18.582975,18.107079,17.463797,16.239592,15.770258,16.170668,16.324924,15.537232,16.085335,16.646564,16.610462,16.068924,15.002257,14.27036,14.345847,14.805334,14.336001,14.096412,13.124924,12.47836,12.668719,13.666463,10.850462,10.020103,9.517949,8.982975,9.350565,8.779488,8.438154,8.457847,8.585847,8.178872,8.602257,7.328821,7.059693,7.9097443,7.4043083,7.017026,5.549949,3.4297438,1.5885129,1.4769232,2.4516926,2.28759,2.0151796,2.1136413,2.5107694,1.3751796,0.8960001,1.4736412,2.7602053,3.6660516,7.7357955,8.937026,9.29477,9.38995,8.362667,8.310155,7.269744,6.193231,5.914257,7.141744,8.192,7.90318,7.250052,6.4065647,4.7392826,3.8662567,3.7021542,3.7710772,4.1780515,5.602462,5.408821,4.3618464,2.8980515,1.5458462,0.95835906,0.81394875,0.7778462,1.0043077,1.394872,1.591795,2.878359,3.5610259,4.886975,6.9054365,8.467693,7.384616,7.177847,6.695385,5.35959,3.1540515,2.3072822,3.9089234,5.0543594,5.2742567,6.521436,9.124104,10.985026,11.907283,11.746463,10.404103,5.5138464,2.8455386,2.1169233,2.5337439,2.7864618,4.2272825,5.1167183,6.550975,8.674462,10.679795,9.705027,8.815591,7.8736415,6.8562055,5.8223596,7.256616,8.579283,9.685334,10.315488,10.069334,10.870154,9.691898,8.996103,9.412924,9.750975,8.753231,7.9852314,7.0400004,5.9963083,5.4547696,5.723898,5.681231,5.0576415,3.9844105,2.989949,2.5632823,3.062154,3.006359,2.612513,3.7907696,2.7437952,1.148718,0.20020515,0.101743594,0.06564103,0.049230773,0.098461546,0.12471796,0.10502565,0.06235898,0.108307704,0.059076928,0.055794876,0.13128206,0.19364104,0.17066668,0.23958977,0.24287182,0.17066668,0.15097436,0.190359,0.27569234,0.29210258,0.24287182,0.24287182,0.25928208,0.33476925,0.33805132,0.27241027,0.28225642,0.30194873,0.39384618,0.508718,0.6498462,0.88943595,1.214359,1.5753847,1.785436,1.9364104,2.4155898,3.889231,4.457026,4.926359,5.533539,5.9569235,7.384616,6.9710774,5.865026,4.8640003,4.4077954,5.1856413,5.7140517,6.4000006,7.145026,7.328821,8.684308,9.252103,9.268514,9.019077,8.848411,8.723693,8.67118,8.4512825,8.132924,8.086975,7.8539495,7.4863596,7.1023593,6.7544622,6.413129,5.9930263,5.910975,5.8880005,5.924103,6.2916927,6.2063594,6.436103,7.1122055,7.975385,8.375795,8.326565,8.362667,8.388924,8.310155,8.050873,7.4404106,7.3321033,7.565129,7.857231,7.788308,7.4732313,7.4765134,7.5618467,7.5520005,7.3058467,7.4371285,7.0892315,6.7249236,6.695385,7.243488,7.4896417,7.9294367,8.146052,7.9195905,7.243488,6.9120007,6.619898,6.5247183,6.764308,7.456821,7.7981544,8.36595,8.667898,8.822155,9.573745,11.290257,10.571488,8.034462,4.962462,3.308308,3.8662567,4.4406157,5.142975,6.1538467,7.712821,5.865026,4.4340515,2.8717952,1.4933335,1.4802053,1.1979488,1.7132308,2.3040001,2.9768207,4.453744,5.4974365,5.76,5.0116925,3.6857438,2.8521028,2.7536411,3.5905645,3.2951798,2.0906668,2.4648206,2.3860514,2.0545642,1.9265642,2.0742567,2.1858463,2.0676925,2.0250258,2.03159,2.1530259,2.550154,2.5271797,2.5698464,2.5698464,2.5731285,2.789744,2.4320002,2.1300514,1.9889232,2.048,2.3072822,2.5764105,2.5796926,2.7470772,3.0982566,3.2196925,3.239385,3.318154,3.8071797,4.519385,4.7327185,4.781949,4.345436,3.8596926,3.5446157,3.383795,3.7448208,4.141949,4.4045134,4.525949,4.673641,4.772103,4.6080003,4.5095387,4.5423594,4.4964104,4.279795,4.1485133,4.2535386,4.57518,4.9362054,4.972308,4.785231,4.713026,4.7950773,4.7655387,5.074052,5.287385,5.5532312,6.1407185,7.456821,6.961231,6.170257,5.83877,5.8289237,5.0904617,5.1167183,6.2687182,6.6494365,5.664821,4.023795,5.0116925,6.1538467,7.062975,7.213949,5.9536414,5.8256416,6.2851286,6.6395903,6.5411286,5.98318,5.85518,5.353026,4.824616,4.637539,5.1954875,4.6080003,3.8104618,3.511795,3.5872824,3.0785644,2.7011285,2.8389745,3.0720003,3.0654361,2.5895386,2.1136413,1.8182565,1.6278975,1.529436,1.5753847,1.6410258,2.048,2.3860514,2.5173335,2.5796926,2.1300514,1.8904617,1.8379488,1.8248206,1.5819489,1.5458462,1.3784616,1.3883078,1.6344616,1.8937438,1.6869745,1.5425643,1.3981539,1.2898463,1.3620514,1.9265642,1.8642052,1.6213335,1.4539489,1.4309745,1.5360001,1.3817437,1.4539489,1.9068719,2.5862565,2.789744,3.0687182,3.0720003,2.865231,2.92759,3.4297438,3.7087183,3.7809234,3.7809234,3.9417439,3.5741541,3.5183592,3.8432825,4.4242053,4.9394875,4.778667,4.604718,4.5522056,4.4373336,3.7251284,2.986667,2.740513,2.9078977,3.4691284,4.450462,5.3760004,7.1089234,8.237949,8.162462,7.0892315,7.24677,7.2205133,7.003898,6.685539,6.4295387,3.2000003,3.4822567,3.7940516,3.9647183,4.069744,4.4307694,5.2381544,5.6943593,6.377026,7.282872,7.8539495,7.680001,7.8145647,7.955693,7.765334,6.8594875,7.2172313,8.214975,9.350565,10.066052,9.757539,9.590155,9.701744,10.240001,11.001437,11.428103,12.274873,12.268309,12.045129,11.835078,11.464206,11.264001,11.050668,11.1294365,11.776001,13.233232,15.1466675,17.010874,19.580719,23.315695,28.383183,32.672825,39.19098,47.36985,57.92821,72.86154,74.76842,63.11385,45.83713,29.459694,19.078566,13.420309,8.966565,5.8453336,3.9286156,2.8258464,2.3860514,2.041436,1.8674873,1.8248206,1.7460514,1.8510771,1.8740515,1.7165129,1.3883078,1.014154,0.72861546,0.60389745,0.6695385,0.8795898,1.1191796,0.95835906,0.702359,0.5021539,0.41682056,0.40369233,0.39712822,0.38728207,0.33476925,0.25271797,0.19692309,0.13128206,0.068923086,0.03938462,0.04594872,0.052512825,0.009846155,0.016410258,0.016410258,0.0032820515,0.009846155,0.04266667,0.2231795,0.49887183,0.75487185,0.8336411,0.51856416,0.5218462,0.73517954,1.020718,1.204513,1.2373334,0.6892308,0.31507695,0.33476925,0.42338464,0.90584624,1.591795,2.0578463,2.1989746,2.2482052,2.8488207,3.4691284,3.6660516,3.6135387,4.1058464,3.4166157,2.4516926,2.4648206,3.1245131,2.5009232,2.412308,2.802872,2.605949,1.9889232,2.359795,2.2580514,2.2022567,2.605949,3.564308,4.8672824,4.6145644,4.3027697,3.8859491,3.7415388,4.6834874,5.1987696,5.277539,5.467898,5.723898,5.398975,5.3070774,5.654975,6.1505647,6.5247183,6.5378466,6.550975,7.77518,10.006975,11.9860525,11.388719,11.286975,11.749744,12.179693,11.959796,10.476309,11.195078,10.305642,9.176616,8.3593855,7.5913854,7.958975,8.907488,9.865847,10.315488,9.777231,10.985026,12.100924,12.78359,12.839386,12.2157955,12.340514,12.461949,12.852514,13.673027,14.966155,14.486976,12.86236,11.208206,9.833026,8.228104,8.631796,10.689642,12.452104,13.289026,13.8765135,13.679591,13.026463,12.5374365,12.393026,12.33395,11.713642,11.483898,11.365745,11.008,10.003693,9.206155,9.002667,9.344001,10.161232,11.372309,11.648001,12.117334,12.120616,11.513436,10.663385,9.074872,8.621949,8.155898,7.4371285,7.1122055,6.6822567,6.5247183,6.7774363,7.243488,7.3714876,7.653744,7.13518,6.669129,6.6592827,7.066257,7.6570263,8.152616,8.884514,9.724719,10.105436,9.764103,9.728001,10.328616,11.766154,14.132514,14.788924,13.643488,12.294565,12.163283,14.490257,16.187078,15.402668,15.189335,16.62031,18.809437,18.83241,18.569847,17.821539,17.10277,17.641027,17.58195,17.93641,18.011898,17.716515,17.552412,17.161848,16.269129,16.09518,16.705643,16.99118,16.886156,17.34236,17.404718,17.178257,17.834667,14.818462,13.571283,14.034052,15.307488,15.635694,15.281232,13.515489,12.005745,11.815386,13.413745,11.096616,9.803488,9.061745,8.864821,9.662359,8.687591,8.333129,8.388924,8.434873,7.8637953,8.306872,8.753231,9.908514,10.528821,7.427283,7.4240007,6.245744,5.333334,4.893539,3.8990772,2.1464617,1.270154,0.9714873,0.9517949,0.94523084,1.0929232,1.0929232,1.2964103,2.7700515,7.2992826,12.461949,12.212514,9.856001,7.650462,6.7840004,7.834257,8.854975,9.065026,8.507077,8.04759,8.828718,9.540924,9.714872,8.769642,6.0028725,4.857436,4.332308,4.20759,4.3749747,4.827898,4.2601027,2.7864618,1.5786668,1.2242053,1.7427694,1.8806155,1.7296412,1.4769232,1.2242053,0.99774367,2.0151796,2.802872,4.2338467,6.0225644,6.747898,6.166975,6.957949,6.941539,5.691077,4.522667,3.0194874,3.2295387,3.6036925,3.8629746,4.9887185,7.1515903,9.964309,12.566976,13.51877,10.79795,6.2129235,3.4067695,2.0775387,1.7920002,1.9790771,2.9078977,3.9023592,4.972308,6.1308722,7.4043083,5.874872,5.7731285,6.5411286,7.207385,6.377026,7.194257,7.5520005,7.7325134,7.7357955,7.2861543,8.195283,7.9950776,7.6931286,7.716103,7.9228725,7.1515903,6.931693,6.626462,6.121026,5.8125134,5.924103,5.8256416,5.2742567,4.414359,3.7940516,3.7152824,3.8662567,3.7284105,3.5774362,4.493129,2.1497438,0.7253334,0.14769232,0.14441027,0.21661541,0.17394873,0.21333335,0.2231795,0.17723078,0.118153855,0.118153855,0.098461546,0.098461546,0.118153855,0.13128206,0.16410258,0.24287182,0.25271797,0.20020515,0.190359,0.28225642,0.3446154,0.35774362,0.3314872,0.2855385,0.3249231,0.37415388,0.34789747,0.27241027,0.2986667,0.3314872,0.39056414,0.5218462,0.76800007,1.1716924,1.6443079,1.7526156,1.6902566,1.7526156,2.3696413,3.5413337,3.7776413,4.135385,5.208616,7.1483083,8.5202055,7.7390776,6.436103,5.3169236,4.161641,4.8672824,5.4514875,6.3474874,7.210667,6.918565,8.260923,8.592411,8.536616,8.539898,8.868103,8.4053335,7.9458466,7.581539,7.4075904,7.5421543,7.2369237,7.062975,6.665847,6.121026,5.927385,5.5269747,5.464616,5.7074876,6.0225644,5.9602056,5.940513,6.954667,8.211693,9.032206,8.828718,8.5202055,8.3593855,8.044309,7.6635904,7.7292314,7.958975,8.339693,8.592411,8.539898,8.100103,7.683283,7.5388722,7.53559,7.5388722,7.4043083,7.1909747,6.75118,6.5772314,6.875898,7.568411,7.6701546,8.146052,8.379078,8.027898,7.0498466,6.51159,6.242462,6.436103,7.026872,7.6767187,7.5618467,7.837539,8.277334,8.786052,9.416205,10.30236,9.905231,7.821129,5.297231,5.2480006,4.266667,4.279795,5.2545643,6.7840004,8.080411,7.24677,4.8049235,2.4188719,1.0962052,1.1946667,1.1126155,1.4539489,1.723077,2.1464617,3.6693337,3.6036925,4.020513,3.876103,2.9111798,1.6377437,1.5688206,2.3040001,2.7831798,2.7831798,2.9013336,2.7011285,2.5042052,2.3794873,2.3893335,2.5764105,2.169436,2.103795,1.9593848,1.7920002,2.1431797,2.231795,2.3105643,2.281026,2.2678976,2.605949,2.3072822,2.0841026,1.9429746,1.8904617,1.9003079,2.546872,2.7766156,2.986667,3.2164104,3.1507695,3.2918978,3.6594875,4.128821,4.5522056,4.7392826,4.6966157,4.417641,4.013949,3.629949,3.4789746,3.8367183,4.2272825,4.31918,4.1846156,4.3027697,4.2240005,4.096,4.125539,4.2830772,4.2994876,4.1156926,3.826872,3.7907696,4.1156926,4.647385,4.588308,4.5817437,4.578462,4.578462,4.637539,4.818052,5.110154,5.5762057,6.294975,7.3714876,6.8430777,6.6461544,6.439385,6.009436,5.293949,5.179077,5.8092313,6.452513,6.2884107,4.417641,4.903385,5.907693,6.9087186,7.39118,6.8594875,6.058667,6.091488,6.4065647,6.49518,5.8880005,5.8190775,5.504,4.893539,4.44718,5.149539,4.634257,3.8695388,3.5610259,3.5741541,2.9243078,2.8225644,3.1737437,3.3608208,3.186872,2.878359,2.2613335,1.9003079,1.6246156,1.4375386,1.5195899,1.8445129,2.2449234,2.5764105,2.7700515,2.8422565,2.2908719,1.8248206,1.785436,2.0742567,2.1398976,1.7690258,1.5261539,1.4802053,1.6311796,1.9003079,1.8018463,1.6508719,1.4473847,1.2603078,1.2209232,1.8215386,1.6968206,1.3718976,1.1848207,1.2964103,1.6278975,1.6443079,1.6213335,1.7952822,2.3630772,2.6945643,3.0227695,3.131077,3.062154,3.1376412,3.6036925,3.7743592,3.8629746,4.010667,4.2962055,4.1846156,3.9975388,4.135385,4.6112823,5.037949,4.716308,4.594872,4.781949,4.841026,3.7842054,3.1245131,2.9078977,3.0752823,3.564308,4.2863593,4.7983594,6.5706673,7.7390776,7.64718,6.8463597,7.4371285,7.824411,7.6701546,7.0957956,6.7117953,3.0424619,3.3280003,3.4691284,3.5511796,3.764513,4.417641,4.7491283,5.080616,5.7632823,6.692103,7.318975,7.1483083,7.125334,7.39118,7.6242056,7.0367184,6.948103,7.752206,8.89436,9.741129,9.573745,9.862565,10.180923,10.509129,10.883283,11.405129,12.2847185,12.12718,11.82195,11.631591,11.172104,10.515693,10.295795,10.66995,11.565949,12.678565,15.195899,17.585232,20.594873,24.546463,29.334976,34.661747,42.262978,52.000824,64.17724,79.53724,77.003494,61.47939,41.951183,25.045336,15.015386,10.259693,7.3714876,5.481026,4.1747694,3.4789746,3.4560003,3.2525132,2.8717952,2.4188719,2.1070771,1.913436,1.8674873,1.654154,1.2307693,0.8008206,1.0666667,1.1782565,1.020718,0.7778462,0.9321026,0.6235898,0.45292312,0.34789747,0.27897438,0.26912823,0.3052308,0.37415388,0.3314872,0.19364104,0.12471796,0.09189744,0.055794876,0.032820515,0.026256412,0.032820515,0.055794876,0.04594872,0.03938462,0.059076928,0.108307704,0.059076928,0.20348719,0.446359,0.69907695,0.8763078,0.702359,0.7384616,0.90584624,1.0568206,0.9682052,0.98461545,0.5513847,0.28225642,0.41682056,0.8566154,1.0469744,1.4276924,1.4244103,1.2504616,1.9265642,2.097231,2.7864618,3.2754874,3.5380516,4.2436924,2.8717952,2.5862565,2.605949,2.6354873,2.868513,2.8422565,3.121231,2.7798977,2.1825643,2.9702566,2.4582565,2.5074873,3.3608208,4.7360005,5.8486156,4.7294364,3.5511796,2.8192823,2.8160002,3.623385,4.650667,4.9788723,5.028103,5.0838976,5.293949,5.58277,6.0225644,6.235898,6.377026,7.1154876,6.9021544,9.15036,12.228924,14.486976,14.276924,12.288001,11.395283,11.45436,11.733335,10.896411,11.47077,10.420513,9.419488,9.048616,8.802463,8.034462,8.418462,9.058462,9.373539,9.094564,10.640411,11.533129,12.320822,12.941129,12.727796,12.107488,11.851488,11.631591,11.634872,12.560411,12.507898,12.593232,12.087796,10.912822,9.6295395,9.426052,10.607591,11.989334,13.092104,14.162052,13.472821,12.596514,11.910565,11.844924,12.891898,11.61518,10.745437,10.47959,10.617436,10.5780525,9.911796,9.268514,9.301334,9.813334,9.754257,9.9282055,10.587898,11.057232,11.08677,10.834052,9.120821,8.55959,8.241231,7.788308,7.3419495,6.9677954,6.675693,6.9645133,7.634052,7.788308,7.466667,7.325539,7.1154876,6.885744,6.951385,7.8145647,8.795898,9.944616,10.998155,11.369026,11.113027,10.919386,11.254155,12.425847,14.578873,15.00554,14.106257,13.233232,13.180719,14.201437,16.374155,16.003283,15.415796,15.944206,17.913437,18.264616,18.75036,18.927591,18.84554,19.03918,18.835693,18.586258,18.018463,17.270155,16.905848,16.548103,16.02954,16.341335,17.457232,18.33354,18.176,18.842258,18.468103,17.447386,18.432001,14.749539,13.282462,13.732103,15.16636,16.02954,15.366566,13.154463,11.437949,11.457642,13.676309,11.588924,10.006975,9.055181,8.815591,9.330873,8.661334,8.572719,8.477539,8.329846,8.6580515,8.251078,9.321027,10.630565,11.126155,9.924924,9.124104,6.426257,6.314667,8.969847,10.233437,3.7940516,1.3522053,0.7975385,0.7318975,0.47589746,1.0272821,1.214359,1.1388719,2.3466668,7.830975,13.4400015,12.2617445,8.592411,5.904411,6.8463597,6.7282057,8.871386,10.512411,10.601027,9.80677,9.248821,9.048616,8.828718,8.008205,5.796103,4.6211286,5.2742567,5.540103,4.6900516,3.4789746,2.5600002,1.3554872,0.84348726,1.4408206,3.0194874,4.013949,3.8728209,3.1442053,2.1070771,0.7778462,1.270154,1.6672822,3.1409233,5.3858466,6.619898,5.8092313,7.0498466,7.640616,6.8332314,5.858462,4.263385,2.793026,2.0742567,2.2186668,2.7995899,4.201026,6.0324106,8.01477,9.179898,7.8506675,5.037949,3.1474874,2.225231,2.097231,2.349949,2.4385643,3.370667,5.159385,6.73477,5.933949,3.2164104,2.858667,4.1485133,5.9634876,6.764308,8.740103,8.704,7.4469748,6.121026,6.235898,6.2227697,7.5913854,7.8539495,6.7150774,6.0783596,6.2194877,6.196513,5.920821,5.4875903,5.156103,5.421949,5.405539,4.9854364,4.31918,3.879385,3.4625645,3.7973337,4.2535386,4.2469745,3.2361028,1.2307693,0.3511795,0.101743594,0.13456412,0.25271797,0.2231795,0.21661541,0.20348719,0.17723078,0.16738462,0.118153855,0.098461546,0.09189744,0.098461546,0.12471796,0.18379489,0.23958977,0.24287182,0.20020515,0.20020515,0.37743592,0.37743592,0.38400003,0.4397949,0.46933338,0.47261542,0.4397949,0.36430773,0.29538465,0.3117949,0.36758977,0.41025645,0.52512825,0.75487185,1.1060513,1.8871796,2.0906668,1.9331284,1.8609232,2.5698464,3.249231,3.383795,3.9154875,5.540103,8.73354,9.570462,8.086975,6.665847,5.87159,4.450462,5.0084105,5.211898,5.737026,6.3573337,5.940513,7.059693,7.7948723,8.228104,8.470975,8.648206,7.975385,7.325539,7.1581545,7.3682055,7.273026,6.7938466,7.0498466,6.9021544,6.2555904,6.0619493,6.0717955,5.9503593,5.979898,6.114462,5.9667697,6.229334,7.4043083,8.553026,9.120821,8.92718,8.792616,8.395488,7.762052,7.2664623,7.637334,8.086975,8.379078,8.470975,8.323282,7.893334,7.719385,7.785026,7.8014364,7.7423596,7.837539,7.1548724,6.4656415,6.3343596,6.7610264,7.1844106,7.453539,8.093539,8.392206,8.060719,7.250052,6.488616,6.3376417,6.409847,6.521436,6.692103,6.9349747,7.197539,7.7259493,8.418462,8.841846,9.140513,8.448001,6.636308,4.955898,6.0619493,4.525949,4.1682053,5.208616,6.567385,5.8486156,5.9536414,3.7054362,1.5589745,0.6892308,0.99774367,1.1749744,1.214359,1.3620514,1.7165129,2.2350771,1.9954873,2.6322052,2.6945643,1.8838975,1.0699488,1.3423591,1.6804104,2.3762052,3.1113849,2.92759,2.605949,2.7437952,2.917744,3.0916924,3.6496413,2.6518977,2.231795,1.8445129,1.4900514,1.719795,1.8346668,1.8707694,1.9003079,1.9954873,2.2350771,2.044718,1.9200002,1.8445129,1.847795,1.9790771,2.5862565,2.993231,3.373949,3.7284105,3.892513,3.9253337,4.1058464,4.2962055,4.5095387,4.896821,4.7425647,4.4800005,4.1091285,3.7218463,3.515077,3.6168208,3.889231,4.0434875,4.1091285,4.450462,4.0533338,3.9942567,4.0467696,4.1091285,4.1911798,4.1091285,3.8859491,3.8498464,4.092718,4.4898467,4.4242053,4.522667,4.6276927,4.6802053,4.71959,4.7950773,5.2709746,5.9634876,6.6461544,7.030154,6.9809237,7.171283,7.0925136,6.616616,5.98318,5.6352825,5.910975,6.7314878,7.2237954,5.717334,5.290667,5.8453336,6.5444107,7.026872,7.433847,6.6034875,6.12759,6.0750775,6.2588725,6.23918,6.045539,5.924103,5.293949,4.522667,4.9099493,4.391385,3.6824617,3.314872,3.2065644,2.6617439,2.789744,3.2853336,3.442872,3.186872,3.0654361,2.5271797,2.225231,1.8543591,1.467077,1.4769232,1.8838975,2.3991797,2.8422565,3.0949745,3.0916924,2.5042052,1.910154,1.7657437,2.044718,2.2383592,1.7985642,1.6246156,1.522872,1.4867693,1.7132308,1.8379488,1.7887181,1.654154,1.5031796,1.3686155,1.6246156,1.4408206,1.1946667,1.1520001,1.4572309,1.7657437,1.8445129,1.8281027,1.8838975,2.2088206,2.5271797,2.7963078,2.9111798,2.92759,3.045744,3.4527183,3.5183592,3.6758976,4.0336413,4.381539,4.3684106,4.325744,4.5095387,4.8771286,5.0674877,4.667077,4.601436,4.95918,5.100308,3.6332312,3.2984617,3.2032824,3.318154,3.620103,4.1058464,4.345436,5.691077,6.692103,6.997334,7.3386674,8.316719,9.025641,8.917334,8.093539,7.3025646,2.8849232,3.3575387,3.4198978,3.3444104,3.4921029,4.2929235,4.2436924,4.522667,5.2545643,6.12759,6.3967185,6.3376417,6.1472826,6.426257,7.030154,7.0367184,6.7840004,7.2369237,8.004924,8.795898,9.416205,10.148104,10.620719,10.545232,10.31877,11.040821,11.795693,11.611898,11.286975,11.250873,11.556104,10.820924,10.443488,11.16554,12.678565,13.617231,16.259283,18.97354,22.04554,25.731283,30.293335,37.35631,46.900517,58.8078,72.562874,87.26975,81.86749,63.172928,41.87898,25.032207,16.022976,12.002462,9.6295395,8.224821,7.4010262,7.059693,7.463385,6.9152827,5.72718,4.3618464,3.4330258,2.6289232,2.2711797,1.8642052,1.2996924,0.8795898,1.5786668,1.9954873,1.7099489,1.0469744,1.0929232,0.5907693,0.41025645,0.35774362,0.33805132,0.33476925,0.35446155,0.40697438,0.3249231,0.13784617,0.09189744,0.11158975,0.08205129,0.04266667,0.01969231,0.02297436,0.108307704,0.10502565,0.128,0.18707694,0.20676924,0.07548718,0.08205129,0.101743594,0.17723078,0.512,0.90256417,1.1257436,1.3128207,1.2898463,0.58092314,0.65641034,0.38728207,0.20676924,0.40697438,1.1290257,0.5546667,0.42338464,0.58420515,0.8369231,0.9419488,1.2176411,1.8412309,2.868513,3.82359,3.69559,2.609231,2.8291285,2.412308,1.6508719,3.058872,2.9210258,3.31159,3.1113849,2.678154,3.8531284,2.9965131,2.7700515,3.764513,5.4416413,6.1472826,4.240411,2.8750772,2.3827693,2.7831798,3.767795,3.7087183,4.069744,4.3060517,4.57518,5.7403083,5.4514875,5.287385,5.142975,5.8223596,9.035488,8.470975,9.754257,12.032001,14.119386,14.49354,11.884309,10.361437,10.496001,11.401847,10.722463,10.811078,10.84718,10.857026,10.774975,10.456616,8.910769,8.891078,9.268514,9.524513,9.770667,11.352616,12.140308,12.737642,13.157744,12.816411,12.2617445,11.835078,10.948924,9.993847,10.331899,11.211488,12.251899,12.442257,11.795693,11.352616,11.034257,10.663385,10.735591,11.529847,13.115078,12.560411,12.156719,11.907283,12.117334,13.367796,11.61518,10.148104,9.619693,9.980719,10.476309,10.134975,9.393231,9.019077,8.963283,8.342975,8.697436,9.363693,9.80677,10.115283,10.994873,9.754257,8.789334,8.310155,8.132924,7.6635904,7.2664623,7.026872,7.381334,8.182155,8.681026,7.7357955,7.7292314,7.893334,7.8441033,7.581539,8.267488,9.609847,10.95877,11.851488,11.995898,12.3536415,12.373334,12.57354,13.403898,15.232001,14.355694,13.430155,13.446565,13.99795,13.279181,15.514257,16.07877,15.980309,15.90154,16.20677,16.105026,16.918976,18.028309,18.95713,19.393642,18.894772,18.379488,17.903591,17.352207,16.452925,15.872002,15.891693,16.810667,18.359797,19.721848,19.282053,20.050053,19.344412,17.440823,17.555695,14.897232,13.4629755,13.443283,14.39836,15.254975,14.263796,12.291283,10.929232,11.1064625,13.069129,11.52,10.177642,9.291488,8.881231,8.720411,8.937026,9.330873,8.818872,8.136206,9.829744,8.832001,9.110975,9.347282,9.91836,12.934566,10.515693,6.3179493,6.311385,10.880001,14.792206,5.7829747,2.556718,1.6836925,1.142154,0.3249231,0.76800007,0.9419488,1.0043077,1.9003079,5.3694363,10.581334,9.258667,6.5312824,5.920821,9.334154,6.550975,8.192,10.371283,11.250873,11.021129,8.982975,6.5837955,5.077334,4.568616,4.013949,3.1671798,5.3891287,6.189949,4.332308,1.8313848,1.1749744,0.7220513,0.82379496,1.7985642,3.9220517,5.691077,5.7042055,4.778667,3.3411283,1.4276924,1.2537436,1.3883078,3.3017437,6.672411,9.38995,6.925129,6.7872825,7.276308,7.1647186,5.681231,5.106872,3.446154,2.5435898,2.6715899,2.553436,3.0687182,2.9768207,2.9472823,3.4756925,4.896821,3.2623591,2.3893335,2.487795,3.1671798,3.4133337,3.2853336,3.7120004,6.498462,9.416205,6.2227697,3.7940516,3.498667,4.2141542,5.4153852,7.1844106,10.249847,10.039796,8.12636,6.5805135,7.975385,7.0859494,9.334154,9.961026,7.972103,6.1505647,7.282872,6.816821,5.7764106,4.916513,4.709744,5.3366156,4.923077,4.125539,3.4100516,3.0424619,1.972513,3.3378465,4.8114877,4.604718,1.4605129,0.51856416,0.12143591,0.029538464,0.072205134,0.15097436,0.16082053,0.15097436,0.128,0.12143591,0.15425642,0.098461546,0.055794876,0.04266667,0.068923086,0.15097436,0.190359,0.24287182,0.26584616,0.23958977,0.18707694,0.41682056,0.38400003,0.39712822,0.53825647,0.6629744,0.58092314,0.48902568,0.40369233,0.33805132,0.32820517,0.42338464,0.46276927,0.52512825,0.6432821,0.77128214,1.8904617,2.428718,2.3958976,2.228513,2.7995899,3.0490258,3.3936412,4.348718,6.3245134,9.6295395,9.6295395,7.962257,6.626462,6.0652313,5.146257,5.536821,4.9952826,4.821334,5.156103,4.9985647,5.8289237,7.53559,8.67118,8.772923,8.356103,7.8637953,7.4699492,7.5946674,7.830975,6.9710774,6.669129,7.3452315,7.4896417,6.892308,6.629744,7.213949,7.0793853,6.698667,6.4295387,6.5444107,7.213949,7.8047185,8.182155,8.41518,8.779488,8.937026,8.425026,7.7981544,7.4699492,7.722667,7.574975,7.4929237,7.5421543,7.6701546,7.706257,7.827693,8.15918,8.237949,8.15918,8.598975,7.6668725,6.747898,6.4722056,6.738052,6.7183595,7.0400004,7.5618467,7.7423596,7.50277,7.207385,6.436103,6.488616,6.3376417,5.792821,5.4843082,6.5050263,6.885744,7.2894363,7.7948723,7.893334,7.6307697,6.226052,4.8311796,4.315898,5.287385,4.342154,4.4767184,5.58277,6.1374364,3.2032824,3.259077,1.8904617,0.72861546,0.44964105,0.77128214,1.1126155,1.1191796,1.2964103,1.4834872,0.86317956,1.2307693,1.7690258,1.6278975,0.9616411,0.9189744,1.7296412,1.8182565,2.2088206,2.8750772,2.7470772,2.1464617,2.7241027,3.4198978,3.9680004,4.8771286,3.3378465,2.5829747,2.028308,1.5458462,1.4834872,1.3784616,1.3029745,1.4769232,1.7427694,1.5885129,1.4998976,1.5097437,1.6278975,1.913436,2.4746668,2.7208207,3.2032824,3.7710772,4.3618464,5.0018463,4.663795,4.266667,4.1452312,4.4373336,5.0642056,4.854154,4.4701543,4.06318,3.7054362,3.3936412,3.131077,3.1638978,3.5282054,4.164923,4.926359,4.4077954,4.391385,4.2994876,4.069744,4.1485133,4.2338467,4.2371287,4.2830772,4.342154,4.2469745,4.3027697,4.4865646,4.781949,5.0642056,5.080616,4.9460516,5.5991797,6.5378466,7.200821,6.997334,7.64718,7.716103,7.5618467,7.256616,6.5706673,6.294975,6.6494365,7.522462,8.2215395,7.4732313,6.1078978,6.1013336,6.298257,6.4656415,7.2894363,7.059693,6.482052,6.235898,6.5083084,7.000616,6.7282057,6.629744,5.976616,4.95918,4.6605134,3.9712822,3.436308,3.1245131,2.9604106,2.6978464,2.865231,3.2131286,3.2951798,3.0654361,2.9144619,2.6322052,2.5009232,2.15959,1.6738462,1.5392822,1.8051283,2.4713848,3.05559,3.3017437,3.18359,2.605949,2.1267693,1.8773335,1.8445129,1.8609232,1.5983591,1.5360001,1.463795,1.3883078,1.5556924,1.8707694,1.8838975,1.847795,1.8313848,1.7296412,1.467077,1.276718,1.1815386,1.2635899,1.6738462,1.8018463,1.8740515,1.9659488,2.0808206,2.156308,2.300718,2.484513,2.5895386,2.6584618,2.9046156,3.1638978,3.1442053,3.3641028,3.876103,4.263385,4.1682053,4.2535386,4.529231,4.8836927,5.0871797,4.667077,4.6145644,4.969026,5.097026,3.6693337,3.6496413,3.639795,3.692308,3.8531284,4.138667,4.2994876,5.0477953,5.8847184,6.7610264,8.064001,9.386667,9.964309,9.714872,8.861539,7.9163084,2.7634873,3.2262566,3.239385,3.1671798,3.2918978,3.8301542,3.879385,4.322462,4.850872,5.3103595,5.677949,5.7731285,5.7534366,5.917539,6.2063594,6.196513,6.9776416,7.017026,7.0465646,7.5881033,8.940309,9.124104,9.416205,9.668923,9.895386,10.28595,10.735591,10.299078,9.9282055,9.8363085,9.504821,10.420513,10.843898,11.697231,13.285745,15.287796,17.657436,20.545643,23.341951,26.436926,31.235285,40.316723,52.66708,67.521645,82.44842,93.338264,83.02277,62.381954,42.02667,27.913849,21.346462,18.17272,16.994463,16.95836,17.155283,16.630156,15.960617,13.676309,11.247591,9.232411,7.27959,5.398975,4.086154,2.9505644,1.9790771,1.5261539,1.5491283,1.719795,1.7099489,1.3850257,0.82379496,0.65312827,0.5546667,0.5973334,0.702359,0.64000005,0.5907693,0.45292312,0.2986667,0.16410258,0.029538464,0.029538464,0.013128206,0.013128206,0.032820515,0.04594872,0.032820515,0.24943592,0.41025645,0.35446155,0.06235898,0.18379489,0.37743592,0.45292312,0.52512825,1.0371283,1.4276924,1.4145643,1.4703591,1.4966155,0.82379496,0.82379496,0.5415385,0.27241027,0.14112821,0.09189744,0.24943592,0.45620516,0.9616411,1.394872,0.74830776,1.2964103,1.5622566,3.1540515,5.5991797,6.3310776,4.6605134,2.7766156,2.7044106,3.826872,2.8980515,1.6771283,2.6190772,3.5413337,3.767795,4.135385,3.9384618,2.930872,2.8258464,3.8137438,4.5456414,2.9243078,2.7634873,2.9965131,3.3050258,4.135385,3.5971284,4.342154,5.2512827,5.543385,4.775385,4.6900516,5.940513,7.325539,8.55959,10.269539,9.892103,10.023385,11.332924,12.760616,11.54954,11.063796,11.050668,10.71918,10.039796,9.734565,9.15036,10.502565,11.936821,12.704822,13.167591,10.752001,10.742155,11.864616,13.00677,13.213539,13.505642,13.039591,13.02318,13.403898,12.87877,12.596514,11.411694,10.640411,10.906258,12.114052,12.652308,12.0549755,12.153437,12.806565,11.900719,11.487181,10.768411,10.292514,10.354873,11.001437,11.113027,11.349334,11.995898,12.62277,12.084514,11.047385,10.148104,9.554052,9.403078,9.780514,10.026668,10.095591,9.6754875,8.917334,8.454565,8.612103,9.009232,9.202872,9.238976,9.6295395,9.724719,8.769642,7.8670774,7.466667,7.3714876,7.2960005,7.0859494,7.4469748,8.474257,9.659078,9.084719,8.795898,9.196308,9.947898,9.947898,9.813334,10.328616,11.441232,12.727796,13.413745,13.338258,12.754052,12.35036,12.826258,14.87754,13.620514,12.967385,13.4170265,14.329437,13.899488,13.99795,14.78236,15.461744,15.622565,15.24513,14.244103,14.313026,15.087591,16.160822,17.073233,16.928822,17.056822,17.135592,16.928822,16.282257,14.549335,15.497848,17.23077,18.793028,20.171488,20.378258,19.899078,19.088411,17.716515,14.969437,14.907078,13.722258,12.914873,12.924719,13.108514,12.888617,12.182976,11.290257,10.443488,9.796924,10.161232,9.649232,9.301334,9.317744,9.048616,9.892103,10.450052,9.3078985,7.3747697,7.890052,8.6580515,9.015796,9.449026,9.711591,8.818872,4.9394875,4.854154,6.370462,7.259898,5.293949,4.8804107,4.9952826,4.2371287,2.3762052,0.3511795,0.26584616,0.30851284,0.7122052,2.3926156,6.957949,9.278359,9.875693,9.278359,8.43159,8.713847,7.381334,9.255385,11.667693,12.471796,10.056206,7.4929237,5.1659493,3.8596926,3.255795,1.9364104,2.2055387,2.612513,2.9965131,2.8816411,1.463795,1.5983591,1.1848207,1.0371283,1.7001027,3.4330258,3.7874875,4.0402055,3.3641028,2.3696413,3.1113849,2.5862565,3.636513,6.196513,9.586872,12.527591,8.303591,3.9253337,2.2514873,3.0818465,3.1442053,4.850872,6.2030773,7.0531287,7.2894363,6.8496413,6.5936418,5.979898,5.290667,4.6178465,3.8596926,2.1267693,2.4451284,3.3608208,3.9876926,4.013949,4.8804107,5.4547696,7.2664623,8.54318,4.197744,6.4557953,9.353847,10.660104,10.272821,10.223591,9.882257,9.347282,9.419488,9.95118,9.842873,9.107693,9.849437,10.883283,11.250873,10.236719,10.545232,9.173334,7.4141545,6.3934364,7.066257,7.762052,5.5532312,2.9407182,1.6640002,2.7011285,2.674872,4.309334,5.481026,5.037949,2.793026,0.764718,0.10502565,0.006564103,0.04266667,0.15097436,0.15097436,0.26256412,0.256,0.13128206,0.108307704,0.118153855,0.08533334,0.06235898,0.07548718,0.13784617,0.19692309,0.27897438,0.40697438,0.4660513,0.19692309,0.3314872,0.38400003,0.54482055,0.73517954,0.6268718,0.41682056,0.4135385,0.4135385,0.36758977,0.36758977,0.49887183,0.52512825,0.58092314,0.74830776,1.0535386,2.103795,2.3827693,2.3893335,2.4582565,2.7602053,2.9440002,3.629949,4.8640003,6.5017443,8.224821,7.7981544,8.021334,7.2336416,5.6943593,5.586052,5.976616,4.9362054,4.529231,4.97559,4.670359,4.962462,7.003898,8.119796,7.90318,8.208411,8.684308,8.805744,8.585847,7.837539,6.163693,6.665847,6.99077,7.1089234,7.056411,6.957949,7.496206,7.4371285,7.3025646,7.456821,8.116513,8.690872,8.861539,8.960001,9.048616,8.92718,8.779488,8.513641,8.4283085,8.333129,7.5520005,7.1515903,7.7718983,8.408616,8.681026,8.864821,8.694155,8.661334,8.484103,8.2445135,8.392206,7.5388722,6.820103,6.9054365,7.680001,8.254359,7.765334,6.957949,6.3310776,6.170257,6.560821,5.7796926,5.7403083,6.0685134,6.5444107,7.0957956,7.069539,7.24677,7.6570263,8.050873,7.90318,5.865026,5.402257,5.5729237,5.7403083,5.5696416,4.7392826,5.986462,7.000616,6.5378466,4.4242053,2.7536411,1.1979488,0.49230772,0.5284103,0.380718,0.67610264,0.90256417,1.1224617,1.2800001,1.204513,1.339077,1.2898463,0.92553854,0.5513847,0.9321026,1.3226668,1.401436,1.8576412,2.6256413,2.868513,2.2088206,2.6387694,3.3476925,3.9253337,4.3651285,3.6562054,3.498667,3.2032824,2.4713848,1.3718976,1.2406155,1.1126155,1.2898463,1.5491283,1.1585642,1.2209232,1.3554872,1.6246156,2.1103592,2.9144619,3.6594875,4.1550775,4.332308,4.269949,4.197744,3.7316926,3.5052311,3.6660516,4.06318,4.2568207,4.342154,4.309334,4.125539,3.7710772,3.2361028,2.7470772,2.5042052,2.6223593,3.117949,3.9384618,4.4242053,4.673641,4.5587697,4.2436924,4.197744,4.3290257,4.1714873,4.1550775,4.125539,3.3575387,3.626667,4.0303593,4.6178465,5.228308,5.5072823,5.0215387,5.6385646,6.633026,7.4141545,7.522462,8.720411,8.661334,8.192,7.5585647,6.422975,6.705231,7.141744,7.6964107,8.205129,8.375795,6.7183595,6.009436,5.7042055,5.6418467,6.058667,6.8988724,7.072821,7.4108725,7.817847,7.2927184,7.0137444,6.8496413,6.4000006,5.477744,4.135385,3.3772311,3.6004105,3.6135387,3.2098465,3.1737437,3.370667,3.4625645,3.4198978,3.18359,2.6715899,2.487795,2.166154,1.8937438,1.7099489,1.5261539,1.782154,2.2482052,2.674872,2.8291285,2.487795,2.231795,2.1858463,2.1431797,2.0578463,2.044718,1.6049232,1.3751796,1.6640002,2.1924105,2.1070771,2.2153847,2.281026,2.097231,1.7788719,1.7558975,1.5097437,1.5688206,1.5261539,1.3193847,1.2209232,1.4769232,1.7788719,1.9692309,2.0217438,2.0611284,2.097231,2.3335385,2.609231,2.8914874,3.2951798,3.2229745,3.259077,3.6004105,4.164923,4.59159,4.70318,4.6211286,4.5029745,4.562052,5.0510774,4.6112823,4.5390773,4.709744,4.890257,4.7294364,4.4373336,4.1911798,4.391385,4.821334,4.637539,4.857436,5.225026,5.9503593,6.951385,7.8441033,9.380103,9.537642,9.005949,8.503796,8.759795,2.8717952,2.9833848,3.0293336,3.1343591,3.3608208,3.6824617,3.8498464,4.086154,4.4865646,5.041231,5.651693,5.7796926,5.786257,5.835488,5.989744,6.232616,7.3353853,7.250052,7.0367184,7.3321033,8.356103,8.743385,9.278359,9.724719,9.93477,9.856001,9.898667,9.7903595,9.672206,9.527796,9.189744,10.036513,10.886565,12.156719,14.017642,16.400412,19.226257,20.795078,22.42954,25.442463,31.136824,40.56944,52.68021,64.095184,72.16247,74.95549,62.336006,45.696003,31.950771,23.634052,18.894772,16.295385,15.153232,15.287796,15.911386,15.632411,15.0088215,13.505642,11.83836,10.28595,8.694155,6.5805135,5.3858466,4.2436924,2.917744,1.782154,1.3784616,1.2996924,1.3292309,1.2438976,0.8467693,0.75487185,0.67610264,0.60389745,0.5907693,0.77456415,0.6662565,0.51856416,0.39712822,0.27241027,0.029538464,0.01969231,0.006564103,0.032820515,0.108307704,0.2297436,0.57764107,0.9419488,0.92225647,0.53825647,0.24287182,0.4135385,0.446359,0.41682056,0.54482055,1.1848207,1.8084104,1.8412309,1.7493335,1.6147693,1.1290257,1.3620514,0.77128214,0.26584616,0.14112821,0.09189744,0.190359,0.24943592,0.5316923,0.82379496,0.42994875,0.8336411,1.142154,1.5360001,2.0512822,2.609231,2.5304618,2.6486156,2.4484105,2.0676925,2.3138463,2.6256413,3.9417439,4.322462,3.6430771,3.6102567,3.0162053,3.6562054,4.522667,4.650667,3.117949,3.2623591,3.495385,3.511795,3.2623591,2.9505644,3.2722054,4.6572313,5.6352825,5.586052,4.7392826,5.182359,6.226052,7.824411,9.80677,11.904001,10.735591,11.864616,12.780309,12.704822,12.599796,11.713642,11.18195,9.833026,8.3823595,9.45559,9.15036,10.44677,11.766154,12.727796,14.119386,12.347078,11.34277,12.1468725,13.8765135,13.702565,14.552616,13.843694,12.872206,12.150155,11.388719,10.794667,10.725744,10.925949,11.201642,11.395283,11.286975,11.877745,12.832822,13.666463,13.718975,12.747488,12.032001,11.378873,10.663385,9.816616,10.482873,11.657847,12.960821,13.824001,13.512206,11.703795,11.027693,10.499283,9.921641,9.892103,9.90195,9.537642,9.40636,9.4457445,8.940309,8.661334,8.897642,9.298052,9.6525135,9.895386,9.38995,8.707283,8.103385,7.781744,7.9195905,7.778462,7.5585647,7.6110773,8.073847,8.87795,9.025641,8.507077,8.874667,10.092308,10.522257,10.699488,10.994873,11.58236,12.3536415,12.898462,12.49477,11.920411,11.575796,11.772718,12.727796,12.750771,12.973949,13.328411,13.761642,14.244103,14.408206,15.314053,15.412514,14.539488,13.8765135,13.656616,13.774771,14.024206,14.49354,15.586463,15.691488,15.855591,15.881847,15.826053,16.000002,15.750566,16.866463,17.91672,18.582975,19.659489,20.864002,21.028105,20.128822,18.454975,16.617027,15.881847,13.735386,11.762873,10.722463,10.545232,11.136001,11.401847,11.1983595,10.581334,9.80677,9.803488,9.645949,10.102155,10.679795,9.609847,10.55836,12.22236,10.971898,7.955693,9.084719,9.481847,11.378873,12.2387705,11.437949,10.28595,6.7938466,6.7938466,7.2172313,6.180103,2.9768207,3.3214362,2.7273848,2.425436,2.3696413,1.2406155,0.5316923,0.30851284,0.45292312,1.5491283,4.893539,4.890257,5.6976414,7.9327188,9.432616,5.2709746,4.516103,7.397744,12.842668,17.138874,13.961847,9.4457445,6.5805135,4.667077,3.3017437,2.3663592,5.0051284,5.287385,5.0084105,4.5489235,2.868513,3.7152824,3.2722054,2.5600002,2.3401027,3.114667,5.481026,5.139693,4.066462,3.511795,4.0041027,4.132103,6.685539,10.226872,13.3940525,14.920206,12.511181,9.386667,6.7807183,5.106872,3.948308,4.4373336,3.8498464,3.5282054,4.0434875,5.21518,6.892308,7.75877,8.224821,7.955693,5.8486156,3.4330258,2.3269746,2.228513,2.6847181,3.1113849,4.269949,5.4941545,6.62318,6.564103,3.2918978,5.0838976,7.9458466,10.473026,11.674257,10.981745,9.202872,7.958975,7.686565,8.218257,8.792616,8.461129,9.324308,10.134975,10.535385,11.044104,11.027693,10.469745,9.078155,7.1909747,5.7829747,6.488616,5.674667,4.082872,2.986667,4.1911798,4.4307694,3.879385,3.757949,3.511795,0.81394875,0.20348719,0.01969231,0.026256412,0.072205134,0.10502565,0.06564103,0.098461546,0.118153855,0.08861539,0.04594872,0.07876924,0.072205134,0.055794876,0.055794876,0.08861539,0.16082053,0.23302566,0.28225642,0.27241027,0.15097436,0.23630771,0.3052308,0.48246157,0.71548724,0.77128214,0.61374366,0.6695385,0.67610264,0.5349744,0.32820517,0.43323082,0.45292312,0.5349744,0.71548724,0.892718,1.6804104,1.8740515,2.1267693,2.6322052,3.1048207,3.0818465,3.1671798,4.269949,6.189949,7.637334,7.056411,8.228104,7.712821,5.612308,5.5597954,5.47118,5.1200004,5.4186673,6.091488,5.671385,6.4623594,7.4404106,7.9852314,8.096821,8.392206,8.576,8.6580515,8.257642,7.387898,6.4590774,6.4590774,6.8463597,7.1023593,7.0465646,6.810257,7.0859494,7.318975,7.529026,7.8112826,8.362667,8.572719,9.570462,10.043077,9.53436,8.425026,8.953437,8.950154,8.474257,7.939283,8.113232,7.496206,7.276308,7.207385,7.2927184,7.778462,8.536616,8.881231,9.133949,9.242257,8.78277,7.899898,7.312411,7.1844106,7.3485136,7.328821,7.1909747,6.7840004,6.340924,6.0849237,6.232616,6.4557953,6.9021544,7.026872,6.7085133,6.2523084,6.5805135,7.0432825,7.1089234,6.626462,5.8157954,4.5587697,4.5456414,5.425231,6.5050263,6.7544622,6.9087186,7.4896417,6.928411,5.221744,3.8990772,1.6508719,0.61374366,0.31507695,0.35774362,0.40697438,0.6892308,0.7253334,0.8172308,1.0404103,1.2406155,1.1815386,1.2209232,1.2603078,1.2668719,1.2832822,1.4211283,1.5458462,2.038154,2.6453335,2.4910772,2.0250258,2.1825643,2.6322052,3.1540515,3.6332312,3.0030773,3.249231,3.4264617,2.9669745,1.7033848,1.4605129,1.273436,1.142154,1.0732309,1.0732309,1.1355898,1.2996924,1.723077,2.3860514,3.0720003,3.3476925,3.186872,3.2525132,3.5872824,3.6102567,3.5872824,3.5807183,3.7349746,4.059898,4.4406157,4.338872,4.2305646,3.9351797,3.4625645,3.0030773,2.612513,2.8192823,3.186872,3.5840003,4.204308,4.263385,4.266667,4.1747694,4.06318,4.1222568,4.5029745,4.578462,4.667077,4.6244106,3.8465643,3.636513,3.6791797,4.020513,4.630975,5.398975,4.9887185,5.540103,6.4656415,7.194257,7.1548724,7.9819493,8.5202055,8.533334,7.9097443,6.6560006,6.6625648,7.2861543,7.6570263,7.7456417,8.375795,8.034462,7.3353853,6.669129,6.301539,6.373744,6.9645133,7.273026,7.778462,8.369231,8.342975,7.9163084,7.6143594,6.994052,6.0652313,5.3070774,3.9745643,3.6430771,3.6758976,3.7021542,3.626667,4.007385,3.7152824,3.6627696,3.876103,3.498667,2.7700515,2.2482052,1.9035898,1.7624617,1.8904617,2.2646155,2.5632823,2.8389745,2.9636924,2.6223593,2.2777438,2.034872,1.9232821,1.8149745,1.4211283,1.1191796,1.1651284,1.4539489,1.8084104,1.9954873,2.3991797,2.5731285,2.231795,1.657436,1.6804104,1.5163078,1.5556924,1.5524104,1.4408206,1.3423591,1.5885129,1.8084104,1.9232821,1.975795,2.1202054,2.166154,2.4155898,2.7175386,2.9965131,3.2361028,3.1803079,3.515077,4.141949,4.8311796,5.228308,4.9362054,4.7458467,4.788513,5.0051284,5.172513,5.221744,5.3366156,5.35959,5.156103,4.6080003,4.5489235,4.309334,4.516103,4.9887185,4.7360005,5.034667,5.2512827,6.012718,7.1647186,7.781744,8.694155,9.176616,9.173334,8.605539,7.3682055,2.6715899,2.7306669,2.865231,3.0884104,3.3903592,3.7021542,3.82359,3.9975388,4.2502565,4.640821,5.2611284,5.609026,5.858462,5.9536414,5.943795,5.98318,6.9349747,7.4404106,7.6570263,7.8080006,8.192,8.329846,8.822155,9.301334,9.43918,8.937026,9.042052,9.061745,8.979693,8.904206,9.045334,10.006975,10.587898,12.018872,14.401642,16.695797,19.616821,20.755693,22.048822,25.189745,31.64226,38.081642,48.31508,54.833237,54.908722,50.60267,41.32431,31.944208,24.116514,18.369642,14.076719,11.017847,9.554052,9.068309,8.854975,8.129642,8.024616,7.6143594,7.02359,6.2752824,5.293949,4.0369234,3.5183592,2.9078977,2.0184617,1.2964103,0.9747693,0.764718,0.69579494,0.69907695,0.6071795,0.6235898,0.5481026,0.49230772,0.5481026,0.8008206,0.69251287,0.57764107,0.4201026,0.21989745,0.029538464,0.1148718,0.13128206,0.15753847,0.25928208,0.4955898,0.83035904,1.0666667,0.8598975,0.3511795,0.16082053,0.22646156,0.2100513,0.18707694,0.32820517,0.9288206,1.7296412,1.8445129,1.8642052,1.9856411,2.028308,1.8018463,0.9485129,0.3511795,0.25271797,0.24615386,0.30194873,0.2855385,0.3511795,0.446359,0.27897438,0.41025645,0.8467693,0.8566154,0.5513847,0.88287187,1.0305642,1.4276924,1.8445129,2.172718,2.422154,2.7076926,3.495385,3.5216413,2.8750772,2.9669745,3.1277952,4.2338467,5.0477953,4.84759,3.4198978,3.7448208,3.9975388,3.8104618,3.43959,3.761231,4.2272825,4.9887185,5.172513,5.0215387,5.910975,6.4623594,7.8802056,9.38995,10.633847,11.680821,12.064821,13.282462,13.545027,12.941129,13.449847,12.511181,12.458668,11.273847,9.363693,9.547488,9.110975,10.541949,12.209231,13.449847,14.55918,14.332719,13.37436,13.797745,14.897232,13.157744,13.308719,12.425847,11.52,11.057232,10.935796,10.400822,10.423796,10.824206,11.132719,10.601027,10.377847,10.774975,11.664412,12.770463,13.66318,13.88636,12.576821,11.290257,10.604308,10.144821,11.008,12.432411,13.367796,13.581129,13.6697445,11.680821,11.785847,11.785847,11.001437,10.276103,9.750975,9.31118,9.304616,9.494975,9.055181,8.736821,8.474257,8.579283,8.887795,8.726975,8.260923,8.264206,7.9195905,7.273026,7.2336416,7.506052,7.39118,7.463385,7.79159,7.9491286,8.316719,8.041026,8.474257,9.622975,10.154668,10.210463,10.171078,10.643693,11.552821,12.140308,11.382154,10.604308,10.374565,10.840616,11.74318,12.245335,13.010053,13.410462,13.61395,14.549335,14.424617,14.818462,14.815181,14.116103,13.039591,13.124924,13.722258,14.194873,14.395078,14.674052,14.227694,14.355694,14.562463,14.880821,15.8654375,16.242872,17.900309,19.055592,19.364103,19.895796,20.41108,20.22072,19.085129,17.591797,17.138874,16.610462,13.656616,10.880001,9.465437,9.199591,10.174359,10.791386,10.774975,10.167795,9.32759,9.777231,9.757539,10.394258,11.497026,11.552821,12.186257,13.088821,12.012309,9.892103,10.8307705,11.648001,12.544001,12.294565,11.890873,14.523078,12.3536415,9.284924,8.553026,9.114257,5.671385,3.501949,2.7142565,2.1234872,1.4506668,1.3456411,0.8172308,0.39712822,0.24615386,0.6498462,2.0250258,1.8937438,2.605949,6.51159,10.8996935,8.008205,6.114462,7.5881033,12.33395,17.880617,19.396925,12.987078,8.546462,5.362872,3.4067695,3.3411283,3.9187696,4.634257,5.179077,5.280821,4.7294364,4.699898,3.9548721,3.1573336,3.0326157,4.391385,6.5345645,5.756718,4.076308,2.9833848,3.43959,4.017231,9.189744,13.5089245,14.880821,14.565744,13.968411,10.906258,7.6274877,5.435077,4.6802053,4.6080003,3.8695388,3.2262566,3.0293336,3.2032824,5.2348723,6.419693,7.9294367,9.009232,6.9710774,4.273231,2.8553848,2.225231,2.0808206,2.297436,2.7995899,4.900103,7.276308,8.349539,6.298257,6.088206,7.7948723,9.892103,10.866873,9.229129,7.069539,5.720616,4.9493337,4.8147697,5.6451287,6.235898,7.0531287,7.6110773,7.8539495,8.15918,9.009232,9.95118,9.334154,7.0465646,4.5095387,4.634257,4.9493337,5.21518,5.297231,5.2020516,4.7261543,3.9778464,3.3805132,2.5271797,0.17394873,0.04266667,0.009846155,0.016410258,0.032820515,0.036102567,0.032820515,0.029538464,0.036102567,0.03938462,0.02297436,0.04266667,0.055794876,0.055794876,0.052512825,0.07548718,0.15097436,0.24943592,0.27241027,0.21333335,0.16410258,0.19364104,0.27241027,0.45620516,0.67938465,0.75487185,0.6892308,0.77128214,0.761436,0.5907693,0.35774362,0.43323082,0.51856416,0.5940513,0.6465641,0.6892308,1.394872,1.7099489,2.281026,3.0194874,3.114667,2.8160002,2.8324106,3.820308,5.5007186,6.669129,6.6592827,7.171283,7.059693,6.232616,5.609026,5.3727183,5.8125134,6.245744,6.235898,5.5630774,6.8955903,7.4174366,7.6274877,7.830975,8.155898,8.52677,8.776206,8.41518,7.4075904,6.163693,6.554257,7.145026,7.463385,7.453539,7.4699492,7.6570263,7.7292314,7.762052,7.8670774,8.201847,8.369231,9.383386,10.105436,9.849437,8.392206,8.736821,8.900924,8.4972315,7.8802056,8.12636,7.456821,7.125334,7.0859494,7.387898,8.185436,8.661334,9.229129,9.527796,9.268514,8.241231,8.43159,8.326565,7.9983597,7.571693,7.2237954,6.954667,7.072821,6.8233852,6.242462,6.166975,6.3934364,6.6625648,6.626462,6.3212314,6.160411,6.8332314,6.8529234,6.0291286,4.7950773,4.2141542,3.1967182,3.5052311,4.6966157,6.0225644,6.426257,8.067283,7.712821,6.229334,4.466872,3.245949,1.529436,0.7318975,0.4004103,0.36102566,0.7220513,0.7187693,0.69579494,0.83035904,1.0994873,1.2865642,1.2077949,1.1848207,1.1979488,1.2176411,1.2176411,1.2898463,1.6246156,1.9659488,2.1103592,1.9200002,1.847795,1.8871796,2.1234872,2.537026,2.9735386,2.9833848,3.259077,3.3772311,2.9735386,1.7493335,1.4867693,1.3620514,1.1520001,0.90256417,0.9419488,1.0699488,1.2471796,1.7952822,2.6223593,3.2328207,3.1113849,3.006359,3.249231,3.6758976,3.629949,3.5807183,3.5478978,3.5971284,3.8334363,4.384821,4.1222568,3.9811285,3.698872,3.2754874,2.989949,2.7634873,3.0096412,3.3444104,3.6562054,4.089436,4.056616,4.1058464,4.1813335,4.2469745,4.2962055,4.5456414,4.827898,4.9132314,4.6802053,4.1058464,3.8564105,3.820308,4.0041027,4.44718,5.21518,5.0871797,5.6287184,6.482052,7.1680007,7.066257,7.7390776,8.224821,8.474257,8.372514,7.719385,7.5487185,7.6274877,7.6931286,7.7981544,8.323282,8.339693,8.004924,7.509334,7.030154,6.747898,7.565129,8.1066675,8.585847,8.956718,8.907488,8.533334,8.316719,7.574975,6.377026,5.5532312,4.818052,3.8137438,3.4527183,3.8006158,4.066462,4.4865646,4.069744,3.8038976,3.9548721,4.082872,3.3772311,2.7011285,2.294154,2.172718,2.1300514,2.4385643,2.7733335,2.993231,2.9965131,2.7175386,2.484513,2.1858463,1.9396925,1.6869745,1.1848207,1.0535386,1.1881026,1.3981539,1.5753847,1.6836925,2.0578463,2.162872,1.9364104,1.5622566,1.4539489,1.6049232,1.6344616,1.4802053,1.3095386,1.5195899,1.7624617,1.9528207,1.9823592,1.9331284,2.044718,2.15959,2.5632823,3.1277952,3.5840003,3.5216413,3.5183592,3.9581542,4.519385,4.9460516,5.0674877,4.903385,4.972308,5.152821,5.284103,5.1954875,5.5696416,5.6451287,5.467898,5.1889234,5.0543594,4.6211286,4.3585644,4.585026,5.10359,5.1987696,5.467898,5.979898,6.87918,7.6242056,6.987488,7.77518,8.996103,9.179898,8.27077,7.604513,2.425436,2.5271797,2.6945643,3.0326157,3.4494362,3.6594875,3.948308,4.135385,4.2535386,4.417641,4.827898,5.156103,5.4449234,5.609026,5.6254363,5.5138464,6.2162056,7.0990777,7.765334,7.9983597,7.752206,7.6176414,7.9195905,8.316719,8.553026,8.457847,8.474257,8.3593855,8.257642,8.375795,8.973129,9.888822,10.706052,12.484924,15.136822,17.417847,19.633232,20.978874,22.403284,25.232412,31.17949,34.454975,41.078156,42.89641,37.933952,30.395079,25.544207,21.56636,17.460514,13.298873,10.20718,7.3485136,5.5762057,4.4964104,3.7218463,2.8816411,2.930872,2.9013336,2.8160002,2.6190772,2.176,1.7099489,1.585231,1.401436,1.083077,0.8992821,0.7089231,0.5218462,0.39384618,0.3511795,0.38728207,0.43651286,0.4201026,0.4004103,0.42994875,0.54482055,0.508718,0.4594872,0.32164106,0.13456412,0.04266667,0.12471796,0.16410258,0.23958977,0.40697438,0.6892308,0.90912825,0.95835906,0.65641034,0.19364104,0.0951795,0.072205134,0.04266667,0.03938462,0.15753847,0.52512825,1.1388719,1.3915899,1.6935385,2.1202054,2.4155898,1.585231,0.88287187,0.52512825,0.4955898,0.5349744,0.51856416,0.44307697,0.3708718,0.2986667,0.15425642,0.15425642,0.47917953,0.45292312,0.12143591,0.23958977,0.27897438,0.56451285,1.5458462,2.7602053,2.8553848,2.6912823,3.1376412,3.170462,2.865231,3.4067695,3.6758976,4.5095387,5.077334,4.896821,3.8432825,3.8629746,3.8006158,3.7251284,3.9876926,5.221744,5.149539,5.914257,6.232616,6.3212314,7.9261546,8.218257,9.590155,10.627283,10.94236,11.162257,12.137027,12.895181,12.832822,12.297847,12.599796,11.785847,12.11077,11.920411,10.866873,9.915077,9.31118,10.978462,12.911591,14.086565,14.480412,14.634667,14.14236,14.060308,13.929027,11.766154,11.674257,11.428103,11.076924,10.932513,11.556104,11.18195,10.742155,10.912822,11.372309,10.807796,10.6469755,10.564924,11.329642,12.819694,14.017642,14.63795,12.908309,11.208206,10.630565,10.985026,12.11077,13.190565,13.397334,12.849232,12.642463,11.237744,12.07795,12.803283,12.393026,11.172104,9.911796,9.314463,9.199591,9.212719,8.848411,8.809027,8.03118,7.653744,7.8112826,7.640616,7.4699492,7.778462,7.581539,6.925129,6.892308,7.076103,7.0137444,7.2960005,7.781744,7.578257,7.637334,7.3386674,7.6012316,8.444718,8.963283,8.740103,8.87795,9.521232,10.469745,11.195078,10.381129,9.6,9.649232,10.463181,11.109744,11.930258,12.786873,13.026463,12.980514,13.98154,13.778052,13.558155,13.51877,13.449847,12.704822,13.302155,14.155488,14.513232,14.227694,13.768207,13.111795,13.236514,13.696001,14.457437,15.908104,16.400412,17.897026,19.104822,19.488823,19.26236,18.724104,18.770052,17.870771,16.41354,16.73518,16.210052,13.157744,10.315488,8.887795,8.52677,9.478565,10.049642,10.056206,9.613129,9.107693,9.5835905,9.8592825,10.509129,11.762873,13.505642,13.856822,13.604104,12.786873,11.940104,12.081232,11.831796,11.45436,10.486155,10.571488,15.465027,15.100719,10.617436,9.596719,12.1698475,11.0145645,4.8311796,2.7569232,2.4976413,2.3335385,1.1027694,0.892718,0.48902568,0.256,0.28882053,0.4201026,0.48574364,1.5327181,5.5893335,10.601027,10.443488,7.0859494,6.5969234,9.137232,13.505642,17.115898,13.302155,9.330873,5.943795,3.8531284,3.761231,2.7273848,3.6660516,4.6211286,5.024821,5.6943593,5.924103,4.785231,3.82359,3.82359,4.8082056,6.633026,6.47877,5.175795,3.7710772,3.5478978,3.8990772,8.667898,12.839386,14.007796,12.393026,10.985026,8.569437,6.193231,4.6080003,4.2469745,4.164923,4.2830772,4.0500517,3.436308,2.917744,4.4340515,5.280821,6.987488,8.51036,6.2063594,4.1156926,3.190154,3.045744,3.18359,2.9768207,2.7437952,4.59159,7.030154,8.500513,7.3682055,6.048821,6.3442054,7.9425645,9.186462,7.0498466,6.87918,5.684513,4.4110775,3.8006158,4.388103,5.543385,6.186667,6.413129,6.2096415,5.4514875,6.626462,8.188719,8.093539,6.042257,3.4592824,3.0162053,4.352,6.157129,6.8988724,4.8311796,5.0510774,4.348718,2.9735386,1.339077,0.04594872,0.016410258,0.009846155,0.006564103,0.0032820515,0.013128206,0.016410258,0.009846155,0.013128206,0.02297436,0.02297436,0.02297436,0.04266667,0.049230773,0.04594872,0.068923086,0.118153855,0.2231795,0.25928208,0.21661541,0.20020515,0.20020515,0.27241027,0.41682056,0.5874872,0.69907695,0.7417436,0.78769237,0.7581539,0.636718,0.4660513,0.48902568,0.5481026,0.5677949,0.5677949,0.67282057,1.3784616,2.15959,2.809436,3.062154,2.6223593,2.5993848,2.934154,3.764513,4.84759,5.5696416,6.436103,6.442667,6.485334,6.685539,6.3967185,5.7698464,6.373744,6.774154,6.409847,5.5893335,6.2129235,6.518154,6.744616,7.0498466,7.5191803,7.830975,7.8539495,7.680001,7.325539,6.75118,7.0334363,7.273026,7.581539,8.027898,8.631796,8.487385,8.4053335,8.329846,8.198565,7.9294367,8.070564,8.493949,8.979693,9.065026,8.0377445,8.129642,8.5202055,8.388924,7.785026,7.643898,7.24677,7.13518,7.243488,7.6143594,8.411898,8.720411,9.3768215,9.573745,9.065026,8.185436,8.79918,8.720411,8.264206,7.7292314,7.4010262,6.8233852,7.200821,7.328821,6.8988724,6.521436,6.626462,6.5280004,6.232616,6.0619493,6.6560006,7.643898,6.7282057,5.2676926,4.1682053,3.879385,2.8127182,3.05559,3.945026,4.84759,5.139693,7.059693,6.688821,5.353026,3.8400004,2.412308,2.3466668,1.214359,0.4955898,0.6301539,1.020718,0.81394875,0.6826667,0.81394875,1.1126155,1.2077949,1.270154,1.2012309,1.2373334,1.3784616,1.4080001,1.4080001,1.6836925,1.8281027,1.7263591,1.5721027,1.6311796,1.6968206,1.8806155,2.2153847,2.6486156,3.0260515,3.170462,3.045744,2.5796926,1.6869745,1.5425643,1.5097437,1.2964103,0.9682052,0.955077,1.1651284,1.4375386,1.9692309,2.6584618,3.1113849,2.917744,2.878359,3.1770258,3.6496413,3.767795,3.7120004,3.6463592,3.5741541,3.6036925,3.945026,3.639795,3.5971284,3.5380516,3.367385,3.1803079,3.18359,3.2689233,3.4166157,3.629949,3.9351797,3.82359,3.7415388,3.8137438,4.096,4.588308,4.7655387,5.024821,5.0182567,4.70318,4.3684106,4.1124105,4.135385,4.266667,4.5390773,5.1856413,5.1987696,5.720616,6.521436,7.171283,7.0334363,7.5388722,8.057437,8.461129,8.592411,8.264206,8.03118,7.755488,7.719385,7.9819493,8.388924,8.490667,8.303591,8.011488,7.7423596,7.571693,8.369231,8.605539,8.832001,9.107693,8.999385,8.661334,8.477539,7.8473854,6.7872825,5.901129,5.805949,4.7261543,4.092718,4.210872,4.2568207,4.637539,4.4340515,4.07959,3.9811285,4.522667,4.1550775,3.4002054,2.8225644,2.5698464,2.3926156,2.740513,2.9013336,2.8980515,2.7667694,2.5796926,2.5435898,2.3958976,2.041436,1.5589745,1.1716924,1.148718,1.339077,1.4867693,1.5392822,1.6607181,1.657436,1.6213335,1.6311796,1.6377437,1.4572309,1.719795,1.7591796,1.5327181,1.2964103,1.5983591,1.9987694,2.2186668,2.1858463,2.0578463,2.2383592,2.4320002,2.6978464,3.2623591,3.8564105,3.7120004,3.564308,3.9712822,4.522667,4.95918,5.175795,5.3037953,5.609026,5.802667,5.805949,5.7435904,6.1046157,6.045539,5.691077,5.293949,5.225026,4.6211286,4.388103,4.6572313,5.211898,5.504,5.7534366,6.5903597,7.4469748,7.719385,6.76759,8.034462,9.366975,9.314463,8.113232,7.6898465,2.300718,2.3729234,2.5009232,2.8947694,3.4067695,3.515077,3.9581542,4.1550775,4.2272825,4.3060517,4.525949,4.5095387,4.594872,4.7556925,4.9329233,5.044513,5.586052,6.373744,7.207385,7.6734366,7.1548724,7.003898,7.0367184,7.194257,7.565129,8.372514,8.024616,7.79159,7.7948723,8.178872,9.097847,9.645949,11.119591,13.266052,15.730873,18.057848,19.511797,21.156105,22.665848,24.697437,28.868925,32.04595,35.28862,34.07754,27.703796,19.291899,16.925539,14.690463,11.969642,9.238976,8.083693,6.2916927,4.588308,3.3641028,2.681436,2.2678976,2.0906668,1.7296412,1.4605129,1.3357949,1.1946667,1.024,0.8763078,0.84348726,0.9485129,1.1257436,0.79425645,0.63343596,0.512,0.38400003,0.31507695,0.30851284,0.3511795,0.33476925,0.24615386,0.15425642,0.21333335,0.2231795,0.17723078,0.10502565,0.08533334,0.06235898,0.13128206,0.29538465,0.5284103,0.77128214,0.9517949,0.8566154,0.5415385,0.18707694,0.12471796,0.08205129,0.03938462,0.03938462,0.09189744,0.17394873,0.36430773,0.6826667,1.1585642,1.6443079,1.8084104,0.8008206,0.56451285,0.5973334,0.64000005,0.69907695,0.5874872,0.4955898,0.4004103,0.26912823,0.03938462,0.068923086,0.098461546,0.101743594,0.07876924,0.068923086,0.10502565,0.47261542,1.6213335,3.0030773,3.0949745,2.7569232,3.4560003,3.8629746,3.8006158,4.2436924,3.9122055,4.2272825,4.601436,4.6112823,4.020513,3.69559,3.6036925,4.07959,5.169231,6.629744,6.1308722,7.8802056,9.18318,9.5146675,10.532104,9.938052,10.453334,10.774975,10.601027,10.620719,10.676514,11.113027,11.300103,11.024411,10.509129,10.020103,10.443488,11.224616,11.588924,10.545232,9.921641,11.431385,13.184001,14.165335,14.214565,13.545027,12.977232,12.22236,11.211488,10.118565,10.768411,11.58236,11.795693,11.71036,12.672001,12.491488,11.595488,11.398565,11.907283,11.72677,11.772718,11.579078,12.393026,14.066873,15.064616,14.8939495,13.223386,11.559385,10.873437,11.59877,13.206975,13.482668,12.931283,12.058257,11.372309,10.742155,11.687386,12.822975,13.141335,12.012309,10.44677,9.468719,9.035488,8.881231,8.5202055,8.78277,7.9294367,7.1844106,7.030154,7.200821,7.145026,7.269744,7.2172313,7.062975,7.318975,6.9677954,6.8463597,7.256616,7.8539495,7.6603084,7.273026,6.688821,6.5903597,7.026872,7.4108725,7.131898,7.762052,8.63836,9.472001,10.33518,9.819899,9.360411,9.642668,10.427077,10.55836,11.572514,12.199386,12.189539,11.98277,12.71795,12.763899,12.225642,11.992617,12.235488,12.389745,13.6467705,14.434463,14.306462,13.525334,13.072412,12.822975,13.082257,13.827283,14.959591,16.292105,16.597334,17.11918,17.874052,18.458258,18.054565,17.138874,17.969233,17.463797,15.724309,16.042667,15.025232,12.370052,9.984001,8.641642,7.9819493,8.67118,9.035488,9.081436,8.979693,9.058462,9.29477,10.04636,10.6469755,11.592206,14.532925,15.107284,14.339283,13.896206,13.938873,13.111795,10.059488,9.642668,9.301334,9.3768215,13.124924,12.914873,9.82318,9.849437,13.35795,15.107284,6.695385,2.5009232,2.8225644,4.529231,1.0601027,0.78769237,0.54482055,0.48902568,0.5513847,0.46276927,0.29210258,1.8937438,4.644103,7.5585647,9.284924,6.6133337,5.0051284,5.356308,7.062975,8.01477,9.009232,7.755488,5.85518,4.3060517,3.5314875,2.7864618,3.498667,4.1058464,4.594872,6.47877,9.780514,9.468719,8.595693,8.264206,7.6209235,7.5487185,7.312411,6.695385,5.6943593,4.5128207,4.414359,6.0028725,8.966565,11.526565,10.427077,6.1341543,4.962462,4.578462,4.0008206,3.6168208,3.3509746,4.325744,4.8377438,4.493129,4.1747694,4.9821544,5.464616,6.4590774,7.0925136,4.7491283,3.761231,3.3017437,3.9614363,5.110154,4.9132314,4.650667,5.2512827,6.229334,6.997334,6.8463597,4.923077,4.076308,5.2053337,6.961231,5.756718,7.9983597,7.1844106,6.114462,5.7534366,5.2545643,6.36718,6.7282057,6.633026,6.0061545,4.378257,4.97559,5.8814363,5.72718,4.4898467,3.4888208,3.1934361,5.0116925,6.7117953,6.5772314,3.4034874,5.3136415,4.4012313,2.1497438,0.13456412,0.0,0.0,0.0,0.0,0.0032820515,0.02297436,0.0032820515,0.009846155,0.02297436,0.029538464,0.029538464,0.01969231,0.029538464,0.036102567,0.036102567,0.059076928,0.072205134,0.15097436,0.21661541,0.23630771,0.2297436,0.2297436,0.27569234,0.34789747,0.45620516,0.636718,0.7778462,0.77456415,0.7253334,0.65969235,0.571077,0.56123084,0.52512825,0.512,0.5940513,0.8598975,1.5721027,2.809436,3.1638978,2.5435898,2.1989746,2.7733335,3.387077,3.9975388,4.4898467,4.6966157,6.2720003,6.488616,6.4295387,6.6592827,7.2270775,6.4065647,6.518154,6.695385,6.4722056,5.792821,4.9788723,5.175795,5.618872,6.0061545,6.488616,6.626462,6.3474874,6.488616,7.1844106,7.890052,7.4436927,7.131898,7.50277,8.493949,9.442462,9.002667,8.887795,8.795898,8.500513,7.860513,7.8408213,7.5618467,7.5454364,7.7292314,7.463385,7.5487185,8.064001,8.152616,7.6012316,6.872616,6.8332314,7.059693,7.2303596,7.4207187,8.086975,8.717129,9.370257,9.403078,8.914052,8.723693,9.045334,8.681026,8.136206,7.6635904,7.259898,6.6527185,7.0859494,7.5946674,7.6143594,6.961231,6.9677954,6.8004107,6.409847,6.23918,7.24677,8.185436,6.6461544,5.074052,4.384821,3.9745643,3.117949,3.6660516,4.1714873,4.1878977,4.3027697,5.346462,5.5105643,4.84759,3.508513,1.7526156,2.937436,1.4408206,0.6859488,1.3751796,1.4966155,1.0108719,0.7318975,0.77456415,1.017436,1.1027694,1.3522053,1.3357949,1.5425643,1.9265642,1.9331284,1.7952822,1.7362052,1.7132308,1.6672822,1.5064616,1.4309745,1.591795,1.8281027,2.100513,2.477949,2.740513,2.8225644,2.5796926,2.097231,1.7001027,1.657436,1.6672822,1.4572309,1.1191796,1.1027694,1.3653334,1.782154,2.1924105,2.5042052,2.6912823,2.7634873,2.7437952,2.986667,3.4789746,3.8301542,3.82359,3.7776413,3.6463592,3.4822567,3.4527183,3.2164104,3.3312824,3.5314875,3.623385,3.4756925,3.623385,3.5216413,3.446154,3.5314875,3.767795,3.7054362,3.3903592,3.3476925,3.8596926,4.9788723,5.1265645,5.225026,5.1265645,4.8804107,4.716308,4.378257,4.450462,4.673641,4.9362054,5.2709746,5.2414365,5.720616,6.498462,7.1515903,7.0334363,7.312411,7.890052,8.310155,8.356103,8.064001,7.9458466,7.7259493,7.7357955,8.034462,8.395488,8.648206,8.438154,8.264206,8.356103,8.67118,9.058462,8.576,8.457847,8.868103,8.884514,8.454565,7.972103,7.5979495,7.253334,6.626462,6.5411286,5.9963083,5.474462,5.0904617,4.588308,4.647385,4.7589746,4.5062566,4.1813335,4.772103,4.788513,4.1846156,3.4330258,2.858667,2.6453335,3.062154,2.8947694,2.5698464,2.349949,2.3072822,2.3860514,2.4976413,2.15959,1.4998976,1.2668719,1.2406155,1.4769232,1.595077,1.585231,1.8149745,1.4178462,1.3029745,1.5130258,1.8182565,1.6935385,1.785436,1.9167181,1.8543591,1.6640002,1.7427694,2.3040001,2.5304618,2.4516926,2.3433847,2.7142565,2.934154,2.9801028,3.3969233,4.0041027,3.892513,3.3903592,3.6463592,4.31918,5.10359,5.720616,6.0258465,6.3442054,6.3868723,6.311385,6.7216415,6.7610264,6.5969234,6.180103,5.622154,5.182359,4.824616,4.59159,4.7392826,5.1889234,5.5138464,6.009436,6.872616,7.4141545,7.39118,7.000616,9.032206,9.8363085,9.511385,8.513641,7.640616,2.349949,2.2153847,2.2908719,2.537026,2.917744,3.4166157,3.186872,3.2656412,3.508513,3.8662567,4.378257,3.95159,3.9286156,3.945026,4.1058464,4.95918,5.421949,6.052103,6.7971287,7.387898,7.3386674,7.5585647,7.2303596,6.875898,6.9054365,7.6143594,7.0531287,7.315693,7.755488,8.36595,9.780514,9.645949,10.794667,12.563693,14.506668,16.374155,18.91118,20.122257,20.98872,22.278566,24.536617,33.972515,38.1079,36.83118,29.935593,17.106052,13.784616,11.142565,8.681026,6.6428723,5.9963083,4.850872,3.9581542,3.0654361,2.3269746,2.3040001,2.3040001,1.9298463,1.4342566,1.0469744,0.9616411,0.8992821,0.86646163,1.024,1.467077,2.2121027,1.2832822,0.81394875,0.636718,0.55794877,0.3511795,0.26584616,0.21661541,0.19364104,0.16738462,0.108307704,0.14441027,0.17066668,0.18379489,0.18379489,0.18379489,0.108307704,0.28225642,0.49887183,0.6629744,0.80738467,1.1126155,0.90584624,0.5152821,0.19692309,0.13784617,0.07548718,0.032820515,0.009846155,0.0032820515,0.016410258,0.08861539,0.14441027,0.20348719,0.2855385,0.380718,0.17394873,0.16738462,0.19692309,0.2100513,0.25928208,0.101743594,0.098461546,0.1148718,0.08861539,0.016410258,0.016410258,0.016410258,0.026256412,0.04594872,0.04594872,0.068923086,0.52512825,1.5458462,2.5928206,2.4713848,2.4976413,3.7382567,4.768821,4.647385,2.9144619,2.9505644,3.062154,2.9505644,3.114667,4.8377438,3.9089234,5.2611284,6.665847,7.3353853,7.936001,8.667898,11.195078,12.383181,12.179693,13.594257,10.9226675,9.980719,9.711591,9.472001,9.032206,8.874667,10.144821,11.047385,10.791386,9.5835905,9.862565,10.8307705,11.221334,11.034257,11.536411,10.998155,11.057232,12.015591,13.495796,14.434463,13.715693,11.254155,9.593436,9.350565,9.216001,10.948924,11.703795,12.068104,12.452104,13.062565,13.292309,12.609642,12.104206,12.009027,11.703795,12.373334,12.642463,13.266052,14.293334,15.074463,14.660924,13.413745,12.002462,11.122872,11.490462,13.712411,12.865642,11.552821,11.113027,11.628308,10.676514,10.502565,10.978462,11.585642,11.414975,11.155693,9.691898,8.868103,8.910769,8.421744,8.507077,8.585847,7.9130263,6.885744,7.020308,6.3967185,6.4590774,6.8562055,7.3419495,7.781744,7.5388722,7.322257,7.3386674,7.4765134,7.2927184,7.1122055,6.7249236,6.482052,6.419693,6.2851286,6.701949,7.0793853,7.9294367,9.153642,10.056206,9.957745,10.006975,9.9282055,9.862565,10.374565,10.8996935,11.32636,11.592206,11.753027,11.946668,12.228924,11.969642,11.323078,10.778257,11.168821,12.425847,13.272616,13.308719,12.977232,13.548308,13.75836,14.395078,15.543797,16.807386,17.319386,17.234053,16.800821,16.544823,16.955078,18.49436,18.6519,19.085129,17.920002,15.849027,16.128002,14.601848,11.88759,9.645949,8.300308,7.020308,7.532308,7.768616,7.8802056,7.9950776,8.241231,9.570462,10.617436,10.866873,11.247591,14.129231,15.924514,15.878566,16.190361,16.820515,15.501129,9.718155,11.218052,12.852514,12.612924,13.627078,8.073847,6.701949,9.07159,12.593232,12.544001,8.4283085,3.4625645,2.481231,4.3290257,1.8773335,0.764718,0.571077,0.79097444,1.0010257,0.8533334,0.39056414,1.5753847,2.044718,2.044718,4.4242053,8.15918,7.2172313,6.193231,5.8518977,3.1442053,2.156308,3.2000003,3.9909747,3.82359,3.5544617,3.006359,3.3641028,4.066462,5.674667,9.872411,19.698874,23.857233,24.523489,23.414156,21.802668,13.147899,7.6898465,5.5302567,5.3792825,4.562052,5.1954875,5.428513,6.6002054,8.986258,11.795693,6.2523084,5.179077,5.5630774,5.8256416,5.8125134,3.8596926,4.4242053,5.35959,5.467898,4.516103,5.041231,5.904411,5.8880005,5.297231,5.979898,5.333334,3.9745643,3.820308,5.0838976,6.2555904,7.3419495,7.312411,7.7390776,9.199591,11.277129,6.0619493,4.5423594,3.8071797,3.5216413,5.8912826,5.7665644,5.83877,6.948103,7.75877,4.7294364,5.5597954,5.546667,5.3760004,5.074052,4.013949,4.1124105,3.8596926,3.0687182,2.937436,6.088206,7.456821,8.208411,6.6461544,3.6102567,2.487795,3.8432825,3.1934361,1.5392822,0.036102567,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.02297436,0.029538464,0.029538464,0.029538464,0.02297436,0.02297436,0.032820515,0.04594872,0.068923086,0.12143591,0.20020515,0.26584616,0.2297436,0.23958977,0.24287182,0.26256412,0.3314872,0.5021539,0.7122052,0.761436,0.67610264,0.5349744,0.47261542,0.571077,0.61374366,0.7220513,0.90912825,1.0666667,1.7394873,2.5665643,2.281026,1.5885129,3.190154,3.56759,3.7087183,4.06318,4.5390773,4.5029745,6.124308,6.5936418,6.5706673,6.38359,6.042257,6.675693,6.294975,5.618872,5.1200004,5.034667,4.388103,4.6933336,5.1265645,5.2545643,5.034667,5.927385,6.488616,7.1122055,7.6570263,7.460103,6.803693,7.131898,7.906462,8.562873,8.513641,8.759795,8.507077,7.9458466,7.604513,8.362667,8.008205,7.7259493,7.7259493,7.8670774,7.6603084,7.830975,7.8637953,7.906462,7.6176414,6.163693,5.920821,6.5903597,6.9645133,7.062975,8.149334,9.002667,9.636104,9.393231,8.615385,8.651488,9.616411,9.718155,8.999385,7.6767187,6.1505647,6.380308,7.1614366,7.5421543,7.240206,6.669129,6.0225644,6.5903597,6.921847,6.770872,7.125334,6.9809237,6.5312824,5.113436,3.131077,2.044718,2.4976413,5.5204105,6.813539,5.914257,6.196513,7.02359,6.3343596,5.35959,4.240411,2.044718,0.9944616,0.5218462,1.4080001,2.9243078,2.8389745,1.3489232,1.0601027,1.0535386,1.0272821,1.2964103,1.5786668,1.6935385,1.9331284,2.2482052,2.2744617,2.028308,1.7657437,1.6082052,1.5425643,1.4342566,1.3981539,1.5819489,1.7624617,1.8445129,1.8313848,1.9298463,2.2547693,2.3040001,2.0545642,1.9692309,1.6508719,1.6082052,1.4178462,1.1126155,1.1749744,1.4178462,1.8379488,2.2022567,2.3630772,2.228513,2.678154,3.2328207,3.7185643,3.9876926,3.892513,3.6102567,3.511795,3.4625645,3.4756925,3.7087183,3.5610259,3.6529233,3.7021542,3.6594875,3.7087183,3.623385,3.4100516,3.2000003,3.121231,3.2820516,3.9384618,3.9318976,4.1025643,4.7327185,5.540103,5.2578464,5.4153852,5.421949,5.179077,5.080616,4.7622566,4.7294364,5.2611284,5.8453336,5.172513,5.172513,5.622154,6.416411,7.1680007,7.2172313,7.387898,7.194257,7.210667,7.5881033,8.024616,8.320001,8.064001,7.824411,7.7981544,7.7981544,8.28718,8.536616,8.644924,8.805744,9.291488,9.32759,8.595693,8.3593855,8.809027,9.078155,8.395488,7.0432825,6.6822567,7.3091288,7.24677,6.3442054,6.23918,6.2129235,6.0652313,6.1046157,5.077334,5.041231,4.8836927,4.466872,4.637539,4.8082056,4.8607183,4.2502565,3.1967182,2.6715899,2.7569232,2.6223593,2.297436,2.038154,2.3204105,2.172718,2.4188719,2.3105643,1.7657437,1.3883078,1.2668719,1.4178462,1.4867693,1.4145643,1.4506668,1.3161026,1.3456411,1.5786668,1.8412309,1.7558975,1.7165129,2.156308,2.5173335,2.5731285,2.425436,2.6945643,2.7175386,2.5928206,2.5796926,3.0654361,3.2000003,3.8104618,4.647385,5.1987696,4.699898,3.7973337,3.7907696,4.4734364,5.4153852,5.9667697,6.11118,6.232616,5.986462,5.8912826,7.3091288,6.954667,6.8496413,6.5805135,6.1341543,5.8912826,5.8157954,5.293949,4.7950773,4.7327185,5.477744,6.882462,7.2336416,7.3058467,7.1581545,6.1341543,8.477539,9.110975,9.373539,9.632821,9.278359,1.8248206,1.8970258,1.9790771,2.1070771,2.28759,2.5140514,2.740513,2.9144619,3.1277952,3.446154,3.892513,4.0500517,4.0533338,4.1714873,4.5128207,5.044513,5.7140517,6.012718,6.166975,6.2884107,6.373744,6.419693,6.294975,6.5903597,7.282872,7.7357955,7.1844106,7.2303596,7.433847,7.8408213,8.963283,9.416205,9.911796,11.1983595,13.656616,17.312822,19.275488,19.367386,20.54236,24.100105,29.686155,33.713234,38.728207,38.18667,29.879797,15.944206,11.588924,8.937026,7.072821,5.786257,5.5696416,4.7458467,3.9351797,3.062154,2.300718,2.0611284,1.8051283,1.5491283,1.276718,1.0502565,1.020718,0.9517949,0.84348726,0.92225647,1.1585642,1.2471796,0.6826667,0.48574364,0.4004103,0.34133336,0.38728207,0.44964105,0.4594872,0.4201026,0.39384618,0.49887183,0.41682056,0.32820517,0.256,0.20020515,0.12143591,0.07876924,0.14112821,0.30194873,0.5021539,0.6498462,0.9747693,0.8172308,0.4660513,0.20348719,0.30851284,0.13128206,0.04266667,0.009846155,0.016410258,0.07548718,0.20676924,0.23958977,0.23302566,0.21661541,0.19692309,0.108307704,0.118153855,0.16738462,0.20676924,0.18707694,0.0951795,0.052512825,0.036102567,0.029538464,0.016410258,0.006564103,0.009846155,0.02297436,0.036102567,0.04594872,0.36430773,2.1858463,3.2689233,3.0326157,2.5698464,3.7842054,3.948308,3.6168208,3.387077,3.879385,3.9154875,4.2436924,3.8859491,3.570872,5.7534366,4.8049235,7.0531287,8.4972315,8.211693,8.349539,10.272821,10.827488,11.523283,12.701539,13.522053,11.904001,10.893129,10.328616,10.364718,11.487181,11.162257,10.9915905,10.962052,10.873437,10.338462,9.7903595,10.886565,11.9171295,12.406155,13.121642,12.507898,12.918155,13.013334,13.059283,14.946463,14.060308,12.3306675,11.493745,11.661129,11.303386,13.584412,14.401642,14.956308,15.327181,14.454155,16.111591,16.246155,15.235283,14.001232,13.99795,13.850258,14.080001,14.345847,14.391796,14.050463,13.206975,12.393026,11.533129,10.902975,11.122872,12.672001,11.644719,10.84718,11.32636,12.347078,11.756309,11.52,11.369026,11.369026,11.900719,11.644719,10.906258,10.197334,9.764103,9.557334,8.851693,8.621949,8.080411,7.3091288,7.240206,6.6067696,6.62318,7.0498466,7.6734366,8.320001,8.914052,8.454565,8.057437,7.90318,7.2205133,6.928411,6.636308,6.439385,6.298257,6.0192823,6.422975,6.813539,8.01477,9.852718,11.16554,10.364718,10.282667,10.427077,10.423796,10.010257,9.498257,9.760821,10.433641,11.23118,11.936821,11.835078,11.664412,11.690667,11.956513,12.281437,13.000206,13.53518,13.328411,12.786873,13.292309,14.427898,15.182771,16.167385,17.188105,17.234053,16.718771,16.384,16.420103,17.201233,19.288616,20.000822,20.627693,19.078566,15.973744,14.614976,13.656616,11.72677,9.915077,8.644924,7.6668725,6.8004107,7.0925136,7.2894363,7.269744,8.03118,9.088,9.964309,10.692924,11.753027,14.057027,16.154257,17.010874,15.753847,13.489232,13.292309,13.718975,13.4629755,13.525334,13.732103,12.721231,8.546462,6.6034875,5.8518977,6.163693,8.333129,7.643898,3.6529233,2.2613335,3.748103,2.7798977,1.5819489,0.8730257,0.73517954,1.024,1.3686155,1.0108719,0.93866676,1.1126155,1.5885129,2.5337439,3.6430771,5.6320004,7.3682055,7.4929237,4.414359,2.993231,2.8750772,3.006359,3.1277952,3.7874875,4.1058464,3.8596926,4.076308,5.21518,7.1876926,12.747488,18.277744,22.281847,24.477541,25.796925,20.109129,13.121642,7.4765134,4.273231,3.0851285,3.1442053,4.388103,5.3398976,6.567385,10.683078,9.078155,7.3616414,7.5421543,8.641642,6.705231,6.012718,5.5007186,5.172513,5.0084105,4.9427695,4.0434875,4.3290257,4.4045134,4.2240005,5.10359,7.2861543,9.196308,9.997129,9.055181,5.9503593,7.125334,6.9776416,7.4699492,8.65477,8.687591,5.720616,5.0609236,5.074052,5.3924108,6.892308,4.2896414,6.764308,8.674462,8.277334,7.719385,8.208411,7.3485136,6.308103,5.353026,3.8432825,5.9503593,5.221744,3.8432825,4.886975,12.314258,8.310155,6.196513,5.930667,6.2129235,4.5128207,3.9154875,2.0808206,0.6465641,0.14441027,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.006564103,0.006564103,0.016410258,0.02297436,0.029538464,0.03938462,0.068923086,0.08533334,0.09189744,0.13128206,0.20676924,0.27897438,0.24943592,0.29538465,0.34789747,0.39056414,0.45620516,0.48574364,0.52512825,0.5546667,0.5677949,0.54482055,0.54482055,0.6826667,0.79097444,0.82379496,0.8369231,1.3718976,2.1267693,2.1234872,1.8084104,3.05559,3.5413337,3.501949,3.5840003,4.020513,4.647385,5.8912826,6.688821,6.803693,6.4000006,6.0783596,6.304821,6.1046157,5.799385,5.5532312,5.3891287,4.926359,4.8311796,4.890257,4.9394875,4.8771286,4.8804107,4.9854364,5.421949,6.1374364,6.7905645,6.738052,7.240206,7.50277,7.3321033,7.1483083,7.860513,7.896616,7.637334,7.4371285,7.6176414,7.8769236,7.896616,7.6668725,7.2861543,6.951385,7.640616,7.817847,7.8080006,7.6242056,6.9809237,6.298257,6.3901544,7.0137444,7.8670774,8.612103,8.694155,9.209436,9.777231,10.079181,9.872411,9.780514,9.468719,8.937026,8.188719,7.197539,7.8703594,7.752206,7.581539,7.512616,7.0957956,6.5083084,6.665847,6.9152827,7.131898,7.762052,8.044309,8.201847,6.6625648,3.945026,2.6420515,3.7087183,4.6769233,4.821334,4.4340515,4.7917953,5.405539,5.211898,4.601436,3.5413337,1.5688206,0.6268718,0.35446155,0.6892308,1.1815386,1.0075898,0.8369231,0.8763078,0.9682052,1.1684103,1.7624617,1.9429746,2.1103592,2.297436,2.4188719,2.2383592,2.0709746,1.7690258,1.522872,1.4309745,1.4966155,1.4473847,1.5721027,1.6672822,1.6705642,1.6475899,1.9396925,1.913436,1.8937438,2.0020514,2.1530259,1.6672822,1.5327181,1.4736412,1.4802053,1.785436,2.0873847,2.4615386,2.5928206,2.422154,2.1300514,2.2482052,2.7766156,3.383795,3.7973337,3.8071797,3.5446157,3.5610259,3.5183592,3.3378465,3.2196925,3.7284105,3.7120004,3.5249233,3.370667,3.2918978,3.2951798,3.242667,3.3476925,3.5872824,3.69559,3.8662567,4.2338467,4.8147697,5.284103,4.9788723,5.284103,5.579488,5.648411,5.467898,5.21518,5.10359,5.290667,5.83877,6.2162056,5.2709746,5.142975,5.927385,6.872616,7.456821,7.387898,7.3353853,7.0892315,6.8693337,7.062975,8.234667,8.457847,8.375795,7.9524107,7.4929237,7.637334,7.50277,7.4043083,7.8441033,8.746667,9.488411,9.301334,9.317744,9.133949,8.625232,7.955693,7.975385,7.276308,7.0137444,7.312411,7.273026,6.62318,6.747898,6.5050263,6.038975,6.8004107,6.8496413,6.5083084,6.1505647,5.7632823,4.955898,5.1856413,5.0182567,4.650667,4.07959,3.0851285,3.0424619,2.8324106,2.3696413,1.8674873,1.8543591,2.1103592,2.3630772,2.4484105,2.3269746,2.097231,1.847795,1.7558975,1.7591796,1.6902566,1.2800001,1.0765129,1.1913847,1.4933335,1.8051283,1.913436,2.0217438,2.3466668,2.5600002,2.5698464,2.5107694,2.7798977,2.6322052,2.4484105,2.4615386,2.7733335,2.92759,3.5577438,4.57518,5.35959,4.7622566,3.9253337,3.8990772,4.5489235,5.549949,6.380308,6.685539,6.9677954,6.931693,6.931693,7.955693,7.4830775,7.1581545,7.0892315,7.02359,6.340924,5.8289237,5.579488,5.398975,5.280821,5.3792825,6.3934364,7.3353853,7.6570263,7.318975,6.7938466,8.178872,8.710565,9.019077,9.252103,9.094564,1.5458462,1.6475899,1.8051283,1.972513,2.1202054,2.2350771,2.4943593,2.6912823,2.861949,3.0884104,3.495385,3.761231,3.7973337,3.9647183,4.4110775,5.074052,5.927385,5.9963083,5.940513,6.0291286,6.1538467,6.4754877,6.629744,6.9842057,7.4896417,7.6767187,6.9710774,6.8266673,6.954667,7.3353853,8.208411,8.5661545,9.344001,10.850462,13.292309,16.777847,18.49436,19.167181,22.025848,26.768412,29.554874,33.270157,40.18872,39.824413,29.77477,15.727591,10.587898,7.965539,6.242462,4.97559,4.893539,4.1517954,3.4822567,2.8488207,2.3302567,2.1169233,1.595077,1.2242053,1.0633847,1.020718,0.86317956,0.8992821,0.86974365,0.892718,0.8992821,0.6498462,0.35774362,0.318359,0.3314872,0.3314872,0.40697438,0.42994875,0.41025645,0.35774362,0.318359,0.34789747,0.38400003,0.32820517,0.256,0.18707694,0.08861539,0.059076928,0.108307704,0.24943592,0.446359,0.6301539,0.8763078,0.75487185,0.446359,0.20348719,0.34133336,0.20676924,0.0951795,0.032820515,0.059076928,0.2297436,0.28882053,0.40369233,0.48574364,0.46933338,0.318359,0.118153855,0.08205129,0.13784617,0.20676924,0.21333335,0.20676924,0.17723078,0.13128206,0.07548718,0.02297436,0.01969231,0.032820515,0.04594872,0.06235898,0.118153855,1.2274873,2.8225644,3.43959,3.2918978,4.2601027,5.1298466,5.2348723,4.6178465,3.9253337,4.414359,4.594872,5.034667,5.0904617,5.2348723,7.017026,7.785026,9.127385,9.40636,8.94359,10.000411,10.624001,11.808822,12.47836,12.790154,14.12595,12.947693,11.58236,10.902975,11.109744,11.716924,11.670976,11.434668,10.880001,10.535385,11.588924,10.072617,10.400822,11.753027,13.197129,13.702565,12.76718,13.095386,13.722258,14.168616,14.424617,13.689437,13.436719,13.13477,12.84595,13.236514,15.763694,16.86318,17.030565,16.548103,15.524104,17.414566,17.112617,16.105026,15.346873,15.258258,15.087591,14.857847,14.78236,14.788924,14.5263605,13.492514,12.438975,11.746463,11.648001,12.202667,13.157744,12.33395,12.068104,12.950975,13.827283,12.983796,12.232206,11.638155,11.313231,11.418258,11.608616,11.0375395,10.233437,9.718155,9.980719,9.275078,8.838565,8.539898,8.2215395,7.6964107,7.069539,6.9382567,7.381334,8.323282,9.5606165,9.93477,9.330873,8.730257,8.3823595,7.824411,7.13518,6.6527185,6.521436,6.5247183,6.0980515,6.2818465,6.7577443,7.8802056,9.4916935,10.9226675,10.509129,10.210463,10.305642,10.660104,10.7158985,9.449026,9.140513,9.537642,10.345026,11.254155,11.352616,11.155693,11.572514,12.737642,13.994668,13.88636,13.548308,12.967385,12.507898,12.898462,14.224411,14.956308,15.832617,16.682669,16.433231,16.009848,16.180513,16.361027,16.66954,17.939693,19.40677,20.004105,18.41231,15.241847,13.019898,12.947693,11.670976,9.974154,8.579283,8.129642,6.5345645,6.7216415,7.1844106,7.640616,9.061745,9.977437,10.308924,11.283693,12.980514,14.313026,16.46277,18.409027,17.814976,15.885129,17.345642,17.250463,15.724309,14.070155,13.036308,12.826258,10.06277,7.958975,6.170257,5.3202057,7.003898,8.743385,5.6451287,5.3694363,8.36595,7.88677,4.7392826,3.6529233,2.8356924,1.7985642,1.339077,1.3554872,1.0108719,0.9419488,1.5885129,3.2131286,4.332308,4.161641,4.785231,6.0619493,5.618872,5.074052,4.194462,3.6036925,3.498667,3.6726158,4.6112823,5.3037953,5.4383593,5.32677,5.8945646,8.182155,11.753027,15.107284,17.536001,19.140924,17.040411,12.619488,8.054154,4.5489235,2.359795,2.3630772,3.0358977,3.387077,4.007385,7.066257,10.039796,8.582564,8.103385,9.288206,8.109949,7.6143594,6.5017443,5.481026,4.916513,4.8114877,4.647385,4.414359,4.2436924,4.1911798,4.2338467,4.8771286,8.267488,11.644719,12.452104,8.326565,6.7840004,6.2588725,6.7117953,7.3321033,6.5411286,5.533539,6.5247183,7.171283,7.0826674,7.8473854,6.7117953,7.8736415,8.434873,7.9327188,8.369231,7.824411,6.0947695,4.850872,4.4438977,3.9286156,4.4373336,4.8836927,4.7425647,5.4186673,10.217027,4.84759,3.1474874,3.9286156,5.2644105,4.453744,4.699898,2.4451284,0.6629744,0.24287182,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.013128206,0.036102567,0.055794876,0.06564103,0.06564103,0.072205134,0.09189744,0.14112821,0.22646156,0.3446154,0.2855385,0.3314872,0.3708718,0.3708718,0.3708718,0.32820517,0.36102566,0.4397949,0.5349744,0.62030774,0.65312827,0.7122052,0.69907695,0.65312827,0.7318975,1.1881026,1.6968206,2.0086155,2.225231,2.7831798,3.436308,3.245949,3.0982566,3.495385,4.5390773,5.3398976,6.1538467,6.2818465,5.7764106,5.428513,5.3825645,5.408821,5.228308,4.9821544,5.2315903,4.6244106,4.529231,4.6966157,4.8607183,4.7622566,4.6966157,4.9099493,5.280821,5.8157954,6.633026,6.669129,6.5280004,6.2687182,6.180103,6.7610264,7.496206,7.719385,7.6110773,7.427283,7.522462,7.8506675,8.011488,7.965539,7.6012316,6.738052,7.3714876,7.7292314,8.103385,8.379078,8.027898,7.4929237,7.50277,7.88677,8.375795,8.608821,8.644924,9.508103,10.240001,10.538668,10.755282,9.997129,9.265231,8.700719,8.247795,7.6274877,7.6898465,7.5454364,7.9294367,8.4283085,7.4863596,7.27959,7.4765134,7.7357955,8.136206,9.18318,8.576,7.5585647,6.4000006,5.1922054,3.8367183,4.0402055,4.768821,5.0051284,4.5587697,4.073026,5.425231,6.114462,5.1856413,2.9243078,0.8467693,0.35446155,0.21989745,0.27897438,0.36430773,0.30194873,0.46933338,0.55794877,0.7450257,1.0732309,1.463795,1.8510771,2.2449234,2.5435898,2.6486156,2.4484105,2.044718,1.6869745,1.3981539,1.2603078,1.401436,1.4605129,1.4802053,1.4506668,1.4244103,1.5097437,1.8149745,1.9659488,2.1333334,2.2908719,2.2055387,1.6311796,1.5130258,1.5425643,1.6672822,2.0841026,2.3368206,2.412308,2.2186668,1.8937438,1.8215386,2.15959,2.6945643,3.186872,3.5249233,3.7284105,3.8596926,3.7185643,3.4789746,3.2951798,3.308308,3.5314875,3.373949,3.1737437,3.0949745,3.1245131,3.245949,3.245949,3.383795,3.5610259,3.314872,3.817026,4.4077954,5.077334,5.543385,5.2480006,5.4153852,5.533539,5.651693,5.674667,5.3694363,5.61559,6.048821,6.3868723,6.314667,5.467898,5.4186673,6.088206,6.806975,7.253334,7.4404106,7.1844106,7.0826674,6.9710774,7.13518,8.3134365,8.681026,8.809027,8.598975,8.218257,8.093539,7.653744,7.1909747,7.6110773,8.802463,9.636104,9.40636,9.386667,9.206155,8.720411,7.9786673,7.939283,7.210667,6.8004107,6.9087186,6.931693,6.226052,6.7150774,7.062975,6.9349747,7.0104623,7.312411,7.24677,7.194257,7.0925136,6.409847,6.314667,5.8978467,5.366154,4.6572313,3.436308,2.9669745,2.989949,2.681436,2.0217438,1.8116925,1.9692309,2.1398976,2.1825643,2.103795,2.0545642,1.8018463,1.5786668,1.4441026,1.3456411,1.1454359,1.0699488,1.3554872,1.6640002,1.8904617,2.1464617,2.2908719,2.537026,2.5862565,2.4746668,2.5435898,2.7963078,2.5107694,2.2711797,2.3466668,2.681436,3.062154,3.5577438,4.3027697,4.8771286,4.33559,3.7152824,3.7349746,4.276513,5.208616,6.373744,6.7314878,6.8266673,6.9120007,7.13518,7.5585647,7.53559,7.5585647,7.755488,7.7948723,6.885744,5.9536414,5.5630774,5.612308,5.970052,6.4722056,6.774154,7.2927184,7.9195905,8.178872,7.204103,8.090257,8.553026,8.822155,8.897642,8.553026,1.4802053,1.5885129,1.7362052,1.913436,2.0939488,2.2022567,2.4976413,2.7011285,2.7634873,2.8324106,3.239385,3.4002054,3.495385,3.7809234,4.338872,5.110154,5.8256416,5.927385,6.0160003,6.229334,6.2129235,6.6494365,7.02359,7.3419495,7.50277,7.2861543,6.9021544,6.8365135,6.87918,7.1483083,8.086975,8.28718,9.288206,10.860309,12.875488,15.307488,17.434258,19.534771,24.33313,29.922464,29.77477,32.630157,41.813335,42.496002,31.16636,15.625848,9.938052,7.3452315,6.058667,5.110154,4.3716927,3.367385,2.789744,2.4615386,2.2219489,1.9364104,1.3915899,1.1224617,1.0371283,1.0043077,0.86317956,0.8992821,0.9682052,0.92553854,0.72861546,0.4594872,0.2986667,0.3052308,0.33805132,0.35774362,0.40697438,0.39712822,0.3117949,0.25271797,0.23958977,0.21989745,0.29210258,0.25928208,0.19692309,0.13456412,0.068923086,0.049230773,0.0951795,0.23630771,0.48902568,0.84348726,0.9878975,0.83035904,0.5316923,0.27897438,0.28225642,0.190359,0.09189744,0.072205134,0.21333335,0.6071795,0.5349744,0.6826667,0.97805136,1.1716924,0.8369231,0.318359,0.15425642,0.13784617,0.15753847,0.190359,0.27897438,0.36102566,0.36102566,0.26256412,0.108307704,0.055794876,0.072205134,0.0951795,0.2297436,0.7417436,2.2744617,3.4921029,4.082872,4.7950773,7.4207187,7.138462,6.7840004,5.904411,4.818052,4.6145644,4.9821544,5.4843082,6.3442054,7.8112826,10.171078,11.063796,10.617436,10.226872,10.870154,13.138052,12.609642,13.446565,13.925745,14.037334,15.481437,13.853539,12.166565,11.516719,11.667693,11.057232,10.978462,11.208206,10.939077,10.518975,11.451077,10.909539,11.008,11.884309,12.973949,13.019898,12.566976,13.059283,13.978257,14.569027,13.833847,13.764924,14.332719,14.447591,14.145642,14.592001,16.515284,17.64431,17.61477,16.57436,15.176207,15.58318,15.323898,15.16636,15.350155,15.589745,15.832617,15.711181,15.37313,14.943181,14.532925,14.391796,13.499078,12.970668,13.115078,13.4170265,14.221129,13.751796,13.499078,13.912617,14.41477,13.797745,13.072412,12.274873,11.559385,11.162257,11.290257,10.692924,9.984001,9.668923,10.144821,10.102155,9.737847,9.4457445,9.15036,8.3134365,7.6274877,7.574975,8.146052,9.304616,11.008,11.011283,10.266257,9.511385,9.032206,8.661334,8.096821,7.2992826,7.026872,7.0826674,6.3179493,6.3179493,7.00718,8.109949,9.317744,10.276103,10.052924,10.000411,10.33518,10.985026,11.588924,10.023385,9.235693,9.432616,10.240001,10.71918,10.469745,10.354873,11.316514,13.35795,15.540514,14.7790785,13.856822,12.832822,12.137027,12.570257,13.538463,13.827283,14.352411,15.018668,14.726565,14.198155,14.867694,15.563488,15.95077,16.515284,18.034874,18.008617,16.406975,13.948719,12.097642,12.626052,11.82195,10.305642,8.907488,8.648206,7.1581545,7.397744,8.116513,9.005949,10.676514,11.428103,11.9860525,13.190565,14.851283,15.740719,17.70995,18.497643,18.002052,17.703386,20.683489,17.404718,16.341335,14.6642065,12.278154,11.825232,10.469745,10.801231,10.522257,9.409642,9.304616,9.747693,7.1876926,7.460103,10.496001,10.328616,6.11118,4.8836927,3.948308,2.4484105,1.3686155,1.3751796,1.024,1.148718,2.1858463,4.1485133,5.9536414,4.601436,3.5872824,4.210872,5.546667,6.088206,5.1200004,4.027077,3.4002054,3.0424619,3.5380516,5.4908724,6.449231,5.9963083,5.733744,6.1997952,8.569437,10.807796,12.114052,12.901745,12.27159,10.584617,8.395488,5.8781543,2.858667,2.4648206,2.484513,2.5238976,2.6584618,3.4264617,7.5913854,7.5881033,7.13518,7.53559,7.6701546,7.0531287,6.180103,5.691077,5.5532312,5.0674877,4.5423594,4.0992823,4.450462,5.0904617,4.2929235,2.868513,4.8771286,8.690872,11.559385,9.622975,5.920821,5.5138464,6.7774363,7.5388722,5.093744,4.7950773,6.294975,7.387898,7.6996927,8.674462,9.225847,8.438154,7.653744,7.4240007,7.512616,5.9503593,4.5390773,4.2207184,4.630975,4.092718,2.6486156,3.9318976,4.562052,4.2994876,6.0258465,2.878359,2.028308,2.3991797,3.1737437,3.8104618,4.1025643,2.1530259,0.57764107,0.18707694,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.009846155,0.029538464,0.055794876,0.068923086,0.049230773,0.06235898,0.08861539,0.14112821,0.21989745,0.32164106,0.3249231,0.37743592,0.39712822,0.36758977,0.3314872,0.3249231,0.32820517,0.36102566,0.43323082,0.571077,0.6892308,0.7515898,0.65641034,0.56123084,0.88615394,1.0568206,1.6640002,2.3335385,2.7995899,2.8750772,3.1409233,2.9538465,2.865231,3.2065644,4.066462,4.4800005,5.2545643,5.4449234,5.077334,5.142975,4.919795,5.0674877,4.926359,4.644103,5.156103,4.9132314,5.0182567,5.034667,4.890257,4.886975,4.896821,5.356308,5.605744,5.687795,6.3277955,6.3376417,5.8190775,5.4613338,5.681231,6.633026,7.653744,8.093539,7.9524107,7.4830775,7.210667,7.427283,7.4863596,7.574975,7.515898,6.764308,7.0400004,7.3583593,7.890052,8.4283085,8.372514,8.198565,8.5891285,8.979693,9.160206,9.26195,9.370257,10.14154,10.696206,10.827488,10.9915905,10.121847,9.242257,8.553026,8.103385,7.7718983,7.460103,7.64718,8.454565,9.061745,7.6996927,7.857231,7.965539,8.172308,8.78277,10.269539,9.101129,6.5345645,4.906667,4.6539493,4.2994876,4.7950773,5.7107697,6.3507695,6.4032826,5.933949,6.2818465,6.442667,5.0838976,2.4549747,0.40697438,0.21661541,0.14441027,0.14112821,0.16082053,0.13784617,0.256,0.318359,0.48574364,0.761436,1.020718,1.5721027,2.044718,2.4320002,2.6518977,2.5764105,2.0644104,1.7394873,1.4473847,1.214359,1.2406155,1.3029745,1.332513,1.3161026,1.2964103,1.3817437,1.6672822,2.0906668,2.3893335,2.3893335,2.0053334,1.6082052,1.5885129,1.6672822,1.8182565,2.281026,2.3958976,2.284308,1.9200002,1.585231,1.8773335,2.3302567,2.7569232,3.1343591,3.4166157,3.5282054,3.6890259,3.5347695,3.3903592,3.3936412,3.508513,3.387077,3.2131286,3.1048207,3.1015387,3.1737437,3.2853336,3.2295387,3.2623591,3.3641028,3.2525132,3.8695388,4.637539,5.2644105,5.5729237,5.5007186,5.5926156,5.681231,5.8125134,5.8978467,5.72718,6.183385,6.5837955,6.6461544,6.3245134,5.792821,5.723898,6.2129235,6.701949,7.0137444,7.3485136,7.1056414,7.2172313,7.4830775,7.9130263,8.746667,9.222565,9.199591,8.94359,8.602257,8.208411,7.75877,7.2664623,7.578257,8.55959,9.107693,9.432616,9.219283,8.78277,8.254359,7.574975,7.387898,6.918565,6.547693,6.5050263,6.8397956,5.989744,6.3376417,7.207385,7.8539495,7.4797955,7.4765134,7.716103,8.057437,8.103385,7.213949,6.633026,6.38359,5.933949,5.077334,3.9318976,3.0818465,2.9243078,2.6683078,2.1398976,1.782154,1.7033848,1.7657437,1.8116925,1.7788719,1.7066668,1.5655385,1.463795,1.3522053,1.2438976,1.2176411,1.3062565,1.6147693,1.8674873,2.0020514,2.1825643,2.3729234,2.5600002,2.5764105,2.4943593,2.6289232,2.8816411,2.605949,2.353231,2.409026,2.7864618,3.249231,3.6332312,4.1025643,4.44718,4.086154,3.5544617,3.7284105,4.3027697,5.172513,6.416411,6.7610264,6.8463597,7.2270775,7.830975,7.962257,7.77518,7.8441033,8.090257,8.146052,7.3485136,6.2752824,6.2227697,6.436103,6.7085133,7.387898,7.3419495,7.5454364,8.283898,8.881231,7.719385,8.234667,8.635077,8.743385,8.503796,7.9819493,1.5064616,1.7165129,1.7624617,1.847795,2.028308,2.2186668,2.5173335,2.7470772,2.7634873,2.7208207,3.0884104,3.131077,3.2623591,3.639795,4.2240005,4.7655387,5.280821,5.687795,6.1374364,6.49518,6.3343596,6.6002054,7.1483083,7.5520005,7.568411,7.1548724,7.256616,7.3058467,7.273026,7.463385,8.546462,8.907488,9.760821,11.021129,12.540719,14.080001,16.505438,20.073027,26.059488,31.757132,30.464003,33.024002,44.356926,46.086567,33.4638,15.37313,9.426052,6.813539,6.048821,5.61559,3.948308,2.5862565,2.0676925,1.9659488,1.8904617,1.5097437,1.204513,1.211077,1.1651284,1.0338463,1.1290257,1.0962052,1.1323078,0.97805136,0.6826667,0.6071795,0.54482055,0.508718,0.47917953,0.47917953,0.574359,0.5907693,0.40369233,0.29538465,0.3117949,0.26256412,0.2297436,0.17066668,0.118153855,0.07876924,0.06564103,0.049230773,0.072205134,0.21989745,0.5284103,0.99774367,1.1454359,0.9353847,0.62030774,0.3446154,0.16738462,0.08861539,0.032820515,0.09189744,0.3446154,0.88943595,0.77456415,0.94523084,1.4539489,1.9200002,1.4998976,0.7187693,0.34133336,0.16410258,0.08533334,0.11158975,0.24615386,0.4266667,0.50543594,0.42994875,0.22646156,0.1148718,0.118153855,0.16738462,0.5546667,1.9593848,3.3411283,4.4832826,5.3103595,6.567385,9.796924,8.39877,7.4896417,6.5411286,5.586052,5.2053337,5.907693,6.166975,7.2992826,9.777231,13.236514,12.5374365,11.503591,11.936821,14.011078,16.246155,15.409232,14.992412,15.225437,15.868719,16.213335,14.250668,12.386462,11.667693,11.631591,10.289231,10.108719,10.765129,11.1294365,10.79795,10.102155,11.739899,12.235488,12.209231,12.002462,11.690667,12.412719,13.548308,14.191591,14.165335,14.03077,14.890668,15.205745,15.681643,16.265848,16.134565,16.630156,16.86318,16.646564,15.780104,14.060308,12.248616,12.583385,13.482668,14.28677,15.264822,15.671796,16.213335,15.763694,14.460719,13.692719,14.710155,14.6182575,14.519796,14.598565,14.112822,15.104001,15.130258,14.546052,13.899488,13.935591,14.089848,14.024206,13.361232,12.310975,11.690667,11.293539,10.627283,10.118565,10.036513,10.466462,11.07036,11.0375395,10.70277,10.134975,9.140513,8.411898,8.513641,9.173334,10.331899,12.137027,12.176412,11.408411,10.604308,10.006975,9.321027,9.15036,8.218257,7.7423596,7.6668725,6.675693,6.564103,7.4174366,8.651488,9.642668,9.718155,9.488411,9.947898,10.735591,11.579078,12.314258,10.820924,9.80677,10.039796,11.011283,10.935796,9.993847,9.947898,11.355898,13.896206,16.36431,15.346873,14.313026,13.016617,11.96636,12.425847,12.63918,12.35036,12.501334,13.010053,12.793437,12.1238985,13.157744,14.546052,15.504412,15.809642,16.554668,15.668514,14.112822,12.731078,12.235488,12.655591,12.22236,11.175385,10.013539,9.481847,8.723693,9.163487,10.115283,11.286975,12.773745,13.617231,15.619284,17.142155,17.723078,18.07754,19.446156,17.47036,15.875283,16.626873,19.945026,15.136822,15.616001,15.360002,12.616206,9.90195,9.271795,12.832822,15.012104,14.316309,13.328411,10.9456415,7.643898,6.7544622,8.467693,9.829744,5.2676926,3.751385,3.249231,2.6256413,1.6311796,1.273436,0.8598975,1.270154,2.5173335,3.7448208,6.170257,6.0258465,4.4964104,3.1671798,4.020513,5.146257,4.8804107,3.7973337,2.6584618,2.422154,1.8215386,3.9614363,5.901129,6.416411,5.979898,5.668103,8.01477,9.898667,10.246565,10.013539,8.989539,8.707283,8.395488,7.250052,4.4340515,2.8553848,2.5206156,2.7602053,2.8324106,1.9003079,4.0500517,5.4449234,5.405539,4.716308,5.618872,5.0051284,4.7491283,5.4153852,6.436103,6.088206,4.1124105,3.5577438,4.5095387,5.805949,5.0576415,3.4888208,2.4615386,3.8334363,6.8529234,8.146052,4.7261543,4.8082056,6.994052,8.36595,4.5029745,3.7120004,4.4832826,5.904411,7.4797955,9.156924,9.590155,8.320001,7.716103,7.817847,6.36718,4.453744,3.8071797,4.535795,5.425231,3.9286156,2.2383592,3.4034874,3.7284105,2.7241027,3.1081028,3.058872,2.4024618,1.6147693,1.4408206,2.8882053,1.9922053,0.86317956,0.16410258,0.01969231,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.02297436,0.036102567,0.026256412,0.06564103,0.072205134,0.10502565,0.16410258,0.21333335,0.32164106,0.39384618,0.41682056,0.39384618,0.35446155,0.39712822,0.36102566,0.32820517,0.34133336,0.41682056,0.571077,0.77456415,0.7122052,0.57764107,1.0732309,1.0633847,2.1825643,3.0194874,3.1376412,3.1048207,2.681436,2.6912823,2.9243078,3.2032824,3.3772311,3.6791797,4.388103,4.706462,4.6605134,5.1167183,4.821334,5.149539,5.2578464,5.100308,5.464616,5.868308,6.0225644,5.6418467,5.0642056,5.2578464,5.1626673,5.7632823,5.927385,5.671385,6.121026,6.0816417,5.7731285,5.7665644,6.262154,7.072821,8.569437,9.065026,8.641642,7.6701546,6.8266673,6.685539,6.4065647,6.416411,6.6822567,6.7314878,6.688821,6.744616,7.1122055,7.6734366,7.975385,8.034462,8.795898,9.383386,9.573745,9.80677,10.269539,10.732308,11.047385,11.034257,10.453334,9.7214365,9.130668,8.4512825,7.8080006,7.6668725,7.6012316,8.080411,8.805744,9.088,7.8670774,8.070564,7.9097443,8.001641,8.815591,10.673231,9.521232,6.0061545,3.5446157,3.255795,3.9647183,5.7698464,6.554257,7.1581545,8.083693,9.504821,7.75877,6.3868723,4.70318,2.6256413,0.67282057,0.27241027,0.13784617,0.18051283,0.256,0.16082053,0.27569234,0.35446155,0.4004103,0.50543594,0.8467693,1.401436,1.7427694,2.0742567,2.4024618,2.5435898,2.2383592,1.9364104,1.6114873,1.2964103,1.083077,1.0469744,1.1946667,1.3029745,1.3095386,1.3193847,1.6836925,2.1792822,2.3860514,2.1924105,1.7985642,1.6869745,1.7460514,1.8543591,2.028308,2.412308,2.4024618,2.281026,1.9331284,1.657436,2.166154,2.5632823,2.865231,3.2000003,3.4592824,3.2820516,3.1015387,3.121231,3.2262566,3.3378465,3.4231799,3.3280003,3.3247182,3.3280003,3.314872,3.3247182,3.2886157,3.1442053,3.117949,3.3312824,3.8137438,4.017231,4.8377438,5.428513,5.549949,5.5762057,5.8125134,6.0291286,6.124308,6.1505647,6.308103,6.695385,6.764308,6.5903597,6.304821,6.0783596,6.012718,6.5083084,6.921847,7.076103,7.240206,7.2172313,7.525744,8.15918,8.884514,9.216001,9.586872,9.229129,8.713847,8.267488,7.765334,7.5191803,7.456821,7.7325134,8.149334,8.152616,9.281642,8.914052,8.044309,7.213949,6.488616,6.3179493,6.6527185,6.6002054,6.314667,6.9809237,6.2785645,6.2194877,7.1548724,8.41518,8.339693,7.8047185,7.9885135,8.372514,8.3134365,7.0400004,6.0324106,6.196513,6.121026,5.3727183,4.4898467,3.508513,2.8816411,2.5271797,2.2219489,1.6443079,1.4112822,1.3489232,1.4736412,1.6180514,1.4145643,1.3817437,1.4998976,1.5327181,1.4506668,1.4145643,1.6213335,1.7624617,1.9167181,2.0578463,2.0184617,2.284308,2.5074873,2.6289232,2.6912823,2.809436,3.0720003,2.9801028,2.8192823,2.8160002,3.1606157,3.3641028,3.5741541,3.9220517,4.240411,4.082872,3.515077,3.9187696,4.6802053,5.540103,6.5772314,6.9645133,7.328821,8.001641,8.812308,9.078155,8.41518,8.188719,8.044309,7.8145647,7.525744,6.6527185,7.3025646,7.765334,7.709539,8.185436,8.188719,8.241231,8.740103,9.248821,8.500513,8.582564,8.677744,8.470975,7.9983597,7.643898,1.4342566,1.8871796,1.8970258,1.8116925,1.8773335,2.2416413,2.0217438,2.353231,2.674872,2.806154,2.930872,2.989949,2.986667,3.1540515,3.373949,3.2032824,4.266667,5.110154,5.865026,6.445949,6.5312824,6.7249236,7.581539,8.1066675,8.195283,8.621949,8.096821,7.581539,7.6734366,8.3364105,8.910769,9.898667,10.5780525,11.565949,13.078976,14.923489,15.668514,19.96472,25.511387,29.023182,26.213745,36.919796,49.99549,49.604927,33.94954,15.274668,9.475283,6.7085133,5.402257,4.4373336,3.1442053,1.8970258,1.5425643,1.4605129,1.3883078,1.3883078,1.3161026,1.2504616,1.1651284,1.1651284,1.4966155,1.6311796,1.332513,0.9747693,0.79097444,0.8992821,1.1684103,1.0633847,0.93866676,1.0010257,1.2832822,1.3193847,0.92553854,0.6498462,0.5546667,0.21333335,0.14112821,0.10502565,0.098461546,0.10502565,0.09189744,0.055794876,0.072205134,0.19692309,0.36430773,0.4135385,0.86317956,0.764718,0.44964105,0.15425642,0.04594872,0.032820515,0.013128206,0.02297436,0.108307704,0.28882053,0.4594872,0.8598975,1.3686155,1.7591796,1.7099489,1.2077949,0.58092314,0.18379489,0.101743594,0.13784617,0.12471796,0.15753847,0.190359,0.20020515,0.21333335,0.190359,0.16410258,0.23302566,0.95835906,3.387077,4.4865646,5.3005133,5.3202057,5.2414365,6.987488,5.4613338,5.9503593,6.5378466,6.744616,7.5388722,9.03877,8.15918,7.496206,8.339693,10.696206,9.793642,12.586668,15.694771,17.073233,16.036104,14.500104,15.632411,16.403694,15.530668,13.505642,13.6008215,11.585642,10.289231,10.243283,9.642668,10.535385,11.270565,11.286975,10.601027,9.796924,11.247591,11.493745,11.35918,11.264001,11.21477,12.521027,14.55918,15.360002,15.031796,15.776822,17.096207,16.676104,17.401438,19.35754,19.820309,18.635489,16.20677,14.657642,14.486976,14.572309,12.301129,12.199386,12.737642,13.410462,14.739694,14.03077,14.742975,14.431181,13.108514,13.22995,13.193847,13.935591,14.690463,14.916924,14.283488,15.24513,16.128002,15.744001,14.362258,13.702565,14.191591,14.634667,14.529642,13.827283,12.924719,12.593232,11.723488,10.975181,10.771693,11.323078,11.30995,11.674257,11.979488,11.72677,10.361437,9.849437,9.554052,9.829744,10.807796,12.406155,13.088821,12.737642,12.242052,11.503591,9.429334,8.576,8.169026,7.9327188,7.6898465,7.384616,7.020308,7.5946674,8.815591,9.83959,9.278359,10.144821,10.453334,11.178667,12.373334,13.167591,11.753027,10.620719,10.663385,11.670976,12.327386,11.851488,11.405129,12.228924,14.263796,16.144411,15.2155905,14.086565,13.115078,12.547283,12.511181,11.670976,11.513436,11.989334,12.560411,12.20595,12.3766165,13.810873,15.136822,15.652103,15.333745,15.153232,14.237539,13.124924,12.550565,13.443283,12.809847,12.852514,12.632616,11.861334,10.909539,10.873437,11.37559,12.675283,14.447591,15.776822,17.69354,22.117744,24.041027,22.373745,19.958155,19.908924,17.289848,14.943181,14.306462,15.379693,15.258258,15.80636,16.06236,14.601848,9.537642,7.6570263,9.43918,11.349334,12.475078,14.5263605,14.854566,7.962257,4.0303593,6.633026,12.711386,5.47118,2.6289232,2.225231,2.4976413,1.8609232,1.4966155,1.0666667,0.74830776,0.7187693,1.1454359,4.588308,4.8082056,3.8006158,2.7241027,1.9068719,2.7503593,3.9680004,3.698872,2.4352822,3.0227695,2.3138463,2.0086155,3.0949745,4.965744,5.4153852,4.1091285,4.3618464,5.5630774,6.485334,5.2644105,5.228308,5.9602056,6.7216415,6.961231,6.301539,2.7142565,1.5885129,2.3269746,3.7809234,4.2568207,5.5762057,5.546667,4.571898,3.7251284,4.775385,4.44718,3.879385,4.4832826,6.235898,7.6734366,6.442667,5.208616,4.342154,4.201026,5.142975,6.436103,4.197744,2.5665643,3.006359,4.2896414,3.9811285,3.9154875,4.70318,5.664821,4.821334,3.3936412,3.9811285,5.7796926,7.8112826,8.910769,7.128616,8.001641,9.947898,10.541949,6.5017443,5.536821,3.3903592,2.7864618,3.5872824,2.793026,3.4264617,4.2830772,4.31918,3.3378465,1.9823592,0.90912825,0.38400003,0.38400003,0.6662565,0.764718,0.20020515,0.02297436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.052512825,0.06235898,0.072205134,0.10502565,0.15097436,0.20020515,0.25928208,0.32164106,0.36758977,0.36758977,0.29210258,0.256,0.32820517,0.42994875,0.32164106,0.3446154,0.67282057,0.7581539,0.5973334,0.7318975,1.4998976,3.1770258,3.495385,2.4943593,2.5173335,2.2121027,2.5665643,3.0982566,3.3411283,2.8521028,3.6726158,4.086154,4.453744,4.6539493,4.1058464,3.8859491,4.9362054,5.907693,6.235898,6.1505647,6.2096415,5.7665644,5.5007186,5.5893335,5.720616,5.3431797,5.907693,6.4032826,6.62318,7.171283,6.87918,6.87918,7.312411,8.195283,9.429334,10.699488,10.604308,9.5606165,8.231385,7.522462,6.2785645,5.5269747,5.3694363,5.720616,6.3179493,6.3901544,6.189949,6.5444107,7.3747697,7.706257,7.509334,7.755488,7.8834877,7.7423596,7.584821,9.609847,10.893129,11.188514,10.512411,9.170052,8.060719,8.267488,8.04759,7.1909747,7.020308,7.325539,7.8047185,8.395488,8.78277,8.392206,8.0377445,7.9130263,8.011488,8.720411,10.817642,9.120821,5.8125134,4.46359,5.0642056,4.013949,5.221744,5.477744,5.024821,5.7468724,11.152411,10.226872,8.914052,6.892308,4.345436,1.9528207,0.5973334,0.18707694,0.2297436,0.3446154,0.25928208,0.6859488,0.8566154,0.8205129,0.7975385,1.1749744,1.6640002,1.847795,1.9593848,2.1530259,2.5337439,2.6551797,2.0808206,1.5819489,1.339077,0.9616411,0.9747693,1.1684103,1.2964103,1.3292309,1.463795,2.1103592,2.3269746,2.2186668,2.041436,2.2121027,1.9561027,1.9200002,2.097231,2.3368206,2.349949,2.412308,2.225231,1.9003079,1.6672822,1.8609232,2.5206156,3.0424619,3.3345644,3.3936412,3.2951798,3.1245131,3.1474874,2.8849232,2.484513,2.7175386,3.0227695,3.308308,3.3936412,3.3247182,3.370667,3.2000003,3.0654361,3.2689233,3.826872,4.4865646,4.1813335,4.663795,5.297231,5.76,6.0258465,6.1374364,6.183385,6.1997952,6.3573337,6.941539,7.026872,6.7577443,6.426257,6.1768208,5.979898,6.482052,7.2927184,7.7325134,7.643898,7.4010262,7.571693,8.008205,8.549745,8.897642,8.605539,8.556309,8.408616,8.1755905,7.824411,7.2631803,7.312411,8.04759,8.4512825,8.247795,7.9195905,8.982975,8.2215395,7.1548724,6.416411,5.7665644,5.5958977,6.8529234,7.13518,6.3474874,6.7150774,7.00718,7.3714876,8.008205,8.756514,9.110975,8.241231,7.7325134,7.384616,7.125334,7.003898,5.868308,5.904411,5.924103,5.4547696,4.7458467,3.9384618,3.5282054,3.2032824,2.6584618,1.5721027,1.3259488,1.1027694,1.1749744,1.4506668,1.4506668,1.2898463,1.2964103,1.273436,1.2307693,1.3883078,1.7066668,1.591795,1.6902566,2.0053334,1.9068719,2.225231,2.7076926,2.9801028,3.006359,3.0654361,3.2984617,3.495385,3.629949,3.748103,3.9680004,3.515077,3.1376412,3.3575387,3.9253337,3.8137438,3.3641028,3.9647183,4.8738465,5.720616,6.514872,7.2369237,7.8637953,8.182155,8.346257,8.89436,9.189744,9.143796,8.001641,6.560821,7.171283,6.7085133,7.315693,8.3823595,9.478565,10.345026,10.174359,9.216001,9.094564,9.7673855,9.537642,9.02236,8.100103,7.4108725,7.2894363,7.765334,1.8740515,2.0118976,1.9528207,1.8642052,1.8445129,1.9364104,1.8445129,2.0512822,2.356513,2.674872,3.0523078,3.0851285,3.1081028,3.2098465,3.3969233,3.6069746,4.210872,4.6966157,4.9493337,5.0904617,5.467898,5.868308,6.482052,7.1187696,7.6110773,7.8047185,7.250052,7.4141545,7.525744,7.6635904,8.763078,9.636104,10.857026,12.566976,14.496821,15.960617,18.005335,21.704206,23.985233,24.612104,26.190771,41.22257,47.425644,40.274055,23.952412,11.378873,8.316719,6.0324106,4.414359,3.2787695,2.3860514,2.1070771,1.8248206,1.5753847,1.3850257,1.2668719,1.1355898,1.1290257,1.2012309,1.2964103,1.3718976,1.1946667,0.9321026,0.6695385,0.49887183,0.508718,0.8369231,0.7089231,0.53825647,0.5349744,0.7089231,0.7450257,0.61374366,0.42338464,0.24615386,0.128,0.0951795,0.06564103,0.06564103,0.09189744,0.128,0.052512825,0.06235898,0.13456412,0.39384618,1.0962052,1.9856411,1.4867693,0.7089231,0.2231795,0.04594872,0.02297436,0.02297436,0.098461546,0.26912823,0.508718,0.5349744,0.72861546,1.0108719,1.2537436,1.2832822,1.0732309,0.56123084,0.21333335,0.18707694,0.3314872,0.7417436,0.46933338,0.380718,0.54482055,0.22646156,1.1782565,2.2383592,2.8816411,3.1442053,3.629949,3.6168208,3.515077,3.442872,3.7842054,5.2053337,5.5269747,5.297231,5.4482055,6.1505647,6.816821,8.953437,8.759795,9.028924,10.331899,11.0375395,11.188514,11.999181,14.037334,16.01641,14.792206,15.264822,16.787693,16.807386,15.396104,15.225437,13.771488,11.936821,10.8996935,10.837335,10.912822,11.559385,11.434668,11.753027,12.209231,11.004719,10.505847,10.6469755,10.742155,10.971898,12.386462,13.682873,15.0088215,15.9343605,16.292105,16.167385,17.165129,18.15631,18.06113,16.922258,15.891693,14.647796,13.873232,14.063591,14.7561035,14.55918,12.964104,12.291283,12.47836,13.74195,16.594053,15.809642,14.106257,13.220103,13.177437,12.314258,12.678565,13.065847,13.495796,13.761642,13.4400015,14.004514,14.683899,14.844719,14.444309,14.020925,14.011078,14.217847,14.437745,14.49354,14.25395,14.034052,13.298873,12.281437,11.178667,10.174359,11.1294365,12.416001,13.226667,13.069129,11.753027,10.134975,9.580308,10.036513,11.109744,12.064821,11.779283,12.396309,12.826258,12.448821,11.113027,9.488411,8.65477,8.438154,8.536616,8.533334,7.8441033,8.362667,9.435898,10.161232,9.373539,10.748719,12.744206,14.168616,14.897232,15.8654375,13.873232,11.881026,10.722463,10.70277,11.595488,12.176412,12.025436,12.78359,14.139078,13.860104,13.558155,13.039591,13.249642,13.840411,13.157744,11.467488,11.510155,12.107488,12.642463,13.062565,14.158771,14.588719,15.346873,16.210052,15.737437,17.585232,16.905848,15.494565,14.575591,14.821745,13.971693,13.46954,13.216822,12.806565,11.533129,13.039591,14.49354,16.603899,18.691284,18.694565,20.319181,32.57108,37.00513,29.56472,20.60472,18.97354,16.689232,15.783386,16.275694,16.200207,14.083283,12.675283,11.690667,11.323078,12.235488,9.212719,9.91836,9.816616,8.67118,10.535385,13.843694,9.826463,5.4843082,4.8672824,9.061745,6.012718,4.821334,5.077334,5.146257,2.166154,1.8871796,1.5392822,1.2274873,1.1552821,1.6311796,2.487795,2.793026,4.1813335,6.0192823,5.3858466,4.33559,3.7382567,2.9505644,2.0873847,2.0086155,1.6213335,1.8018463,2.5928206,3.5511796,3.7218463,3.0785644,3.5544617,4.1747694,4.886975,6.557539,5.4974365,4.896821,4.5587697,4.414359,4.5062566,3.7021542,3.6463592,4.269949,4.857436,4.023795,5.0215387,5.1265645,4.640821,4.128821,4.397949,6.117744,5.7501545,4.7261543,4.1222568,4.6244106,4.630975,5.4514875,5.540103,4.8836927,4.9821544,4.9788723,4.1058464,3.6036925,3.7907696,4.066462,5.6385646,5.1889234,4.663795,4.827898,5.2742567,4.3027697,4.381539,5.546667,7.604513,10.118565,7.9852314,7.9491286,8.730257,8.704,5.914257,7.0793853,6.1013336,6.2687182,6.941539,3.5478978,3.5971284,4.0336413,4.3290257,4.0434875,2.8258464,2.0250258,1.6049232,1.1946667,0.6892308,0.24943592,0.068923086,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.0032820515,0.01969231,0.04594872,0.07876924,0.128,0.22646156,0.20676924,0.22646156,0.256,0.28225642,0.28225642,0.31507695,0.33476925,0.3446154,0.3314872,0.27241027,0.3052308,0.5316923,0.69579494,0.76800007,0.9517949,1.8281027,2.806154,2.934154,2.5042052,3.05559,2.6223593,2.8291285,2.8422565,2.5271797,2.4516926,3.0720003,3.498667,3.9876926,4.4373336,4.384821,4.457026,5.681231,7.2861543,8.251078,7.2960005,6.5870776,6.4557953,6.4754877,6.301539,5.674667,5.0609236,5.0609236,5.405539,5.8781543,6.3277955,6.806975,7.030154,7.3616414,7.768616,7.817847,9.058462,9.147078,8.641642,8.073847,7.962257,7.1548724,6.675693,6.626462,6.997334,7.683283,7.8834877,7.634052,7.325539,7.0957956,6.8397956,7.1122055,7.6274877,7.6176414,7.312411,7.9261546,8.730257,9.284924,9.764103,9.9282055,9.133949,8.297027,8.146052,8.044309,7.7292314,7.325539,8.116513,8.185436,7.936001,7.75877,8.001641,6.9645133,7.2172313,7.939283,8.214975,7.0334363,6.8693337,7.0432825,8.766359,10.115283,6.038975,6.2720003,7.2861543,8.369231,9.209436,9.921641,10.820924,8.828718,6.163693,4.7360005,6.1505647,1.5655385,0.26584616,0.32164106,0.571077,0.60061544,1.0469744,1.1355898,1.1881026,1.4080001,1.8937438,1.6705642,1.847795,2.038154,2.1300514,2.2646155,2.3958976,2.0808206,1.6672822,1.3292309,1.0601027,1.1684103,1.1618463,1.2471796,1.4506668,1.6246156,1.8806155,1.9331284,2.0217438,2.1431797,2.028308,1.7624617,1.9593848,2.2055387,2.3433847,2.4713848,2.0644104,1.8412309,1.9462565,2.2416413,2.300718,2.6289232,2.9505644,2.8750772,2.6683078,3.2361028,2.9078977,2.917744,3.0752823,3.3050258,3.6430771,3.7349746,3.6069746,3.4198978,3.2886157,3.2984617,3.2951798,3.0687182,3.495385,4.5489235,5.3169236,4.571898,4.4307694,4.6276927,4.893539,4.9788723,5.3891287,5.76,6.189949,6.5805135,6.6494365,6.99077,7.0137444,6.8332314,6.521436,6.1407185,6.5247183,7.2237954,7.8112826,8.096821,8.146052,7.965539,8.152616,8.484103,8.713847,8.556309,9.005949,9.019077,8.425026,7.5552826,7.2270775,6.8463597,7.253334,7.827693,8.201847,8.274052,8.493949,7.893334,6.9809237,6.242462,6.1341543,5.671385,5.917539,6.1013336,6.163693,6.764308,7.056411,7.2894363,7.9819493,8.996103,9.524513,9.301334,8.477539,7.860513,7.634052,7.3452315,6.11118,6.045539,5.8125134,5.0838976,4.5128207,4.07959,3.626667,3.245949,2.802872,1.9495386,1.4145643,1.2471796,1.339077,1.4998976,1.4605129,1.332513,1.3817437,1.4375386,1.4703591,1.6213335,1.7329233,1.7001027,1.8116925,2.034872,2.0053334,2.284308,2.7175386,3.0523078,3.239385,3.4560003,3.3969233,3.314872,3.501949,3.9942567,4.565334,3.8498464,3.4133337,3.4034874,3.6529233,3.6791797,4.0008206,4.5095387,5.0674877,5.7042055,6.626462,7.6668725,8.51036,9.147078,9.504821,9.409642,8.628513,7.939283,7.13518,6.6592827,7.6110773,7.79159,8.320001,9.097847,9.957745,10.637129,10.44677,9.330873,9.110975,9.911796,10.148104,8.969847,8.297027,7.9195905,7.7948723,8.034462,1.8543591,1.910154,1.8871796,1.8904617,1.910154,1.8149745,2.041436,2.2777438,2.5764105,2.9407182,3.3280003,3.186872,3.117949,3.170462,3.383795,3.8006158,4.1485133,4.525949,4.57518,4.397949,4.571898,5.287385,6.163693,6.8529234,7.4108725,8.283898,7.6570263,7.8769236,7.8408213,7.6242056,8.500513,9.399796,11.313231,14.086565,17.08636,19.177027,23.16472,24.267488,23.903181,25.298054,33.47036,42.151386,38.11775,26.742155,14.283488,7.8802056,6.1308722,4.588308,3.3509746,2.4681027,1.9331284,1.8576412,1.6213335,1.3850257,1.1881026,0.9616411,0.9321026,1.0469744,1.2635899,1.4145643,1.204513,0.97805136,0.7581539,0.60389745,0.5546667,0.6301539,0.92225647,0.9189744,0.7450257,0.57764107,0.6301539,0.71548724,0.6432821,0.49230772,0.3314872,0.23630771,0.20348719,0.14441027,0.190359,0.27569234,0.128,0.16738462,0.23302566,0.56123084,1.2471796,2.2449234,2.6157951,1.913436,0.9714873,0.2986667,0.072205134,0.032820515,0.016410258,0.072205134,0.19692309,0.3446154,0.5021539,0.88943595,1.3456411,1.6344616,1.4408206,0.90912825,0.71548724,0.571077,0.43323082,0.46276927,0.8533334,0.8369231,0.77128214,0.7778462,0.7318975,2.0086155,2.7273848,3.0227695,3.1606157,3.5282054,3.2361028,2.993231,3.3378465,4.07959,4.3027697,5.671385,5.58277,5.549949,6.3868723,8.231385,9.330873,9.741129,10.571488,11.392001,10.236719,11.332924,11.191795,11.9171295,13.656616,14.598565,15.14995,16.147694,16.498873,15.8884115,14.775796,12.691693,12.232206,12.084514,11.841642,11.999181,11.772718,10.66995,10.476309,11.224616,11.204924,10.561642,10.919386,11.290257,11.355898,11.500309,13.66318,15.382976,16.771284,17.499899,16.768002,16.292105,17.778873,18.179283,16.679386,14.697027,14.129231,14.313026,14.401642,14.093129,13.640206,13.019898,12.603078,13.285745,14.897232,16.200207,15.832617,14.7561035,14.171899,14.290052,14.329437,14.36554,13.676309,13.249642,13.275898,13.11836,13.59754,14.500104,14.706873,14.208001,14.099693,13.912617,13.7386675,13.850258,14.158771,14.194873,14.181745,13.840411,13.010053,11.82195,10.692924,11.099898,12.35036,13.778052,14.303181,12.448821,10.469745,10.039796,10.325335,10.640411,10.459898,10.738873,11.864616,12.504617,12.3076935,11.894155,10.820924,10.089026,9.6525135,9.32759,8.792616,8.500513,9.15036,10.151385,10.614155,9.353847,11.10318,13.692719,15.540514,16.315079,16.935387,14.8709755,12.563693,10.8307705,10.167795,10.755282,11.618463,11.296822,11.74318,13.052719,13.472821,13.489232,12.507898,12.120616,12.35036,11.644719,11.0145645,11.88759,12.711386,13.069129,13.676309,14.907078,15.29436,16.200207,17.476925,17.476925,20.227283,19.18031,17.240616,16.187078,16.659693,15.960617,14.296617,13.289026,13.036308,12.12718,15.087591,18.248207,21.16595,22.436104,19.689028,23.811283,47.025234,56.37908,43.52985,24.740105,21.11672,17.184822,15.038361,14.815181,14.680616,13.036308,13.3251295,12.435693,10.486155,10.811078,8.976411,9.199591,8.756514,7.5585647,8.155898,12.668719,12.724514,8.67118,3.95159,5.1167183,5.356308,6.121026,6.560821,5.924103,3.5610259,2.5009232,1.9528207,1.6443079,1.4867693,1.5819489,2.1989746,2.5107694,3.757949,5.733744,6.7971287,5.4449234,3.9253337,2.5009232,1.5327181,1.4703591,1.4309745,1.8281027,2.0906668,2.1333334,2.3729234,2.0775387,2.225231,2.425436,2.8455386,4.2371287,4.082872,4.1025643,4.197744,3.9712822,2.7503593,3.2262566,4.1156926,4.70318,4.70318,4.269949,4.1091285,4.2240005,4.6178465,5.402257,6.7938466,7.2927184,6.8397956,5.6352825,4.315898,3.9614363,4.4832826,5.3136415,5.658257,5.2742567,4.4767184,4.6900516,3.9253337,3.7021542,4.210872,4.315898,5.3136415,5.5762057,5.546667,5.2644105,4.3716927,3.501949,3.3509746,4.128821,5.756718,7.8408213,5.428513,4.788513,5.543385,6.4557953,5.428513,6.166975,6.741334,8.195283,8.861539,4.388103,3.5577438,4.2830772,4.598154,3.9647183,3.3017437,2.0775387,1.4703591,1.0305642,0.5481026,0.049230773,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.0,0.006564103,0.009846155,0.006564103,0.0032820515,0.0,0.013128206,0.036102567,0.07548718,0.128,0.20676924,0.21333335,0.24615386,0.24615386,0.22646156,0.27897438,0.35446155,0.34789747,0.36102566,0.4201026,0.4594872,0.380718,0.41025645,0.52512825,0.7318975,1.0535386,2.284308,2.674872,2.6912823,2.7044106,3.0162053,2.6387694,2.8192823,2.7208207,2.353231,2.5698464,3.0687182,3.2361028,3.639795,4.279795,4.601436,4.7983594,5.8223596,7.1089234,7.899898,7.253334,6.803693,6.7117953,6.6625648,6.3967185,5.733744,4.857436,4.9362054,5.428513,6.0324106,6.685539,7.066257,7.2960005,7.712821,8.136206,7.899898,8.776206,8.818872,8.362667,7.8408213,7.788308,7.0498466,6.7577443,6.9120007,7.2927184,7.466667,8.050873,7.8769236,7.5552826,7.3353853,7.1154876,6.9809237,7.1122055,7.1548724,7.181129,7.6996927,8.310155,9.380103,9.882257,9.55077,8.868103,8.539898,8.060719,7.5618467,7.1581545,6.941539,7.565129,7.6077952,7.397744,7.2336416,7.4010262,6.633026,7.1154876,8.027898,8.41518,7.204103,7.6964107,7.0432825,7.4830775,8.513641,6.892308,8.251078,9.833026,11.542975,11.926975,8.165744,8.1755905,6.3474874,4.7950773,4.279795,4.20759,1.6475899,0.6301539,0.4660513,0.6104616,0.6498462,1.1027694,1.2340513,1.332513,1.5064616,1.6804104,1.5360001,1.723077,2.0250258,2.2022567,2.0053334,2.1891284,2.1234872,1.9232821,1.6836925,1.467077,1.4933335,1.3029745,1.3029745,1.5425643,1.7165129,1.8838975,1.9462565,2.0512822,2.1333334,1.9298463,1.910154,2.1858463,2.4320002,2.4713848,2.2908719,2.1267693,1.8510771,1.719795,1.7690258,1.8149745,2.0906668,2.7076926,2.989949,3.0194874,3.639795,3.2229745,3.114667,3.3214362,3.6627696,3.764513,3.56759,3.4330258,3.3214362,3.2098465,3.114667,2.9636924,2.9144619,3.6463592,4.768821,4.8377438,4.342154,4.266667,4.457026,4.7327185,4.8804107,5.0543594,5.6418467,6.226052,6.5312824,6.413129,6.5805135,6.6494365,6.744616,6.820103,6.6560006,6.5050263,6.7610264,7.3550773,7.9950776,8.1755905,8.03118,8.192,8.362667,8.464411,8.635077,9.012513,9.009232,8.438154,7.6110773,7.3353853,7.125334,6.9021544,7.1909747,7.9491286,8.546462,8.887795,8.864821,8.329846,7.581539,7.3780518,6.803693,6.4722056,6.4000006,6.5247183,6.692103,7.1844106,7.5618467,8.080411,8.704,9.078155,9.019077,8.3823595,8.004924,7.893334,7.256616,5.786257,5.737026,5.7468724,5.32677,4.886975,4.4996924,3.945026,3.3017437,2.6420515,2.0545642,1.5031796,1.4178462,1.5721027,1.7033848,1.5392822,1.401436,1.404718,1.4112822,1.4244103,1.5885129,1.522872,1.5885129,1.782154,2.0184617,2.1300514,2.3335385,2.7634873,3.0982566,3.3280003,3.7284105,3.6168208,3.5413337,3.8367183,4.3749747,4.5587697,3.895795,3.6758976,3.6791797,3.8432825,4.279795,4.667077,4.923077,5.2545643,5.8486156,6.872616,7.8637953,8.723693,9.472001,9.91836,9.691898,8.766359,7.8834877,7.240206,7.1089234,7.830975,8.385642,8.818872,9.488411,10.315488,10.765129,10.161232,9.048616,8.769642,9.435898,9.95118,8.651488,8.119796,8.008205,7.9950776,7.781744,2.0742567,2.0939488,2.1431797,2.172718,2.1267693,1.9364104,2.2547693,2.4943593,2.809436,3.2229745,3.623385,3.2886157,3.2361028,3.2820516,3.4231799,3.8531284,4.1485133,4.4996924,4.535795,4.342154,4.457026,5.287385,6.186667,6.744616,7.1876926,8.36595,8.064001,8.14277,7.9917955,7.7718983,8.425026,8.999385,11.017847,14.575591,19.127796,23.48636,28.150156,26.41395,25.783796,30.693747,42.509132,40.868107,28.711388,16.28554,8.828718,6.5805135,5.074052,3.7710772,2.7700515,2.097231,1.7296412,1.585231,1.4276924,1.3128207,1.1946667,0.9485129,0.9878975,1.1290257,1.2603078,1.2865642,1.1093334,0.8960001,0.702359,0.60389745,0.636718,0.7975385,1.0962052,1.1913847,1.0108719,0.7187693,0.702359,0.82379496,0.83035904,0.7187693,0.56451285,0.48574364,0.571077,0.4135385,0.33805132,0.36102566,0.17723078,0.44964105,0.8041026,1.3915899,2.1792822,2.9472823,2.9636924,2.1891284,1.1946667,0.41025645,0.12143591,0.098461546,0.1148718,0.13784617,0.16410258,0.19364104,0.42338464,0.9321026,1.6902566,2.3302567,2.1366155,1.270154,1.1060513,1.1257436,1.0732309,0.96492314,0.9714873,1.0699488,1.1224617,1.1355898,1.2570257,2.2613335,3.05559,3.4067695,3.442872,3.6627696,3.5938463,3.2328207,3.5446157,4.276513,3.9680004,5.07077,5.1922054,5.35959,6.2588725,8.247795,8.480822,9.035488,9.645949,9.777231,8.625232,10.390975,10.262975,10.322052,11.382154,12.983796,14.336001,15.100719,15.497848,15.376411,14.234258,12.225642,12.005745,11.762873,11.185231,11.474052,11.008,10.171078,10.217027,10.9915905,10.955488,10.94236,11.513436,11.930258,11.884309,11.500309,14.03077,15.484719,16.640001,17.394873,16.75159,16.646564,17.552412,17.959387,17.106052,14.979283,14.897232,14.575591,13.699283,12.616206,12.340514,12.196103,12.609642,13.718975,14.844719,14.470565,14.788924,14.7331295,14.831591,15.350155,16.292105,15.970463,14.503386,13.558155,13.53518,13.590976,14.027489,14.54277,14.683899,14.490257,14.506668,13.860104,13.082257,12.859077,13.24636,13.686155,13.909334,13.90277,13.472821,12.635899,11.621744,11.201642,12.160001,13.817437,14.769232,12.875488,10.535385,10.203898,10.197334,9.833026,9.432616,9.714872,10.9456415,11.687386,11.684103,11.867898,12.153437,11.608616,11.034257,10.660104,10.134975,9.90195,10.328616,11.07036,11.52,10.794667,12.340514,14.352411,15.763694,16.377438,16.896002,15.136822,12.895181,11.024411,10.066052,10.272821,11.218052,10.7848215,11.109744,12.580104,13.814155,14.073437,12.842668,11.670976,11.1064625,10.706052,11.145847,12.685129,13.430155,13.433437,14.697027,15.753847,15.90154,16.20349,16.840206,17.129026,19.977848,19.99754,18.582975,17.28,17.811693,16.817232,14.7561035,13.243078,12.78359,12.800001,16.521847,20.67036,23.798155,24.431591,21.093744,29.732105,63.993443,79.23529,62.221134,31.130259,25.022362,18.947283,15.136822,14.224411,15.241847,13.640206,13.846975,13.35795,11.405129,8.940309,8.211693,8.503796,8.155898,7.0859494,6.7938466,10.154668,12.041847,9.163487,3.6758976,3.190154,4.059898,5.684513,6.3376417,5.687795,4.818052,3.1967182,2.2678976,1.9954873,2.034872,1.7526156,2.4516926,3.0096412,3.6496413,4.6933336,6.5706673,5.835488,4.381539,2.6256413,1.214359,1.024,1.1257436,1.5458462,1.6902566,1.5195899,1.5425643,1.3259488,1.2898463,1.3029745,1.5097437,2.3138463,3.2098465,3.8006158,3.8564105,3.2787695,2.097231,2.5665643,3.5741541,4.342154,4.5587697,4.378257,4.096,4.9329233,6.0980515,7.1548724,8.021334,7.200821,6.491898,5.5926156,4.7983594,5.0182567,5.349744,5.536821,5.61559,5.4449234,4.7327185,6.245744,6.0291286,5.5269747,5.2578464,4.821334,4.824616,6.698667,7.8834877,7.2270775,4.9854364,3.2295387,2.7503593,3.5807183,5.113436,6.1013336,4.1813335,3.508513,4.201026,5.3366156,4.95918,5.139693,5.9634876,7.6077952,8.4512825,5.097026,4.269949,4.8640003,4.7458467,3.6824617,3.3214362,1.6180514,0.9714873,0.65641034,0.3249231,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.02297436,0.029538464,0.029538464,0.01969231,0.009846155,0.0,0.006564103,0.013128206,0.032820515,0.06564103,0.108307704,0.15753847,0.17723078,0.22646156,0.24287182,0.23302566,0.28882053,0.3314872,0.3249231,0.38728207,0.508718,0.5284103,0.45292312,0.4135385,0.49887183,0.7384616,1.1093334,2.556718,2.6617439,2.6486156,2.8553848,2.7602053,2.5435898,2.6912823,2.6026669,2.3794873,2.8192823,3.0720003,3.2656412,3.826872,4.644103,5.0543594,5.0018463,5.4416413,6.193231,6.8299494,6.6428723,6.4689236,6.491898,6.432821,6.193231,5.85518,5.0904617,5.221744,5.733744,6.2916927,6.764308,7.1187696,7.2369237,7.584821,8.096821,8.155898,8.841846,9.032206,8.477539,7.5913854,7.453539,7.0498466,6.8463597,7.1023593,7.522462,7.24677,7.6996927,7.650462,7.509334,7.4240007,7.256616,7.0531287,6.99077,7.1089234,7.322257,7.4371285,7.857231,8.763078,9.143796,8.838565,8.539898,8.28718,7.568411,6.806975,6.419693,6.813539,6.9349747,7.069539,7.030154,6.892308,6.99077,6.564103,7.076103,8.096821,8.815591,8.027898,8.086975,6.948103,6.521436,6.997334,6.8693337,8.369231,8.887795,9.954462,10.568206,7.177847,7.0104623,5.6287184,4.6178465,3.9253337,1.8576412,1.2898463,0.7220513,0.48902568,0.6268718,0.88287187,1.1585642,1.2865642,1.4080001,1.5031796,1.4080001,1.4572309,1.7099489,2.0578463,2.2350771,1.8281027,2.1366155,2.166154,2.0808206,1.9987694,1.9922053,1.7788719,1.4769232,1.3653334,1.467077,1.5655385,2.048,2.1792822,2.1989746,2.156308,1.9167181,2.0841026,2.231795,2.3696413,2.428718,2.2613335,2.103795,1.8543591,1.6377437,1.5655385,1.7558975,1.9298463,2.6157951,3.0687182,3.1803079,3.495385,3.2328207,3.259077,3.515077,3.754667,3.5446157,3.436308,3.3444104,3.2951798,3.2295387,2.993231,2.8160002,3.0358977,3.9351797,4.900103,4.4406157,4.4077954,4.3585644,4.493129,4.788513,4.9788723,5.2480006,5.805949,6.2884107,6.488616,6.3376417,6.2523084,6.311385,6.7610264,7.3386674,7.273026,6.626462,6.47877,6.931693,7.653744,7.8834877,8.070564,8.352821,8.4972315,8.585847,8.996103,9.114257,8.841846,8.395488,7.9819493,7.788308,7.6176414,7.059693,6.9809237,7.6931286,8.953437,9.399796,9.875693,9.659078,8.848411,8.362667,7.8408213,7.4108725,7.3091288,7.4075904,7.204103,7.565129,7.955693,8.155898,8.195283,8.339693,8.523488,8.119796,7.857231,7.6996927,6.8496413,5.861744,5.924103,6.0652313,5.8912826,5.5565133,4.962462,4.457026,3.7809234,2.9571285,2.284308,1.8313848,1.7263591,1.8773335,2.0808206,2.0086155,1.529436,1.3981539,1.4441026,1.5491283,1.6344616,1.3817437,1.4375386,1.7099489,2.0808206,2.422154,2.3827693,2.7503593,3.1277952,3.4100516,3.7842054,3.6627696,3.626667,3.9417439,4.391385,4.2962055,3.8564105,3.7316926,3.817026,4.1911798,5.113436,5.10359,5.0477953,5.32677,6.0750775,7.1909747,8.113232,8.802463,9.321027,9.6065645,9.4916935,9.097847,8.2215395,7.6570263,7.6734366,8.050873,8.487385,8.756514,9.301334,10.079181,10.564924,9.4457445,8.470975,8.211693,8.710565,9.468719,8.503796,8.136206,8.152616,8.188719,7.752206,2.5665643,2.4976413,2.5337439,2.5042052,2.3696413,2.1858463,2.3171284,2.537026,2.930872,3.4724104,4.013949,3.570872,3.5774362,3.5807183,3.5741541,3.9876926,4.2994876,4.578462,4.6211286,4.5587697,4.850872,5.5269747,6.0717955,6.439385,6.803693,7.5487185,7.7981544,7.9294367,7.8506675,7.817847,8.4283085,8.507077,10.197334,14.011078,19.872822,27.122873,30.897234,28.205952,29.745234,38.048824,47.481438,36.709747,21.507284,11.050668,7.6635904,6.8233852,5.093744,3.7021542,2.6912823,2.048,1.7033848,1.5097437,1.4539489,1.4375386,1.3784616,1.2242053,1.2373334,1.2931283,1.204513,1.0371283,1.1323078,0.8598975,0.7122052,0.65969235,0.6859488,0.76800007,1.1684103,1.2832822,1.148718,0.90584624,0.80738467,0.92225647,0.9878975,0.8992821,0.71548724,0.6826667,0.8730257,0.67610264,0.4397949,0.36430773,0.46933338,1.024,1.7165129,2.3466668,2.7864618,2.9801028,2.9997952,2.2350771,1.2570257,0.48246157,0.15753847,0.16738462,0.29210258,0.3511795,0.30851284,0.28225642,0.47261542,0.86974365,1.7624617,2.789744,2.9505644,1.9954873,1.595077,1.6935385,2.044718,2.2022567,2.0020514,2.100513,2.3466668,2.5764105,2.609231,2.8521028,4.1583595,4.9887185,4.850872,4.3027697,4.594872,3.7349746,3.4198978,3.882667,3.882667,3.620103,3.7349746,4.194462,4.9526157,5.943795,6.1013336,6.47877,6.747898,6.8627696,7.056411,8.592411,8.845129,8.996103,9.540924,10.262975,12.908309,13.820719,13.764924,13.436719,13.449847,11.96636,10.850462,9.849437,9.189744,9.603283,9.780514,10.361437,11.319796,11.969642,10.962052,11.385437,11.74318,12.032001,12.33395,12.803283,14.55918,14.923489,15.376411,16.210052,16.518566,18.051283,17.841232,17.542566,17.270155,15.616001,15.130258,13.689437,12.196103,11.35918,11.67754,11.621744,12.806565,13.794462,13.804309,12.714667,13.46954,13.774771,14.506668,15.698052,16.55795,16.452925,14.815181,13.853539,14.083283,14.306462,14.34913,14.181745,14.575591,15.258258,14.890668,13.853539,12.763899,12.245335,12.47836,13.200411,13.656616,13.909334,13.814155,13.302155,12.373334,11.497026,12.288001,13.682873,14.421334,13.075693,10.538668,10.102155,9.800206,9.189744,9.353847,8.874667,9.816616,10.752001,11.34277,12.337232,13.53518,12.859077,12.087796,12.005745,12.402873,11.992617,11.825232,12.209231,12.937847,13.289026,14.588719,15.425642,15.625848,15.563488,16.15754,15.015386,13.210258,11.444513,10.276103,10.144821,11.034257,10.902975,11.533129,13.15118,14.437745,15.00554,13.961847,12.557129,11.52,11.047385,11.444513,12.875488,13.298873,13.252924,15.829334,16.935387,16.610462,15.563488,14.70359,15.136822,17.066668,18.914463,18.976822,17.736206,17.83795,16.420103,15.159796,13.879796,13.088821,13.988104,17.942976,21.815796,24.293745,24.786053,23.424002,35.99426,78.785645,101.169235,83.74811,38.3639,30.030771,22.14072,17.184822,16.088617,18.202257,15.80636,13.968411,13.344822,12.547283,8.149334,7.821129,8.162462,7.7292314,6.547693,6.11118,6.9152827,8.155898,6.954667,4.023795,3.6758976,3.245949,4.309334,5.156103,5.2447186,5.1987696,3.5478978,2.3991797,2.2153847,2.605949,2.3204105,2.4681027,3.239385,3.8465643,4.2994876,5.3924108,5.3431797,4.6769233,3.1376412,1.3095386,0.63343596,0.6826667,0.97805136,1.3784616,1.5753847,1.0994873,0.88287187,0.90256417,1.0633847,1.4441026,2.3204105,3.8071797,4.2962055,3.5314875,2.3105643,2.4648206,2.3958976,2.7602053,3.6168208,4.493129,4.3618464,4.9920006,6.445949,7.643898,7.860513,6.744616,5.9470773,4.9460516,4.279795,4.4898467,6.11118,6.0619493,5.8453336,5.5269747,5.353026,5.717334,8.064001,8.871386,8.310155,6.8955903,5.4875903,4.8738465,7.7357955,9.481847,8.608821,6.705231,4.4734364,3.9286156,4.7360005,5.901129,5.7435904,5.3103595,5.1265645,5.3694363,5.5630774,4.5817437,5.2512827,4.7655387,4.9493337,5.7632823,5.3136415,5.5597954,5.3398976,4.571898,3.6102567,3.2328207,1.1979488,0.6170257,0.39384618,0.108307704,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.01969231,0.052512825,0.12471796,0.10502565,0.06564103,0.026256412,0.006564103,0.013128206,0.013128206,0.032820515,0.052512825,0.072205134,0.108307704,0.108307704,0.15753847,0.21333335,0.25271797,0.27569234,0.26256412,0.2986667,0.39712822,0.48574364,0.41025645,0.47589746,0.53825647,0.65312827,0.8533334,1.1224617,2.609231,2.8225644,2.809436,2.868513,2.546872,2.4320002,2.5731285,2.5173335,2.3991797,2.92759,2.8980515,3.4888208,4.44718,5.32677,5.4843082,5.097026,5.0576415,5.536821,6.157129,5.9995904,5.8912826,6.23918,6.2818465,5.9470773,5.861744,5.5696416,5.579488,5.9963083,6.5706673,6.692103,7.207385,7.1548724,7.269744,7.6701546,7.860513,8.408616,9.002667,8.562873,7.387898,7.1581545,7.3025646,7.030154,7.1614366,7.6110773,7.384616,7.4207187,7.5454364,7.512616,7.282872,7.017026,7.076103,7.200821,7.312411,7.3386674,7.1844106,7.171283,7.1187696,7.322257,7.752206,8.054154,7.680001,6.918565,6.183385,6.0258465,7.125334,6.6034875,6.7544622,6.7774363,6.5706673,6.7216415,6.47877,6.9809237,8.034462,8.897642,8.260923,6.744616,6.5936418,7.177847,7.680001,7.0990777,7.4141545,5.8518977,5.330052,6.2720003,6.6100516,7.463385,6.5247183,5.21518,3.882667,1.8018463,1.3554872,0.67282057,0.37415388,0.63343596,1.1946667,1.214359,1.2635899,1.3784616,1.4736412,1.3292309,1.467077,1.7985642,2.1103592,2.172718,1.7526156,2.2121027,2.2022567,2.0611284,2.048,2.3401027,1.9003079,1.6016412,1.3915899,1.2898463,1.3883078,2.225231,2.3893335,2.3269746,2.231795,2.0118976,2.2153847,2.162872,2.1300514,2.225231,2.359795,1.9692309,1.8346668,1.8149745,1.8904617,2.15959,2.297436,2.6322052,2.858667,2.8947694,2.8914874,2.9078977,3.1803079,3.511795,3.6529233,3.318154,3.5971284,3.4822567,3.387077,3.3378465,2.986667,2.9997952,3.511795,4.332308,4.9788723,4.6802053,4.844308,4.601436,4.5095387,4.709744,4.893539,5.681231,6.0750775,6.308103,6.439385,6.3474874,6.1472826,6.3245134,7.0367184,7.7981544,7.4863596,6.8988724,6.626462,6.87918,7.460103,7.77518,8.349539,8.772923,8.996103,9.170052,9.639385,9.449026,8.828718,8.461129,8.467693,8.39877,7.939283,7.3649235,6.9743595,7.273026,8.966565,9.590155,10.161232,10.06277,9.3768215,8.910769,8.470975,8.090257,8.129642,8.4512825,8.4053335,8.320001,8.477539,8.342975,7.9163084,7.752206,8.201847,8.01477,7.680001,7.2664623,6.416411,6.5739493,6.701949,6.73477,6.636308,6.4000006,5.5072823,5.169231,4.634257,3.748103,2.9440002,2.3401027,2.0775387,2.15959,2.4484105,2.674872,1.8215386,1.4834872,1.6311796,1.9429746,1.8018463,1.4375386,1.3784616,1.6804104,2.2482052,2.8324106,2.4648206,2.737231,3.2131286,3.6004105,3.7448208,3.570872,3.56759,3.7776413,4.0434875,4.007385,3.8006158,3.6168208,3.754667,4.4012313,5.6287184,5.2414365,5.0609236,5.4416413,6.4000006,7.5913854,8.65477,9.110975,9.238976,9.235693,9.235693,9.225847,8.218257,7.6668725,7.906462,8.162462,8.303591,8.375795,8.730257,9.43918,10.269539,8.825437,7.9950776,7.8145647,8.198565,8.956718,8.41518,8.293744,8.395488,8.434873,8.04759,2.7011285,2.4582565,2.2121027,2.176,2.294154,2.2580514,2.2350771,2.612513,3.2164104,3.95159,4.8049235,4.4045134,4.1189747,3.8695388,3.8531284,4.562052,4.709744,4.7917953,4.6145644,4.3651285,4.6080003,4.9985647,5.297231,5.799385,6.3901544,6.560821,6.7807183,7.50277,7.7981544,7.64718,7.965539,8.257642,10.243283,13.906053,19.51836,27.648003,30.25067,30.998978,35.52821,42.23344,42.28267,27.181952,14.444309,8.060719,7.056411,5.4941545,3.9318976,3.2098465,2.6190772,1.9954873,1.7394873,1.654154,1.6311796,1.4933335,1.2832822,1.2964103,1.2603078,1.270154,1.2077949,1.1323078,1.2668719,0.79097444,0.77128214,0.90584624,0.9156924,0.5481026,1.0732309,1.214359,1.3489232,1.4441026,1.0535386,1.1257436,0.9419488,0.73517954,0.5973334,0.48902568,0.36758977,0.45620516,0.508718,0.64000005,1.3128207,2.0808206,2.6223593,2.9440002,3.0260515,2.806154,2.477949,1.7624617,0.95835906,0.32820517,0.12143591,0.108307704,0.39056414,0.6170257,0.67282057,0.67282057,0.93866676,1.1454359,1.6738462,2.487795,3.0982566,2.231795,1.8215386,2.048,2.9604106,4.4865646,5.2414365,5.989744,6.5083084,6.7577443,6.882462,6.038975,6.4590774,6.931693,6.6822567,5.402257,5.792821,3.9942567,3.1540515,3.7710772,3.7218463,1.9298463,2.048,2.176,2.038154,2.989949,3.2853336,3.7973337,5.3398976,7.1548724,6.8955903,6.23918,6.1013336,6.449231,7.466667,9.567181,10.886565,11.250873,11.1983595,10.873437,10.056206,9.238976,8.418462,8.260923,8.579283,8.346257,9.275078,10.870154,11.713642,11.707078,12.084514,11.864616,11.050668,11.398565,12.803283,13.289026,13.22995,13.105232,13.88636,15.67836,17.716515,18.008617,17.385027,17.007591,16.836924,15.638975,13.35795,12.668719,12.363488,12.248616,13.154463,13.810873,14.726565,15.002257,14.250668,12.603078,12.763899,13.3251295,14.27036,15.094155,14.8020525,16.032822,14.391796,13.420309,13.915898,13.915898,12.672001,13.174155,14.63795,15.609437,13.961847,13.948719,13.899488,13.4859495,12.868924,12.711386,13.443283,14.165335,14.03077,13.243078,13.046155,12.117334,12.95754,13.843694,13.820719,12.711386,11.1983595,10.535385,9.931488,9.268514,9.110975,8.815591,9.035488,10.072617,12.228924,15.793232,15.474873,13.994668,12.36677,11.720206,13.305437,13.745232,13.131488,13.459693,14.634667,14.450873,16.987898,17.24718,16.246155,15.097437,14.998976,14.792206,13.971693,12.360206,10.545232,9.888822,10.131693,10.925949,12.317539,14.060308,15.609437,16.597334,15.333745,14.152206,13.377642,11.352616,10.266257,10.341744,10.732308,11.946668,15.852309,17.769028,17.83795,16.196924,14.477129,15.809642,15.064616,16.085335,17.135592,17.398155,16.984617,16.482462,16.705643,16.406975,15.783386,16.479181,21.06749,23.7719,24.835283,24.976412,25.38995,36.877132,83.49211,116.30606,106.39098,44.84595,36.141953,26.899694,20.97231,19.27877,19.790771,17.811693,17.05354,15.107284,11.529847,7.8441033,8.356103,7.604513,6.9021544,6.5903597,6.0258465,5.356308,6.4689236,6.4623594,5.152821,5.080616,4.630975,4.4077954,4.8344617,5.356308,4.4406157,2.8291285,2.1891284,2.176,2.4910772,2.868513,1.9528207,2.0644104,3.2229745,4.5390773,4.197744,3.9023592,4.076308,3.3575387,1.7460514,0.6104616,0.65969235,0.7253334,1.014154,1.2340513,0.6104616,0.65969235,0.48902568,1.2077949,2.6354873,3.2951798,5.5171285,5.989744,4.9788723,3.3575387,2.6256413,2.7700515,2.5796926,2.6715899,3.3969233,4.8377438,5.546667,5.07077,4.778667,4.841026,4.2436924,4.5095387,3.3411283,2.6715899,3.2295387,4.5456414,4.9493337,4.9329233,4.71959,4.8640003,6.2555904,6.3179493,6.99077,7.8473854,8.0377445,6.3179493,5.0609236,5.421949,5.412103,4.9362054,5.8125134,6.961231,7.716103,7.2205133,5.6943593,4.4242053,6.2063594,6.678975,6.5772314,6.0225644,4.532513,6.669129,4.4832826,2.048,1.7985642,4.532513,6.1078978,5.0182567,4.0402055,4.013949,3.8301542,1.3751796,0.43323082,0.128,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01969231,0.101743594,0.32164106,0.32164106,0.2100513,0.0951795,0.02297436,0.0,0.013128206,0.032820515,0.032820515,0.02297436,0.04594872,0.0951795,0.098461546,0.108307704,0.15097436,0.21333335,0.24943592,0.3052308,0.33476925,0.33476925,0.33476925,0.48246157,0.6662565,0.83035904,0.9517949,1.0371283,2.7109745,3.3936412,3.3017437,2.8291285,2.546872,2.2055387,2.5698464,2.6683078,2.4385643,2.7306669,2.7798977,3.7710772,4.8836927,5.47118,5.080616,5.044513,5.668103,6.301539,6.452513,5.7665644,6.11118,6.892308,6.806975,5.874872,5.4482055,5.546667,5.6254363,6.3212314,7.4863596,8.195283,8.326565,8.113232,8.12636,8.129642,7.0793853,6.7872825,7.75877,8.021334,7.269744,6.8660517,6.987488,6.3967185,6.1341543,6.49518,7.020308,7.581539,8.01477,7.9294367,7.4436927,7.1876926,6.6133337,6.8266673,6.806975,6.439385,6.5017443,6.340924,6.229334,6.370462,6.73477,7.066257,7.4929237,7.0400004,6.294975,6.052103,7.3091288,6.0652313,6.0652313,6.2785645,6.245744,6.088206,6.2851286,7.128616,7.7948723,8.139488,8.713847,4.598154,4.522667,6.1472826,8.01477,9.55077,9.760821,7.762052,5.717334,4.6572313,4.4865646,5.0838976,4.57518,3.9154875,3.6102567,3.7087183,3.1343591,1.3062565,0.26912823,0.49887183,0.8992821,0.9616411,0.9682052,1.0272821,1.1224617,1.0994873,1.4408206,1.7263591,1.9659488,2.044718,1.7394873,2.28759,2.2711797,1.9790771,1.7788719,2.1202054,1.7657437,1.6246156,1.4112822,1.2800001,1.8149745,2.1956925,2.2711797,2.2646155,2.2678976,2.2416413,2.487795,2.4943593,2.3401027,2.1530259,2.0906668,2.1530259,2.156308,2.0841026,1.9396925,1.7690258,2.4549747,2.3696413,2.4713848,2.9144619,3.0358977,3.0227695,3.0129232,3.1277952,3.3050258,3.2820516,3.6463592,3.5905645,3.4822567,3.3772311,3.0358977,3.1967182,4.059898,4.571898,4.670359,5.280821,4.8771286,4.59159,4.3684106,4.2962055,4.637539,5.6385646,6.1013336,6.173539,6.091488,6.163693,6.091488,6.695385,7.2992826,7.3747697,6.547693,7.131898,7.1220517,7.3058467,7.88677,8.484103,9.107693,9.517949,9.764103,9.980719,10.420513,9.764103,9.140513,8.792616,8.704,8.605539,7.8736415,7.0400004,6.308103,6.1472826,7.2927184,9.330873,9.475283,9.268514,9.42277,9.826463,9.242257,8.326565,8.185436,8.953437,9.796924,9.5146675,9.353847,9.042052,8.457847,7.6307697,7.6898465,8.064001,7.9524107,7.2369237,6.4557953,7.430565,7.3452315,7.315693,7.571693,7.460103,6.4590774,6.117744,5.330052,4.240411,4.2272825,2.665026,2.1989746,2.2186668,2.4188719,2.8225644,2.4549747,1.8445129,1.9035898,2.3729234,1.8018463,1.654154,1.5064616,1.7690258,2.4418464,3.1113849,2.6486156,2.917744,3.4921029,3.9647183,3.95159,3.7185643,3.892513,3.9647183,3.8367183,3.8006158,3.6529233,3.6069746,3.7349746,4.1878977,5.1889234,5.211898,5.4941545,6.0356927,6.8955903,8.178872,9.67877,10.092308,10.14154,10.151385,10.039796,8.868103,7.138462,6.5050263,7.138462,7.7357955,8.247795,8.2215395,8.441437,9.242257,10.512411,9.206155,8.323282,8.169026,8.480822,8.408616,7.748924,7.9130263,8.339693,8.546462,8.132924,2.6157951,2.6256413,2.4451284,2.3204105,2.3072822,2.2711797,2.3630772,2.5961027,3.0030773,3.5577438,4.1485133,4.4964104,4.240411,4.073026,4.325744,4.965744,4.5456414,4.4800005,4.5554876,4.565334,4.2896414,4.896821,5.402257,5.9667697,6.304821,5.6943593,5.8157954,6.229334,6.416411,6.377026,6.6461544,7.1548724,9.517949,13.856822,20.804924,31.494566,31.701336,33.368618,39.11549,44.514465,38.1079,20.43077,11.398565,7.9228725,6.9152827,5.284103,3.5380516,2.7864618,2.3072822,1.8937438,1.8609232,1.7362052,1.522872,1.3620514,1.3128207,1.332513,1.394872,1.404718,2.1792822,3.1442053,2.3401027,1.3357949,0.9616411,0.9485129,1.1585642,1.5753847,1.3883078,1.2471796,1.1749744,1.1323078,1.017436,1.020718,0.827077,0.7187693,0.7384616,0.69579494,0.7187693,0.7581539,1.0666667,1.6738462,2.3729234,3.3378465,3.5478978,3.6004105,3.7251284,3.761231,2.5993848,1.3423591,0.4955898,0.17394873,0.072205134,0.06235898,0.29210258,0.5349744,0.6629744,0.63343596,0.86317956,1.214359,1.4933335,1.9003079,2.986667,3.4691284,3.4855387,4.2994876,6.009436,7.525744,9.337437,11.907283,14.418053,16.449642,17.975796,17.184822,15.55036,13.61395,11.661129,9.734565,8.815591,7.4765134,6.439385,5.664821,4.3585644,3.3936412,3.3772311,3.826872,4.1156926,3.4658465,3.8662567,4.818052,5.720616,6.1997952,6.091488,6.0685134,6.0750775,6.62318,7.4469748,7.515898,8.356103,10.213744,10.7848215,10.085744,10.469745,9.974154,8.681026,8.54318,9.268514,8.333129,9.865847,11.073642,11.648001,11.861334,12.560411,13.590976,13.771488,12.980514,11.96636,12.337232,13.039591,13.6237955,14.851283,16.584206,17.811693,17.54913,17.227488,17.552412,18.153027,17.58195,15.00554,14.102976,13.755078,13.456411,13.3251295,13.699283,14.697027,15.241847,14.772514,13.249642,13.945437,14.592001,15.074463,14.982565,13.604104,14.388514,13.99795,13.338258,13.059283,13.538463,13.610668,13.6008215,13.929027,14.598565,15.205745,13.778052,13.236514,12.868924,12.652308,13.236514,13.702565,14.089848,13.804309,13.036308,12.754052,12.655591,12.685129,12.632616,12.626052,13.138052,12.885334,12.36677,12.091078,11.628308,9.632821,9.6065645,9.83959,10.456616,11.953232,15.195899,16.331488,15.287796,14.122667,13.784616,14.112822,14.112822,14.355694,14.683899,14.946463,14.998976,16.44636,16.180513,15.1466675,14.257232,14.41477,14.342566,14.641232,14.145642,12.780309,11.536411,11.398565,11.746463,12.868924,14.677335,16.695797,17.411283,15.704617,13.833847,12.36677,10.194052,10.082462,9.787078,9.655796,10.509129,13.643488,15.287796,16.8599,17.043694,16.502155,17.870771,18.395899,19.222977,19.344412,18.720821,18.277744,18.38277,18.12677,17.88718,18.448412,21.008411,27.346054,29.029745,27.871181,26.246567,27.0999,35.245953,70.51816,106.9555,113.624626,54.63631,41.9479,33.81826,27.369028,22.147284,20.132105,20.079592,18.011898,14.49354,10.709334,8.477539,7.768616,7.7981544,7.177847,6.2162056,6.892308,4.962462,5.8420515,6.2752824,5.077334,3.1277952,2.5206156,3.6660516,5.8945646,7.0957956,3.7185643,2.8816411,2.4681027,2.5600002,3.2656412,4.7360005,4.5423594,3.6693337,3.7218463,4.5128207,4.073026,3.7710772,3.0720003,2.2580514,1.4605129,0.6465641,0.48246157,0.4004103,0.43323082,0.51856416,0.512,1.5097437,1.0765129,0.77128214,1.1782565,1.9167181,2.8192823,3.2787695,2.6453335,1.404718,1.1585642,1.5589745,1.7099489,2.2908719,3.620103,5.668103,5.7698464,6.2818465,6.416411,5.8420515,4.6572313,4.279795,3.9253337,3.5413337,3.5249233,4.706462,6.232616,6.2096415,6.009436,6.2227697,6.6461544,5.917539,5.398975,5.07077,4.900103,4.841026,4.1091285,3.367385,3.0851285,3.9253337,6.7183595,11.136001,10.538668,8.569437,6.49518,3.2032824,4.2535386,5.504,6.557539,7.131898,7.059693,6.636308,4.713026,3.242667,2.8947694,3.0424619,3.2886157,2.3204105,1.719795,1.9561027,2.3893335,2.231795,0.9321026,0.055794876,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.118153855,0.45620516,0.48246157,0.36102566,0.19364104,0.06564103,0.013128206,0.02297436,0.029538464,0.036102567,0.04266667,0.059076928,0.08861539,0.09189744,0.108307704,0.14112821,0.15097436,0.17066668,0.21333335,0.27241027,0.3511795,0.45620516,0.56451285,0.6662565,0.7581539,0.9747693,1.5885129,3.629949,3.4756925,2.9111798,2.681436,2.487795,2.7503593,2.612513,2.4713848,2.5928206,3.1081028,3.4724104,3.948308,4.6145644,5.2315903,5.2414365,5.3103595,5.602462,5.937231,6.2851286,6.744616,6.3540516,7.0334363,7.213949,6.6461544,6.373744,5.8486156,5.792821,6.6560006,8.034462,8.694155,7.9294367,7.778462,7.962257,8.093539,7.6767187,7.131898,7.936001,8.546462,8.349539,7.683283,6.5280004,5.8190775,5.5138464,5.7009234,6.616616,7.5881033,7.712821,7.427283,7.131898,7.197539,7.026872,6.5936418,6.124308,5.8092313,5.792821,5.9963083,5.8125134,5.786257,6.038975,6.2720003,7.1581545,7.026872,6.445949,6.0192823,6.370462,6.3934364,6.314667,6.0356927,5.805949,6.2227697,6.301539,6.619898,9.084719,11.32636,6.675693,4.9329233,3.31159,2.6157951,3.4625645,6.2818465,6.6527185,6.564103,6.550975,6.11118,3.7054362,3.629949,2.9571285,2.7963078,3.2525132,3.4264617,3.6824617,1.9954873,0.73517954,0.69907695,1.1191796,0.8992821,1.4408206,1.6475899,1.3193847,1.148718,1.1979488,1.3817437,1.6246156,1.785436,1.6672822,1.9331284,1.9298463,1.785436,1.7329233,2.1333334,1.7788719,1.6443079,1.5753847,1.595077,1.8773335,2.3040001,2.2383592,2.0676925,2.038154,2.2678976,2.4320002,2.5238976,2.550154,2.5304618,2.4681027,2.5206156,2.4713848,2.3762052,2.3072822,2.3794873,2.809436,2.8225644,2.740513,2.6453335,2.3762052,2.9604106,2.7470772,2.8291285,3.446154,3.9876926,3.817026,3.5347695,3.3247182,3.2984617,3.4625645,3.7776413,4.0008206,4.1747694,4.460308,5.110154,5.0871797,4.7458467,4.4800005,4.562052,5.1265645,5.4449234,5.346462,5.3760004,5.681231,6.0192823,5.9930263,6.186667,6.439385,6.7544622,7.3025646,8.054154,7.9261546,7.9097443,8.162462,8.008205,8.454565,9.225847,10.056206,10.683078,10.850462,9.701744,9.258667,9.156924,9.248821,9.5835905,9.366975,9.170052,8.789334,8.2904625,8.01477,9.025641,9.954462,10.157949,9.688616,9.301334,8.470975,8.0377445,8.119796,8.874667,10.466462,10.167795,9.232411,8.549745,8.198565,7.4469748,7.653744,7.785026,7.568411,6.99077,6.294975,7.076103,7.6603084,8.293744,8.832001,8.730257,7.4174366,7.0400004,6.308103,5.4482055,6.229334,4.3716927,2.8389745,2.2777438,2.553436,2.7602053,2.5895386,2.2547693,2.0250258,1.9626669,1.8970258,1.654154,2.1267693,2.7175386,3.121231,3.3312824,3.0818465,3.3772311,3.8432825,4.1550775,4.023795,4.2929235,4.4767184,4.384821,4.1911798,4.457026,4.056616,3.8531284,3.826872,4.0369234,4.637539,5.4449234,5.9503593,6.9120007,8.280616,9.193027,9.412924,9.885539,9.875693,9.370257,9.065026,8.917334,7.6767187,6.9349747,6.9021544,6.4065647,7.5421543,8.293744,8.910769,9.53436,10.20718,9.281642,8.667898,8.395488,8.339693,8.237949,8.192,8.277334,8.392206,8.3134365,7.6931286,2.300718,2.3302567,2.3630772,2.284308,2.1858463,2.3827693,2.4188719,2.3762052,2.6190772,3.1671798,3.7087183,4.332308,4.5062566,4.6112823,4.785231,4.9099493,4.7458467,5.097026,5.3760004,5.284103,4.8049235,5.100308,5.5991797,6.2523084,6.5969234,5.7698464,5.861744,6.180103,6.3540516,6.298257,6.189949,6.810257,9.281642,14.844719,22.741335,30.194874,28.199387,32.180515,38.97108,41.941338,30.98585,15.402668,8.920616,6.6494365,5.4383593,3.879385,2.7011285,2.2186668,2.1431797,2.2022567,2.176,2.1792822,2.034872,1.9396925,1.9298463,1.8740515,1.6508719,1.6738462,2.0578463,2.546872,2.537026,2.0512822,1.847795,1.7624617,1.7263591,1.7657437,2.176,2.0841026,1.8248206,1.5327181,1.1257436,0.99774367,0.827077,0.77128214,0.8336411,0.8763078,0.7318975,0.6498462,0.85005134,1.3357949,1.8904617,2.6518977,2.6683078,2.5271797,2.4549747,2.294154,1.5721027,0.761436,0.24287182,0.08533334,0.032820515,0.049230773,0.14769232,0.23958977,0.3511795,0.6071795,1.1191796,1.6705642,1.972513,2.294154,3.4724104,4.466872,4.598154,5.024821,6.048821,7.1220517,9.255385,10.476309,11.592206,12.924719,14.306462,14.923489,14.700309,13.696001,12.3306675,11.385437,11.641437,11.437949,10.532104,8.937026,6.925129,4.9427695,4.273231,4.4865646,4.821334,4.1813335,4.2502565,5.1298466,5.796103,5.924103,5.907693,6.547693,6.163693,6.170257,7.0334363,8.257642,10.390975,11.096616,10.568206,9.665642,9.924924,9.626257,8.835282,9.232411,10.322052,9.429334,10.637129,10.955488,11.546257,12.389745,12.278154,12.681848,12.865642,12.501334,11.956513,12.2847185,12.199386,12.714667,13.692719,15.379693,18.405745,17.906874,18.008617,18.517334,18.838976,17.985641,15.944206,14.464001,13.7386675,13.869949,14.87754,15.123693,15.491283,15.717745,15.281232,13.403898,14.454155,15.271386,15.061335,13.984821,13.177437,13.167591,13.650052,13.824001,13.587693,13.525334,13.489232,13.636924,13.958565,14.634667,16.039387,14.148924,13.367796,12.914873,12.78359,13.74195,13.948719,13.699283,12.895181,11.976206,11.910565,12.137027,12.86236,13.062565,12.754052,12.987078,13.633642,13.384206,13.223386,12.921437,11.047385,10.541949,10.282667,10.213744,10.857026,13.315283,14.831591,14.959591,15.025232,15.415796,15.61272,15.274668,14.946463,14.749539,14.818462,15.300924,16.436514,16.170668,15.379693,15.1466675,16.764719,15.484719,15.816206,15.652103,14.431181,13.11836,13.026463,13.259488,14.135796,15.570052,17.076513,17.322668,15.428925,13.778052,12.872206,11.323078,10.44677,9.173334,8.553026,9.301334,11.818667,13.906053,15.816206,16.39713,16.489027,18.898052,20.079592,21.270975,21.280823,20.292925,19.85313,19.75795,19.643078,20.358566,22.30154,25.416206,31.14667,31.67508,29.705849,28.146873,30.099695,36.58503,57.97744,88.65806,104.8517,64.68267,49.138874,41.40308,34.330257,26.446772,21.930668,21.572926,18.809437,14.864411,11.126155,9.140513,7.532308,7.827693,7.8145647,6.948103,6.340924,7.1187696,6.669129,6.3442054,5.805949,3.0162053,2.2646155,2.9571285,4.44718,5.4482055,4.0336413,3.0227695,2.225231,2.4648206,3.7185643,5.110154,5.32677,4.778667,4.670359,5.10359,5.077334,4.2962055,3.308308,2.546872,1.9528207,0.98461545,0.5907693,0.318359,0.18051283,0.16738462,0.23302566,0.7187693,0.54482055,0.39056414,0.83035904,2.349949,2.9965131,2.9538465,2.3794873,1.6180514,1.1881026,1.2832822,1.3128207,1.8806155,3.245949,5.32677,6.1472826,7.5520005,7.578257,5.986462,4.240411,4.4996924,4.322462,4.017231,4.135385,5.4514875,7.315693,8.52677,7.8506675,6.1374364,6.314667,5.927385,4.9821544,4.7360005,5.097026,4.6080003,4.2502565,3.6890259,3.761231,4.6080003,5.661539,8.730257,8.434873,7.181129,5.976616,4.4373336,4.33559,4.969026,5.477744,5.504,5.1626673,4.972308,4.699898,4.3618464,3.8137438,2.7437952,2.231795,1.6410258,1.4966155,1.7723079,1.8740515,1.2209232,0.43651286,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.013128206,0.12143591,0.48902568,0.4660513,0.52512825,0.43651286,0.20348719,0.06235898,0.04266667,0.04594872,0.068923086,0.10502565,0.12471796,0.12143591,0.12471796,0.12471796,0.118153855,0.118153855,0.14441027,0.22646156,0.3249231,0.41025645,0.47917953,0.5907693,0.67938465,0.83035904,1.2274873,2.162872,3.2000003,2.930872,2.6486156,2.6880002,2.4451284,2.8521028,2.7569232,2.6847181,2.9440002,3.6430771,3.8137438,4.059898,4.7983594,5.681231,5.5991797,5.4186673,5.2709746,5.5171285,6.0783596,6.4590774,6.3376417,6.698667,6.672411,6.2162056,6.0849237,5.6352825,5.671385,6.1440005,6.925129,7.8112826,7.315693,7.0957956,7.13518,7.2369237,7.030154,6.9710774,7.5946674,8.195283,8.14277,6.892308,6.0717955,5.907693,5.9963083,6.3376417,7.328821,8.763078,8.490667,7.906462,7.6274877,7.50277,6.8594875,6.1997952,5.9930263,6.196513,6.245744,6.1440005,5.9930263,6.042257,6.3179493,6.6133337,7.637334,7.204103,6.3442054,5.7468724,5.76,5.609026,5.602462,5.7632823,6.0192823,6.193231,5.9470773,6.7971287,8.277334,8.618668,4.7261543,4.466872,3.623385,3.0030773,3.3312824,5.2611284,5.113436,4.9132314,4.6276927,3.9647183,2.3729234,2.1891284,2.605949,3.314872,4.0434875,4.585026,4.5489235,4.338872,3.4002054,2.048,1.4572309,0.7056411,1.2504616,1.6180514,1.4375386,1.4441026,1.3456411,1.3915899,1.5491283,1.7001027,1.6475899,1.7394873,1.8379488,1.7690258,1.6705642,1.9987694,1.8576412,1.6278975,1.5556924,1.6443079,1.6344616,1.7591796,1.785436,1.7788719,1.8674873,2.228513,2.4188719,2.6551797,2.7470772,2.6912823,2.681436,2.7667694,2.546872,2.5074873,2.7011285,2.7241027,2.8849232,2.7995899,2.678154,2.6486156,2.7437952,3.3444104,3.186872,3.3378465,3.9844105,4.450462,3.7940516,3.3247182,3.1442053,3.2525132,3.5511796,3.636513,3.7382567,3.9942567,4.4307694,4.965744,5.1265645,4.9788723,4.926359,5.2053337,5.87159,5.8289237,5.4974365,5.346462,5.543385,5.943795,6.114462,6.298257,6.498462,6.7610264,7.1909747,7.765334,8.054154,8.162462,8.067283,7.6143594,8.119796,8.87795,9.783795,10.5780525,10.873437,10.049642,9.750975,9.626257,9.626257,10.000411,10.253129,10.243283,9.7903595,9.015796,8.323282,9.005949,9.961026,10.161232,9.521232,8.914052,8.3593855,8.585847,8.989539,9.412924,10.14154,10.187488,9.32759,8.746667,8.549745,7.765334,8.077128,8.228104,8.027898,7.4797955,6.7872825,7.1614366,7.9491286,8.700719,9.107693,9.002667,7.5881033,6.885744,6.23918,5.72718,6.160411,4.7950773,3.2853336,2.5698464,2.7273848,2.9669745,2.6912823,2.4451284,2.1431797,1.8970258,1.9954873,2.034872,2.7569232,3.626667,4.135385,3.8006158,3.31159,3.4888208,3.95159,4.4373336,4.775385,5.077334,5.031385,4.8640003,4.781949,4.962462,4.5128207,3.948308,3.5741541,3.6562054,4.4274874,5.979898,7.0826674,8.39877,9.77395,10.279386,10.210463,10.469745,10.19077,9.452309,9.268514,9.334154,8.385642,7.762052,7.6012316,6.8693337,7.768616,8.185436,8.641642,9.291488,9.938052,9.475283,9.32759,9.032206,8.579283,8.43159,8.454565,8.743385,8.986258,8.897642,8.234667,2.294154,2.1956925,2.2646155,2.2186668,2.166154,2.5961027,2.481231,2.297436,2.4451284,2.92759,3.367385,3.9778464,4.4865646,4.84759,4.9920006,4.8377438,4.9788723,5.431795,5.7665644,5.7698464,5.4547696,5.208616,5.72718,6.4689236,6.774154,5.8880005,6.048821,6.2030773,6.49518,6.8004107,6.7249236,7.4207187,10.70277,17.302977,24.91077,28.179695,24.067284,29.879797,36.358566,35.84985,22.298258,11.477334,7.53559,5.9470773,4.4110775,2.8717952,2.1366155,1.8313848,2.0611284,2.5074873,2.4320002,2.5042052,2.5173335,2.4681027,2.3302567,2.038154,1.6836925,1.5983591,1.5327181,1.5819489,2.169436,2.15959,2.2449234,2.3302567,2.3204105,2.1202054,2.7864618,2.6322052,2.2744617,1.9167181,1.3522053,1.0305642,0.8598975,0.7844103,0.77128214,0.7975385,0.6170257,0.50543594,0.58092314,0.8566154,1.2307693,1.6508719,1.5360001,1.3226668,1.1520001,0.8730257,0.62030774,0.32820517,0.12471796,0.03938462,0.02297436,0.049230773,0.055794876,0.06235898,0.16082053,0.5415385,1.332513,2.0808206,2.5206156,2.8455386,3.7218463,4.8377438,5.0609236,4.962462,5.028103,5.664821,8.257642,8.989539,8.848411,8.615385,8.851693,10.358154,11.382154,11.697231,11.32636,10.555078,10.9686165,11.1064625,10.423796,9.032206,7.6931286,6.6592827,6.1472826,6.183385,6.12759,4.663795,5.1954875,6.370462,6.961231,6.885744,7.213949,7.936001,7.13518,7.253334,8.917334,10.948924,12.225642,11.539693,10.79795,10.614155,10.315488,9.878975,9.344001,9.639385,10.466462,10.30236,10.857026,10.840616,11.565949,12.727796,12.386462,12.258463,12.084514,12.265027,12.672001,12.668719,11.769437,11.897437,13.08554,15.448617,19.157335,18.632206,18.409027,18.638771,18.888206,18.14318,16.603899,14.969437,14.470565,15.432206,17.283283,16.551386,16.193642,16.210052,16.085335,14.769232,15.399385,15.816206,15.16636,13.912617,13.853539,13.778052,14.316309,14.746258,14.7790785,14.588719,14.185027,14.362258,14.76595,15.504412,17.138874,15.209026,14.089848,13.522053,13.436719,13.961847,13.781334,13.1872835,12.248616,11.369026,11.306667,11.451077,12.619488,13.184001,12.875488,12.793437,13.650052,14.057027,14.063591,13.587693,12.425847,11.500309,10.860309,10.253129,10.19077,11.972924,13.751796,14.641232,15.140103,15.579899,16.114874,15.425642,14.769232,14.460719,14.706873,15.619284,16.617027,16.469334,15.980309,16.082052,17.821539,16.771284,17.152,17.03713,15.937642,14.792206,14.500104,14.523078,14.660924,15.081027,16.315079,16.643284,15.793232,14.936617,14.395078,13.640206,11.401847,9.337437,8.27077,8.635077,10.459898,11.999181,14.224411,15.209026,15.465027,17.93641,19.744822,20.93949,21.750156,22.137438,21.809233,21.947079,22.422976,23.945848,26.486156,29.269335,33.444103,34.31713,32.531696,30.706875,33.42441,39.821133,51.20657,70.347496,85.29723,69.4318,54.465645,46.21785,38.422977,29.673027,23.42072,21.431797,19.14749,15.780104,11.936821,9.580308,8.123077,7.785026,7.9852314,7.768616,5.8223596,7.2303596,6.304821,5.5269747,5.179077,3.3509746,2.5173335,2.422154,2.793026,3.2886157,3.515077,2.8849232,2.1202054,2.425436,3.8498464,5.277539,5.5729237,5.5105643,5.4580517,5.4875903,5.3727183,4.516103,3.6496413,3.062154,2.5600002,1.467077,0.8566154,0.4201026,0.3314872,0.4660513,0.41025645,0.67610264,0.5349744,0.4201026,0.9682052,3.0096412,3.515077,2.858667,2.3072822,2.15959,1.723077,1.6935385,1.4473847,1.5983591,2.4188719,3.82359,4.818052,6.445949,6.619898,5.2414365,4.2272825,4.7524104,4.266667,4.273231,4.9788723,5.3103595,6.242462,7.427283,7.250052,6.170257,6.7183595,6.0291286,4.9526157,4.9394875,5.61559,4.785231,4.263385,3.882667,3.8104618,3.9942567,4.1550775,5.1232824,5.2742567,4.7392826,4.138667,4.59159,4.9132314,4.7491283,4.2141542,3.5249233,3.0030773,3.6529233,4.384821,4.919795,5.0116925,4.457026,2.3236926,1.401436,1.3193847,1.4966155,1.1355898,0.256,0.013128206,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0,0.006564103,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.013128206,0.098461546,0.3708718,0.42338464,0.6465641,0.7089231,0.5284103,0.24287182,0.16738462,0.14441027,0.16082053,0.19692309,0.21661541,0.18379489,0.15425642,0.12143591,0.098461546,0.118153855,0.15097436,0.27241027,0.39384618,0.45620516,0.45620516,0.5973334,0.7318975,0.9714873,1.4998976,2.5600002,2.5337439,2.3696413,2.477949,2.6912823,2.281026,2.609231,2.8914874,3.114667,3.3575387,3.7776413,3.8301542,3.9909747,4.7294364,5.7107697,5.802667,5.3070774,4.9821544,5.297231,6.0061545,6.1341543,6.157129,6.2063594,5.9995904,5.6418467,5.6320004,5.3760004,5.366154,5.3398976,5.481026,6.432821,6.4754877,6.445949,6.4590774,6.47877,6.298257,6.931693,7.456821,7.821129,7.781744,6.892308,6.2884107,6.2096415,6.675693,7.574975,8.677744,9.961026,9.278359,8.372514,7.9425645,7.6570263,6.5936418,6.2030773,6.377026,6.764308,6.7971287,6.3868723,5.9930263,5.8978467,6.157129,6.5936418,7.5388722,7.00718,6.045539,5.32677,5.172513,4.9788723,5.0510774,5.674667,6.49518,6.5280004,5.8781543,7.13518,7.6996927,6.564103,4.31918,4.1189747,4.240411,4.709744,5.349744,5.756718,5.691077,4.31918,3.0851285,2.4155898,1.719795,1.4539489,2.8258464,4.2896414,5.398975,6.816821,4.772103,5.2512827,5.7764106,5.1987696,3.7120004,1.2865642,1.1388719,1.3981539,1.3620514,1.4998976,1.4834872,1.5425643,1.6836925,1.7920002,1.6475899,1.6443079,1.8018463,1.7624617,1.6114873,1.8707694,1.8740515,1.6672822,1.5885129,1.657436,1.5819489,1.3915899,1.463795,1.6246156,1.8412309,2.2153847,2.3926156,2.5862565,2.6880002,2.6978464,2.737231,2.8816411,2.5206156,2.5042052,2.858667,2.7864618,2.809436,2.7076926,2.6354873,2.7175386,3.0654361,3.7316926,3.876103,4.076308,4.4373336,4.601436,4.013949,3.4822567,3.2000003,3.2328207,3.498667,3.6332312,3.945026,4.3585644,4.7622566,5.0084105,5.211898,5.093744,5.1265645,5.5007186,6.1341543,5.7829747,5.5105643,5.4416413,5.654975,6.189949,6.485334,6.695385,6.928411,7.145026,7.1581545,7.430565,7.7981544,8.027898,8.004924,7.7292314,8.113232,8.4972315,9.229129,10.200616,10.860309,10.850462,10.745437,10.624001,10.581334,10.752001,10.9686165,10.7158985,10.098872,9.344001,8.786052,9.025641,9.55077,9.82318,9.632821,9.127385,8.868103,9.301334,9.688616,9.787078,9.865847,10.230155,9.42277,8.736821,8.51036,8.12636,8.710565,8.736821,8.667898,8.562873,8.093539,8.018052,8.257642,8.467693,8.549745,8.631796,7.3353853,6.3540516,5.8190775,5.6320004,5.47118,4.6769233,3.498667,2.7470772,2.7044106,3.1442053,3.0030773,2.7536411,2.3958976,2.0808206,2.1234872,2.3696413,3.1409233,4.059898,4.5817437,4.020513,3.3805132,3.4330258,3.8498464,4.457026,5.2512827,5.612308,5.5269747,5.3366156,5.221744,5.1954875,4.716308,3.82359,3.2656412,3.4888208,4.634257,6.5280004,8.004924,9.399796,10.59118,11.017847,11.040821,11.113027,10.745437,10.059488,9.77395,9.8363085,8.891078,8.385642,8.4053335,7.686565,8.444718,8.280616,8.36595,8.966565,9.462154,9.199591,9.396514,9.298052,8.874667,8.815591,8.730257,9.16677,9.432616,9.212719,8.562873,2.6387694,2.4057438,2.3171284,2.2482052,2.284308,2.7142565,2.556718,2.4648206,2.5632823,2.8225644,3.0752823,3.5577438,4.076308,4.532513,4.8147697,4.772103,5.024821,5.208616,5.4908724,5.7796926,5.737026,5.228308,5.799385,6.4754877,6.6002054,5.8420515,6.242462,6.0750775,6.4722056,7.4371285,7.857231,8.874667,13.705847,20.594873,26.584618,27.536413,21.287386,26.863592,31.67508,28.261745,14.293334,8.51036,6.9382567,5.9602056,4.2469745,2.733949,2.028308,1.6738462,1.9200002,2.4549747,2.3860514,2.4943593,2.550154,2.4582565,2.1825643,1.7526156,1.529436,1.332513,1.2307693,1.2931283,1.595077,1.585231,1.782154,2.100513,2.3794873,2.3630772,2.5928206,2.4188719,2.172718,1.9790771,1.7460514,1.3161026,1.1158975,0.92553854,0.6859488,0.5152821,0.47917953,0.44964105,0.5021539,0.65969235,0.8763078,1.0338463,0.8566154,0.67938465,0.58420515,0.40369233,0.24287182,0.16082053,0.08861539,0.02297436,0.02297436,0.052512825,0.08205129,0.1148718,0.19692309,0.42994875,1.2274873,2.028308,2.678154,3.1770258,3.6660516,4.6769233,5.208616,5.1232824,4.8082056,5.1889234,8.146052,10.889847,11.828514,10.94236,9.760821,11.352616,12.2847185,12.914873,12.898462,11.1983595,10.010257,9.07159,7.8441033,6.518154,6.0225644,7.634052,8.195283,8.536616,8.073847,4.772103,6.5378466,8.234667,8.67118,8.342975,9.4457445,9.6754875,9.097847,10.125129,12.553847,13.558155,12.517745,11.812103,11.844924,12.09436,11.090053,10.624001,9.987283,9.728001,10.056206,10.84718,11.116308,11.61518,12.337232,13.056001,13.354668,13.699283,13.082257,12.980514,13.426873,13.02318,11.736616,11.529847,13.305437,16.518566,19.167181,19.193438,18.110361,17.650873,18.176,18.678156,17.67713,16.44636,16.426668,17.778873,19.380514,17.430975,16.758156,16.869745,17.217642,17.220924,17.23077,16.777847,16.019693,15.471591,16.003283,16.256,16.144411,16.019693,16.068924,16.305231,15.908104,15.904821,16.019693,16.49231,18.080822,16.59077,15.268104,14.690463,14.690463,14.372104,13.755078,12.980514,12.2387705,11.723488,11.608616,11.490462,12.202667,12.675283,12.609642,12.488206,12.987078,14.201437,14.608412,13.978257,13.387488,12.645744,12.235488,11.457642,10.748719,11.661129,13.83713,14.923489,15.084309,14.831591,15.028514,14.401642,14.621539,14.841437,15.015386,15.898257,16.633438,16.610462,16.433231,16.512001,17.060104,17.706669,18.36308,18.241642,17.227488,15.868719,15.330462,15.29436,14.546052,13.653335,14.953027,15.927796,16.738462,16.70236,16.036104,15.852309,13.184001,10.683078,9.127385,8.822155,9.6,9.636104,12.002462,13.676309,14.194873,15.652103,17.778873,19.154053,21.077335,23.102362,23.026873,24.218258,25.465437,27.2279,29.528618,31.947489,34.983387,37.408825,36.558773,34.241642,36.755695,43.736618,50.980106,58.36144,64.436516,66.43529,55.85067,47.5438,39.702976,31.684925,24.001642,21.07077,19.324718,16.485744,12.626052,10.157949,9.255385,7.7423596,7.4075904,7.653744,5.474462,5.2480006,5.0674877,4.31918,3.31159,3.2984617,2.4746668,2.1398976,2.0939488,2.169436,2.2383592,2.5435898,2.3827693,2.6354873,3.692308,5.4547696,5.691077,5.8125134,5.7829747,5.4875903,4.7261543,4.8311796,3.9712822,3.318154,2.9538465,1.8740515,1.1158975,0.5907693,0.6498462,1.1158975,1.2898463,2.300718,2.0512822,1.5753847,1.7296412,3.1737437,3.7809234,2.737231,2.1070771,2.3105643,2.1202054,2.1267693,1.719795,1.6607181,2.2088206,3.1277952,3.6562054,5.0084105,5.546667,5.142975,5.169231,5.208616,4.0992823,4.2994876,5.4514875,4.388103,4.1124105,4.1878977,5.218462,6.806975,7.5454364,6.1440005,5.3924108,5.2053337,5.169231,4.5390773,3.6627696,3.114667,2.5698464,2.2744617,3.0358977,3.0227695,3.3050258,2.8553848,2.100513,2.9078977,4.535795,4.2174363,3.242667,2.484513,2.412308,3.2361028,3.9122055,4.969026,6.3179493,7.273026,3.117949,1.148718,0.67282057,0.7450257,0.15097436,0.029538464,0.0,0.0,0.0032820515,0.0,0.013128206,0.006564103,0.0,0.0032820515,0.006564103,0.0032820515,0.0032820515,0.0032820515,0.0032820515,0.0,0.0,0.0,0.009846155,0.059076928,0.190359,0.4397949,0.7384616,0.9485129,0.9288206,0.5481026,0.37415388,0.28882053,0.27241027,0.30194873,0.35774362,0.26584616,0.18051283,0.118153855,0.101743594,0.15097436,0.17723078,0.318359,0.4266667,0.45292312,0.44964105,0.60389745,0.7778462,1.0502565,1.5786668,2.5895386,2.2646155,2.1530259,2.3827693,2.6486156,2.2153847,2.4024618,3.006359,3.4888208,3.6135387,3.4494362,3.6036925,3.8400004,4.4701543,5.3398976,5.8486156,5.156103,4.9329233,5.366154,6.0685134,6.0685134,5.920821,5.786257,5.6352825,5.5105643,5.5302567,5.2578464,5.0674877,4.772103,4.647385,5.4547696,5.933949,6.1046157,6.0816417,5.989744,5.9602056,7.0432825,7.5520005,7.719385,7.785026,8.011488,7.3452315,6.9842057,7.571693,8.923898,10.020103,10.240001,9.110975,8.096821,7.6964107,7.4404106,6.485334,6.445949,6.7282057,6.954667,6.9710774,6.377026,5.674667,5.346462,5.504,5.907693,6.7314878,6.554257,5.901129,5.211898,4.857436,4.972308,5.0543594,5.8157954,6.9349747,7.072821,6.2227697,7.2960005,7.8637953,6.987488,5.2315903,4.2830772,4.71959,5.933949,7.030154,6.8004107,7.4765134,4.850872,3.1113849,3.1081028,2.3335385,1.9692309,3.170462,4.7294364,6.5411286,9.616411,5.0609236,4.394667,6.091488,8.034462,7.499488,3.2098465,1.6377437,1.2176411,1.1257436,1.2635899,1.4473847,1.7427694,1.9889232,2.0217438,1.6475899,1.6147693,1.785436,1.7657437,1.6082052,1.8084104,1.8740515,1.7624617,1.6804104,1.719795,1.8346668,1.5031796,1.4769232,1.6344616,1.9003079,2.225231,2.2711797,2.2908719,2.4484105,2.678154,2.6683078,2.789744,2.4681027,2.4155898,2.6847181,2.6584618,2.7011285,2.7142565,2.733949,2.858667,3.2196925,4.0434875,4.4701543,4.6867695,4.7917953,4.8114877,4.6244106,4.023795,3.4756925,3.2754874,3.5478978,4.073026,4.532513,4.890257,5.097026,5.093744,5.2315903,4.962462,4.9854364,5.435077,5.8945646,5.4186673,5.297231,5.4482055,5.8518977,6.557539,6.918565,7.0892315,7.3058467,7.5520005,7.5618467,7.604513,7.506052,7.6209235,7.9294367,8.024616,8.241231,8.310155,8.92718,10.102155,11.149129,11.674257,11.684103,11.690667,11.805539,11.759591,11.54954,10.8537445,10.043077,9.366975,8.976411,8.841846,9.074872,9.701744,10.289231,9.941334,9.711591,9.862565,9.892103,9.77395,9.96759,10.315488,9.347282,8.310155,7.8802056,8.182155,9.143796,8.940309,9.07159,9.688616,9.616411,9.238976,8.65477,8.083693,7.77518,8.018052,6.7774363,5.7468724,5.356308,5.3792825,4.926359,4.519385,3.5610259,2.7273848,2.5304618,3.2820516,3.5872824,3.4133337,2.9538465,2.4582565,2.2383592,2.5009232,3.2623591,3.9844105,4.2929235,3.9778464,3.442872,3.4330258,3.7316926,4.2863593,5.1954875,5.83877,6.012718,5.7764106,5.346462,5.0838976,4.6145644,3.6463592,3.2032824,3.767795,5.277539,7.030154,8.4972315,9.747693,10.712616,11.204924,11.369026,11.388719,11.090053,10.522257,9.954462,10.033232,9.058462,8.648206,8.881231,8.300308,8.992821,8.704,8.569437,8.841846,8.891078,8.585847,8.864821,9.078155,9.058462,9.091283,8.923898,9.334154,9.40636,8.92718,8.392206,2.8849232,2.6880002,2.5665643,2.4681027,2.3827693,2.3335385,2.5796926,2.7503593,2.7437952,2.674872,2.868513,3.2722054,3.4921029,3.8334363,4.2469745,4.332308,4.7622566,5.077334,5.3891287,5.5893335,5.3727183,5.5663595,5.989744,6.193231,6.121026,6.1341543,7.0137444,6.482052,6.6822567,7.9195905,8.651488,10.752001,16.961643,23.003899,26.706053,27.999182,19.515078,21.4679,24.454565,21.897848,10.056206,6.8332314,5.973334,5.2644105,3.9680004,2.806154,2.0151796,1.5425643,1.5097437,1.7526156,1.8018463,2.1924105,1.9593848,1.6902566,1.6410258,1.7394873,1.6049232,1.6738462,1.6968206,1.5458462,1.204513,0.9616411,0.8992821,0.98461545,1.079795,0.94523084,1.0305642,1.6114873,1.8740515,1.8543591,2.4418464,2.2449234,2.0676925,1.6475899,0.9911796,0.380718,0.29538465,0.35774362,0.380718,0.3511795,0.4135385,0.571077,0.48246157,0.3708718,0.318359,0.24287182,0.21989745,0.18707694,0.118153855,0.036102567,0.0,0.098461546,0.26912823,0.2986667,0.2231795,0.32164106,0.6498462,1.1257436,2.1103592,3.3476925,3.9811285,4.5554876,5.835488,6.7872825,7.141744,7.384616,9.288206,15.753847,20.965746,22.311386,20.368412,22.567387,23.299284,23.414156,22.931694,21.024822,18.497643,15.314053,11.273847,7.0826674,4.348718,5.973334,7.4141545,8.766359,8.753231,4.699898,7.177847,8.474257,8.408616,8.224821,10.604308,10.384411,11.483898,13.154463,14.181745,12.86236,13.364513,14.815181,14.211283,11.431385,9.245539,9.941334,9.8592825,10.121847,11.053949,12.176412,13.334975,14.762668,14.9628725,14.293334,14.953027,16.626873,15.396104,13.761642,12.937847,12.86236,11.021129,10.807796,12.22236,14.677335,16.984617,18.960411,17.814976,16.30195,16.44636,19.5479,20.096,19.328001,18.405745,18.22195,19.393642,18.185848,18.021746,18.202257,18.428719,18.78318,19.712002,18.809437,17.946259,18.23836,20.020514,19.285336,18.435284,17.591797,17.027283,17.135592,17.19795,17.440823,17.014154,16.384,17.348925,17.42113,16.827078,16.49231,16.518566,16.190361,15.360002,13.722258,12.685129,12.721231,13.367796,13.170873,12.983796,12.852514,12.511181,11.414975,11.572514,12.993642,14.116103,14.352411,14.083283,14.424617,15.2155905,14.677335,12.84595,11.54954,13.797745,15.37313,16.003283,15.323898,12.895181,13.712411,16.242872,17.145437,16.091898,15.763694,16.128002,16.420103,16.682669,17.033848,17.670565,18.756924,19.22954,18.996513,17.723078,14.831591,15.074463,16.026258,15.432206,13.830565,14.5263605,15.980309,16.827078,16.896002,16.498873,16.449642,16.20349,13.197129,10.906258,10.187488,9.245539,8.598975,9.4457445,11.221334,13.174155,14.358975,15.323898,19.042463,21.11672,20.841026,21.195488,23.781746,25.593437,27.2279,29.348104,32.66954,36.26995,39.240208,40.01477,39.36821,40.40534,46.946465,53.51713,56.461132,56.02134,56.352825,52.358566,47.36985,41.74113,34.68144,24.247797,24.198566,20.246977,15.894976,13.016617,11.85477,9.878975,7.7357955,6.370462,5.5958977,4.1189747,5.671385,6.2490263,4.8640003,2.5895386,2.5796926,1.8838975,2.1202054,2.3762052,2.3236926,2.2121027,2.5173335,2.806154,2.9505644,3.3280003,4.8082056,5.208616,5.4843082,5.677949,5.543385,4.532513,7.0104623,5.175795,3.498667,3.131077,1.9232821,1.1651284,0.6465641,0.5907693,1.2176411,2.7306669,5.0510774,5.4547696,4.9132314,4.017231,2.989949,5.152821,4.2535386,3.0030773,2.4615386,2.0611284,1.4998976,1.3029745,2.353231,4.6178465,7.1548724,8.2904625,9.764103,10.039796,8.795898,6.928411,6.633026,4.775385,3.9154875,4.4012313,4.3651285,5.0838976,5.796103,6.7544622,7.4699492,6.7150774,6.445949,7.2664623,6.5017443,4.1846156,3.0358977,2.7175386,2.2383592,2.3466668,2.8291285,2.487795,2.4746668,3.1573336,3.0851285,2.1136413,1.4178462,1.8346668,2.422154,2.6486156,2.5862565,2.9144619,2.878359,3.6463592,5.110154,6.931693,8.530052,4.3552823,1.5524104,0.571077,0.6892308,0.029538464,0.006564103,0.0,0.006564103,0.013128206,0.0,0.013128206,0.006564103,0.006564103,0.01969231,0.029538464,0.01969231,0.016410258,0.016410258,0.013128206,0.0,0.0,0.0,0.006564103,0.04266667,0.15097436,0.5316923,0.9288206,1.1355898,1.086359,0.8533334,0.512,0.33476925,0.2986667,0.39384618,0.6268718,0.3708718,0.23958977,0.18051283,0.16082053,0.19692309,0.24615386,0.37743592,0.4266667,0.4135385,0.5349744,0.62030774,0.69579494,0.8730257,1.2832822,2.0742567,2.550154,2.3762052,2.359795,2.6683078,2.8389745,2.8980515,3.1967182,3.436308,3.4231799,3.0818465,3.2656412,3.9056413,4.827898,5.7140517,6.1046157,5.3825645,5.2020516,5.612308,6.1078978,5.6320004,5.7632823,5.5696416,5.6418467,5.933949,5.737026,5.1987696,5.0477953,4.9329233,4.9788723,5.7829747,6.7216415,6.262154,5.4875903,5.179077,5.8125134,6.7282057,7.240206,7.634052,8.04759,8.500513,8.92718,9.196308,9.649232,10.240001,10.545232,8.858257,7.1023593,6.6002054,7.1220517,6.8660517,6.5870776,6.038975,5.98318,6.482052,6.8955903,5.835488,5.549949,5.612308,5.664821,5.431795,6.3245134,6.6461544,6.5739493,6.2129235,5.61559,5.2480006,5.293949,6.0947695,7.1220517,6.987488,6.5870776,7.13518,7.4765134,6.987488,5.586052,4.8049235,5.405539,5.674667,5.664821,7.200821,8.1066675,5.146257,3.948308,5.106872,4.164923,4.1517954,3.4625645,3.8301542,6.514872,12.314258,7.7981544,4.1583595,3.2984617,5.668103,10.269539,6.705231,3.0490258,1.0699488,0.92225647,1.1290257,1.3128207,2.0184617,2.4582565,2.294154,1.6475899,1.6836925,1.913436,1.9364104,1.7624617,1.785436,2.0545642,1.8084104,1.6311796,1.7723079,2.1530259,1.8707694,1.6738462,1.6607181,1.847795,2.1530259,1.9429746,2.0020514,2.4057438,2.8258464,2.5337439,2.3630772,2.3926156,2.3302567,2.2416413,2.546872,2.6715899,2.737231,2.8947694,3.2820516,4.013949,4.562052,4.7458467,5.044513,5.533539,5.874872,5.47118,4.46359,3.6529233,3.4756925,4.013949,4.673641,4.6539493,4.519385,4.5554876,4.775385,4.7261543,4.532513,4.9099493,5.7009234,5.858462,5.9569235,5.723898,5.602462,5.8256416,6.422975,7.0104623,7.256616,7.3353853,7.512616,8.149334,8.208411,7.6110773,7.240206,7.318975,7.4174366,8.100103,8.756514,9.672206,10.8537445,12.038565,11.634872,11.34277,11.490462,11.9171295,11.979488,11.625027,10.729027,9.498257,8.254359,7.460103,8.205129,9.179898,10.387693,11.30995,10.893129,10.371283,10.30236,10.059488,9.711591,10.039796,9.833026,8.976411,7.9327188,7.27959,7.706257,8.805744,8.766359,9.097847,9.921641,9.993847,9.665642,9.225847,8.5661545,7.8703594,7.6143594,5.805949,4.972308,4.781949,4.827898,4.6080003,4.585026,3.6529233,2.7175386,2.5271797,3.6627696,4.2962055,4.529231,4.0402055,3.0326157,2.228513,2.556718,3.3345644,3.7743592,3.820308,4.1517954,3.761231,3.7349746,3.9680004,4.4012313,5.034667,6.11118,6.626462,6.2030773,5.182359,4.6080003,4.414359,3.8038976,3.6890259,4.519385,6.301539,7.643898,9.032206,10.197334,10.889847,10.86359,11.145847,11.178667,10.689642,9.882257,9.429334,9.429334,8.999385,8.828718,9.009232,9.032206,8.740103,9.317744,9.501539,9.035488,8.681026,8.474257,8.625232,8.923898,9.104411,8.835282,8.63836,8.976411,8.937026,8.464411,8.329846,2.3236926,2.166154,2.1267693,2.284308,2.5632823,2.7503593,2.7602053,2.930872,2.9538465,2.8947694,3.1967182,3.5610259,3.501949,3.82359,4.414359,4.2371287,4.6145644,4.7524104,4.890257,5.100308,5.2611284,5.4482055,5.7009234,5.7403083,5.7764106,6.51159,6.688821,6.0849237,6.4754877,8.004924,9.176616,14.391796,21.7239,29.19713,33.217644,28.586668,18.313848,21.044514,24.448002,21.428514,10.105436,6.3245134,5.1265645,4.6867695,4.0500517,3.1245131,2.300718,1.8379488,1.6935385,1.6640002,1.3620514,1.8018463,1.8576412,1.7952822,1.7493335,1.7394873,1.6049232,1.5327181,1.529436,1.529436,1.4145643,1.1191796,1.2964103,1.3915899,1.2898463,1.3128207,1.3981539,1.3915899,1.211077,1.0108719,1.1979488,1.4211283,1.2832822,1.024,0.7450257,0.41682056,0.4201026,0.36430773,0.3117949,0.318359,0.44964105,0.44964105,0.39056414,0.3052308,0.21989745,0.14769232,0.11158975,0.10502565,0.072205134,0.016410258,0.0,0.01969231,0.15753847,0.29538465,0.3511795,0.27241027,0.43651286,0.7384616,1.2307693,1.9035898,2.665026,3.764513,5.4482055,6.961231,7.79159,7.6668725,7.4108725,9.02236,13.653335,19.190155,20.23713,18.057848,16.94195,17.752617,20.020514,21.953642,22.455797,21.146257,17.88718,13.472821,9.645949,7.899898,6.265436,5.211898,4.713026,4.2371287,5.0051284,6.5706673,7.9491286,8.73354,9.091283,7.532308,9.02236,11.437949,13.331694,13.938873,17.378464,18.107079,15.904821,12.068104,9.393231,9.170052,9.547488,10.450052,11.59877,12.504617,12.09436,13.866668,15.205745,15.530668,16.295385,17.362053,15.698052,14.217847,14.066873,14.608412,13.449847,13.046155,14.043899,15.547078,15.140103,18.435284,17.85436,16.662975,16.603899,17.900309,18.379488,17.952822,17.299694,16.99118,17.490053,18.097233,18.320412,18.405745,18.579693,19.03918,20.096,20.020514,19.91877,20.361847,21.412104,20.384823,19.052309,18.392616,18.635489,19.236105,19.265642,18.500925,17.746052,17.72636,19.06872,18.615797,18.225233,18.103796,18.090668,17.654156,16.531694,15.481437,14.884104,14.78236,14.8939495,15.126975,15.156514,14.86113,13.909334,11.756309,11.270565,11.923694,13.144616,14.299898,14.693745,13.728822,14.775796,15.796514,15.51754,13.443283,15.084309,15.366566,15.839181,16.088617,13.748514,13.892924,16.187078,17.85436,17.867489,16.981335,17.739489,18.724104,18.999796,18.875078,19.892515,19.40677,19.075283,19.009642,18.399181,15.514257,15.074463,16.475899,17.001026,16.193642,15.845745,15.520822,16.531694,17.473642,17.539284,16.521847,16.649847,15.527386,14.385232,13.249642,10.932513,9.941334,8.769642,8.513641,9.954462,13.541744,12.386462,13.548308,16.62359,19.922052,20.46359,22.806976,24.914053,25.698463,26.134975,29.252926,31.93436,35.245953,39.486362,43.49703,44.65231,48.725338,54.3278,56.69744,54.3278,48.964928,46.10626,43.8318,40.34626,34.3959,25.24554,21.51713,17.746052,14.585437,12.179693,10.171078,10.440206,8.172308,5.914257,5.07077,5.8781543,5.7009234,5.4153852,4.6112823,3.442872,2.6387694,2.0118976,2.5764105,3.006359,2.8291285,2.3958976,3.0227695,3.045744,3.0260515,3.4133337,4.5390773,5.1659493,5.4974365,5.3070774,4.713026,4.1780515,5.651693,4.5390773,3.4658465,3.0785644,2.0578463,1.5360001,1.1684103,0.8369231,0.90584624,2.2416413,6.380308,9.429334,11.303386,12.107488,12.156719,7.532308,4.7327185,3.2722054,2.7470772,2.8521028,1.9987694,1.6344616,1.7132308,2.2416413,3.2886157,8.201847,10.240001,9.747693,7.7390776,5.8912826,6.5739493,8.1755905,8.293744,6.9021544,6.3277955,5.612308,4.5456414,4.345436,4.7524104,4.0041027,5.1922054,6.3967185,6.1013336,4.70318,4.5128207,4.8705645,3.8400004,3.2196925,3.1507695,2.097231,2.8553848,3.0424619,2.681436,2.1070771,1.9692309,1.9626669,1.4736412,0.9321026,0.72861546,1.204513,2.681436,3.9680004,4.378257,3.7284105,2.3302567,1.5425643,1.1323078,0.8205129,0.45292312,0.01969231,0.0032820515,0.006564103,0.009846155,0.0032820515,0.0,0.0032820515,0.0,0.0,0.009846155,0.029538464,0.009846155,0.009846155,0.01969231,0.02297436,0.0,0.009846155,0.0032820515,0.006564103,0.026256412,0.06564103,0.41682056,0.7975385,0.9124103,0.8533334,1.1093334,0.7975385,0.5907693,0.48246157,0.4660513,0.5513847,0.35446155,0.30851284,0.26912823,0.20676924,0.17394873,0.18379489,0.21661541,0.24287182,0.2986667,0.49887183,0.64000005,0.702359,1.0305642,1.6836925,2.428718,2.3794873,2.8127182,2.9013336,2.6223593,2.7536411,3.0293336,3.3214362,3.2787695,2.9505644,2.8127182,3.1343591,3.6758976,4.5095387,5.3070774,5.346462,4.8705645,5.3234878,5.7501545,5.7632823,5.5204105,5.3924108,5.3070774,5.3103595,5.182359,4.4307694,3.9712822,4.0008206,4.3618464,4.9887185,5.8814363,6.5280004,6.770872,6.803693,6.9054365,7.4141545,7.430565,7.755488,8.297027,8.805744,8.87795,10.213744,10.226872,9.485129,8.838565,9.4457445,8.188719,7.213949,7.1122055,7.640616,7.6964107,6.232616,6.1768208,6.2916927,6.124308,5.9930263,5.5269747,5.7665644,5.970052,5.9569235,6.114462,5.7074876,5.677949,6.0980515,6.449231,5.6287184,5.037949,5.3924108,6.196513,6.7971287,6.3901544,6.0356927,7.1680007,7.9885135,7.515898,5.586052,4.850872,6.2063594,7.059693,6.770872,6.629744,6.340924,4.164923,3.058872,3.9187696,5.605744,5.691077,4.417641,4.588308,5.730462,4.0992823,7.9819493,8.4053335,6.616616,5.0084105,7.1187696,7.755488,5.6254363,2.8455386,0.98461545,1.0568206,1.5327181,1.9593848,2.1333334,2.1103592,2.1858463,1.8510771,1.9200002,1.9298463,1.7690258,1.6738462,1.9823592,1.9626669,1.9889232,2.1234872,2.103795,1.7920002,1.6246156,1.5097437,1.5655385,2.1136413,2.2482052,2.428718,2.5600002,2.487795,2.0217438,2.2022567,2.2022567,2.169436,2.176,2.2186668,2.8488207,3.239385,3.6496413,4.164923,4.71959,4.7425647,4.457026,4.7655387,5.5630774,5.7403083,5.142975,4.3060517,3.8367183,3.9122055,4.2929235,4.9427695,5.031385,4.667077,4.2436924,4.4340515,4.315898,4.9329233,5.668103,6.009436,5.543385,5.5532312,5.540103,5.4908724,5.6320004,6.422975,7.2631803,7.7357955,7.785026,7.768616,8.454565,8.388924,7.640616,7.1548724,7.3616414,8.172308,8.864821,10.387693,11.753027,12.530872,12.855796,12.688411,12.360206,12.481642,12.800001,12.199386,11.346052,10.7158985,10.010257,9.147078,8.254359,8.500513,8.736821,9.465437,10.509129,10.9915905,11.132719,10.86359,10.551796,10.450052,10.712616,9.977437,8.861539,7.7259493,7.0498466,7.4371285,8.224821,7.837539,7.8112826,8.438154,8.772923,8.533334,8.772923,8.553026,7.857231,7.6012316,6.2818465,5.4449234,4.972308,4.7392826,4.6080003,4.6605134,3.9253337,3.1638978,3.1113849,4.4800005,4.598154,4.7950773,4.2272825,3.0162053,2.2383592,2.7634873,3.3444104,3.6102567,3.7316926,4.394667,3.7874875,3.7251284,4.0303593,4.5522056,5.156103,5.8125134,6.180103,5.8978467,5.2709746,5.2414365,5.037949,4.522667,4.598154,5.405539,6.3376417,7.8080006,8.871386,9.777231,10.676514,11.608616,12.475078,12.668719,12.137027,11.099898,10.052924,10.256411,9.921641,9.3078985,8.822155,9.032206,9.199591,9.708308,9.813334,9.468719,9.32759,8.585847,8.454565,8.736821,9.03877,8.763078,8.264206,8.385642,8.2904625,7.7948723,7.3682055,2.3729234,2.2711797,2.2744617,2.353231,2.487795,2.6880002,2.5665643,2.5862565,2.6322052,2.7831798,3.3280003,3.6069746,3.6562054,3.9220517,4.2830772,4.0467696,4.6112823,4.7228723,4.8738465,5.293949,5.9667697,5.4547696,5.4514875,5.425231,5.3202057,5.5532312,5.7074876,5.504,6.301539,8.41518,11.109744,17.867489,24.966566,30.903797,32.36431,24.25436,18.582975,24.086977,27.625029,22.86277,10.262975,6.7314878,5.3169236,4.670359,4.0336413,3.239385,2.5074873,2.0053334,1.7329233,1.6410258,1.654154,2.172718,2.0545642,1.782154,1.6508719,1.7755898,1.8116925,1.6836925,1.4703591,1.2865642,1.2898463,1.1093334,1.1782565,1.2209232,1.1782565,1.211077,1.2176411,1.0929232,1.0305642,1.1355898,1.4244103,1.7985642,1.913436,1.7394873,1.4244103,1.2800001,0.8992821,0.62030774,0.49230772,0.48246157,0.4660513,0.4004103,0.35446155,0.29538465,0.21661541,0.15097436,0.10502565,0.07548718,0.049230773,0.02297436,0.009846155,0.009846155,0.07548718,0.18379489,0.29538465,0.37743592,0.44307697,0.5973334,0.8533334,1.2438976,1.8412309,3.1376412,4.854154,6.2129235,6.820103,6.665847,6.173539,6.3245134,8.195283,11.001437,12.091078,11.411694,10.65354,11.053949,13.00677,16.06236,17.171694,17.02072,15.176207,12.166565,9.468719,8.280616,6.012718,4.279795,3.876103,4.7622566,5.330052,6.99077,7.8703594,7.8473854,8.556309,7.939283,9.009232,10.151385,10.761847,11.247591,14.053744,15.337027,14.844719,13.141335,11.628308,10.41395,10.220308,10.778257,11.605334,12.012309,12.048411,13.715693,15.189335,15.763694,15.855591,14.8939495,14.759386,15.133539,15.556924,15.402668,14.86113,14.677335,15.520822,16.584206,15.586463,17.234053,17.51959,16.961643,16.515284,17.56882,18.648617,18.921026,18.766771,18.251488,17.122463,18.084105,18.487797,18.491077,18.602669,19.698874,20.178053,20.033642,19.91549,20.135386,20.680206,20.657232,20.184616,19.98113,20.26995,20.775387,20.558771,20.178053,19.56759,19.252514,20.342155,20.729437,20.299488,19.734976,19.154053,18.103796,16.928822,15.993437,15.386257,15.291079,15.970463,16.134565,16.36431,16.229744,15.225437,12.757335,11.539693,11.910565,13.184001,14.549335,15.074463,14.821745,15.514257,16.118155,16.006565,14.959591,15.570052,15.940925,17.033848,17.926565,15.819489,15.451899,17.650873,20.20431,21.441643,20.263386,20.201027,20.486567,20.722874,20.854155,21.159386,19.652925,19.111385,19.062155,18.65518,16.682669,15.684924,16.361027,16.764719,16.324924,15.852309,16.262566,17.09949,18.228514,18.579693,16.164104,15.894976,15.504412,15.241847,14.946463,14.080001,12.018872,10.597744,9.816616,9.885539,11.241027,10.19077,10.660104,13.8075905,18.44513,21.03795,22.895592,24.625233,25.071592,25.097849,27.582361,27.867899,30.152208,35.121235,41.248825,44.790157,50.07754,54.587082,54.961235,50.737236,44.3438,41.199593,39.67344,38.009438,34.530464,27.631592,21.559797,17.542566,15.189335,13.380924,10.272821,9.872411,8.54318,6.7216415,5.149539,4.890257,5.720616,5.3005133,4.522667,3.6824617,2.4910772,2.422154,2.9538465,3.2689233,3.1540515,2.9997952,3.4231799,3.3017437,3.2229745,3.5478978,4.414359,5.0477953,5.540103,5.658257,5.287385,4.417641,5.405539,4.673641,3.7152824,3.1442053,2.6945643,2.0906668,1.8182565,1.4375386,1.0896411,1.4998976,4.4406157,6.7577443,10.082462,14.36554,17.847795,13.147899,7.4797955,3.4822567,1.9954873,2.034872,1.6213335,2.425436,2.9111798,2.7273848,2.6945643,6.340924,6.931693,6.806975,6.8299494,6.370462,6.157129,7.282872,7.634052,6.7117953,5.622154,4.955898,4.089436,4.568616,5.7403083,4.7458467,5.0149746,5.3924108,5.2644105,4.8836927,5.3858466,4.8049235,4.0369234,3.7349746,3.8662567,3.7120004,3.373949,2.868513,2.678154,3.0654361,4.092718,3.2951798,1.7427694,0.5677949,0.2986667,0.8336411,1.8838975,2.740513,2.8980515,2.15959,0.64000005,0.50543594,0.48902568,0.40369233,0.20348719,0.02297436,0.0032820515,0.009846155,0.01969231,0.026256412,0.026256412,0.013128206,0.013128206,0.02297436,0.029538464,0.029538464,0.01969231,0.02297436,0.026256412,0.029538464,0.026256412,0.026256412,0.016410258,0.013128206,0.029538464,0.08205129,0.702359,1.0962052,1.1585642,1.017436,1.0371283,1.1290257,0.9419488,0.75487185,0.6892308,0.7089231,0.4955898,0.36102566,0.28225642,0.23302566,0.17723078,0.16082053,0.17723078,0.21661541,0.29210258,0.45292312,0.54482055,0.702359,1.1520001,1.7985642,2.225231,1.9462565,2.284308,2.5140514,2.5337439,2.858667,3.1442053,3.131077,2.9046156,2.6322052,2.5435898,3.0326157,3.5380516,4.017231,4.348718,4.342154,4.5423594,5.1922054,5.651693,5.654975,5.3103595,5.4580517,5.691077,5.717334,5.540103,5.4416413,4.9952826,4.962462,5.2578464,5.799385,6.5083084,7.3550773,7.640616,7.6898465,7.821129,8.372514,8.4053335,8.63836,8.897642,8.953437,8.533334,9.298052,9.613129,9.288206,8.726975,8.940309,8.15918,7.460103,7.1154876,7.2894363,8.03118,6.8233852,6.436103,6.3573337,6.2162056,5.786257,5.586052,5.579488,5.5565133,5.5663595,5.910975,5.648411,5.8880005,6.1472826,6.0225644,5.182359,4.7392826,4.890257,5.4383593,5.9930263,5.9569235,5.9667697,6.73477,7.5585647,7.8145647,6.9776416,6.87918,8.14277,7.6668725,5.6943593,5.805949,6.370462,4.890257,3.2886157,3.5249233,7.5946674,6.2916927,5.756718,6.442667,7.1023593,4.7917953,9.468719,11.67754,10.023385,6.377026,5.874872,7.975385,7.7981544,5.651693,2.6847181,0.88287187,1.2832822,1.6278975,1.7394873,1.7296412,1.972513,1.7132308,1.7591796,1.7755898,1.6771283,1.6311796,1.8576412,2.0020514,2.2121027,2.3893335,2.162872,1.7657437,1.595077,1.5360001,1.6213335,2.03159,1.9232821,2.1169233,2.412308,2.5862565,2.3958976,2.3040001,2.169436,2.297436,2.5600002,2.412308,2.868513,3.4855387,3.8859491,4.0041027,4.092718,4.7228723,4.466872,4.532513,5.041231,5.0215387,4.4242053,4.194462,4.31918,4.630975,4.8114877,5.2676926,5.182359,4.709744,4.2568207,4.466872,4.6572313,5.4383593,6.0947695,6.235898,5.8190775,5.691077,5.605744,5.865026,6.373744,6.6527185,6.685539,6.944821,7.240206,7.5946674,8.254359,7.958975,7.6964107,7.837539,8.631796,10.220308,10.834052,11.313231,11.959796,12.58995,12.530872,12.73436,12.570257,12.1698475,11.670976,11.218052,10.79795,10.637129,10.476309,10.134975,9.504821,8.904206,8.848411,9.275078,10.092308,11.18195,11.434668,10.978462,10.561642,10.410667,10.240001,9.819899,8.697436,7.6012316,7.030154,7.269744,8.15918,7.9294367,7.778462,8.123077,8.605539,8.254359,8.237949,8.057437,7.565129,6.948103,6.413129,5.8978467,5.3070774,4.7950773,4.772103,4.640821,4.3749747,3.9778464,3.8104618,4.59159,4.6539493,4.706462,4.2240005,3.2328207,2.3171284,3.0720003,3.5380516,3.6594875,3.7776413,4.601436,4.2272825,4.1550775,4.309334,4.6244106,5.031385,5.612308,6.0028725,6.1505647,6.1407185,6.2063594,5.8157954,5.412103,5.4514875,6.0160003,6.7971287,8.136206,9.209436,10.171078,11.149129,12.225642,12.360206,12.071385,11.369026,10.689642,10.9226675,11.21477,10.79795,10.138257,9.6525135,9.711591,9.750975,10.102155,9.980719,9.442462,9.409642,8.726975,8.329846,8.320001,8.493949,8.323282,7.821129,7.8145647,7.6701546,7.204103,6.6592827,2.4484105,2.4910772,2.5829747,2.5632823,2.4681027,2.5107694,2.4057438,2.422154,2.4713848,2.6387694,3.1803079,3.5183592,3.6693337,3.8400004,3.9876926,3.8465643,4.522667,4.6900516,4.9296412,5.4941545,6.2851286,5.5958977,5.5236926,5.4613338,5.172513,4.7983594,4.965744,5.3005133,6.308103,8.4053335,11.910565,19.081848,25.366976,29.846977,29.797747,20.70318,18.766771,24.484104,26.548515,20.657232,9.488411,7.1647186,5.910975,5.1987696,4.647385,4.017231,3.2820516,2.7044106,2.2088206,1.9265642,2.1924105,2.6387694,2.2186668,1.7099489,1.5195899,1.6738462,1.8051283,1.6640002,1.4539489,1.332513,1.401436,1.3915899,1.3915899,1.3522053,1.3161026,1.4375386,1.4572309,1.1979488,1.0732309,1.2471796,1.6508719,2.1464617,2.3893335,2.228513,1.8510771,1.7657437,1.2176411,0.8992821,0.7844103,0.7384616,0.508718,0.36102566,0.2986667,0.25928208,0.22646156,0.2297436,0.16410258,0.10502565,0.059076928,0.026256412,0.016410258,0.016410258,0.036102567,0.08861539,0.18707694,0.34133336,0.40369233,0.5284103,0.7417436,1.0601027,1.4736412,2.5928206,4.076308,5.1364107,5.467898,5.2611284,4.9427695,4.775385,4.7556925,4.9952826,5.6943593,6.744616,7.276308,7.571693,8.39877,11.044104,11.871181,12.091078,11.35918,9.852718,8.267488,7.433847,5.799385,4.388103,4.0303593,5.3891287,6.5280004,7.8112826,8.3364105,8.362667,9.301334,9.498257,9.449026,9.527796,9.783795,9.924924,11.109744,12.258463,13.177437,13.51877,12.780309,10.9915905,10.138257,10.387693,11.152411,11.067078,11.707078,13.105232,15.051488,16.800821,17.079796,15.530668,16.357744,17.250463,17.293129,16.951796,16.31836,16.259283,16.928822,17.696821,17.14872,16.938667,17.834667,17.844515,17.046976,17.56882,19.528206,20.210873,20.384823,19.968002,18.021746,18.149744,18.793028,19.18031,19.324718,20.033642,20.184616,20.184616,19.984411,19.738258,19.767796,20.30277,20.824617,21.11672,21.3399,22.009438,21.75672,21.809233,21.50072,21.074053,21.67795,22.409847,22.078362,21.3399,20.296207,18.5239,17.03713,15.803078,15.172924,15.468308,16.978052,17.191385,17.631182,17.772308,16.984617,14.503386,12.672001,13.000206,14.375385,15.750566,16.118155,15.737437,16.052513,16.239592,16.187078,16.472616,16.49231,17.263592,18.822565,19.938463,18.113642,17.306257,18.947283,21.868309,24.287182,23.785027,23.04,22.4919,22.498463,22.816822,22.6199,20.457027,19.396925,18.891489,18.41231,17.463797,16.46277,16.39713,16.580925,16.577642,16.183796,17.214361,17.729643,17.920002,17.83795,17.385027,16.38072,16.039387,16.118155,16.36431,16.508718,13.856822,12.576821,11.414975,10.19077,9.80677,8.461129,8.822155,11.204924,15.120412,19.305027,20.59159,22.038977,23.033438,23.870361,25.744411,24.287182,25.734566,30.178463,36.273235,41.252106,48.256004,52.237133,51.17703,46.23426,41.750977,38.751183,36.975594,36.164925,34.917747,30.70031,24.18872,19.478975,16.439796,14.211283,11.1983595,9.990565,9.042052,7.4830775,5.4482055,4.1124105,5.0084105,5.0084105,4.7491283,4.1189747,2.2646155,2.733949,3.2886157,3.370667,3.1048207,3.31159,3.5347695,3.5347695,3.5905645,3.8695388,4.4406157,5.044513,5.5597954,5.874872,5.786257,5.0116925,5.661539,5.4613338,4.4242053,3.2262566,3.2065644,2.5961027,2.294154,1.8937438,1.3850257,1.1618463,2.0545642,2.9111798,5.7698464,10.948924,17.05354,16.311796,11.362462,5.989744,2.4385643,1.4178462,1.3357949,2.878359,4.2272825,4.453744,3.511795,4.5390773,4.273231,5.3924108,7.243488,5.8420515,6.49518,7.0367184,6.87918,5.986462,4.850872,4.7556925,4.5522056,5.408821,6.47877,4.9099493,5.3398976,5.4449234,5.353026,5.2676926,5.4580517,4.4734364,3.9811285,3.9876926,4.269949,4.3651285,4.1091285,3.8990772,3.757949,3.9417439,4.9460516,3.4002054,1.723077,0.67282057,0.5218462,1.0469744,1.1848207,1.5556924,1.6246156,1.1881026,0.39712822,0.19692309,0.08861539,0.055794876,0.052512825,0.02297436,0.0032820515,0.013128206,0.029538464,0.03938462,0.032820515,0.013128206,0.02297436,0.032820515,0.03938462,0.036102567,0.036102567,0.03938462,0.049230773,0.055794876,0.052512825,0.04594872,0.03938462,0.036102567,0.055794876,0.14441027,0.7844103,1.1979488,1.2996924,1.1618463,1.024,1.3981539,1.273436,1.0929232,1.020718,0.92225647,0.62030774,0.41682056,0.30194873,0.24287182,0.17723078,0.15753847,0.17394873,0.21989745,0.29210258,0.37743592,0.4660513,0.7778462,1.2373334,1.723077,2.0841026,1.8412309,1.8445129,1.910154,2.0545642,2.5173335,2.9604106,3.0194874,2.9046156,2.7831798,2.802872,3.1015387,3.446154,3.7185643,3.8498464,3.82359,4.535795,5.080616,5.4908724,5.7107697,5.5597954,5.986462,6.3179493,6.2884107,6.117744,6.485334,6.189949,5.9995904,6.117744,6.564103,7.181129,7.8112826,7.8473854,7.7948723,8.041026,8.858257,9.094564,9.147078,9.07159,8.779488,8.024616,8.198565,8.786052,9.084719,8.992821,9.032206,8.536616,7.8441033,7.276308,7.13518,7.702975,6.9087186,6.5247183,6.363898,6.189949,5.7074876,5.546667,5.280821,5.0904617,5.152821,5.654975,5.622154,5.85518,5.730462,5.146257,4.522667,4.4077954,4.4701543,4.95918,5.674667,5.979898,6.114462,6.3212314,7.069539,8.123077,8.556309,9.668923,10.364718,8.464411,5.4613338,6.491898,6.957949,6.518154,5.658257,5.691077,8.736821,7.765334,7.1515903,7.4765134,8.119796,7.269744,9.291488,11.867898,11.319796,7.680001,4.70318,6.547693,8.14277,7.683283,4.844308,0.77128214,1.014154,1.2603078,1.3292309,1.3259488,1.6344616,1.7001027,1.7985642,1.8051283,1.7558975,1.8445129,2.0184617,2.1267693,2.2449234,2.2908719,2.0118976,1.6082052,1.4769232,1.4867693,1.6016412,1.8740515,1.7099489,1.8445129,2.2416413,2.6518977,2.5961027,2.3696413,2.1464617,2.2711797,2.6256413,2.6256413,2.8914874,3.6168208,4.0467696,3.9811285,3.8038976,4.460308,4.414359,4.4110775,4.598154,4.5128207,4.2601027,4.388103,4.6834874,4.955898,5.037949,5.080616,5.0182567,4.6769233,4.2929235,4.5423594,5.1987696,5.786257,6.196513,6.3606157,6.245744,6.160411,6.0258465,6.2490263,6.6592827,6.482052,6.157129,6.340924,6.9710774,7.899898,8.87795,8.690872,8.996103,9.475283,10.177642,11.513436,12.173129,12.2387705,12.448821,12.773745,12.402873,12.672001,12.616206,12.06154,11.234463,10.761847,10.59118,10.581334,10.594462,10.522257,10.292514,9.465437,9.344001,9.609847,10.194052,11.280411,11.756309,11.559385,11.185231,10.742155,9.93477,9.596719,8.740103,7.890052,7.3419495,7.1647186,7.6996927,8.01477,8.109949,8.205129,8.746667,8.605539,8.165744,7.8080006,7.4863596,6.7282057,6.6461544,6.308103,5.5729237,4.8049235,4.8705645,4.466872,4.568616,4.571898,4.4242053,4.6178465,4.8672824,4.772103,4.345436,3.6004105,2.553436,3.4198978,3.8498464,3.9548721,4.082872,4.8344617,4.768821,4.670359,4.647385,4.772103,5.0674877,5.540103,6.048821,6.5411286,6.872616,6.806975,6.3901544,6.0816417,6.1341543,6.6067696,7.3747697,8.615385,9.875693,10.7848215,11.506873,12.744206,12.248616,11.306667,10.515693,10.450052,11.641437,12.032001,11.641437,11.139283,10.893129,10.9686165,10.94236,10.768411,10.134975,9.255385,8.864821,8.434873,8.100103,7.8802056,7.702975,7.430565,7.1647186,7.0432825,6.7938466,6.4000006,6.1046157,2.4484105,2.5895386,2.7306669,2.737231,2.605949,2.477949,2.4582565,2.5895386,2.6157951,2.6026669,2.917744,3.3444104,3.4888208,3.5905645,3.7054362,3.7251284,4.312616,4.578462,4.9920006,5.5729237,5.924103,5.668103,5.7731285,5.691077,5.2611284,4.706462,4.7622566,5.412103,6.235898,7.5979495,10.627283,17.129026,22.6199,27.040823,27.716925,19.350975,18.727386,22.501745,22.170258,15.858873,8.349539,7.525744,6.560821,5.8814363,5.4974365,5.0051284,4.417641,3.8432825,3.0818465,2.4024618,2.540308,2.7536411,2.172718,1.6344616,1.467077,1.5064616,1.5655385,1.4211283,1.4080001,1.5786668,1.7066668,1.8838975,1.8970258,1.8379488,1.8084104,1.9200002,1.9856411,1.529436,1.1191796,1.0535386,1.3718976,1.847795,1.9889232,1.8346668,1.5589745,1.4736412,1.1158975,1.0010257,0.98461545,0.8960001,0.53825647,0.31507695,0.2297436,0.21661541,0.23958977,0.28882053,0.2100513,0.13784617,0.07548718,0.029538464,0.01969231,0.016410258,0.02297436,0.049230773,0.0951795,0.15097436,0.26584616,0.47917953,0.79425645,1.1881026,1.6246156,2.425436,3.5905645,4.522667,4.8836927,4.6211286,4.1452312,3.6496413,3.3805132,3.5183592,4.1517954,5.0543594,6.5345645,7.2992826,7.64718,9.468719,10.144821,10.276103,10.246565,9.813334,8.113232,6.0783596,5.169231,4.4800005,4.2371287,5.7764106,7.3780518,8.195283,9.160206,10.292514,10.692924,10.699488,9.596719,9.6065645,10.880001,11.510155,11.831796,11.85477,12.580104,13.571283,12.964104,11.277129,9.888822,9.586872,10.138257,10.299078,11.122872,11.999181,14.322873,17.345642,18.166155,18.484514,19.702156,19.93518,19.236105,19.59713,18.481232,18.09395,18.307283,18.786463,18.963694,18.04472,18.852104,19.226257,18.582975,17.923283,20.171488,20.50954,20.706463,20.890259,19.554462,18.563284,19.403488,20.43077,20.74913,20.22072,20.217438,20.483284,20.522669,20.217438,19.83672,19.908924,20.814772,21.494156,21.822361,22.596926,22.488617,22.482054,22.4919,22.62318,23.174566,23.23036,22.90872,22.212925,20.975592,18.86195,17.089642,15.599591,15.218873,16.170668,18.090668,18.556719,18.894772,19.167181,18.793028,16.554668,14.572309,14.772514,16.06236,17.371899,17.650873,16.118155,16.111591,16.466053,16.932104,18.159592,18.070976,18.999796,20.598156,21.730463,20.46031,19.183592,19.705437,22.275284,25.498259,26.368002,25.488413,24.566156,24.175592,24.201847,23.867079,21.62872,19.958155,18.881643,18.28431,17.903591,17.306257,17.05354,17.257027,17.611488,17.371899,18.189129,18.330257,17.010874,16.039387,19.826874,18.130053,17.660719,17.496616,17.319386,17.391592,15.186052,13.702565,11.923694,10.033232,9.412924,7.210667,7.282872,8.618668,11.030975,15.143386,16.039387,17.191385,18.776617,20.74913,22.836515,21.799387,22.852924,26.384413,31.501131,36.050053,43.25744,47.156517,46.099697,41.96431,40.15262,38.53785,36.65395,35.859695,35.61354,33.48349,27.825233,22.478771,17.988924,14.716719,12.84595,11.542975,9.885539,7.79159,5.658257,4.3716927,3.8465643,4.3027697,4.818052,4.4012313,2.0151796,2.861949,3.498667,3.4100516,2.92759,3.2131286,3.4034874,3.6726158,3.9909747,4.338872,4.673641,5.2742567,5.6385646,5.8157954,5.8486156,5.7632823,5.8092313,6.9054365,5.9995904,3.5446157,3.4822567,2.9013336,2.484513,2.0250258,1.5589745,1.3423591,0.82379496,0.892718,1.9495386,4.775385,10.515693,14.083283,13.210258,9.196308,4.3027697,1.7657437,1.4834872,2.7142565,4.667077,5.914257,4.4077954,4.0402055,3.9089234,5.7403083,7.6668725,4.2338467,6.997334,7.781744,7.0826674,5.7665644,5.0642056,5.353026,5.4974365,5.792821,5.7501545,4.086154,5.930667,6.009436,5.7632823,5.658257,5.1954875,4.594872,4.082872,3.9318976,3.95159,3.501949,4.8738465,5.412103,4.844308,3.7710772,3.698872,2.0184617,1.086359,0.7450257,0.8533334,1.2898463,0.9189744,0.9747693,0.8402052,0.41682056,0.15097436,0.06564103,0.026256412,0.013128206,0.013128206,0.013128206,0.0032820515,0.016410258,0.032820515,0.036102567,0.01969231,0.009846155,0.01969231,0.029538464,0.029538464,0.04266667,0.04266667,0.052512825,0.068923086,0.08205129,0.072205134,0.128,0.12471796,0.108307704,0.128,0.25271797,0.5874872,1.0108719,1.214359,1.1848207,1.1946667,1.5458462,1.467077,1.3718976,1.3357949,1.0732309,0.7778462,0.5481026,0.380718,0.26256412,0.18379489,0.16082053,0.16410258,0.20020515,0.25928208,0.3052308,0.46276927,0.9288206,1.3095386,1.6049232,2.2219489,2.1300514,1.782154,1.4506668,1.3915899,1.8313848,2.4943593,2.989949,3.2164104,3.2754874,3.4658465,3.3345644,3.5413337,3.8728209,4.1156926,4.0303593,4.8672824,5.2020516,5.408821,5.674667,6.0028725,6.422975,6.6133337,6.567385,6.4656415,6.6592827,6.5312824,6.298257,6.4295387,6.994052,7.64718,7.571693,7.3747697,7.387898,7.860513,8.950154,9.147078,9.065026,8.920616,8.628513,7.8047185,7.8703594,8.3823595,8.871386,9.186462,9.488411,9.15036,8.3593855,7.712821,7.4108725,7.2303596,6.5870776,6.51159,6.38359,5.976616,5.47118,5.2447186,4.9460516,4.7983594,4.9821544,5.6287184,5.3924108,5.1954875,4.821334,4.345436,4.1156926,4.2141542,4.3618464,4.9788723,5.8847184,6.3245134,6.183385,6.0685134,6.810257,8.3364105,9.655796,11.877745,11.703795,9.18318,6.4722056,7.8080006,7.53559,7.8769236,8.342975,8.828718,9.622975,10.86359,9.639385,8.201847,7.6931286,8.123077,7.8145647,9.737847,10.532104,8.539898,3.8334363,4.2535386,6.3868723,7.6570263,6.189949,0.81066674,0.8992821,0.9911796,1.024,1.1126155,1.5556924,1.8412309,2.0250258,2.048,2.0020514,2.1300514,2.3040001,2.2744617,2.1497438,1.9593848,1.6508719,1.404718,1.3357949,1.3522053,1.4408206,1.6935385,1.7526156,1.8871796,2.3040001,2.7536411,2.556718,2.3269746,2.1234872,2.1070771,2.3040001,2.6026669,2.9505644,3.570872,4.059898,4.2436924,4.1846156,4.0992823,4.2535386,4.3618464,4.348718,4.3618464,4.6572313,4.70318,4.6539493,4.644103,4.781949,4.4077954,4.5456414,4.457026,4.210872,4.644103,5.5893335,5.8912826,6.1407185,6.485334,6.62318,6.6527185,6.560821,6.426257,6.2523084,5.9602056,6.0061545,6.3573337,7.3780518,8.923898,10.338462,10.440206,11.23118,11.651283,11.572514,11.782565,12.599796,13.003489,13.200411,13.131488,12.4685135,12.458668,12.383181,12.1468725,11.697231,11.040821,10.778257,10.676514,10.551796,10.43036,10.545232,10.029949,9.987283,10.240001,10.676514,11.237744,12.182976,12.57354,12.3766165,11.628308,10.450052,9.718155,9.176616,8.621949,7.975385,7.2894363,6.9809237,7.748924,8.300308,8.434873,9.051898,9.521232,8.868103,8.192,7.79159,7.1647186,7.1909747,6.7282057,5.8453336,4.9920006,5.024821,4.4438977,4.522667,4.7950773,4.9821544,5.0018463,5.3103595,5.034667,4.59159,4.0303593,3.0326157,3.8498464,4.342154,4.5456414,4.6605134,5.0674877,5.146257,5.07077,5.0051284,5.07077,5.35959,5.622154,6.2555904,6.9152827,7.259898,6.9743595,6.6034875,6.419693,6.629744,7.1909747,7.8145647,9.117539,10.601027,11.319796,11.638155,13.233232,12.619488,11.2672825,10.512411,10.857026,11.953232,12.445539,12.3306675,12.130463,12.160001,12.507898,12.488206,11.497026,10.233437,9.074872,8.067283,7.827693,7.7259493,7.39118,6.8004107,6.2851286,6.3277955,6.1505647,5.85518,5.6352825,5.796103,2.7766156,2.605949,2.5074873,2.612513,2.806154,2.7470772,2.6978464,2.7044106,2.674872,2.674872,2.930872,3.0654361,3.2886157,3.498667,3.6529233,3.8006158,4.141949,4.57518,5.3136415,5.9602056,5.5072823,5.2644105,5.6320004,5.5893335,5.0116925,4.670359,4.8049235,5.156103,5.425231,5.986462,7.90318,12.288001,17.447386,22.78072,24.84513,17.348925,19.74154,24.805746,23.824411,16.111591,9.032206,8.5202055,7.200821,5.933949,5.0674877,4.457026,4.84759,4.588308,3.6824617,2.612513,2.3204105,2.2711797,1.910154,1.6311796,1.5688206,1.6180514,1.4703591,1.332513,1.2668719,1.3259488,1.5721027,1.975795,1.7723079,1.913436,2.284308,1.723077,1.5655385,1.2504616,1.0010257,0.9321026,1.0535386,0.892718,0.8172308,0.8041026,0.81394875,0.7778462,0.5940513,0.7515898,0.8172308,0.65969235,0.4266667,0.29210258,0.25928208,0.28882053,0.30194873,0.16738462,0.108307704,0.055794876,0.029538464,0.029538464,0.029538464,0.01969231,0.016410258,0.026256412,0.052512825,0.07548718,0.16082053,0.5316923,1.024,1.6246156,2.4418464,3.3214362,4.345436,5.35959,6.0980515,6.196513,5.2315903,4.384821,4.007385,4.017231,3.9056413,4.2240005,5.0084105,5.973334,7.125334,8.772923,9.957745,10.282667,11.250873,11.88759,8.713847,5.3202057,4.0402055,4.0467696,4.8114877,6.117744,7.0465646,8.4053335,9.813334,10.8767185,11.168821,10.607591,9.974154,10.243283,11.707078,13.978257,15.100719,14.355694,14.240822,15.186052,15.563488,14.697027,12.402873,9.691898,8.28718,10.604308,11.88759,11.529847,11.949949,13.016617,12.038565,15.872002,19.43959,21.192207,21.428514,22.308104,21.612309,20.230566,19.472412,19.731693,20.476719,19.938463,19.639797,20.256823,21.011694,19.669334,20.266668,19.216412,19.249231,20.545643,20.752413,19.83672,20.368412,21.428514,22.075079,21.333336,20.233849,19.620104,20.25354,21.48431,21.241438,20.434053,20.854155,21.7239,22.242464,21.605745,21.313643,21.02154,21.412104,22.675694,24.507078,23.699694,22.44595,20.992002,19.498669,18.021746,17.06995,16.20677,16.49559,17.897026,19.288616,19.764515,19.012924,18.927591,19.328001,17.959387,16.725334,16.354464,16.800821,17.713232,18.432001,17.211079,16.521847,16.810667,18.100513,20.004105,19.505232,20.33231,21.930668,23.40431,23.512617,21.609028,20.886976,22.59036,25.80677,27.464207,26.489437,25.593437,24.825438,24.050873,22.964514,21.828924,20.795078,20.073027,19.590565,18.966976,18.464823,18.550156,18.527182,18.399181,18.875078,19.826874,19.534771,17.641027,16.420103,20.76554,18.727386,18.54031,17.703386,16.354464,17.257027,16.426668,14.306462,12.281437,10.535385,8.057437,6.774154,6.0783596,7.1220517,9.636104,11.933539,12.993642,12.849232,12.99036,14.683899,18.966976,21.395695,21.435078,23.919592,29.128208,32.790977,37.82236,41.137234,41.298054,39.223797,38.22277,38.990772,38.44267,37.74031,36.89026,34.727386,29.430157,24.562874,20.424206,17.398155,15.944206,14.224411,11.303386,8.129642,5.5532312,4.332308,3.515077,3.623385,3.629949,3.0030773,1.7099489,3.0162053,3.3772311,3.383795,3.3247182,3.190154,3.31159,3.5971284,4.1058464,4.7327185,5.2348723,5.805949,5.986462,6.0717955,6.23918,6.5444107,5.2512827,9.15036,9.094564,4.6178465,3.9220517,2.9702566,2.4648206,1.9823592,1.5392822,1.5885129,1.1355898,1.214359,1.2832822,1.4966155,2.7175386,6.2818465,7.8112826,7.568411,5.805949,2.793026,1.7657437,2.15959,3.9614363,5.723898,4.578462,5.5302567,4.6867695,4.1517954,4.332308,3.95159,5.3694363,5.2742567,5.395693,5.9667697,5.720616,5.805949,5.930667,5.58277,5.0642056,5.477744,6.882462,4.8147697,3.8990772,5.100308,5.720616,4.6605134,4.027077,3.370667,2.793026,2.9768207,5.1987696,4.6900516,3.0851285,1.6968206,1.5261539,1.0371283,0.65969235,0.65969235,0.9747693,1.204513,1.0601027,0.51856416,0.15425642,0.101743594,0.07548718,0.03938462,0.02297436,0.009846155,0.0,0.0,0.0,0.009846155,0.03938462,0.06564103,0.029538464,0.029538464,0.029538464,0.02297436,0.01969231,0.029538464,0.029538464,0.03938462,0.04594872,0.06235898,0.12143591,0.39056414,0.33805132,0.25271797,0.28882053,0.47261542,0.58420515,0.9485129,1.2176411,1.3029745,1.3883078,1.5360001,1.3981539,1.3718976,1.4276924,1.0994873,1.2209232,0.88615394,0.5316923,0.34133336,0.24287182,0.18379489,0.16738462,0.18051283,0.21989745,0.3052308,0.49887183,1.0436924,1.4112822,1.6607181,2.4418464,2.3794873,1.6147693,1.1552821,1.3062565,1.6475899,2.0873847,2.6354873,3.131077,3.501949,3.7842054,3.564308,4.1517954,4.650667,4.7524104,4.716308,5.421949,5.717334,5.481026,5.110154,5.540103,5.6352825,5.8256416,6.2162056,6.5969234,6.439385,6.048821,6.1440005,6.6560006,7.3682055,7.90318,7.3780518,7.2303596,7.351795,7.765334,8.621949,8.438154,8.713847,8.986258,8.900924,8.195283,8.195283,8.247795,8.63836,9.304616,9.842873,9.915077,8.989539,7.9885135,7.509334,7.827693,7.499488,6.8562055,6.380308,5.9963083,5.080616,4.824616,4.4307694,4.4307694,4.919795,5.5532312,5.0182567,4.5522056,4.3716927,4.4701543,4.6539493,4.457026,4.33559,4.7950773,5.723898,6.409847,5.858462,5.76,6.4656415,8.021334,10.131693,12.012309,10.660104,8.297027,6.514872,6.2720003,8.224821,7.430565,6.6560006,7.9852314,12.832822,15.284514,15.616001,11.556104,6.1341543,7.6603084,8.746667,8.92718,9.908514,10.289231,5.5532312,3.501949,3.4297438,4.8049235,5.3398976,1.0075898,0.8598975,0.84348726,1.0010257,1.3489232,1.8609232,1.7624617,2.0151796,2.2022567,2.1530259,1.9232821,2.0578463,2.1267693,2.1136413,1.9331284,1.4178462,1.5031796,1.4244103,1.3522053,1.401436,1.6311796,1.585231,2.028308,2.8356924,3.508513,3.2032824,2.3368206,2.2383592,2.2580514,2.1989746,2.3335385,2.9440002,3.062154,3.3608208,3.9154875,4.197744,3.9647183,4.2436924,4.2207184,3.8859491,4.0434875,4.6900516,4.4964104,4.086154,3.9023592,4.197744,3.892513,3.8596926,3.82359,3.9975388,5.097026,5.671385,5.8420515,6.23918,6.8430777,6.987488,6.7577443,6.633026,6.426257,6.1078978,5.8125134,5.9963083,6.416411,7.9819493,10.230155,11.352616,11.168821,12.570257,13.315283,12.895181,12.527591,13.380924,12.58995,12.015591,12.005745,11.382154,11.126155,10.998155,10.889847,10.7848215,10.771693,10.870154,11.076924,11.017847,10.801231,11.030975,10.226872,10.482873,10.9226675,11.126155,11.139283,12.409437,13.056001,12.937847,12.304411,11.779283,10.765129,10.102155,9.498257,8.805744,8.011488,7.194257,7.4830775,8.241231,9.101129,9.980719,11.10318,10.420513,9.268514,8.326565,7.6307697,7.9950776,7.2894363,6.47877,5.989744,5.720616,5.2447186,4.7228723,4.9362054,5.733744,6.0258465,5.720616,5.0871797,4.647385,4.4012313,3.8137438,4.535795,5.1987696,5.5007186,5.408821,5.1889234,5.152821,5.32677,5.4547696,5.504,5.674667,5.87159,6.560821,7.384616,7.8408213,7.27959,6.498462,6.5870776,7.0498466,7.5454364,7.890052,9.416205,11.0145645,11.776001,12.120616,13.794462,12.977232,11.828514,11.090053,11.08677,11.733335,12.199386,12.616206,12.937847,13.266052,13.840411,13.252924,11.605334,10.049642,8.933744,7.7981544,7.6274877,7.273026,6.5936418,5.786257,5.3727183,5.5302567,5.5138464,5.546667,5.720616,6.0258465,2.7175386,2.5731285,2.412308,2.3729234,2.425436,2.3433847,2.481231,2.5698464,2.5238976,2.4648206,2.7208207,2.9046156,3.0982566,3.2328207,3.3280003,3.495385,3.945026,4.529231,5.290667,5.9995904,6.1440005,5.586052,5.4514875,5.356308,5.1856413,5.097026,5.0642056,5.802667,6.36718,6.685539,7.5388722,10.085744,14.785643,18.454975,18.766771,14.260514,22.580515,27.877747,25.639387,16.95836,8.5202055,7.3550773,6.2752824,5.2644105,4.391385,3.820308,4.5423594,4.453744,3.692308,2.7076926,2.2580514,2.2580514,1.9331284,1.5688206,1.3653334,1.4342566,1.6672822,1.4506668,1.3193847,1.4178462,1.4867693,1.4900514,1.3029745,1.1913847,1.1782565,1.0765129,0.9878975,0.8730257,0.86317956,0.9517949,1.0043077,0.9616411,0.827077,0.7384616,0.702359,0.6071795,0.4135385,0.5513847,0.7417436,0.7515898,0.40369233,0.39712822,0.39384618,0.3249231,0.20020515,0.0951795,0.08205129,0.036102567,0.016410258,0.032820515,0.04266667,0.01969231,0.016410258,0.04266667,0.0951795,0.15097436,0.27241027,0.65969235,1.1388719,1.7887181,2.930872,4.1780515,5.546667,7.02359,8.257642,8.549745,7.7325134,7.312411,7.026872,6.76759,6.5805135,6.770872,7.141744,7.194257,7.325539,8.848411,10.305642,11.58236,14.076719,15.852309,11.654565,7.138462,5.3891287,4.7589746,4.562052,5.0576415,5.5926156,7.565129,9.337437,10.184206,10.289231,10.33518,12.186257,12.343796,10.8307705,11.204924,12.49477,13.617231,13.607386,13.403898,15.832617,14.624822,12.412719,9.829744,8.231385,9.701744,11.441232,11.047385,11.286975,12.576821,12.967385,16.17395,18.642054,20.65067,22.144001,22.711796,21.343182,20.719591,20.608002,20.709745,20.673643,21.504002,22.035694,22.636309,22.86277,21.461334,20.86072,19.728413,20.227283,21.91754,21.753437,23.299284,23.542156,23.22708,22.800411,22.419695,21.152822,20.036924,20.12554,21.156105,21.546669,21.792822,22.340925,22.961233,23.273027,22.71836,23.54872,23.059694,22.15713,21.897848,23.506054,24.516926,23.217232,21.14954,19.242668,17.824821,17.273438,16.790976,17.010874,17.91672,18.858667,19.383797,19.18031,18.855387,18.51077,17.739489,17.641027,17.673847,17.355488,17.165129,18.579693,18.619078,17.956104,17.312822,17.54913,19.685745,21.208616,22.583797,23.499489,24.33313,26.161232,23.88677,23.40759,24.218258,25.744411,27.3559,27.707079,27.414976,25.993849,23.978668,22.94154,23.082668,22.400002,21.947079,21.809233,21.077335,20.480001,19.669334,19.127796,19.127796,19.728413,20.768822,20.946053,19.003078,16.505438,17.811693,17.132309,18.609232,18.875078,18.228514,20.627693,19.43631,17.194668,14.454155,11.746463,9.570462,7.936001,7.4010262,7.9524107,9.609847,12.432411,11.667693,9.908514,9.468719,11.539693,16.196924,19.88595,21.257847,25.314463,31.337029,32.902565,34.054565,38.869335,41.728004,41.18318,39.968822,38.1998,39.476517,40.63508,38.87918,31.786669,27.88431,25.895386,23.187695,19.528206,17.06995,13.774771,10.203898,7.1154876,5.0674877,4.4438977,2.6190772,2.2547693,2.6289232,2.9965131,2.612513,3.4100516,3.5282054,3.7054362,4.0402055,3.9811285,3.7907696,4.0369234,4.5489235,5.110154,5.464616,6.3901544,6.7544622,6.738052,6.514872,6.2523084,5.730462,7.0826674,7.0859494,5.293949,4.0303593,2.8750772,2.1956925,1.7723079,1.4342566,1.0732309,0.76800007,0.9156924,0.8533334,0.65312827,1.0929232,1.9429746,2.7733335,3.5741541,3.9023592,2.878359,2.0676925,1.7591796,3.0326157,4.972308,4.663795,5.8781543,5.2480006,4.4274874,4.493129,5.940513,5.786257,4.066462,3.564308,4.384821,3.9647183,4.9985647,4.5423594,4.0041027,4.644103,7.578257,6.7938466,5.1922054,5.080616,6.3212314,6.3212314,5.277539,5.2381544,5.2315903,4.604718,2.9997952,4.138667,4.0402055,2.681436,0.95835906,0.7089231,0.40369233,0.761436,0.9616411,0.79425645,0.65641034,0.47917953,0.2855385,0.16082053,0.118153855,0.06564103,0.016410258,0.0032820515,0.0032820515,0.0,0.0,0.0,0.009846155,0.01969231,0.026256412,0.01969231,0.029538464,0.029538464,0.029538464,0.032820515,0.055794876,0.04594872,0.04594872,0.04594872,0.052512825,0.072205134,0.20348719,0.21333335,0.37415388,0.6465641,0.69251287,0.7056411,0.81394875,0.8172308,0.8041026,1.1454359,1.3095386,1.3686155,1.4112822,1.4145643,1.2209232,1.2242053,0.9353847,0.6826667,0.5677949,0.45292312,0.3314872,0.24287182,0.19692309,0.2231795,0.36758977,0.47261542,0.892718,1.1848207,1.463795,2.3794873,1.8806155,1.4867693,1.273436,1.2340513,1.2832822,1.3883078,1.7952822,2.2186668,2.550154,2.8816411,3.8038976,4.2272825,4.2305646,4.069744,4.1911798,5.464616,6.2687182,6.2490263,5.7042055,5.5762057,5.6451287,6.2129235,7.072821,7.785026,7.683283,7.4108725,7.7259493,7.965539,7.821129,7.3419495,7.3058467,7.328821,7.6077952,8.04759,8.267488,7.604513,7.6734366,7.955693,8.041026,7.6077952,7.6274877,8.448001,8.786052,8.5891285,9.048616,10.138257,10.220308,9.258667,7.9458466,7.719385,6.5083084,5.648411,5.412103,5.4186673,4.630975,4.1485133,4.086154,4.388103,4.818052,4.955898,4.84759,4.5128207,4.164923,4.056616,4.4832826,4.5128207,4.4832826,4.9296412,5.674667,5.8223596,5.9470773,5.832206,6.2227697,7.4896417,9.632821,10.807796,10.341744,9.137232,7.210667,3.69559,7.4174366,7.6209235,5.6352825,4.0533338,6.741334,11.82195,17.115898,15.268104,7.9458466,5.8289237,10.771693,11.191795,10.518975,9.03877,3.882667,3.0129232,2.7208207,3.9647183,5.0609236,1.7033848,1.4309745,1.079795,1.0929232,1.4867693,1.8740515,1.8346668,1.910154,1.9462565,1.9429746,2.03159,1.9331284,1.913436,1.7362052,1.4276924,1.2832822,1.3686155,1.394872,1.4867693,1.6180514,1.595077,1.595077,2.1792822,2.9013336,3.3509746,3.1442053,2.412308,2.2022567,2.3105643,2.6026669,3.0293336,3.0162053,3.4133337,4.066462,4.532513,4.1091285,3.7120004,3.9876926,4.1682053,4.0303593,3.895795,4.086154,4.161641,3.9876926,3.6332312,3.3772311,3.2689233,3.2656412,3.4921029,4.1846156,5.681231,5.737026,6.1472826,6.629744,7.00718,7.1844106,6.308103,6.0028725,6.048821,6.232616,6.3507695,6.485334,7.3714876,9.209436,11.290257,11.976206,12.865642,13.643488,12.62277,10.745437,11.54954,12.524308,12.770463,12.616206,12.242052,11.687386,10.857026,11.030975,11.418258,11.644719,11.749744,12.432411,12.465232,12.009027,11.447796,11.385437,11.1064625,11.152411,11.411694,11.487181,10.686359,11.625027,12.504617,12.616206,12.189539,12.3766165,11.490462,10.988309,10.374565,9.508103,8.595693,8.228104,8.182155,8.320001,8.884514,10.502565,12.173129,12.258463,11.539693,10.459898,9.130668,8.63836,7.899898,7.328821,6.9710774,6.5280004,6.2752824,5.7534366,5.536821,5.83877,6.5017443,6.1013336,5.346462,4.7261543,4.460308,4.5095387,5.425231,6.045539,6.193231,5.858462,5.1889234,5.142975,5.796103,6.3540516,6.6527185,7.1647186,7.39118,8.241231,9.124104,9.186462,7.315693,6.426257,6.6625648,7.312411,7.9819493,8.595693,10.043077,11.506873,12.425847,12.852514,13.4400015,13.305437,12.416001,11.608616,11.319796,11.588924,12.570257,13.00677,13.505642,14.25395,15.025232,13.840411,11.766154,10.20718,9.278359,7.8080006,7.24677,6.4065647,5.5269747,4.8836927,4.8082056,4.4110775,4.7622566,5.097026,5.2742567,5.7829747,2.8192823,2.8389745,2.6880002,2.6322052,2.6715899,2.5271797,2.4549747,2.356513,2.2646155,2.2350771,2.359795,2.540308,2.7667694,2.9505644,3.0523078,3.062154,3.8367183,4.4800005,5.3431797,6.2227697,6.3376417,5.805949,5.2644105,5.0018463,5.0149746,5.0116925,4.9362054,6.012718,6.6461544,6.7905645,7.9327188,10.66995,16.144411,18.520617,16.790976,14.79877,21.950361,24.726976,20.644104,11.979488,5.7665644,5.907693,5.720616,5.208616,4.525949,4.010667,4.2305646,3.6791797,2.7963078,2.0086155,1.7493335,1.782154,1.591795,1.273436,1.0502565,1.2800001,1.7755898,1.6147693,1.4933335,1.6410258,1.8116925,1.9200002,1.7952822,1.6147693,1.4375386,1.1979488,0.8763078,0.73517954,0.78769237,0.9124103,0.8467693,0.76800007,0.90256417,0.90584624,0.7515898,0.7384616,0.7187693,0.84348726,0.9714873,0.93866676,0.56123084,0.38728207,0.32820517,0.27241027,0.18051283,0.06564103,0.07548718,0.052512825,0.032820515,0.032820515,0.036102567,0.055794876,0.06235898,0.08533334,0.16082053,0.3314872,0.4004103,0.5546667,1.1454359,2.1792822,3.3345644,4.420923,5.3202057,6.232616,6.961231,6.9152827,6.6034875,6.554257,6.3376417,5.907693,5.58277,6.422975,6.705231,6.449231,6.0258465,6.183385,8.155898,11.277129,13.50236,13.778052,12.068104,9.938052,8.172308,6.5247183,5.156103,4.634257,5.4843082,7.315693,9.363693,10.581334,9.632821,7.965539,8.933744,9.7673855,10.049642,11.703795,11.021129,12.944411,13.863386,13.131488,13.062565,12.675283,11.372309,9.337437,7.6635904,8.349539,10.696206,11.116308,11.785847,13.351386,14.920206,18.592821,21.444925,24.067284,26.36472,27.572515,24.986258,24.795898,24.694157,23.680002,22.058668,21.661541,22.600206,23.827694,24.356104,23.240208,21.654976,21.123283,21.592617,22.327797,21.940514,24.33313,25.478565,25.107695,23.814566,23.046566,22.193232,20.499695,19.951591,20.824617,21.704206,22.317951,22.931694,24.119797,25.24554,24.451284,25.416206,24.730259,23.611078,23.14831,24.326567,24.77949,23.430567,21.139694,18.944002,18.06113,17.70995,17.10277,16.846771,17.204514,18.09395,19.173744,19.577436,19.242668,18.33354,17.237335,16.745028,16.804104,17.06995,17.532719,18.507488,18.802874,18.182566,17.408,17.283283,18.681437,21.668104,24.146053,25.1799,25.22913,26.148104,25.80677,25.655796,25.99713,26.873438,28.071386,28.980515,28.82954,27.323078,25.219284,24.326567,24.562874,24.710566,25.209438,25.744411,25.212719,24.457848,22.560822,21.195488,20.801643,20.59159,22.226053,21.861746,19.429745,16.692514,17.211079,15.675078,16.30195,17.801847,20.004105,23.857233,23.98195,22.393438,19.190155,15.126975,11.605334,9.202872,8.572719,8.201847,8.044309,9.527796,9.494975,7.450257,6.5936418,8.421744,12.737642,17.877335,21.202053,25.439182,29.88308,30.401644,31.780106,36.519386,40.8878,43.254158,44.130466,40.66462,41.153645,41.796925,39.542156,32.09518,27.795694,25.61313,22.57395,18.261335,14.805334,11.828514,8.749949,6.121026,4.46359,4.2863593,2.4484105,1.913436,2.3466668,3.0096412,2.7569232,3.7185643,3.764513,3.9417439,4.4406157,4.565334,4.5456414,4.8607183,5.3169236,5.8157954,6.3277955,7.197539,7.7259493,7.9885135,7.7390776,6.426257,5.8847184,6.12759,6.2851286,5.8912826,4.890257,3.2131286,2.2908719,1.785436,1.3817437,0.8008206,0.5907693,0.64000005,0.62030774,0.85005134,2.28759,2.487795,2.3401027,2.3072822,2.353231,1.9364104,1.5458462,1.2406155,1.7591796,2.8291285,3.1540515,4.6933336,4.6966157,4.1222568,3.8334363,4.6178465,4.9099493,3.8498464,4.073026,5.405539,4.8607183,5.346462,4.5817437,4.420923,5.6352825,7.9195905,5.277539,6.0685134,6.62318,5.943795,5.681231,4.7261543,4.6769233,4.775385,4.417641,3.1442053,3.9351797,3.8629746,2.6289232,0.9124103,0.35774362,0.3052308,0.6826667,0.761436,0.45620516,0.33476925,0.2855385,0.27897438,0.23302566,0.13784617,0.06235898,0.013128206,0.0,0.0032820515,0.009846155,0.009846155,0.009846155,0.01969231,0.03938462,0.059076928,0.052512825,0.08533334,0.08205129,0.06564103,0.049230773,0.04266667,0.03938462,0.049230773,0.059076928,0.059076928,0.04266667,0.10502565,0.15097436,0.38728207,0.67610264,0.56451285,0.7417436,0.8598975,0.8467693,0.8598975,1.2832822,1.5425643,1.6935385,1.4900514,1.1093334,1.142154,1.0666667,0.8533334,0.7778462,0.85005134,0.82379496,0.5940513,0.3314872,0.19364104,0.2297436,0.380718,0.43651286,0.79097444,1.1651284,1.5360001,2.1366155,1.5031796,1.3423591,1.2471796,1.1191796,1.1520001,1.1782565,1.4080001,1.7558975,2.169436,2.6289232,3.43959,4.2207184,4.6539493,4.778667,4.965744,5.6254363,6.2818465,6.491898,6.2555904,5.979898,6.245744,6.872616,7.5979495,8.155898,8.28718,7.890052,7.50277,7.2960005,7.269744,7.240206,7.6176414,7.5979495,7.5552826,7.755488,8.352821,7.512616,7.39118,7.512616,7.5913854,7.5618467,7.8441033,8.205129,8.1755905,7.906462,8.198565,8.753231,9.081436,8.763078,7.8080006,6.675693,6.2063594,5.5958977,5.3760004,5.32677,4.4996924,4.056616,4.096,4.2469745,4.4045134,4.7228723,4.6572313,4.5029745,4.164923,3.8564105,4.1091285,4.4077954,4.6211286,4.9887185,5.47118,5.7403083,6.6494365,6.380308,6.2720003,7.145026,9.324308,10.522257,10.581334,9.944616,8.2445135,4.279795,6.36718,6.7117953,5.9470773,4.7294364,3.7448208,9.980719,15.330462,15.763694,12.166565,10.331899,13.282462,11.565949,8.461129,5.61559,3.0424619,3.3345644,4.059898,5.2578464,5.5597954,2.2055387,1.8642052,1.4506668,1.2996924,1.4867693,1.8116925,1.8018463,1.8576412,1.8740515,1.8609232,1.9495386,1.8346668,1.6738462,1.404718,1.1454359,1.214359,1.3062565,1.3029745,1.4473847,1.6607181,1.522872,1.6804104,2.1858463,2.7831798,3.1737437,3.0260515,2.7208207,2.4352822,2.3958976,2.665026,3.1507695,3.058872,3.186872,3.4921029,3.7382567,3.4756925,3.5282054,3.9745643,4.132103,3.9220517,3.8596926,3.9351797,3.9712822,3.7743592,3.383795,3.0818465,3.2689233,3.5774362,4.266667,5.2315903,6.012718,5.9536414,5.924103,5.8092313,5.654975,5.677949,5.3202057,5.6385646,6.180103,6.547693,6.4032826,6.928411,8.864821,11.122872,12.760616,12.99036,13.725539,13.794462,13.00677,12.084514,12.672001,12.931283,13.00677,12.885334,12.557129,12.022155,11.805539,12.11077,12.251899,12.09436,12.028719,12.714667,12.754052,12.137027,11.365745,11.437949,11.890873,12.455385,12.914873,12.839386,11.58236,12.012309,12.760616,12.806565,12.356924,12.849232,12.498053,12.022155,11.260718,10.28595,9.373539,9.002667,8.815591,8.979693,9.596719,10.699488,11.884309,12.314258,12.268309,11.753027,10.502565,9.452309,8.51036,8.04759,7.9294367,7.53559,7.213949,6.7971287,6.416411,6.3507695,6.997334,6.803693,5.924103,4.9788723,4.5128207,5.0149746,6.0061545,6.5411286,6.4032826,5.7468724,5.0674877,5.0215387,5.7632823,6.49518,6.9809237,7.565129,7.768616,8.779488,9.77395,9.846154,8.001641,7.328821,7.394462,7.9819493,8.805744,9.498257,10.71918,12.018872,13.016617,13.636924,14.139078,13.75836,12.635899,12.153437,12.62277,13.298873,13.764924,13.157744,13.200411,14.234258,15.218873,14.070155,12.402873,10.834052,9.442462,7.77518,7.381334,6.3245134,5.2020516,4.4077954,4.1485133,3.9023592,4.397949,4.8377438,5.07077,5.5663595,2.9472823,3.0391798,2.9768207,2.8882053,2.7766156,2.4910772,2.3926156,2.2383592,2.166154,2.2088206,2.2744617,2.3860514,2.6847181,2.92759,3.0293336,3.05559,3.6660516,4.204308,5.10359,6.0619493,6.0324106,5.8518977,5.464616,5.208616,5.1364107,5.0215387,4.919795,6.045539,6.6100516,6.7282057,8.43159,11.621744,17.165129,18.638771,15.868719,14.913642,20.164925,20.660515,15.38954,7.3321033,3.4264617,4.31918,5.0576415,5.1232824,4.6244106,4.273231,4.1747694,3.0851285,2.041436,1.5622566,1.6311796,1.4703591,1.2865642,1.083077,0.9517949,1.0666667,1.6836925,1.7427694,1.6968206,1.7788719,1.9823592,2.1267693,2.0512822,1.847795,1.5524104,1.1454359,0.86974365,0.77128214,0.8205129,0.8992821,0.761436,0.71548724,0.9419488,1.024,0.9353847,1.020718,1.0338463,1.0075898,0.9714873,0.8730257,0.574359,0.32164106,0.23302566,0.21989745,0.19364104,0.06235898,0.059076928,0.055794876,0.049230773,0.03938462,0.049230773,0.118153855,0.128,0.15097436,0.24943592,0.44964105,0.47917953,0.5940513,1.1815386,2.2383592,3.370667,4.394667,4.9887185,5.428513,5.737026,5.7009234,5.661539,5.861744,5.802667,5.3792825,4.8804107,5.835488,5.973334,5.7009234,5.218462,4.516103,5.5171285,8.264206,10.079181,10.341744,10.512411,10.607591,9.002667,6.8004107,4.9460516,4.2141542,5.0215387,6.7282057,8.500513,9.508103,8.923898,6.5247183,6.1407185,7.030154,8.697436,10.896411,9.872411,11.083488,12.087796,11.690667,9.96759,11.792411,11.437949,9.987283,8.63836,8.690872,10.154668,11.746463,13.433437,14.92677,15.681643,19.498669,23.105642,25.737848,27.136002,27.536413,25.291489,25.826464,26.177643,25.22913,23.719387,22.22277,23.391182,24.94031,25.672207,25.48513,23.62749,22.774155,22.636309,22.662565,22.035694,24.218258,26.157951,26.525541,25.35713,24.041027,23.374771,21.782976,20.722874,20.795078,21.753437,22.757746,23.535591,25.051899,26.561644,25.616413,26.62072,26.272823,25.258669,24.306873,24.178873,24.1559,23.302567,21.451488,19.34113,18.62236,17.85436,17.270155,16.79754,16.679386,17.483488,18.816002,19.531488,19.620104,19.016207,17.608206,15.95077,15.799796,16.584206,17.680412,18.41559,18.881643,18.41231,17.716515,17.375181,17.85436,20.936207,23.91631,25.353848,25.491693,26.246567,27.385439,27.414976,27.569233,28.26831,29.131489,30.31631,30.447592,29.289028,27.680822,27.529848,27.858053,28.754053,29.738668,30.362259,30.194874,29.348104,26.594463,24.034464,22.52472,21.684515,23.489643,22.94154,20.289642,17.08636,16.200207,14.864411,14.464001,16.449642,20.519386,24.628515,26.83077,27.497028,25.83631,21.782976,16.01313,12.553847,10.525539,8.507077,6.8562055,7.709539,8.339693,6.232616,5.1298466,6.442667,9.235693,14.7790785,19.383797,23.095797,25.600002,26.213745,29.111797,33.398155,38.002876,42.515694,47.18934,44.288002,42.289234,40.66462,37.90113,31.478157,26.17436,23.223797,19.561028,14.746258,11.001437,8.973129,6.882462,5.0838976,3.9581542,3.9023592,2.4713848,1.8412309,1.9823592,2.4320002,2.281026,2.989949,3.2853336,3.564308,4.013949,4.601436,4.6933336,5.156103,5.7796926,6.5378466,7.581539,8.369231,8.861539,9.199591,8.950154,7.1220517,6.2884107,6.0160003,6.0356927,5.927385,5.1167183,3.9384618,2.9472823,2.2121027,1.6114873,0.83035904,0.60061544,0.54482055,0.62030774,1.1454359,2.789744,3.131077,2.8455386,2.356513,1.8871796,1.4605129,1.1454359,0.90256417,0.9485129,1.2898463,1.7394873,2.8914874,3.4756925,3.5314875,3.3772311,3.5971284,4.138667,3.8038976,4.2174363,5.346462,5.4843082,6.0225644,5.113436,4.630975,5.3366156,6.882462,4.273231,5.9503593,6.5936418,5.2480006,5.32677,4.604718,4.1780515,4.2830772,4.417641,3.3444104,3.5380516,3.0293336,1.9889232,0.85005134,0.3249231,0.31507695,0.446359,0.40697438,0.20676924,0.15097436,0.17394873,0.24287182,0.21661541,0.10502565,0.04266667,0.009846155,0.0,0.0032820515,0.009846155,0.009846155,0.02297436,0.052512825,0.08861539,0.1148718,0.08205129,0.12143591,0.118153855,0.098461546,0.08205129,0.06235898,0.06564103,0.07548718,0.072205134,0.059076928,0.04266667,0.08533334,0.13128206,0.28225642,0.4660513,0.43651286,0.7515898,0.8402052,0.90912825,1.0469744,1.2176411,1.5491283,1.6771283,1.3751796,0.88943595,0.94523084,0.86646163,0.7515898,0.7581539,0.8795898,0.93866676,0.65312827,0.35774362,0.21989745,0.26912823,0.40697438,0.4955898,0.78769237,1.1158975,1.4211283,1.7591796,1.2898463,1.2307693,1.1881026,1.0601027,1.024,1.1126155,1.2340513,1.4769232,1.8543591,2.297436,3.0424619,4.017231,4.8377438,5.32677,5.5138464,6.038975,6.62318,6.957949,6.889026,6.416411,6.7774363,7.27959,7.686565,7.9917955,8.4283085,8.01477,7.1483083,6.7840004,7.0957956,7.4699492,7.821129,7.6274877,7.39118,7.499488,8.241231,7.4240007,7.194257,7.3091288,7.5552826,7.7456417,7.962257,7.7325134,7.499488,7.5979495,8.237949,8.083693,7.6701546,7.3058467,6.9120007,5.9963083,6.058667,5.5663595,5.208616,4.9920006,4.204308,3.9876926,3.9122055,3.9548721,4.1517954,4.601436,4.2929235,4.2502565,4.082872,3.8137438,3.879385,4.1878977,4.457026,4.8672824,5.4514875,6.0816417,7.328821,6.8332314,6.377026,7.072821,9.3768215,10.8307705,11.510155,10.955488,8.976411,5.6385646,6.0192823,5.986462,6.488616,7.0334363,5.684513,10.5780525,13.400617,14.401642,14.037334,12.964104,11.684103,8.707283,5.546667,3.3509746,2.878359,3.8564105,4.3585644,4.565334,4.164923,2.3335385,2.0578463,1.7001027,1.4703591,1.4408206,1.5688206,1.7066668,1.7427694,1.8609232,2.028308,2.0053334,1.8313848,1.5688206,1.2537436,1.0338463,1.1651284,1.2209232,1.2603078,1.4309745,1.6311796,1.529436,1.7329233,2.425436,3.0851285,3.4034874,3.3017437,3.18359,2.8750772,2.6880002,2.7569232,3.0260515,3.1671798,2.9636924,2.9210258,3.0654361,2.9571285,3.249231,3.7448208,3.895795,3.7349746,3.8531284,3.892513,3.895795,3.6660516,3.2787695,3.0654361,3.3345644,3.8334363,4.7228723,5.651693,5.7632823,5.61559,5.333334,4.9394875,4.588308,4.571898,4.640821,5.3825645,6.1341543,6.5247183,6.49518,8.41518,10.65354,12.402873,13.482668,14.322873,14.680616,14.204719,13.791181,13.804309,14.086565,14.007796,13.692719,13.620514,13.702565,13.272616,13.341539,13.233232,12.839386,12.455385,12.786873,13.449847,13.633642,13.15118,12.343796,12.097642,12.550565,13.459693,14.099693,13.896206,12.42913,12.708103,13.092104,13.013334,12.770463,13.51877,13.361232,12.626052,11.785847,10.988309,10.059488,9.724719,9.53436,9.764103,10.423796,11.254155,11.61518,12.097642,12.36677,12.176412,11.382154,10.033232,9.005949,8.352821,8.004924,7.778462,7.463385,7.2664623,6.9743595,6.764308,7.204103,7.194257,6.452513,5.5762057,5.0838976,5.421949,6.38359,6.738052,6.2785645,5.3858466,5.044513,5.0674877,5.7829747,6.550975,7.145026,7.7292314,7.9425645,8.976411,9.95118,10.171078,9.130668,8.940309,8.891078,9.202872,9.80677,10.345026,11.08677,12.360206,13.515489,14.25395,14.628103,14.03077,13.00677,12.737642,13.4170265,14.244103,14.424617,13.551591,13.216822,13.846975,14.700309,14.050463,12.62277,10.9226675,9.271795,7.824411,7.4207187,6.193231,4.97559,4.194462,3.8662567,3.826872,4.3290257,4.716308,4.900103,5.346462,3.0129232,3.0424619,3.0818465,2.9111798,2.537026,2.162872,2.3269746,2.28759,2.2646155,2.3401027,2.4681027,2.487795,2.7995899,3.0326157,3.1376412,3.3903592,3.442872,3.820308,4.650667,5.5072823,5.412103,5.792821,5.940513,5.8814363,5.668103,5.3792825,5.221744,6.114462,6.5280004,6.698667,8.621949,11.313231,15.707899,16.843489,14.473847,13.075693,18.737232,18.825848,13.63036,6.2588725,2.6157951,3.05559,4.1846156,4.5456414,4.023795,3.8498464,3.9417439,2.7273848,1.782154,1.6869745,2.041436,1.6082052,1.3489232,1.2340513,1.1684103,0.97805136,1.5097437,1.7165129,1.7493335,1.7591796,1.8707694,1.8642052,1.7690258,1.5163078,1.1520001,0.8533334,0.84348726,0.827077,0.84348726,0.86974365,0.8402052,0.9189744,0.9353847,0.9682052,1.0633847,1.2438976,1.148718,0.92553854,0.73517954,0.61374366,0.45620516,0.27241027,0.20676924,0.2100513,0.20020515,0.06564103,0.04266667,0.03938462,0.04266667,0.04594872,0.07548718,0.16082053,0.20676924,0.25928208,0.35446155,0.49887183,0.67938465,1.0010257,1.5261539,2.3269746,3.4855387,4.598154,5.3202057,5.789539,6.114462,6.377026,6.4032826,6.5378466,6.5017443,6.173539,5.618872,5.943795,5.737026,5.4514875,5.175795,4.6211286,3.9745643,4.6966157,6.4656415,8.254359,8.342975,8.815591,7.3747697,5.579488,4.450462,4.4964104,4.841026,6.163693,6.9152827,7.0793853,8.165744,6.701949,5.681231,5.723898,6.741334,7.906462,8.487385,8.372514,8.697436,9.120821,7.830975,11.385437,11.759591,11.18195,10.745437,10.387693,9.82318,12.33395,14.903796,15.842463,14.795488,17.490053,21.56636,23.952412,23.995079,23.460104,23.06954,24.287182,24.953438,24.704002,24.966566,23.683285,25.124104,26.499285,27.001438,27.831797,26.259695,24.464413,23.768618,23.844105,22.711796,24.113234,26.384413,27.670977,27.254156,25.537643,24.713848,23.827694,22.672413,21.72718,22.153849,23.54872,24.513643,25.688618,26.643694,25.888823,26.978464,27.378874,26.505848,24.67118,23.082668,23.368206,23.286156,22.186668,20.417643,19.328001,17.621334,17.30954,17.02072,16.571077,16.94195,18.198977,19.072002,19.764515,19.905643,18.550156,16.180513,15.744001,16.387283,17.473642,18.579693,19.236105,18.881643,18.304,17.992207,18.139898,20.214155,22.800411,24.484104,25.370258,27.083488,28.360207,28.389746,28.416002,28.931284,29.659899,30.84472,31.556925,31.271387,30.723284,31.921234,33.09949,34.32041,34.980106,35.01621,34.917747,34.287594,31.314054,27.588924,24.474258,23.115488,24.25108,23.870361,21.54995,17.942976,14.7790785,14.857847,14.211283,15.67836,19.38708,22.757746,26.512413,29.929028,31.304207,29.075695,21.815796,17.473642,13.000206,8.966565,6.688821,8.198565,8.2215395,6.0947695,5.0051284,5.7632823,6.810257,11.319796,15.921232,19.098257,20.617847,21.553232,25.69518,29.590977,33.444103,38.422977,46.664207,46.303185,41.744415,37.270977,33.61149,27.940105,22.390156,19.081848,15.133539,10.338462,7.1483083,5.901129,4.84759,4.0992823,3.6890259,3.564308,2.556718,1.8281027,1.5589745,1.6443079,1.6902566,1.8576412,2.4057438,2.7798977,3.0785644,4.0369234,4.2240005,4.8672824,5.8453336,7.125334,8.772923,9.77395,10.20718,10.279386,9.813334,8.241231,7.1581545,6.518154,6.0324106,5.4514875,4.5489235,4.414359,3.498667,2.6157951,2.0250258,1.4211283,1.1158975,0.8369231,0.8402052,1.2077949,1.8445129,2.284308,2.5731285,2.5895386,2.284308,1.6869745,1.1158975,0.79097444,0.7253334,0.8566154,1.0338463,1.3554872,2.2580514,3.0194874,3.43959,3.8432825,3.7415388,3.501949,3.442872,3.9581542,5.5302567,6.2523084,5.159385,3.895795,3.5905645,4.850872,4.07959,4.8311796,5.2053337,4.923077,5.3070774,5.2053337,4.532513,4.588308,4.896821,3.1967182,2.4385643,1.522872,0.90256417,0.63343596,0.36758977,0.38400003,0.23958977,0.13128206,0.101743594,0.049230773,0.052512825,0.11158975,0.10502565,0.032820515,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.036102567,0.0951795,0.14441027,0.15425642,0.108307704,0.11158975,0.10502565,0.101743594,0.108307704,0.10502565,0.11158975,0.108307704,0.08861539,0.06564103,0.07548718,0.1148718,0.128,0.14441027,0.20676924,0.380718,0.69907695,0.7056411,0.84348726,1.083077,0.90256417,1.1979488,1.2242053,1.0896411,0.90256417,0.761436,0.6629744,0.60389745,0.6071795,0.6662565,0.76800007,0.47917953,0.30851284,0.26584616,0.32820517,0.4397949,0.5907693,0.81394875,0.9616411,1.0732309,1.3587693,1.1979488,1.1716924,1.1454359,1.0502565,0.8533334,1.0338463,1.1388719,1.270154,1.4867693,1.7887181,2.6978464,3.495385,4.2994876,5.0051284,5.293949,6.380308,7.177847,7.571693,7.4929237,6.9382567,7.076103,7.3649235,7.5487185,7.716103,8.293744,8.034462,7.351795,7.1581545,7.5388722,7.752206,7.7259493,7.3747697,7.1876926,7.3649235,7.821129,7.256616,7.0104623,7.2369237,7.6996927,7.8047185,7.709539,7.397744,7.213949,7.5388722,8.795898,8.421744,6.9776416,5.9536414,5.796103,5.920821,5.684513,5.142975,4.6966157,4.388103,3.9056413,3.8038976,3.5183592,3.620103,4.086154,4.3060517,3.7021542,3.6824617,3.7743592,3.7809234,3.7940516,3.9187696,4.096,4.663795,5.579488,6.409847,7.529026,6.9120007,6.514872,7.387898,9.665642,11.411694,12.763899,11.930258,9.019077,6.058667,6.308103,5.917539,6.747898,8.809027,10.28595,11.441232,11.877745,11.989334,11.74318,10.696206,6.491898,4.2502565,3.2000003,2.865231,3.0523078,4.7491283,3.3444104,1.8313848,1.5261539,2.0545642,1.9692309,1.7657437,1.5327181,1.3489232,1.2832822,1.6344616,1.6180514,1.8215386,2.2153847,2.1497438,1.8609232,1.591795,1.276718,1.0338463,1.1355898,1.1027694,1.2635899,1.4539489,1.5786668,1.5885129,1.785436,2.806154,3.6069746,3.8137438,3.7251284,3.564308,3.2951798,3.0818465,2.9571285,2.8160002,3.186872,2.9243078,2.8225644,2.9801028,2.806154,2.989949,3.3969233,3.5840003,3.5774362,3.8531284,3.9384618,3.9548721,3.7087183,3.2853336,3.0785644,3.2229745,3.6627696,4.4307694,5.1889234,5.2447186,5.024821,4.827898,4.640821,4.516103,4.5456414,4.647385,5.4580517,6.1407185,6.5411286,7.194257,10.384411,11.9860525,12.678565,13.410462,15.409232,15.786668,15.27795,14.834873,14.834873,15.107284,15.323898,14.87754,14.78236,15.090873,14.867694,14.651078,13.984821,13.193847,12.914873,14.10954,15.235283,15.497848,15.156514,14.460719,13.653335,13.492514,14.306462,14.907078,14.651078,13.410462,13.607386,13.620514,13.587693,13.755078,14.454155,14.034052,12.954257,12.160001,11.716924,10.811078,10.597744,10.371283,10.486155,11.116308,12.2617445,12.104206,12.507898,12.57354,12.1468725,11.828514,10.404103,9.396514,8.342975,7.4174366,7.4436927,7.325539,7.3353853,7.128616,6.820103,6.9842057,7.066257,6.7544622,6.3868723,6.091488,5.796103,6.49518,6.626462,6.012718,5.1626673,5.2414365,5.346462,5.9963083,6.774154,7.463385,8.073847,8.434873,9.360411,10.102155,10.328616,10.118565,10.387693,10.496001,10.630565,10.840616,11.0375395,11.264001,12.524308,13.787898,14.470565,14.444309,14.152206,13.564719,13.22995,13.361232,13.817437,14.244103,14.119386,13.797745,13.604104,13.846975,13.761642,12.189539,10.387693,8.986258,7.9983597,7.128616,5.717334,4.6211286,4.135385,3.9811285,3.9811285,4.4242053,4.6539493,4.663795,5.110154,2.9768207,2.937436,2.9669745,2.733949,2.3236926,2.2121027,2.5435898,2.477949,2.3302567,2.3105643,2.5173335,2.5173335,2.6289232,2.737231,2.9013336,3.3411283,3.3542566,3.7973337,4.5095387,5.093744,4.896821,5.83877,6.0717955,6.1407185,6.186667,5.9667697,5.76,6.373744,6.5903597,6.6560006,8.316719,8.92718,11.881026,13.528616,12.612924,10.269539,18.36308,20.22072,16.321642,9.084719,2.8849232,2.8849232,3.4067695,3.186872,2.2646155,1.9823592,2.3860514,1.910154,1.6738462,1.9922053,2.3958976,2.1267693,2.041436,1.8642052,1.5885129,1.463795,1.5885129,1.3620514,1.3686155,1.6640002,1.785436,1.7985642,1.5622566,1.2209232,0.9878975,1.1585642,0.90256417,0.67282057,0.5513847,0.6432821,1.083077,1.1815386,0.97805136,0.76800007,0.7811283,1.1585642,1.1224617,0.9485129,0.761436,0.6301539,0.58092314,0.33476925,0.28225642,0.25271797,0.17723078,0.09189744,0.06564103,0.04266667,0.02297436,0.026256412,0.07548718,0.11158975,0.31507695,0.43651286,0.47589746,0.67282057,1.4145643,1.847795,2.5928206,3.7415388,4.850872,5.681231,6.5411286,7.24677,7.6242056,7.4765134,7.9885135,7.450257,6.747898,6.314667,6.117744,5.937231,5.330052,4.7622566,4.4373336,4.3027697,4.6802053,5.98318,7.4240007,8.2445135,7.719385,7.000616,5.668103,5.3727183,6.377026,7.5388722,7.939283,7.2992826,6.370462,6.1046157,7.6307697,6.8496413,5.353026,4.529231,4.781949,5.540103,6.5411286,6.73477,7.450257,8.15918,6.5017443,7.3321033,8.470975,9.941334,11.096616,10.620719,9.202872,11.641437,13.551591,13.610668,13.548308,13.403898,17.48677,20.995283,22.997335,26.427078,27.19836,27.746464,26.368002,24.22154,25.344002,25.235695,27.16554,28.435694,28.514463,29.052721,27.539694,26.420515,26.505848,26.811079,24.566156,25.078156,27.779284,29.459694,28.918156,26.978464,26.233438,25.75426,25.27836,24.641644,23.78831,24.81231,25.6919,26.04636,25.924925,25.80349,26.41395,27.204926,26.676516,24.963284,23.863796,24.20513,24.080412,23.079386,21.415386,19.912207,17.398155,17.109335,17.040411,16.439796,15.793232,17.391592,18.907898,19.70872,19.492104,18.294155,17.378464,16.722052,16.810667,17.772308,19.347694,19.505232,18.858667,18.681437,19.396925,20.568617,21.861746,23.732515,25.11754,25.947899,27.145847,28.205952,28.18954,27.858053,27.792412,28.366772,28.816412,30.129232,31.556925,33.16513,35.826874,38.94154,39.955696,39.94913,39.43385,38.36062,38.629745,36.4439,32.43323,27.913849,24.887796,24.605541,23.335386,21.792822,19.685745,15.730873,15.488001,14.959591,15.258258,16.984617,20.217438,23.318975,26.932514,30.076721,30.605131,25.222567,20.93949,14.529642,9.147078,6.9152827,8.940309,7.3058467,5.973334,5.3070774,5.602462,7.0793853,9.557334,12.934566,16.259283,18.379488,17.913437,22.711796,25.990566,28.724516,32.8238,41.124107,43.27057,38.452515,32.246155,26.962053,21.651693,18.17272,14.36554,10.305642,6.5969234,4.3651285,3.4002054,3.186872,3.4067695,3.7218463,3.7842054,2.9407182,2.2186668,1.9495386,2.0217438,1.8609232,2.556718,2.540308,2.5337439,2.793026,3.0982566,3.9778464,4.7622566,5.940513,7.565129,9.26195,10.994873,11.894155,11.674257,10.607591,9.521232,8.362667,7.466667,6.3376417,5.0510774,4.2568207,3.43959,2.4484105,1.9396925,2.1792822,3.0194874,2.7536411,1.7887181,1.2274873,1.3193847,1.463795,1.5622566,1.7526156,2.1530259,2.3958976,1.6016412,1.0404103,0.67938465,0.5284103,0.5349744,0.5940513,0.9353847,1.9462565,2.989949,3.6332312,3.6463592,2.8521028,2.9013336,3.3280003,4.4438977,7.325539,5.3234878,3.69559,2.9440002,2.802872,2.228513,3.3509746,4.1714873,4.8311796,5.0642056,4.197744,5.504,5.481026,5.077334,4.2436924,1.9364104,0.69251287,0.45620516,0.6268718,0.67282057,0.12143591,0.84348726,0.43651286,0.03938462,0.02297436,0.0,0.013128206,0.016410258,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.036102567,0.108307704,0.15097436,0.15425642,0.16738462,0.0951795,0.06564103,0.06235898,0.06564103,0.09189744,0.07876924,0.0951795,0.118153855,0.13784617,0.13784617,0.13784617,0.118153855,0.15097436,0.2100513,0.19692309,0.4660513,0.6071795,0.7187693,0.8172308,0.8533334,0.90256417,0.8336411,0.92553854,1.0666667,0.74830776,0.40697438,0.26584616,0.3446154,0.5481026,0.67282057,0.34133336,0.23958977,0.27241027,0.35446155,0.4266667,0.49887183,0.67282057,0.7844103,0.8566154,1.1126155,1.1027694,1.1520001,1.1290257,0.9878975,0.79425645,0.96492314,1.079795,1.1782565,1.3259488,1.6180514,2.0086155,2.5074873,3.1540515,3.9286156,4.7458467,5.8814363,6.8496413,7.4436927,7.709539,7.965539,7.4765134,7.529026,7.719385,7.8802056,8.086975,7.90318,7.8112826,7.752206,7.6898465,7.6307697,7.460103,7.1515903,6.892308,6.918565,7.4929237,7.5881033,7.394462,7.394462,7.5585647,7.3386674,7.4141545,7.7423596,7.522462,7.1483083,8.208411,8.001641,6.9152827,6.0356927,5.723898,5.61559,4.8344617,4.637539,4.457026,4.2240005,4.394667,3.7842054,3.4297438,3.5216413,3.7940516,3.5249233,2.937436,2.9472823,3.2361028,3.511795,3.5249233,3.7185643,4.0434875,4.6605134,5.431795,5.920821,6.9809237,6.633026,6.87918,8.237949,9.750975,11.946668,13.4859495,12.160001,8.241231,4.4701543,6.157129,6.1538467,6.7840004,8.746667,11.139283,7.39118,8.743385,8.805744,6.422975,5.691077,3.3247182,2.8127182,2.4484105,2.0644104,3.0523078,6.944821,3.570872,1.0666667,1.6278975,1.4802053,1.6508719,1.7591796,1.5195899,1.148718,1.3423591,1.7329233,1.7132308,1.7066668,1.8445129,1.9528207,1.7329233,1.5688206,1.3259488,1.086359,1.1585642,1.0502565,1.1946667,1.3784616,1.4900514,1.5261539,2.0250258,2.7634873,3.3280003,3.5183592,3.370667,3.446154,3.2984617,3.18359,3.0358977,2.487795,2.7175386,2.8422565,2.865231,2.8455386,2.868513,3.1507695,3.5872824,3.6463592,3.4756925,3.892513,4.3552823,4.204308,3.7415388,3.2262566,2.8849232,3.0194874,3.2820516,3.9351797,4.8311796,5.4153852,5.4908724,5.152821,4.9854364,5.044513,4.8377438,5.2512827,6.4722056,7.3714876,7.899898,9.110975,10.610872,11.59877,12.498053,13.627078,15.212309,16.226463,16.65313,16.52513,16.15754,16.144411,16.643284,16.275694,15.494565,14.808617,14.769232,14.759386,14.516514,13.8765135,13.522053,14.998976,17.503181,17.42113,16.646564,16.108309,15.776822,15.556924,16.216616,16.571077,16.36431,16.265848,15.350155,15.304206,15.714462,16.003283,15.442053,14.867694,13.873232,13.170873,12.826258,12.251899,11.812103,11.244308,11.234463,11.979488,13.213539,13.446565,13.824001,13.446565,12.511181,12.3306675,11.011283,9.810052,8.474257,7.4436927,7.857231,8.004924,7.9491286,7.351795,6.5083084,6.363898,6.669129,6.8365135,6.951385,6.8562055,6.1505647,6.1374364,6.124308,5.874872,5.546667,5.7074876,5.681231,6.1341543,6.9645133,7.9163084,8.576,9.357129,10.164514,10.505847,10.328616,10.010257,10.180923,10.755282,11.424822,11.844924,11.611898,11.85477,12.714667,13.587693,14.066873,13.932309,14.480412,13.866668,13.348104,13.341539,13.426873,13.988104,14.230975,14.204719,13.883078,13.138052,13.065847,11.516719,10.069334,9.196308,8.254359,6.6428723,5.142975,4.325744,4.164923,4.0434875,4.128821,4.5062566,4.5489235,4.378257,4.8672824,3.1967182,3.0424619,3.0162053,2.7963078,2.3794873,2.103795,2.1989746,2.1924105,2.2022567,2.2646155,2.3466668,2.4746668,2.7044106,2.8291285,2.8849232,3.1573336,3.4724104,3.9417439,4.529231,5.077334,5.3005133,5.7632823,5.664821,5.85518,6.3310776,6.245744,6.038975,6.186667,6.3967185,6.816821,8.04759,8.36595,10.902975,12.35036,12.396309,13.722258,24.208412,24.257643,18.028309,9.668923,3.31159,3.114667,3.121231,2.7503593,1.9561027,1.2274873,1.2012309,1.0272821,1.1388719,1.522872,1.7001027,1.6180514,1.6738462,1.657436,1.5786668,1.6607181,1.5589745,1.5163078,1.6804104,1.8970258,1.7362052,1.7493335,1.8281027,1.7690258,1.5195899,1.1716924,1.1881026,0.90256417,0.761436,0.892718,1.1093334,1.0305642,1.014154,1.0732309,1.1881026,1.3423591,1.1191796,0.8992821,0.7417436,0.6268718,0.46933338,0.4594872,0.3511795,0.24943592,0.190359,0.10502565,0.098461546,0.049230773,0.016410258,0.02297436,0.052512825,0.118153855,0.25271797,0.380718,0.58092314,1.0994873,2.2055387,2.868513,3.6594875,4.7392826,5.8420515,6.7085133,7.8408213,8.612103,8.884514,8.989539,9.074872,8.786052,8.516924,8.356103,8.070564,7.6635904,6.872616,6.2588725,6.665847,9.196308,11.421539,10.059488,9.291488,9.980719,9.662359,8.776206,7.936001,7.75877,8.441437,9.747693,10.745437,10.259693,9.002667,7.8145647,7.6898465,6.810257,5.366154,4.076308,3.5380516,4.197744,4.640821,5.284103,6.422975,7.2369237,5.792821,5.8912826,7.2303596,8.421744,9.110975,9.974154,10.889847,10.962052,10.8537445,11.063796,11.890873,12.806565,15.501129,18.907898,23.033438,28.954258,29.860106,28.232206,26.837336,26.666668,26.919386,25.189745,26.870155,28.035284,27.979488,29.200413,28.084515,28.465233,28.544003,27.349335,24.713848,24.982977,25.491693,26.646976,27.874464,27.6119,25.091284,24.218258,24.582565,25.472002,25.875694,25.70831,26.341745,26.689644,26.817642,27.926977,26.807796,27.044106,26.597746,25.091284,23.814566,23.532309,22.849644,22.002874,20.919796,19.193438,16.932104,16.758156,16.78113,16.288822,15.721026,15.287796,16.347898,17.604925,18.162872,17.513027,17.283283,17.51959,17.91672,18.372925,18.970259,18.01518,18.159592,18.944002,20.040207,21.251284,22.994053,24.677746,25.097849,24.641644,25.291489,26.118567,26.640411,26.535387,25.961027,25.557335,25.728003,27.414976,29.952002,33.155285,37.3399,40.36595,41.7838,41.389954,40.165745,40.300312,40.786053,39.348515,35.462566,30.532925,27.913849,26.489437,24.01149,21.648413,19.157335,14.890668,16.226463,16.17395,16.311796,17.332514,19.032618,20.073027,23.40759,27.398565,29.312002,25.294771,20.729437,14.828309,10.148104,7.899898,7.9524107,6.6002054,6.8233852,6.413129,5.618872,7.1548724,8.43159,11.753027,14.9628725,16.561232,15.717745,19.19672,22.357334,25.222567,28.176413,31.954054,33.184822,29.93231,24.546463,19.301744,16.403694,12.514462,9.42277,6.2227697,3.308308,2.3729234,2.2121027,2.0644104,2.3794873,3.2131286,4.2601027,3.1048207,2.1267693,1.6902566,1.8773335,2.5206156,3.4789746,2.9997952,2.7536411,3.4166157,4.6605134,4.7491283,4.8607183,5.8880005,7.817847,9.750975,11.894155,13.095386,13.289026,12.42913,10.473026,8.651488,7.1515903,5.664821,4.2830772,3.4888208,2.8258464,2.1300514,1.719795,1.591795,1.4112822,1.6672822,1.6935385,1.7066668,1.8149745,2.0020514,2.1497438,2.5764105,2.678154,2.3794873,2.1530259,2.097231,1.4112822,0.71548724,0.3708718,0.4594872,0.764718,1.2570257,1.7296412,2.0184617,2.0118976,2.0578463,2.9604106,3.6463592,3.7710772,3.7218463,7.8539495,6.9776416,6.4590774,6.6560006,2.8980515,5.8978467,4.9887185,4.2962055,5.2644105,6.672411,4.8344617,3.2886157,2.3204105,1.7132308,0.75487185,0.318359,0.24615386,0.36430773,0.41025645,0.036102567,0.17066668,0.0951795,0.01969231,0.016410258,0.013128206,0.0032820515,0.0032820515,0.006564103,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.036102567,0.118153855,0.18051283,0.22646156,0.3249231,0.3117949,0.2855385,0.20348719,0.12471796,0.17723078,0.16410258,0.13456412,0.17394873,0.23630771,0.13784617,0.108307704,0.11158975,0.14769232,0.17723078,0.12471796,0.27569234,0.52512825,0.72861546,0.827077,0.8533334,0.6104616,0.57764107,0.67938465,0.7417436,0.49230772,0.4135385,0.4266667,0.47589746,0.49887183,0.4266667,0.27241027,0.2231795,0.24615386,0.2986667,0.35446155,0.34789747,0.512,0.6826667,0.8402052,1.0765129,0.9878975,1.0338463,1.0404103,0.9321026,0.7581539,0.9682052,1.2176411,1.4309745,1.5786668,1.6672822,1.8018463,2.15959,2.6683078,3.308308,4.086154,5.671385,6.8266673,7.456821,7.755488,8.198565,7.5520005,6.941539,6.9382567,7.5191803,8.086975,7.4732313,7.384616,7.397744,7.3452315,7.325539,7.0957956,6.7282057,6.436103,6.3507695,6.5017443,7.020308,6.7544622,6.665847,6.9809237,7.181129,7.3616414,8.113232,8.326565,7.9195905,7.830975,7.7981544,7.1023593,6.377026,5.8092313,5.113436,4.8607183,4.5029745,4.3060517,4.2305646,3.9417439,3.6660516,3.570872,3.6036925,3.6726158,3.6463592,3.255795,3.2196925,3.3017437,3.367385,3.3903592,3.8695388,4.4110775,5.0510774,5.6352825,5.8092313,6.432821,6.4065647,6.918565,8.392206,10.482873,12.3766165,12.806565,11.789129,9.216001,4.84759,5.21518,7.0104623,8.356103,8.6580515,8.598975,6.2687182,7.709539,7.240206,4.7458467,5.7042055,4.781949,3.190154,2.1202054,1.9692309,2.3302567,5.346462,2.8717952,1.4572309,2.353231,1.4933335,1.5360001,1.6475899,1.467077,1.1913847,1.5622566,1.5721027,1.595077,1.6869745,1.7329233,1.4539489,1.6738462,1.5885129,1.3981539,1.2964103,1.4769232,1.522872,1.5392822,1.591795,1.6082052,1.3915899,2.0184617,2.3926156,2.7208207,2.9735386,2.8947694,3.4592824,3.5347695,3.4789746,3.4264617,3.318154,3.1967182,3.3476925,3.0326157,2.5206156,3.1015387,3.31159,3.5347695,3.5413337,3.4034874,3.4756925,3.754667,3.7776413,3.6594875,3.5347695,3.5544617,3.4264617,3.5478978,3.6496413,3.7152824,3.9876926,4.5587697,4.969026,5.2381544,5.2676926,4.824616,5.346462,6.9677954,8.303591,9.094564,10.197334,11.969642,13.167591,13.830565,14.470565,16.068924,16.945232,17.316103,17.58195,17.690258,17.11918,17.785437,16.925539,16.587488,17.270155,17.906874,16.800821,16.551386,16.183796,15.625848,15.694771,16.95836,17.667284,17.795284,17.381744,16.534975,16.33477,17.004309,17.385027,17.381744,17.985641,16.925539,16.331488,16.636719,17.237335,16.49231,15.527386,14.726565,13.912617,13.2562065,13.279181,13.443283,13.203693,12.99036,13.259488,14.470565,15.212309,14.9628725,13.915898,12.724514,12.511181,11.506873,10.473026,9.508103,8.809027,8.687591,8.697436,8.953437,8.408616,7.174565,6.521436,6.885744,7.315693,7.4765134,7.253334,6.7610264,5.907693,5.5171285,5.5926156,5.9503593,6.2063594,6.426257,6.7282057,7.4207187,8.39877,9.137232,10.220308,10.929232,11.30995,11.365745,11.047385,10.965334,11.313231,12.07795,12.816411,12.675283,13.239796,13.879796,14.01436,13.702565,13.627078,14.332719,14.234258,14.03077,13.952001,13.745232,13.778052,13.574565,13.298873,12.983796,12.504617,11.835078,11.191795,10.233437,9.025641,8.04759,6.629744,5.5532312,4.7261543,4.197744,4.1517954,3.761231,3.8498464,4.073026,4.33559,4.7950773,2.5173335,2.6289232,2.5993848,2.4582565,2.2416413,1.975795,1.9003079,2.048,2.1956925,2.28759,2.4320002,2.540308,2.7864618,2.8882053,2.8455386,2.937436,3.387077,3.9909747,4.565334,5.07077,5.612308,5.684513,5.901129,6.242462,6.488616,6.235898,6.4754877,6.7314878,6.8693337,7.174565,8.356103,9.009232,10.555078,11.513436,12.780309,17.6279,27.503592,25.51467,17.066668,7.781744,3.501949,3.570872,3.508513,2.92759,1.9232821,1.0666667,1.0568206,0.9189744,0.9124103,1.083077,1.2406155,1.0502565,1.142154,1.211077,1.2307693,1.4605129,1.3915899,1.4802053,1.6640002,1.8018463,1.6771283,1.7427694,2.1825643,2.3860514,2.0808206,1.339077,1.1191796,0.92225647,0.8172308,0.8172308,0.892718,1.1027694,1.1257436,1.0962052,1.1060513,1.1946667,1.1093334,1.014154,0.8172308,0.5973334,0.5874872,0.6465641,0.4955898,0.3052308,0.16082053,0.06235898,0.052512825,0.036102567,0.02297436,0.026256412,0.026256412,0.08533334,0.19692309,0.33805132,0.69251287,1.6278975,2.6978464,3.2951798,3.9745643,4.923077,5.940513,7.0990777,7.77518,8.786052,10.279386,11.739899,12.074668,12.3076935,12.626052,12.836103,12.3306675,11.2672825,10.364718,9.655796,9.472001,10.459898,14.089848,13.019898,10.781539,9.32759,9.028924,9.370257,8.854975,8.743385,9.435898,10.463181,11.172104,11.040821,10.364718,9.570462,9.225847,8.966565,7.8539495,5.7042055,3.7185643,4.457026,4.1156926,3.8465643,4.4734364,5.546667,5.3398976,4.962462,5.474462,5.9602056,6.485334,8.090257,11.076924,11.933539,11.382154,10.738873,11.913847,13.062565,15.205745,17.142155,19.22954,23.40759,26.77826,29.321848,29.843695,28.793438,28.274874,26.341745,27.034258,28.612925,30.148926,31.524105,29.266054,28.855797,28.85908,28.245335,26.397541,25.924925,25.642668,26.482874,27.785849,27.323078,25.284925,24.119797,24.244514,25.028925,24.805746,25.701746,27.211489,28.084515,28.120617,28.17313,27.72349,27.759592,26.922668,25.232412,24.106668,23.299284,22.764309,22.127592,20.95918,18.766771,16.728617,16.003283,15.8654375,15.75713,15.281232,14.260514,14.503386,15.655386,16.836924,16.66954,16.02954,16.597334,17.736206,18.819284,19.232822,18.130053,18.395899,19.19672,20.115694,21.139694,23.213951,24.871386,25.222567,24.149336,22.327797,23.578259,24.451284,25.088001,25.531078,25.72472,25.96431,27.053951,29.216824,32.39713,36.28308,40.39221,42.643696,42.706055,41.58031,41.609848,41.83303,40.576004,37.300514,33.00103,30.208002,28.215797,25.176617,22.38031,19.849848,16.354464,16.521847,16.600616,17.09949,18.087385,19.213129,20.565334,23.341951,26.345028,27.421541,23.483078,19.495386,14.621539,10.791386,8.65477,7.5881033,6.76759,7.253334,7.250052,6.7314878,7.456821,8.01477,10.9456415,14.670771,17.174976,16.009848,17.043694,18.78318,21.287386,23.913027,25.334156,25.573746,21.546669,16.544823,12.731078,11.155693,8.687591,6.452513,4.0336413,1.8740515,1.273436,1.6902566,1.6738462,1.9035898,2.5238976,3.1540515,2.5993848,1.9167181,1.585231,1.9429746,3.190154,3.826872,3.314872,3.006359,3.4756925,4.529231,4.345436,4.647385,5.76,7.581539,9.570462,11.004719,11.657847,11.713642,11.07036,9.373539,7.9195905,6.452513,4.972308,3.564308,2.3893335,1.8182565,1.7755898,1.595077,1.1618463,0.90584624,0.9747693,1.3456411,1.5327181,1.5556924,1.972513,2.048,2.3860514,2.6387694,2.6387694,2.409026,1.8674873,1.3817437,0.85005134,0.4004103,0.41682056,0.6662565,0.97805136,1.3128207,1.6082052,1.785436,1.4769232,2.5698464,3.5446157,4.0041027,4.673641,8.211693,6.5805135,5.024821,4.6112823,2.2350771,3.6004105,2.937436,2.5107694,3.2131286,4.57518,3.1442053,1.9528207,1.083077,0.56451285,0.36758977,0.15753847,0.098461546,0.15097436,0.190359,0.016410258,0.0032820515,0.0032820515,0.006564103,0.006564103,0.016410258,0.0032820515,0.0,0.0032820515,0.026256412,0.101743594,0.101743594,0.03938462,0.0,0.0,0.0,0.029538464,0.14441027,0.18707694,0.17723078,0.28225642,0.27569234,0.27897438,0.28225642,0.27897438,0.28882053,0.32164106,0.24287182,0.20676924,0.21989745,0.16410258,0.15097436,0.17066668,0.16738462,0.13128206,0.108307704,0.20676924,0.39712822,0.5940513,0.69251287,0.56123084,0.4135385,0.380718,0.39056414,0.380718,0.318359,0.3708718,0.44964105,0.46276927,0.39384618,0.30194873,0.2297436,0.19692309,0.2100513,0.25271797,0.28225642,0.32164106,0.47589746,0.64000005,0.8008206,1.0404103,0.88615394,0.85005134,0.8566154,0.82379496,0.67282057,1.0404103,1.2504616,1.3489232,1.4112822,1.5491283,1.9528207,2.3269746,2.7569232,3.2722054,3.8564105,5.2381544,6.5870776,7.4765134,7.778462,7.6603084,7.1876926,6.813539,6.921847,7.427283,7.748924,7.2336416,7.0137444,6.885744,6.8627696,7.200821,7.273026,6.882462,6.616616,6.62318,6.62318,7.0334363,6.705231,6.557539,6.9152827,7.53559,8.182155,8.579283,8.572719,8.293744,8.155898,7.650462,7.463385,6.9809237,6.0816417,5.146257,4.7655387,4.4373336,4.1813335,3.8564105,3.1606157,3.3608208,3.4625645,3.4330258,3.3017437,3.1540515,2.8356924,2.8849232,2.993231,3.121231,3.511795,4.2962055,4.598154,4.923077,5.330052,5.435077,5.661539,6.311385,7.2237954,8.516924,10.57477,11.697231,11.71036,10.788103,8.841846,5.5105643,5.2414365,6.9842057,7.906462,7.50277,7.6077952,6.180103,7.1056414,6.5903597,4.7589746,5.661539,4.9821544,3.114667,1.8806155,2.03159,3.249231,5.58277,3.131077,1.4966155,2.0578463,1.972513,1.7132308,1.7362052,1.5688206,1.339077,1.7920002,1.4933335,1.4900514,1.6410258,1.7001027,1.3357949,1.5786668,1.4145643,1.3850257,1.5458462,1.4736412,1.4933335,1.5327181,1.5655385,1.5753847,1.5491283,2.0709746,2.2646155,2.4713848,2.7044106,2.6584618,3.4133337,3.3050258,3.18359,3.2623591,3.0949745,2.733949,3.0030773,2.917744,2.5796926,3.1671798,3.2820516,3.4756925,3.7382567,3.7940516,3.0687182,3.0162053,3.2328207,3.245949,3.0982566,3.3378465,3.626667,3.8564105,3.945026,3.9154875,3.9056413,4.71959,5.3037953,5.405539,5.2676926,5.654975,6.5936418,7.8047185,9.242257,10.752001,12.097642,13.069129,13.732103,14.355694,15.307488,17.024002,17.900309,17.585232,17.250463,17.385027,17.811693,17.877335,17.394873,17.660719,18.665028,19.104822,17.739489,17.26031,17.61477,18.28431,18.258053,18.697847,19.075283,19.009642,18.658463,18.727386,17.956104,18.225233,18.546873,18.694565,19.213129,18.582975,17.194668,16.745028,17.266872,17.112617,16.357744,15.337027,14.79877,14.831591,14.8709755,14.486976,14.135796,13.801026,13.994668,15.737437,16.31836,16.006565,14.805334,13.289026,12.586668,12.265027,11.946668,11.323078,10.476309,9.875693,9.603283,9.465437,8.694155,7.397744,6.5903597,6.951385,7.653744,7.955693,7.785026,7.762052,6.0652313,5.4416413,5.691077,6.380308,6.8463597,7.017026,7.4929237,8.211693,8.953437,9.350565,10.525539,11.227899,11.815386,12.160001,11.634872,11.483898,11.667693,12.173129,12.793437,13.141335,13.561437,14.093129,14.273643,14.063591,13.843694,14.500104,14.552616,14.523078,14.490257,14.099693,13.994668,13.338258,12.770463,12.340514,11.529847,10.998155,10.709334,9.957745,8.707283,7.5913854,6.1308722,5.4416413,5.149539,4.9427695,4.565334,4.007385,3.748103,3.8301542,4.089436,4.1452312,2.4516926,2.546872,2.5140514,2.409026,2.2744617,2.1398976,2.038154,2.100513,2.15959,2.2383592,2.5435898,2.733949,2.9078977,2.937436,2.8422565,2.793026,3.2065644,3.8859491,4.532513,5.093744,5.7468724,5.8157954,6.2818465,6.5312824,6.416411,6.242462,6.8332314,6.951385,7.0498466,7.50277,8.576,9.865847,11.08677,11.805539,13.35795,18.835693,25.590157,21.96677,13.476104,5.5762057,3.6660516,3.4921029,3.058872,2.3335385,1.4834872,0.892718,1.020718,1.0404103,0.9944616,0.9714873,1.1257436,0.8763078,0.8598975,0.90256417,0.9616411,1.1093334,1.1651284,1.3292309,1.5589745,1.7690258,1.8051283,1.8642052,2.1103592,2.2088206,1.9626669,1.3226668,1.0469744,1.0633847,0.9682052,0.71548724,0.636718,0.892718,0.92553854,0.9353847,0.9911796,1.014154,1.1684103,1.1126155,0.90912825,0.69907695,0.72861546,0.6826667,0.5349744,0.3314872,0.13784617,0.04266667,0.029538464,0.036102567,0.055794876,0.07548718,0.08205129,0.072205134,0.15097436,0.33805132,0.78769237,1.785436,2.7700515,3.4921029,4.378257,5.504,6.626462,7.778462,8.539898,10.174359,12.793437,15.366566,15.986873,16.019693,16.141129,16.20349,15.238565,13.75836,12.452104,11.546257,11.113027,11.063796,14.001232,14.106257,12.163283,9.613129,8.546462,9.462154,9.068309,8.973129,9.757539,10.988309,11.35918,11.405129,11.234463,10.988309,10.807796,10.617436,9.235693,6.7544622,4.2568207,3.8498464,3.373949,2.8291285,2.8980515,3.5938463,4.266667,3.9647183,4.0041027,4.3618464,5.225026,6.9743595,9.3768215,11.989334,13.049437,13.033027,14.641232,16.200207,18.54359,19.715284,19.928617,21.563078,22.948105,25.878977,27.841642,28.245335,28.402874,26.866875,27.221336,29.607388,32.741745,33.893745,31.291079,29.866669,29.256207,28.882053,27.959797,26.505848,26.305643,27.293541,28.52431,28.160002,27.158976,25.67549,24.946875,25.088001,25.097849,26.34831,28.104208,29.512207,30.034054,29.449848,28.793438,28.074669,26.873438,25.353848,24.293745,23.43713,23.072823,22.475489,21.10031,18.60595,17.165129,16.216616,16.02954,16.082052,15.084309,14.099693,14.066873,14.697027,15.501129,15.803078,14.844719,15.205745,16.666258,18.33354,18.638771,17.723078,18.107079,18.822565,19.442873,20.059898,22.002874,23.056412,23.102362,21.973335,19.452719,21.392412,22.698668,24.01477,25.478565,26.702772,27.076925,27.19508,28.406157,30.913643,33.792004,38.03898,40.98626,42.289234,42.423798,42.702774,42.108723,40.615387,37.970055,34.579697,31.510977,29.056002,25.888823,23.05313,20.647387,17.801847,16.833643,17.286566,18.189129,19.045746,19.85313,21.50072,23.072823,24.664618,24.864822,20.762259,17.664001,14.070155,11.546257,10.043077,7.8802056,6.7577443,7.6734366,8.342975,8.054154,7.6701546,7.817847,9.911796,13.883078,17.634462,17.033848,16.597334,16.262566,18.070976,21.11672,21.54995,20.913233,16.259283,11.500309,8.598975,7.584821,6.0685134,4.466872,2.92759,1.6640002,0.9747693,1.273436,1.3883078,1.5261539,1.7099489,1.7920002,1.7329233,1.4211283,1.332513,1.913436,3.6036925,3.9680004,3.564308,3.1409233,3.1081028,3.5413337,3.511795,4.082872,5.2676926,6.810257,8.192,8.375795,8.323282,8.172308,7.7718983,6.695385,5.786257,4.71959,3.7809234,2.8816411,1.5360001,1.2570257,1.4769232,1.3686155,0.8960001,0.79097444,0.7089231,0.9878975,1.1946667,1.3193847,1.7591796,1.5786668,1.6508719,1.910154,2.1103592,1.8281027,1.2176411,1.1126155,0.9682052,0.67938465,0.58420515,0.5940513,0.84348726,1.1224617,1.3653334,1.657436,1.2800001,1.9298463,2.6453335,3.501949,5.5991797,6.170257,4.453744,3.5511796,3.5938463,1.7263591,1.6508719,1.4605129,1.4900514,1.8740515,2.546872,1.6738462,1.0043077,0.49230772,0.18379489,0.20020515,0.07548718,0.049230773,0.072205134,0.08205129,0.009846155,0.0032820515,0.0,0.0,0.0032820515,0.009846155,0.0032820515,0.0,0.0,0.01969231,0.101743594,0.101743594,0.059076928,0.01969231,0.0,0.0,0.01969231,0.108307704,0.13784617,0.1148718,0.19692309,0.24615386,0.27897438,0.30194873,0.30194873,0.27897438,0.34789747,0.3446154,0.3052308,0.25928208,0.23302566,0.25271797,0.22646156,0.17394873,0.13128206,0.13784617,0.19692309,0.29538465,0.446359,0.5546667,0.39712822,0.4004103,0.32820517,0.24615386,0.2231795,0.33476925,0.33476925,0.380718,0.3708718,0.2986667,0.23958977,0.23958977,0.20676924,0.20020515,0.2231795,0.23302566,0.28225642,0.4266667,0.574359,0.7187693,0.9353847,0.8369231,0.7253334,0.67282057,0.6662565,0.5940513,0.9911796,1.2668719,1.3883078,1.4178462,1.5327181,2.0020514,2.3958976,2.8291285,3.314872,3.761231,4.772103,5.8223596,6.6625648,7.0826674,6.9021544,6.8332314,6.9349747,7.174565,7.39118,7.27959,7.24677,7.056411,6.885744,6.925129,7.384616,7.568411,7.2205133,6.8660517,6.76759,6.928411,7.197539,6.8332314,6.816821,7.381334,8.041026,8.562873,8.316719,7.7981544,7.456821,7.7357955,7.453539,7.4830775,7.1187696,6.232616,5.2676926,4.8344617,4.466872,4.141949,3.7316926,2.9965131,3.2164104,3.4658465,3.5774362,3.4822567,3.2098465,2.9833848,2.9604106,2.986667,3.1507695,3.7743592,4.4012313,4.33559,4.381539,4.7491283,5.0642056,5.362872,6.8233852,8.004924,8.648206,9.665642,10.95877,10.676514,9.29477,7.273026,5.07077,5.651693,6.514872,6.5903597,6.498462,8.54318,7.171283,7.0334363,5.9930263,4.2863593,4.4964104,4.125539,3.3312824,2.8455386,3.255795,5.0215387,6.678975,3.6102567,1.4441026,1.719795,1.8674873,1.7755898,1.9265642,1.782154,1.4998976,1.9265642,1.7591796,1.6475899,1.6804104,1.7493335,1.5392822,1.585231,1.4211283,1.5589745,1.8773335,1.6213335,1.5556924,1.5753847,1.5589745,1.5491283,1.7329233,2.0939488,2.169436,2.3696413,2.7208207,2.8914874,3.3575387,3.2328207,3.062154,3.0194874,2.930872,2.5928206,2.868513,2.993231,2.9505644,3.4560003,3.495385,3.5183592,3.6627696,3.5971284,2.5337439,2.3729234,2.6847181,2.809436,2.7733335,3.3017437,3.9417439,4.1583595,4.266667,4.414359,4.5587697,5.346462,5.8092313,5.9569235,6.088206,6.803693,7.4075904,8.41518,10.006975,11.98277,13.764924,14.221129,14.444309,15.113848,16.374155,17.821539,18.432001,17.719797,17.270155,17.680412,18.582975,18.084105,18.376207,18.884924,19.324718,19.689028,19.032618,18.68472,19.213129,20.171488,20.115694,19.669334,19.593847,19.465847,19.442873,20.279797,19.222977,18.802874,18.81272,19.06872,19.416616,18.838976,17.270155,16.482462,16.800821,17.06995,16.66954,16.164104,16.479181,17.224207,16.695797,15.386257,14.713437,14.322873,14.624822,16.78113,17.027283,16.49559,15.435489,14.162052,13.072412,13.00677,13.02318,12.626052,11.749744,10.778257,10.374565,9.665642,8.530052,7.194257,6.242462,7.0826674,7.824411,8.054154,7.830975,7.6767187,6.0652313,5.5236926,5.858462,6.6428723,7.2237954,7.194257,7.8802056,8.700719,9.3078985,9.590155,10.71918,11.716924,12.534155,12.852514,12.068104,11.841642,12.06154,12.389745,12.701539,13.092104,13.292309,13.909334,14.240822,14.12595,13.922462,14.677335,14.841437,14.742975,14.539488,14.227694,14.14236,13.410462,12.790154,12.212514,10.79795,10.512411,10.180923,9.481847,8.4053335,7.2336416,5.8518977,5.3234878,5.280821,5.297231,4.8836927,4.4438977,3.95159,3.7251284,3.7087183,3.4658465,3.045744,2.878359,2.8389745,2.740513,2.5993848,2.6486156,2.5304618,2.3236926,2.166154,2.2022567,2.556718,2.8849232,2.9604106,2.917744,2.8488207,2.793026,3.0916924,3.6726158,4.3716927,5.0576415,5.618872,5.9634876,6.4623594,6.5280004,6.2851286,6.567385,7.1548724,6.8266673,6.944821,7.7718983,8.454565,10.407386,11.963078,12.471796,13.033027,16.489027,19.5479,15.363283,8.851693,3.9220517,3.4560003,2.802872,2.0217438,1.4605129,1.1848207,0.9878975,1.0535386,1.2406155,1.2898463,1.204513,1.2438976,1.0633847,0.92553854,0.892718,0.93866676,0.9517949,1.0896411,1.2964103,1.6082052,1.9331284,2.0644104,2.0578463,1.7723079,1.5261539,1.3817437,1.1520001,1.1060513,1.2438976,1.0994873,0.69251287,0.508718,0.46933338,0.512,0.7187693,0.9616411,0.92553854,1.2504616,1.1520001,1.020718,0.955077,0.74830776,0.5349744,0.43323082,0.318359,0.17066668,0.08205129,0.049230773,0.049230773,0.08205129,0.128,0.15753847,0.07876924,0.118153855,0.34133336,0.8008206,1.5392822,2.5304618,3.5249233,4.841026,6.4623594,8.011488,8.960001,10.371283,12.540719,15.402668,18.520617,19.403488,18.710976,17.910154,17.240616,15.711181,14.309745,12.498053,11.35918,11.254155,11.818667,12.842668,13.59754,13.052719,11.260718,9.360411,9.6,9.225847,9.252103,10.023385,11.218052,11.204924,11.011283,10.952206,11.063796,11.113027,10.210463,8.418462,6.6034875,4.8672824,2.540308,2.3302567,2.2153847,2.0118976,1.972513,2.802872,2.9505644,3.1376412,3.8301542,5.034667,6.3179493,6.816821,10.512411,13.873232,15.95077,18.41231,20.614565,23.729233,25.478565,25.550772,25.59672,21.48759,19.610258,20.949335,24.280617,26.2039,25.96431,26.978464,30.0439,33.847797,34.989952,33.22421,31.448618,29.952002,28.944412,28.553848,26.679796,26.906258,28.248617,29.709131,30.267078,30.244104,28.517746,26.752003,26.0759,27.076925,27.536413,28.655592,30.313028,31.766977,31.668516,29.659899,27.946669,26.627285,25.501541,24.06072,23.584822,23.315695,22.724924,21.395695,19.016207,18.04472,17.38831,17.385027,17.348925,15.556924,14.680616,14.772514,14.841437,14.726565,15.117129,14.293334,14.214565,15.27795,16.761436,16.843489,16.210052,16.889437,17.69354,18.090668,18.20554,19.462566,19.620104,19.11795,18.22195,17.030565,19.291899,20.854155,22.390156,24.241232,26.427078,27.181952,26.663387,27.073643,28.842669,30.657644,33.851078,37.316925,40.277336,42.436928,43.979492,42.486156,40.297028,37.782978,34.993233,31.668516,28.629335,25.859283,23.299284,20.8279,18.264616,17.014154,17.929848,18.960411,19.40677,19.899078,21.376001,21.707489,22.38031,22.46236,18.625643,16.311796,13.59754,12.025436,11.099898,8.27077,6.4065647,7.890052,9.025641,8.4972315,7.3649235,7.640616,8.779488,12.337232,16.840206,17.778873,17.188105,15.081027,15.924514,19.19672,19.383797,18.688002,14.769232,10.433641,7.433847,6.482052,4.6572313,3.3476925,2.7306669,2.4713848,1.7263591,1.2307693,1.2012309,1.1946667,1.0404103,0.86974365,0.8730257,0.8172308,0.95835906,1.7033848,3.6069746,4.089436,3.8334363,3.2787695,2.7700515,2.5665643,2.7241027,3.245949,4.312616,5.504,5.8190775,4.95918,4.525949,4.3290257,4.1156926,3.564308,2.930872,2.3794873,2.2121027,2.1103592,1.142154,1.270154,1.3161026,1.1651284,0.88943595,0.7515898,0.81394875,0.8467693,1.0075898,1.2898463,1.5360001,1.0535386,0.92225647,1.0010257,1.0732309,0.86646163,0.86974365,0.97805136,1.0896411,1.0962052,0.9156924,0.5546667,0.6859488,0.85005134,0.9616411,1.2931283,1.4276924,1.3915899,1.4473847,2.2121027,4.644103,3.9056413,3.2032824,3.8038976,4.522667,1.7165129,1.591795,1.5655385,1.7165129,1.9495386,1.9561027,0.86646163,0.3117949,0.128,0.1148718,0.052512825,0.02297436,0.068923086,0.0951795,0.06564103,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.036102567,0.036102567,0.0,0.0,0.013128206,0.03938462,0.06564103,0.098461546,0.15425642,0.28882053,0.34133336,0.29538465,0.20676924,0.190359,0.27569234,0.37743592,0.39056414,0.32820517,0.2986667,0.33476925,0.27897438,0.22646156,0.2100513,0.190359,0.20020515,0.23958977,0.3446154,0.4594872,0.42994875,0.46933338,0.3511795,0.24943592,0.27241027,0.4594872,0.318359,0.29538465,0.29210258,0.256,0.21333335,0.27897438,0.24943592,0.21661541,0.21333335,0.21333335,0.2297436,0.3511795,0.48574364,0.61374366,0.8041026,0.827077,0.6859488,0.56123084,0.5284103,0.5415385,0.79097444,1.1815386,1.463795,1.5721027,1.6311796,1.8904617,2.2449234,2.6715899,3.1573336,3.6726158,4.397949,4.778667,5.2611284,5.8945646,6.3442054,6.770872,7.076103,7.1876926,7.0859494,6.7807183,7.243488,7.3025646,7.2894363,7.3485136,7.456821,7.5618467,7.351795,6.9152827,6.5903597,6.9645133,7.0367184,6.75118,7.069539,7.9163084,8.182155,8.1066675,7.4797955,6.6428723,6.1538467,6.7872825,7.259898,7.1056414,6.665847,6.0685134,5.2348723,4.9099493,4.4274874,4.07959,3.8564105,3.4625645,3.3312824,3.5544617,3.9318976,4.201026,4.0434875,3.8301542,3.6168208,3.442872,3.4855387,4.0533338,4.2174363,3.817026,3.698872,4.125539,4.7622566,5.4186673,7.387898,8.641642,8.621949,8.228104,10.180923,9.842873,8.073847,5.868308,4.348718,6.482052,7.003898,6.6002054,6.741334,9.685334,8.339693,6.816821,4.9821544,3.387077,3.255795,3.1474874,3.9548721,4.4800005,4.8377438,6.4590774,7.460103,3.8137438,1.4473847,1.7099489,1.3653334,1.6705642,2.038154,1.9429746,1.5885129,1.910154,2.2186668,2.0578463,1.9068719,1.9035898,1.8445129,1.6968206,1.5753847,1.7788719,2.1103592,1.8806155,1.7788719,1.7001027,1.6114873,1.6049232,1.8937438,2.044718,2.041436,2.2580514,2.7437952,3.239385,3.1803079,3.2623591,3.1015387,2.8291285,3.0949745,2.937436,3.1048207,3.2229745,3.3280003,3.8531284,3.889231,3.6332312,3.308308,2.878359,2.034872,2.0020514,2.225231,2.4648206,2.7831798,3.5446157,4.164923,4.322462,4.493129,4.8672824,5.346462,6.0980515,6.436103,6.8233852,7.3091288,7.5191803,7.3485136,8.700719,10.633847,12.665437,14.772514,15.120412,15.268104,16.141129,17.618053,18.533745,18.553438,18.06113,18.090668,18.71754,19.072002,18.615797,19.695591,20.345438,20.276514,20.847591,21.057642,21.031385,21.18236,21.369438,20.906668,19.718565,19.544617,19.695591,19.971283,20.644104,19.862976,18.901335,18.435284,18.553438,18.773335,18.176,17.263592,16.79754,16.866463,16.873028,16.531694,16.964924,18.25477,19.442873,18.54031,16.646564,15.579899,15.117129,15.543797,17.67713,17.673847,16.692514,15.842463,15.31077,14.368821,13.804309,13.522053,13.144616,12.435693,11.306667,10.965334,9.800206,8.231385,6.698667,5.661539,7.243488,7.77518,7.6635904,7.1909747,6.514872,5.930667,5.648411,5.976616,6.744616,7.322257,7.1023593,7.968821,8.960001,9.642668,10.089026,11.293539,12.691693,13.51877,13.443283,12.557129,12.416001,12.645744,12.891898,12.964104,12.832822,12.868924,13.548308,13.860104,13.689437,13.801026,14.667488,14.933334,14.578873,14.017642,14.086565,13.909334,13.50236,13.128206,12.4685135,10.620719,10.30236,9.714872,8.953437,8.03118,6.8693337,5.796103,5.2315903,5.037949,5.028103,4.969026,4.7360005,4.1714873,3.639795,3.2853336,3.0358977,2.8980515,2.9472823,2.934154,2.9702566,3.1015387,3.2951798,2.8553848,2.6190772,2.5206156,2.4976413,2.4713848,2.6420515,2.6945643,2.7076926,2.7667694,2.9768207,3.255795,3.508513,4.0533338,4.775385,5.142975,5.5072823,6.2588725,6.6133337,6.688821,7.506052,7.752206,7.381334,7.522462,8.15918,8.149334,10.59118,11.88759,11.21477,10.020103,12.009027,14.168616,11.241027,6.3507695,2.3794873,1.9528207,2.1103592,2.3991797,2.6847181,2.7963078,2.5009232,2.0020514,1.7296412,1.6082052,1.5130258,1.2832822,1.0994873,1.1454359,1.1323078,1.1093334,1.463795,1.5130258,1.7723079,2.034872,2.176,2.1530259,2.1136413,1.9954873,1.7624617,1.467077,1.2373334,1.211077,0.95835906,0.7318975,0.6432821,0.65641034,0.44964105,0.45292312,0.5973334,0.79097444,0.8992821,1.2176411,1.1946667,1.2504616,1.2603078,0.56451285,0.3314872,0.28225642,0.31507695,0.31507695,0.16738462,0.059076928,0.029538464,0.04266667,0.06235898,0.06235898,0.049230773,0.08205129,0.24615386,0.6235898,1.2832822,2.3433847,3.1409233,4.4832826,6.5444107,8.864821,10.148104,11.529847,13.00677,15.104001,18.875078,20.50954,19.941746,18.57313,17.05354,15.258258,14.257232,12.596514,11.352616,10.988309,11.369026,12.675283,12.826258,12.416001,11.789129,11.030975,10.19077,9.961026,10.551796,11.096616,9.642668,8.349539,7.4141545,7.4141545,8.205129,8.92718,7.351795,6.774154,6.688821,6.055385,3.2951798,2.3926156,1.5622566,1.1520001,1.3718976,2.28759,2.5928206,2.7241027,2.9571285,3.3017437,3.508513,5.8518977,8.854975,11.949949,15.113848,18.875078,21.060925,25.258669,28.097643,28.576822,28.074669,23.634052,19.088411,16.935387,17.80513,20.476719,23.870361,25.846155,28.494772,31.937643,34.31713,32.974773,31.22872,29.581131,28.445541,28.153439,27.762875,28.242054,29.338259,30.706875,31.891695,33.29313,31.704618,29.105232,27.090054,26.870155,27.493746,28.36349,29.889643,31.520823,31.753849,29.971695,28.547285,27.32636,25.816618,23.194258,23.108925,23.32554,23.207386,22.360617,20.614565,18.58954,18.110361,18.41559,18.46154,16.938667,15.973744,15.419078,15.461744,15.668514,14.982565,14.276924,14.116103,14.299898,14.572309,14.634667,14.549335,15.415796,16.183796,16.384,16.128002,16.324924,16.610462,16.410257,15.616001,14.601848,15.9343605,16.79754,17.857643,19.72513,22.934977,24.960001,24.97313,25.27836,26.446772,27.313232,29.902771,34.182568,38.560825,42.354874,45.82072,44.370056,40.818874,37.372723,34.43857,30.654362,26.883284,25.455591,23.299284,20.073027,18.14318,16.288822,16.866463,17.611488,17.772308,18.12677,20.483284,21.156105,21.776411,21.920822,19.088411,17.19795,13.912617,10.988309,9.051898,7.5979495,6.439385,7.1023593,7.430565,6.7774363,5.9963083,7.584821,8.411898,11.011283,15.179488,17.975796,17.11918,14.792206,14.372104,15.904821,16.114874,17.371899,15.514257,12.140308,8.946873,7.752206,5.0674877,3.8367183,3.9286156,4.522667,4.1189747,2.6551797,1.7132308,1.2537436,1.0043077,0.44307697,0.4660513,0.62030774,0.8336411,1.4342566,3.1442053,4.194462,4.2174363,3.8071797,3.249231,2.5173335,2.1891284,2.3171284,2.9768207,3.6824617,3.4034874,2.609231,2.3827693,2.2613335,2.038154,1.7690258,1.086359,0.9353847,0.97805136,1.0305642,1.0666667,1.276718,1.3554872,1.404718,1.3357949,0.88615394,1.1520001,1.1651284,1.079795,1.0601027,1.2668719,0.81394875,0.83035904,1.0436924,1.1848207,0.97805136,1.3784616,1.2242053,1.204513,1.3915899,1.2209232,0.63343596,0.42338464,0.47261542,0.7581539,1.3423591,1.6738462,1.4441026,1.3095386,1.6672822,2.6551797,5.9995904,6.1046157,4.394667,2.3269746,1.3718976,1.2996924,1.8051283,2.1333334,1.8576412,0.86974365,0.35774362,0.101743594,0.026256412,0.052512825,0.07548718,0.026256412,0.068923086,0.07548718,0.026256412,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02297436,0.06564103,0.10502565,0.13128206,0.16738462,0.30194873,0.35446155,0.3249231,0.26256412,0.27569234,0.3708718,0.26912823,0.19692309,0.22646156,0.27569234,0.26256412,0.40697438,0.4594872,0.36102566,0.21333335,0.16410258,0.190359,0.256,0.3314872,0.380718,0.3314872,0.2297436,0.2100513,0.30194873,0.4135385,0.28882053,0.3249231,0.34133336,0.2855385,0.21333335,0.24943592,0.23958977,0.2231795,0.21333335,0.21333335,0.2855385,0.3511795,0.43651286,0.571077,0.7778462,0.8041026,0.65312827,0.5481026,0.5415385,0.5021539,0.5874872,0.74830776,0.9616411,1.2406155,1.6180514,1.9462565,2.2580514,2.4484105,2.7306669,3.6463592,4.20759,4.2830772,4.6080003,5.3792825,6.2720003,7.138462,6.9809237,6.449231,6.0717955,6.2555904,6.62318,6.9809237,7.194257,7.0892315,6.4557953,6.8332314,6.882462,6.7774363,6.6822567,6.744616,6.0356927,6.0980515,6.806975,7.5585647,7.27959,7.3386674,7.171283,6.8430777,6.665847,7.200821,7.2631803,6.7282057,6.0685134,5.5007186,4.9887185,4.391385,3.9680004,3.7120004,3.6102567,3.6463592,3.5741541,3.3280003,3.7218463,4.630975,4.95918,4.325744,4.1747694,3.9975388,3.820308,4.210872,4.394667,3.698872,3.3378465,3.7152824,4.4110775,4.896821,6.3934364,7.6635904,8.067283,7.568411,8.349539,8.982975,8.513641,7.1680007,6.363898,8.388924,10.807796,11.132719,9.209436,7.2336416,7.817847,4.9985647,3.4724104,4.342154,5.110154,3.7316926,4.457026,4.59159,4.1780515,5.9963083,6.547693,3.5052311,1.5425643,1.7920002,1.8773335,1.7066668,1.7920002,1.723077,1.5425643,1.7394873,2.300718,2.4582565,2.3926156,2.1956925,1.8904617,1.7952822,1.4572309,1.4966155,1.8313848,1.7099489,1.6836925,1.5589745,1.5360001,1.7362052,2.2121027,1.9331284,1.9528207,2.03159,2.1989746,2.7634873,2.6157951,2.6322052,2.537026,2.4713848,3.0227695,2.8258464,2.9604106,3.0654361,3.18359,3.767795,3.892513,3.629949,3.255795,2.806154,2.0611284,2.034872,1.910154,2.1300514,2.7044106,3.2032824,3.5577438,4.1517954,4.9329233,5.61559,5.674667,6.8955903,7.4404106,7.4043083,7.056411,6.8365135,7.1056414,9.058462,11.37559,13.443283,15.333745,14.821745,14.959591,16.466053,18.678156,19.5479,18.960411,19.042463,18.865232,18.336823,18.202257,18.71754,20.299488,22.022566,23.240208,23.604515,23.092514,22.65272,22.89231,23.348515,22.505028,21.592617,21.609028,21.592617,21.218464,20.8279,20.522669,19.91549,19.170464,18.507488,18.189129,19.055592,19.226257,19.14749,18.81272,17.77559,16.75159,16.777847,18.070976,19.846565,20.309336,18.806156,17.332514,16.643284,17.129026,18.81272,18.691284,17.572104,16.784412,16.699078,16.722052,15.074463,14.28677,13.6467705,12.832822,11.9171295,11.625027,10.187488,8.1066675,6.186667,5.540103,7.1515903,7.433847,6.872616,6.0750775,5.7829747,6.2227697,5.9569235,6.12759,6.9054365,7.4929237,7.2861543,8.461129,9.760821,10.5780525,10.955488,12.786873,14.106257,14.385232,13.804309,13.22995,13.840411,13.489232,13.354668,13.505642,12.895181,12.685129,12.898462,13.15118,13.410462,14.007796,14.385232,14.470565,13.873232,13.157744,13.853539,13.157744,13.15118,13.138052,12.57354,11.047385,10.243283,9.399796,8.4053335,7.2369237,5.9667697,5.2447186,4.709744,4.568616,4.7622566,4.9427695,4.663795,4.069744,3.4133337,2.92759,2.8521028,2.3860514,2.5140514,2.6420515,2.8849232,3.170462,3.245949,2.9833848,2.7175386,2.5993848,2.6387694,2.7044106,2.5829747,2.7733335,2.8389745,2.7011285,2.6453335,3.006359,3.2328207,3.6758976,4.378257,5.106872,5.5991797,6.4557953,7.0367184,7.240206,7.4830775,7.4929237,7.532308,7.634052,7.785026,7.9294367,9.472001,10.272821,10.906258,13.259488,20.54236,19.702156,13.403898,6.564103,2.2153847,1.4769232,1.4309745,2.2219489,3.1507695,3.5610259,2.8553848,2.2777438,2.0086155,1.9265642,1.8871796,1.7329233,1.5097437,1.4506668,1.4408206,1.5491283,2.038154,2.5074873,2.6387694,2.674872,2.7864618,3.05559,2.9210258,2.228513,1.6738462,1.4769232,1.3817437,1.3883078,1.3522053,1.2635899,1.1585642,1.1323078,0.78769237,0.7778462,0.88287187,0.9517949,0.92553854,1.086359,1.083077,1.0010257,0.81394875,0.380718,0.29538465,0.256,0.2297436,0.20348719,0.14441027,0.101743594,0.098461546,0.10502565,0.101743594,0.072205134,0.09189744,0.0951795,0.2100513,0.6268718,1.5983591,3.2164104,4.1813335,5.5926156,7.896616,10.880001,13.000206,14.667488,15.977027,17.152,18.520617,18.428719,17.506462,16.108309,14.959591,15.136822,14.496821,13.850258,12.76718,11.523283,11.113027,11.703795,11.526565,11.116308,10.880001,11.07036,11.35918,12.416001,14.040616,14.65436,11.316514,7.522462,6.157129,5.8420515,5.533539,4.5456414,3.6824617,3.4592824,3.5938463,3.7382567,3.4789746,2.986667,2.1202054,1.3489232,1.0469744,1.4966155,1.2340513,1.7066668,2.038154,2.103795,2.546872,5.10359,8.123077,10.804514,12.629334,13.371078,16.689232,22.311386,28.18954,31.888412,30.628105,27.13272,22.800411,18.898052,16.656412,17.28,20.30277,24.87795,29.508924,32.774567,33.329235,30.257233,28.70154,28.20267,28.527592,29.689438,28.90831,28.192823,28.553848,30.053745,31.806362,31.599592,32.12472,31.520823,29.558157,27.638157,27.178669,27.631592,28.422565,29.088823,29.249643,28.737642,28.291285,27.625029,26.279387,23.59467,23.14831,23.745644,24.185438,23.83754,22.629745,20.903387,19.606976,18.95713,18.661745,17.939693,16.718771,16.02954,16.042667,16.288822,15.655386,14.624822,14.276924,14.326155,14.290052,13.4629755,13.689437,14.024206,14.828309,15.940925,16.689232,15.908104,15.474873,14.834873,13.866668,12.895181,12.973949,13.4170265,14.073437,15.396104,18.441847,20.164925,21.845335,22.340925,22.324514,24.274054,27.408413,32.64657,38.101337,42.817646,46.7758,45.26277,41.4359,37.776413,34.530464,29.689438,23.955694,23.289438,22.439386,19.994259,18.386053,16.354464,15.31077,15.300924,16.456207,18.95713,21.106873,21.362873,21.4679,21.589334,20.309336,19.111385,15.465027,12.370052,10.683078,9.124104,7.768616,7.899898,7.9983597,7.328821,5.910975,7.000616,8.149334,11.349334,15.947489,18.645334,16.823795,13.925745,12.327386,12.33395,12.1698475,15.684924,16.456207,15.616001,14.034052,12.340514,9.508103,7.6931286,7.256616,7.5552826,6.928411,2.9538465,1.404718,1.020718,0.98133343,0.9189744,0.80738467,1.8182565,2.0841026,1.6869745,2.6551797,4.125539,4.8836927,4.709744,3.7809234,2.6880002,2.1136413,1.8904617,2.5271797,3.5938463,3.6824617,2.0217438,1.5130258,1.3981539,1.3226668,1.3193847,0.9189744,0.761436,0.79097444,1.0305642,1.591795,1.6443079,2.0644104,2.0217438,1.4244103,0.9353847,1.211077,1.9298463,2.228513,1.9626669,1.6804104,1.142154,1.2242053,1.1520001,0.7778462,0.5481026,0.6695385,0.5316923,0.5316923,0.78769237,1.1355898,0.81394875,0.47917953,0.318359,0.42338464,0.79425645,1.0633847,1.2603078,1.585231,1.9528207,1.9954873,3.006359,3.6693337,3.2918978,2.1103592,1.276718,2.0906668,2.6190772,2.4615386,1.6640002,0.7220513,1.8215386,1.0896411,0.25928208,0.09189744,0.380718,0.08861539,0.318359,0.3314872,0.036102567,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.0,0.013128206,0.068923086,0.09189744,0.07876924,0.0951795,0.18051283,0.22646156,0.22646156,0.19364104,0.17723078,0.23630771,0.26256412,0.3446154,0.50543594,0.702359,0.86646163,0.7450257,0.61374366,0.5284103,0.3249231,0.24615386,0.23302566,0.26584616,0.32164106,0.380718,0.3511795,0.28225642,0.23958977,0.24287182,0.26584616,0.2986667,0.26912823,0.23302566,0.22646156,0.24943592,0.256,0.26912823,0.29538465,0.3249231,0.33476925,0.3511795,0.35446155,0.43651286,0.60389745,0.8041026,0.76800007,0.78769237,0.7187693,0.571077,0.5152821,0.56123084,0.6301539,0.7811283,1.014154,1.276718,1.4309745,1.5786668,1.7985642,2.225231,3.0720003,3.5282054,3.7021542,3.8990772,4.5128207,6.038975,6.564103,6.7314878,6.701949,6.636308,6.6822567,6.8430777,7.0104623,7.1647186,7.2205133,7.017026,6.633026,6.892308,6.9842057,6.7282057,6.5739493,6.5017443,6.882462,7.584821,8.260923,8.339693,7.785026,7.1483083,6.678975,6.47877,6.518154,6.314667,6.1768208,5.9470773,5.730462,5.8912826,5.5007186,4.673641,3.9417439,3.4921029,3.1474874,3.4921029,3.498667,3.8400004,4.535795,4.923077,4.601436,4.667077,4.397949,3.82359,3.7349746,3.761231,3.2689233,3.0260515,3.2098465,3.4100516,3.9253337,4.903385,6.2096415,7.5618467,8.4972315,7.8112826,7.269744,7.322257,7.3747697,5.789539,6.301539,8.073847,9.475283,9.90195,9.770667,7.1548724,6.2818465,7.0925136,8.001641,5.8814363,5.35959,5.421949,5.2676926,5.277539,6.997334,9.032206,4.7589746,1.522872,1.4703591,1.5360001,1.7755898,1.6607181,1.5130258,1.5064616,1.6902566,1.9003079,1.9364104,1.9889232,2.0118976,1.6968206,1.6672822,1.5031796,1.4966155,1.6738462,1.7952822,1.9068719,1.7952822,1.7460514,1.8445129,1.9692309,2.0184617,2.044718,2.038154,2.162872,2.7241027,2.5009232,2.7175386,2.7831798,2.6223593,2.6912823,2.8192823,3.05559,3.2229745,3.442872,4.1485133,4.161641,3.4855387,2.8389745,2.4746668,2.169436,2.3893335,2.537026,2.7044106,2.9505644,3.314872,3.764513,4.3749747,5.113436,5.8190775,6.1997952,6.485334,6.2720003,6.226052,6.485334,6.675693,8.224821,9.613129,11.349334,13.262771,14.480412,14.562463,15.156514,15.947489,16.889437,18.215385,19.456001,20.565334,21.024822,20.87713,20.742565,20.814772,21.425232,22.800411,24.375797,24.789335,23.739079,22.87918,22.78072,23.220514,23.190975,22.754463,23.40431,23.46995,22.92513,23.40431,22.357334,21.776411,21.353027,20.752413,19.603693,21.858463,22.610052,22.281847,21.097027,19.081848,17.765745,17.184822,17.88718,19.561028,21.041233,20.683489,19.925335,19.012924,18.579693,19.669334,19.672617,19.272207,18.694565,18.07754,17.46708,16.308514,15.284514,14.135796,12.852514,11.674257,11.447796,9.90195,7.8670774,6.3967185,6.7840004,7.5552826,7.2631803,6.449231,5.76,5.9536414,6.921847,6.8463597,6.8266673,7.2270775,7.6767187,7.5552826,8.516924,9.682052,10.66995,11.61518,13.397334,14.168616,13.952001,13.298873,13.289026,14.605129,14.421334,13.883078,13.479385,13.065847,12.681848,12.806565,13.095386,13.35795,13.5548725,14.139078,13.974976,13.269335,12.5374365,12.596514,12.156719,12.209231,12.393026,12.35036,11.74318,10.079181,8.946873,7.7292314,6.445949,5.7829747,5.208616,4.781949,4.4307694,4.2272825,4.3716927,3.95159,3.4592824,3.0785644,2.878359,2.806154,2.3958976,2.3663592,2.5862565,2.806154,2.9636924,3.190154,3.2032824,3.0096412,2.7733335,2.5928206,2.4976413,2.6157951,2.7241027,2.665026,2.537026,2.665026,2.8291285,3.0654361,3.5249233,4.2272825,5.0609236,5.7764106,6.5083084,7.1187696,7.532308,7.722667,7.6668725,7.896616,7.958975,8.109949,9.31118,9.5606165,9.67877,12.084514,17.93313,27.122873,23.794874,15.094155,7.328821,3.2098465,1.8445129,1.0633847,1.1651284,1.6311796,2.0250258,1.9659488,1.9462565,1.9003079,1.9068719,1.8970258,1.6443079,1.5885129,1.6738462,1.7296412,1.8116925,2.1825643,2.5271797,2.5928206,2.6945643,2.9013336,3.0227695,2.8717952,2.2678976,1.8313848,1.7558975,1.8116925,1.5392822,1.4900514,1.4441026,1.3193847,1.1585642,1.1323078,1.1191796,1.0732309,0.99774367,0.9682052,0.9419488,0.8598975,0.79097444,0.7318975,0.5907693,0.50543594,0.40697438,0.30194873,0.20676924,0.15425642,0.108307704,0.07876924,0.06235898,0.055794876,0.049230773,0.059076928,0.06235898,0.24287182,0.79425645,1.9265642,3.6824617,4.9821544,6.705231,9.225847,12.389745,14.339283,15.780104,16.968206,17.72636,17.424412,16.820515,15.799796,14.65436,14.178463,15.691488,16.036104,15.701335,14.41477,12.448821,10.617436,10.226872,10.663385,10.8996935,10.880001,11.526565,12.987078,15.448617,17.545847,17.444103,12.859077,8.109949,6.1505647,5.3202057,4.5817437,3.5314875,2.7733335,2.15959,2.0512822,2.359795,2.5271797,2.546872,2.3171284,1.6869745,0.92553854,0.72861546,0.72861546,1.0272821,1.0502565,0.88943595,1.2865642,3.058872,6.058667,8.769642,10.499283,11.388719,13.751796,18.950565,25.212719,29.814156,29.08554,27.497028,24.546463,20.837746,17.818258,17.752617,21.691078,26.12185,30.605131,33.956104,34.244926,31.08431,29.256207,28.074669,27.30667,27.155695,27.175386,27.808823,28.65231,29.715694,31.419079,31.136824,32.36759,33.08308,31.967182,28.445541,27.874464,28.022156,28.176413,28.084515,27.940105,27.559387,26.729027,26.01354,25.360413,24.100105,24.536617,25.140514,25.212719,24.697437,24.201847,22.934977,21.842052,20.598156,19.324718,18.609232,18.06113,16.925539,16.38072,16.521847,16.38072,15.314053,14.726565,14.280207,13.633642,12.445539,12.84595,13.190565,14.162052,15.868719,17.828104,17.851078,17.42113,15.96718,13.896206,12.593232,11.382154,11.674257,12.452104,13.673027,16.265848,17.942976,19.551182,20.171488,19.908924,19.899078,23.023592,28.947695,35.222977,40.146053,42.77498,40.933746,36.788517,32.863182,29.77477,26.217028,23.089233,23.151592,22.675694,20.775387,19.416616,16.741745,15.402668,15.570052,17.283283,20.447182,20.276514,19.856411,19.797335,20.233849,20.854155,20.355284,18.01518,16.216616,14.841437,11.254155,9.754257,8.513641,8.493949,8.736821,6.3474874,6.747898,8.067283,11.437949,15.586463,16.856617,14.299898,11.332924,9.636104,9.278359,8.723693,11.848206,13.974976,15.645539,16.748308,16.518566,15.665232,13.761642,12.2847185,11.208206,8.992821,4.397949,2.2613335,1.3981539,1.1618463,1.4506668,2.0709746,3.8629746,4.525949,3.754667,3.245949,4.893539,6.3606157,6.432821,5.1298466,3.7185643,2.865231,2.1431797,2.1136413,2.7241027,3.3312824,2.0906668,1.339077,0.955077,0.81394875,0.79425645,0.7581539,0.7089231,0.75487185,0.9714873,1.404718,1.6213335,1.910154,1.7952822,1.3029745,0.955077,1.142154,1.7132308,2.4418464,2.989949,2.937436,2.0906668,1.5031796,1.0075898,0.6104616,0.48902568,0.49230772,0.4201026,0.4266667,0.574359,0.83035904,0.90256417,0.64000005,0.380718,0.35774362,0.7187693,0.955077,1.332513,1.6607181,1.7460514,1.4178462,1.9429746,2.2678976,2.041436,1.4605129,1.2800001,2.169436,1.9692309,1.4408206,1.3850257,2.6453335,1.5261539,0.6268718,0.13456412,0.049230773,0.18379489,0.04266667,0.15097436,0.15753847,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0,0.013128206,0.04266667,0.055794876,0.068923086,0.14112821,0.18379489,0.190359,0.23630771,0.29538465,0.23630771,0.41682056,0.8533334,1.1881026,1.2832822,1.2307693,1.2898463,0.9353847,0.69907695,0.6629744,0.45292312,0.3446154,0.33805132,0.3446154,0.33476925,0.33476925,0.318359,0.27569234,0.24615386,0.23630771,0.2297436,0.27897438,0.23302566,0.20348719,0.2297436,0.2855385,0.2855385,0.28882053,0.3117949,0.34789747,0.36758977,0.31507695,0.28225642,0.29210258,0.39056414,0.65312827,0.6629744,0.8369231,0.8467693,0.65312827,0.51856416,0.69579494,0.69907695,0.6859488,0.764718,0.99774367,0.9189744,1.0075898,1.332513,1.8674873,2.5009232,2.8389745,3.31159,3.7743592,4.457026,5.979898,6.7872825,6.8955903,6.7905645,6.688821,6.5345645,6.7905645,6.672411,6.678975,6.7872825,6.432821,5.8814363,6.4000006,6.9087186,7.062975,7.243488,7.88677,8.408616,8.700719,8.740103,8.595693,7.824411,7.128616,6.5870776,6.2490263,6.163693,5.8092313,5.937231,6.160411,6.232616,6.0717955,5.0149746,4.2863593,3.7842054,3.4658465,3.3312824,3.43959,3.5872824,4.0041027,4.5128207,4.529231,4.3716927,4.457026,4.325744,3.8662567,3.3247182,3.1277952,2.9702566,3.0490258,3.255795,3.1770258,3.570872,4.519385,5.549949,6.5050263,7.5552826,7.181129,7.250052,7.778462,7.8080006,5.425231,6.432821,8.854975,10.095591,9.229129,7.0104623,6.12759,9.645949,10.545232,8.024616,7.499488,7.0498466,5.8223596,5.366154,6.6034875,9.83959,9.69518,6.7249236,3.6004105,1.8543591,1.8806155,1.7591796,1.6147693,1.4933335,1.4998976,1.8149745,1.8806155,1.8248206,1.8904617,1.9856411,1.6738462,1.7001027,1.6311796,1.5885129,1.6607181,1.9167181,1.719795,1.6311796,1.6213335,1.7066668,1.9626669,2.1858463,2.0709746,2.0184617,2.156308,2.359795,2.0053334,2.356513,2.7076926,2.7536411,2.5731285,2.7733335,3.0785644,3.4034874,3.7382567,4.141949,3.5577438,2.8849232,2.5107694,2.4910772,2.5731285,2.7437952,2.9013336,3.0490258,3.2032824,3.3772311,3.9581542,4.4307694,5.044513,5.7731285,6.3245134,6.0356927,5.8256416,5.85518,6.314667,7.433847,9.110975,10.896411,12.576821,13.8075905,14.102976,14.9628725,15.333745,16.049232,17.38831,19.10154,20.43077,21.169233,21.32677,21.195488,21.333336,22.393438,23.269745,24.214975,25.028925,25.074873,24.264208,23.558565,23.151592,23.253336,24.083694,25.422771,25.376822,24.20513,22.99077,23.637335,23.302567,22.951385,22.564104,22.09149,21.431797,23.089233,24.346258,24.864822,24.037745,21.011694,19.121233,18.23836,18.592821,19.91549,21.444925,21.714052,21.428514,20.936207,20.614565,20.844309,20.499695,20.178053,19.64636,18.760206,17.47036,16.390566,15.02195,13.568001,12.150155,10.788103,10.6469755,9.124104,7.3714876,6.4295387,7.2237954,7.529026,7.177847,6.521436,6.0061545,6.160411,7.0104623,7.3058467,7.4732313,7.6701546,7.785026,7.8769236,8.960001,10.266257,11.52,12.950975,13.63036,13.860104,13.636924,13.344822,13.764924,15.356719,14.966155,13.935591,13.131488,12.934566,12.754052,12.865642,13.069129,13.262771,13.433437,13.929027,13.7386675,12.908309,11.956513,11.881026,11.897437,11.808822,11.792411,11.739899,11.2672825,9.77395,8.484103,7.3550773,6.3934364,5.6451287,4.8377438,4.2207184,3.7415388,3.4264617,3.383795,3.0949745,2.9604106,2.9472823,2.9997952,3.058872,2.487795,2.2514873,2.3729234,2.5074873,2.605949,2.9144619,3.186872,3.1048207,2.8127182,2.4516926,2.172718,2.4352822,2.5107694,2.4582565,2.4681027,2.8521028,2.8389745,3.170462,3.623385,4.1878977,5.0904617,6.294975,6.9120007,7.4797955,8.070564,8.2904625,8.211693,8.369231,8.349539,8.625232,10.548513,9.524513,10.121847,13.794462,20.118977,26.794668,20.483284,12.389745,6.5247183,3.8465643,2.2711797,1.0765129,0.53825647,0.47261542,0.69251287,1.0010257,1.2504616,1.3292309,1.467077,1.5885129,1.332513,1.394872,1.5688206,1.7985642,2.0939488,2.5173335,2.4943593,2.6223593,2.7437952,2.7569232,2.6223593,2.5337439,2.1792822,1.910154,1.8313848,1.8116925,1.5688206,1.5688206,1.5556924,1.4342566,1.2865642,1.4703591,1.3817437,1.211077,1.079795,1.0535386,0.90584624,0.77128214,0.84348726,1.079795,1.1848207,0.81394875,0.5874872,0.43323082,0.32820517,0.30194873,0.16410258,0.07548718,0.036102567,0.036102567,0.06564103,0.12143591,0.23958977,0.6268718,1.3489232,2.3269746,3.9154875,5.287385,7.003898,9.278359,11.999181,13.978257,15.688207,16.843489,17.024002,15.668514,15.067899,14.70359,14.834873,15.970463,18.871796,22.239182,20.900105,17.942976,14.969437,12.107488,10.981745,11.739899,12.563693,13.000206,13.948719,15.730873,18.888206,21.284103,20.801643,15.343591,9.921641,7.0892315,5.3398976,4.0500517,3.4822567,3.0490258,2.4943593,2.297436,2.3827693,2.1431797,2.0775387,2.1891284,1.847795,1.0896411,0.5940513,0.5218462,0.49230772,0.3446154,0.21989745,0.5481026,1.2635899,4.194462,7.0104623,8.592411,9.045334,11.0145645,14.565744,19.347694,23.93272,25.819899,26.574772,26.187489,23.758772,20.309336,18.776617,21.635284,25.659079,30.227695,33.90359,34.44513,32.482464,30.782362,29.32513,28.150156,27.349335,26.41067,26.935797,27.680822,28.75077,31.61272,31.507694,32.981335,34.49436,34.38277,30.854567,29.571285,29.101952,28.865643,28.498053,27.82195,27.030977,25.898668,25.419489,25.616413,25.570463,26.308926,26.499285,26.072617,25.16677,24.106668,22.849644,22.606771,22.144001,21.270975,20.844309,20.693335,19.236105,17.956104,17.391592,17.138874,16.52513,15.514257,14.519796,13.545027,12.199386,12.747488,13.289026,14.27036,15.82277,17.769028,18.947283,19.780924,18.927591,16.548103,14.303181,12.517745,12.471796,12.931283,13.853539,16.38072,18.12677,18.422155,18.208822,17.654156,16.137848,19.462566,25.504822,31.363285,35.091694,35.68903,33.119183,29.229952,25.90195,23.899899,22.89231,23.988514,24.451284,23.601233,21.687796,19.882668,17.378464,16.338053,16.649847,18.005335,19.88595,16.873028,16.25272,16.889437,18.290873,20.62113,21.88472,20.847591,19.035898,16.561232,12.084514,10.65354,8.825437,8.621949,9.212719,6.921847,6.8955903,7.8539495,10.643693,13.83713,13.74195,10.505847,7.972103,6.9382567,7.069539,6.9087186,9.619693,10.811078,12.642463,15.182771,16.403694,19.006361,20.581745,19.712002,16.469334,12.3995905,8.247795,5.3924108,3.5216413,2.5304618,2.487795,3.4756925,5.6451287,6.672411,5.9963083,4.8147697,5.9503593,7.522462,7.77518,6.744616,6.2785645,4.6605134,2.8750772,1.8674873,2.0020514,3.045744,2.3269746,1.4506668,1.2176411,1.394872,0.7089231,1.0765129,1.0929232,1.0469744,1.0929232,1.2438976,1.404718,1.5064616,1.4145643,1.1913847,1.083077,1.2832822,1.6147693,2.4976413,3.7087183,4.378257,2.92759,1.5622566,0.7581539,0.53825647,0.4955898,0.5677949,0.7450257,0.7187693,0.51856416,0.512,0.86317956,0.86974365,0.7417436,0.67610264,0.8467693,1.0666667,1.2832822,1.3259488,1.2406155,1.2603078,1.6836925,1.5885129,1.2832822,1.0633847,1.211077,1.4539489,0.9189744,0.45292312,0.75487185,2.3893335,0.6695385,0.101743594,0.009846155,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.01969231,0.04266667,0.026256412,0.026256412,0.072205134,0.13784617,0.13456412,0.20676924,0.256,0.38728207,0.636718,0.98461545,0.9124103,1.3915899,1.8904617,2.3926156,3.4034874,2.917744,2.3663592,1.6147693,0.88287187,0.761436,0.42994875,0.33476925,0.30194873,0.27241027,0.26912823,0.30851284,0.27897438,0.256,0.26256412,0.23958977,0.29210258,0.24287182,0.2297436,0.27241027,0.27569234,0.2855385,0.28882053,0.29210258,0.2986667,0.32820517,0.2986667,0.256,0.2100513,0.24615386,0.5316923,0.62030774,0.8008206,0.8172308,0.67282057,0.63343596,0.7975385,0.7844103,0.6662565,0.57764107,0.7417436,0.7089231,0.8041026,1.1323078,1.6804104,2.3236926,2.540308,3.058872,3.817026,4.841026,6.23918,7.3616414,7.6996927,7.5487185,7.138462,6.633026,6.6494365,6.1505647,5.943795,6.055385,5.7501545,5.6385646,6.0258465,6.564103,7.2237954,8.3134365,9.43918,9.685334,9.429334,9.009232,8.743385,7.88677,7.204103,6.688821,6.2916927,5.933949,5.61559,5.8256416,6.2194877,6.380308,5.805949,4.2601027,3.7973337,3.7349746,3.7152824,3.7120004,3.255795,3.2820516,3.5971284,3.8432825,3.4658465,3.6824617,3.9286156,4.010667,3.7776413,3.121231,2.7963078,2.7602053,2.865231,3.0096412,3.1638978,3.639795,4.332308,5.2053337,6.1407185,6.9382567,6.9743595,7.9130263,8.474257,7.975385,6.3343596,5.9602056,8.372514,9.659078,8.369231,5.5138464,7.0531287,10.748719,10.771693,7.240206,6.2490263,6.183385,5.169231,4.6539493,5.366154,7.312411,9.517949,8.73354,5.398975,1.7985642,2.0578463,1.5819489,1.5031796,1.5097437,1.5327181,1.7558975,1.8215386,1.8149745,1.8576412,1.9200002,1.8149745,1.8642052,1.7723079,1.7001027,1.7165129,1.8018463,1.4178462,1.4211283,1.5327181,1.723077,2.1891284,2.1136413,1.9692309,1.9429746,2.034872,2.048,1.8313848,2.1825643,2.5829747,2.7569232,2.6584618,2.7798977,3.0884104,3.4166157,3.6693337,3.8006158,2.989949,2.5928206,2.4910772,2.5993848,2.8717952,2.934154,3.0654361,3.2295387,3.3247182,3.1540515,3.515077,3.9876926,4.647385,5.3431797,5.687795,5.5236926,5.7796926,6.262154,7.056411,8.546462,9.938052,11.697231,13.144616,14.007796,14.418053,15.560206,16.147694,17.529438,19.813745,21.842052,22.068514,22.186668,22.150566,22.199797,22.846361,24.448002,25.383387,25.80349,25.649233,24.661335,24.58913,24.602259,24.362669,24.132925,24.763079,26.77826,26.26954,24.864822,23.840822,24.100105,23.962257,23.77518,23.338669,22.856207,22.94154,23.433847,24.838566,26.17436,26.006977,22.452515,19.98113,19.081848,19.56759,20.913233,22.249027,22.3639,22.20308,22.226053,22.33108,21.868309,21.234873,20.745848,19.810463,18.330257,16.682669,15.740719,14.355694,12.786873,11.237744,9.865847,9.7214365,8.316719,6.9087186,6.3868723,7.273026,7.4207187,7.128616,6.7085133,6.4557953,6.6625648,7.0925136,7.680001,8.054154,8.083693,7.899898,8.277334,9.432616,10.761847,12.038565,13.410462,13.810873,13.843694,13.538463,13.331694,14.043899,15.445334,14.907078,13.728822,12.839386,12.76718,12.760616,12.944411,13.13477,13.269335,13.39077,13.495796,13.200411,12.416001,11.608616,11.795693,11.864616,11.336206,10.755282,10.322052,9.888822,9.16677,8.260923,7.312411,6.2884107,5.0051284,4.1124105,3.3641028,2.8717952,2.6354873,2.537026,2.3958976,2.6453335,2.9965131,3.2689233,3.3805132,2.556718,2.284308,2.1858463,2.1858463,2.281026,2.540308,2.8816411,2.9144619,2.674872,2.28759,1.9462565,2.1825643,2.300718,2.3466668,2.481231,2.9702566,2.930872,3.4034874,3.7809234,4.1058464,5.093744,6.7905645,7.387898,7.9917955,8.756514,8.900924,8.914052,8.953437,8.759795,8.897642,10.729027,9.097847,11.149129,15.366566,19.488823,20.489847,11.539693,6.3573337,4.1189747,3.4198978,2.284308,1.4473847,0.90912825,0.702359,0.75487185,0.86317956,0.80738467,0.83035904,1.014154,1.2242053,1.1191796,1.1355898,1.2865642,1.6836925,2.2613335,2.7569232,2.4385643,2.6715899,2.7109745,2.3893335,2.1070771,2.1234872,1.9462565,1.8051283,1.7066668,1.4178462,1.4998976,1.6246156,1.6246156,1.5163078,1.5064616,1.6311796,1.4473847,1.2340513,1.1126155,1.0568206,0.90912825,0.8205129,1.0502565,1.4867693,1.657436,1.0043077,0.6859488,0.56451285,0.5415385,0.5513847,0.256,0.13456412,0.08861539,0.07876924,0.128,0.25928208,0.5546667,1.1749744,2.0020514,2.6518977,3.8498464,5.093744,6.557539,8.388924,10.70277,13.4400015,15.691488,16.54154,15.80636,14.053744,13.88636,14.811898,16.538258,19.045746,22.567387,28.688412,26.692924,22.160412,18.067694,14.78236,13.761642,14.54277,15.8654375,17.188105,18.68472,19.90236,22.488617,24.795898,24.559591,18.904617,12.73436,8.759795,5.796103,3.6824617,3.2984617,3.249231,3.1967182,3.1376412,2.9636924,2.4582565,1.9593848,1.9429746,1.8445129,1.4933335,1.1126155,0.6268718,0.256,0.09189744,0.15753847,0.40369233,0.7122052,3.0752823,5.3398976,6.2851286,5.6254363,8.306872,10.381129,13.8765135,18.83241,23.286156,25.032207,26.87672,26.17108,22.905437,19.695591,19.373951,22.86277,27.542976,31.343592,32.74831,33.076515,32.41354,31.602875,31.16308,31.300926,28.425848,26.752003,26.28267,27.572515,31.737438,31.80308,33.46708,35.43631,36.28636,34.464825,32.31508,31.087593,30.46072,29.906054,28.681849,27.67754,26.758566,26.59118,27.11631,27.569233,27.871181,27.40513,26.5879,25.330873,23.059694,21.474463,21.93395,23.194258,24.329847,24.763079,24.30359,22.846361,21.205336,19.790771,18.62236,18.251488,16.820515,15.573335,14.644514,13.062565,13.197129,13.725539,14.5263605,15.491283,16.528412,18.491077,21.30708,22.485334,21.162668,18.087385,16.278976,15.691488,15.258258,15.376411,17.880617,19.577436,18.159592,16.452925,15.461744,14.372104,17.94954,23.424002,27.782566,29.508924,28.57354,25.46872,22.432823,20.427488,20.036924,21.454771,25.363695,25.951181,24.536617,22.117744,19.38708,17.522873,16.722052,16.997746,17.539284,16.692514,12.182976,11.85477,13.348104,15.744001,19.56759,22.85949,22.255592,19.11795,14.916924,11.224616,9.947898,9.048616,8.976411,9.009232,7.253334,6.9743595,7.53559,9.580308,11.638155,10.128411,6.889026,5.3366156,5.031385,5.6418467,6.9152827,9.69518,8.608821,8.641642,10.774975,11.972924,17.821539,24.329847,25.728003,21.661541,17.174976,15.015386,10.758565,7.1515903,5.1626673,3.9712822,4.33559,6.0258465,7.141744,7.0432825,6.3507695,6.3277955,7.197539,7.4797955,7.2960005,8.342975,6.0717955,3.4724104,1.8838975,1.7952822,2.861949,2.6387694,2.034872,2.2449234,2.7766156,1.4769232,1.9856411,1.7952822,1.4473847,1.2373334,1.2373334,1.1093334,1.204513,1.2176411,1.1782565,1.4276924,1.8248206,2.284308,3.170462,4.414359,5.4941545,3.6463592,1.972513,0.92553854,0.5481026,0.45292312,0.6826667,1.0929232,1.024,0.52512825,0.3708718,0.71548724,0.98133343,1.1520001,1.1684103,0.9485129,1.0338463,0.90912825,0.6859488,0.6498462,1.2406155,1.3981539,1.1552821,0.9682052,0.9682052,0.9714873,0.42994875,0.16082053,0.059076928,0.036102567,0.036102567,0.036102567,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.03938462,0.0951795,0.04594872,0.032820515,0.11158975,0.20676924,0.101743594,0.23630771,0.39384618,0.62030774,1.0535386,1.910154,1.401436,1.6213335,2.2777438,3.5314875,5.9995904,5.07077,4.6112823,3.4264617,1.8543591,1.7591796,0.65641034,0.23958977,0.14769232,0.15425642,0.20348719,0.318359,0.318359,0.30194873,0.2986667,0.26912823,0.3117949,0.26584616,0.26912823,0.3117949,0.24287182,0.256,0.26912823,0.25928208,0.24943592,0.2986667,0.34133336,0.31507695,0.26256412,0.26584616,0.4660513,0.5940513,0.67610264,0.6695385,0.6498462,0.80738467,0.80738467,0.82379496,0.7122052,0.5513847,0.6498462,0.8533334,0.94523084,1.1716924,1.6836925,2.5435898,2.7076926,2.9997952,3.889231,5.3202057,6.7117953,7.8769236,8.592411,8.585847,7.958975,7.197539,6.688821,5.9634876,5.5729237,5.5696416,5.5105643,5.8912826,5.986462,6.3310776,7.318975,9.209436,10.180923,9.984001,9.380103,8.835282,8.5202055,7.821129,7.197539,6.7577443,6.36718,5.658257,5.586052,5.7468724,5.9634876,5.9503593,5.2709746,3.8334363,3.564308,3.764513,3.9286156,3.7284105,2.8849232,2.665026,2.7208207,2.7306669,2.3958976,2.9538465,3.4231799,3.623385,3.4855387,3.0654361,2.6486156,2.5337439,2.3991797,2.359795,2.9801028,3.626667,3.9680004,4.9952826,6.567385,7.4043083,7.5520005,8.592411,8.713847,7.8670774,7.7456417,4.4701543,6.058667,7.899898,7.90318,6.4689236,10.151385,9.819899,8.234667,6.3474874,3.2951798,3.7185643,4.0992823,3.8301542,2.7831798,1.2964103,8.024616,9.271795,5.8453336,1.2832822,1.8609232,1.3161026,1.3357949,1.5064616,1.5819489,1.4802053,1.6836925,1.8182565,1.8281027,1.8116925,1.9889232,1.9167181,1.8149745,1.7624617,1.7066668,1.4506668,1.2635899,1.3456411,1.5622566,1.8707694,2.3368206,1.8313848,1.8051283,1.8543591,1.8510771,1.9495386,1.9954873,2.2908719,2.5271797,2.6518977,2.861949,2.9078977,3.1474874,3.31159,3.31159,3.242667,2.7831798,2.7076926,2.6486156,2.5895386,2.8849232,2.9013336,2.9735386,3.1442053,3.239385,2.8717952,2.878359,3.3542566,4.06318,4.6572313,4.6802053,5.1987696,6.163693,7.276308,8.395488,9.547488,10.929232,12.225642,13.210258,13.984821,14.992412,15.986873,17.30954,19.5479,22.370462,24.523489,23.77518,23.67672,23.922874,24.448002,25.442463,26.78154,27.155695,27.044106,26.423798,24.786053,25.570463,26.285952,26.368002,25.790361,25.08472,26.285952,26.112001,25.731283,25.54749,25.173336,24.395489,24.365952,24.047592,23.502771,23.867079,23.545437,24.592413,26.102156,26.420515,23.135181,20.585028,19.88595,20.70318,22.258873,23.345232,22.734772,22.42954,22.728207,23.213951,22.754463,22.032412,21.225027,19.51836,17.174976,15.504412,14.8480015,13.748514,12.173129,10.456616,9.330873,8.864821,7.709539,6.7249236,6.485334,7.2861543,7.3682055,7.138462,6.9710774,7.0531287,7.387898,7.53559,8.136206,8.493949,8.372514,8.008205,8.667898,9.718155,10.8537445,11.936821,13.003489,13.958565,14.027489,13.53518,13.180719,14.043899,14.949745,14.467283,13.50236,12.737642,12.629334,12.609642,12.964104,13.266052,13.318565,13.164309,12.754052,12.2387705,11.703795,11.428103,11.881026,11.513436,10.528821,9.432616,8.608821,8.346257,8.264206,7.972103,7.1187696,5.677949,3.9811285,3.2623591,2.612513,2.2219489,2.1070771,2.1103592,2.15959,2.6420515,3.1934361,3.5872824,3.7218463,2.8389745,2.934154,2.7766156,2.4582565,2.2350771,2.5009232,2.5009232,2.6387694,2.5238976,2.1530259,1.9232821,2.4713848,2.4615386,2.3269746,2.359795,2.7011285,2.7995899,3.2984617,3.5905645,3.8006158,4.775385,6.2785645,6.8627696,7.755488,8.891078,8.92718,9.426052,9.764103,9.242257,8.556309,9.764103,9.081436,11.82195,16.41354,19.318155,15.044924,6.4754877,3.0523078,2.15959,2.028308,1.723077,2.0775387,2.0841026,2.041436,2.0841026,2.1825643,1.6082052,1.5392822,1.4539489,1.2668719,1.3259488,1.1684103,1.3751796,1.6804104,1.8510771,1.6935385,1.522872,1.6443079,1.723077,1.6311796,1.4342566,1.5195899,1.4769232,1.6607181,1.8838975,1.4178462,1.4802053,1.5031796,1.4309745,1.2996924,1.2504616,1.276718,1.1716924,0.98133343,0.78769237,0.702359,0.702359,0.77456415,0.96492314,1.1454359,1.024,0.79097444,0.6498462,0.67282057,0.7844103,0.74830776,0.29538465,0.2297436,0.21661541,0.15097436,0.15097436,0.27569234,0.6268718,1.2307693,1.9561027,2.5173335,3.190154,4.630975,6.3376417,8.480822,11.88759,15.95077,17.562258,17.06995,15.409232,14.112822,15.333745,17.434258,18.894772,19.551182,20.614565,23.190975,24.805746,23.046566,18.517334,14.831591,15.392821,17.161848,19.531488,22.14072,24.887796,25.458874,25.951181,26.95877,27.047386,22.75118,16.305231,11.040821,6.9809237,4.276513,3.190154,2.4582565,2.100513,1.9528207,1.9364104,2.044718,1.9364104,1.9790771,2.0217438,1.9561027,1.723077,1.6278975,0.8041026,0.28225642,0.26912823,0.18379489,1.8313848,2.2416413,2.2383592,2.5009232,3.5872824,6.550975,9.472001,15.209026,22.111181,24.018053,22.344208,23.033438,24.103386,24.139488,22.308104,19.817028,20.420925,22.46236,25.314463,29.4039,33.10277,34.550156,34.097233,33.16841,34.254772,33.010876,29.761642,27.703796,27.966362,29.600822,30.614977,32.295387,34.54359,36.562054,36.880413,36.197746,34.845543,33.17826,31.501131,30.06031,29.974977,29.184002,28.097643,27.460926,28.35036,28.973951,28.048412,26.59118,25.133951,23.742361,22.314669,22.104616,24.116514,27.336206,28.71795,27.556105,26.407387,25.51467,24.480822,22.245745,20.292925,18.937437,18.12349,17.237335,15.074463,13.072412,12.921437,13.59754,14.598565,15.931078,18.274464,22.17354,25.06831,25.570463,23.483078,21.077335,20.201027,19.02277,17.818258,18.966976,20.17477,17.867489,15.481437,14.690463,15.412514,18.20554,22.505028,25.550772,26.351591,25.682053,23.532309,21.366156,20.25354,20.722874,22.734772,24.95672,25.796925,24.520206,21.559797,18.507488,15.77354,14.588719,15.291079,15.960617,12.422565,9.882257,9.659078,10.262975,12.1468725,17.700104,20.630976,19.541334,16.52513,13.019898,9.796924,8.342975,9.737847,11.063796,10.427077,6.9743595,5.9602056,7.4732313,10.105436,11.1294365,6.514872,5.405539,5.474462,4.890257,4.522667,7.965539,9.711591,7.90318,7.2861543,8.297027,7.066257,13.216822,18.81272,21.99631,22.436104,21.300514,24.46113,17.188105,10.656821,8.205129,5.32677,4.07959,3.8498464,4.644103,5.789539,5.937231,4.6539493,4.1583595,4.240411,4.670359,5.218462,4.023795,2.937436,2.1858463,1.910154,2.166154,3.3378465,3.9056413,3.8498464,3.4789746,3.4166157,3.2229745,2.2482052,1.332513,0.88287187,0.86974365,0.77128214,1.086359,1.1848207,1.2077949,2.0742567,2.7831798,3.9220517,5.21518,6.1407185,5.920821,4.9920006,3.9647183,2.4024618,0.76800007,0.4266667,0.69579494,0.7811283,0.7253334,0.6170257,0.58092314,0.5316923,0.6662565,1.024,1.3029745,0.8402052,0.38728207,0.20020515,0.14112821,0.190359,0.45620516,0.51856416,0.3314872,0.3708718,0.60389745,0.51856416,0.16410258,0.029538464,0.0,0.0,0.0,0.0,0.009846155,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.02297436,0.04594872,0.04594872,0.036102567,0.04266667,0.101743594,0.25928208,0.35774362,0.51856416,0.8008206,1.1520001,1.4342566,1.2274873,1.6771283,2.8389745,4.266667,5.034667,5.024821,5.421949,5.3858466,4.8016415,4.2863593,1.3456411,0.28882053,0.08861539,0.118153855,0.16738462,0.23958977,0.37743592,0.40369233,0.318359,0.3052308,0.23302566,0.2231795,0.25928208,0.3052308,0.3052308,0.26912823,0.23302566,0.23302566,0.2855385,0.39712822,0.41025645,0.4201026,0.39056414,0.3314872,0.32164106,0.3708718,0.446359,0.5874872,0.74830776,0.80738467,0.80738467,0.8467693,0.8205129,0.80738467,1.0535386,1.1388719,1.1126155,1.3161026,1.8871796,2.7766156,3.1081028,3.2984617,4.1091285,5.5893335,7.066257,7.955693,8.260923,8.303591,8.198565,7.8441033,7.256616,6.9349747,6.5936418,6.157129,5.7665644,5.5729237,6.0652313,6.954667,8.050873,9.245539,8.930462,8.851693,8.513641,7.752206,6.7150774,6.872616,6.6461544,6.2063594,5.6943593,5.218462,5.546667,5.7042055,5.5565133,5.1232824,4.562052,3.5741541,3.308308,3.3378465,3.2787695,2.7766156,2.3630772,2.2121027,2.176,2.3236926,2.9440002,3.006359,3.239385,3.259077,3.0293336,2.8849232,2.1530259,2.1070771,2.044718,1.9298463,2.3794873,2.6978464,3.5905645,5.0149746,6.7183595,8.27077,9.110975,8.982975,8.52677,7.9524107,7.0498466,3.9614363,5.579488,7.640616,7.8112826,5.677949,13.538463,11.657847,6.9349747,3.895795,4.699898,4.1747694,4.3552823,4.5062566,4.092718,2.7602053,3.2886157,5.98318,5.156103,1.4342566,1.7394873,1.214359,1.2668719,1.5097437,1.6147693,1.2964103,1.785436,1.9429746,1.9068719,1.8445129,1.9528207,1.3915899,1.5983591,1.7099489,1.4506668,1.1454359,1.4867693,1.4441026,1.4933335,1.7165129,1.8018463,1.7165129,1.785436,1.8346668,1.8510771,1.9987694,1.8412309,2.231795,2.5107694,2.605949,3.0227695,3.1934361,3.3280003,3.370667,3.2065644,2.6715899,2.6584618,2.674872,2.4976413,2.297436,2.6387694,2.674872,2.4385643,2.5042052,2.934154,3.249231,3.5314875,3.4822567,3.6529233,4.1091285,4.4242053,5.5958977,7.3649235,8.572719,9.147078,10.085744,12.343796,14.12595,15.018668,15.05477,14.723283,15.983591,17.604925,19.643078,21.851898,23.683285,24.195284,24.431591,25.11754,26.138258,26.564924,27.992617,27.812105,27.339489,27.290258,27.739899,29.023182,29.279182,28.727797,27.418259,25.206156,25.69518,26.22031,26.305643,25.833027,25.03877,24.12308,24.608822,24.90749,24.598976,24.42831,24.037745,24.234669,25.16677,25.747694,23.637335,22.255592,21.828924,22.373745,23.371489,23.7719,22.577232,22.104616,22.347488,23.108925,23.985233,23.11877,21.658258,19.265642,16.49559,14.785643,14.273643,13.2562065,11.644719,9.980719,9.429334,7.965539,7.2861543,7.030154,7.0793853,7.568411,7.2861543,7.2894363,7.6274877,8.034462,7.9491286,8.487385,8.667898,8.667898,8.4972315,7.9950776,8.851693,9.760821,10.676514,11.746463,13.321847,13.797745,13.5778475,13.266052,13.348104,14.191591,14.667488,14.319591,13.525334,12.714667,12.360206,12.2617445,12.905026,13.338258,13.154463,12.481642,11.798975,11.168821,10.962052,11.113027,11.122872,10.256411,9.472001,8.697436,8.054154,7.857231,7.24677,6.738052,5.7796926,4.4307694,3.3575387,2.7470772,2.4385643,2.2186668,2.0644104,2.1366155,2.6617439,3.131077,3.4855387,3.7842054,4.210872,2.6420515,2.5271797,2.678154,2.678154,2.484513,2.428718,2.3302567,2.422154,2.4385643,2.297436,2.0939488,2.3794873,2.3269746,2.2055387,2.2055387,2.4188719,2.5271797,2.986667,3.4494362,3.9614363,4.9460516,5.8518977,6.5378466,7.499488,8.546462,8.828718,9.905231,10.509129,10.098872,9.235693,9.593436,8.802463,10.807796,14.441027,16.502155,11.762873,5.3792825,2.789744,2.0578463,1.972513,2.028308,2.550154,2.8455386,2.8849232,2.8192823,2.9768207,2.4910772,2.1497438,1.7558975,1.3653334,1.2800001,1.404718,1.6804104,1.8051283,1.719795,1.6213335,1.8018463,1.8281027,1.6738462,1.4244103,1.2865642,1.2668719,1.2471796,1.339077,1.4539489,1.3226668,1.529436,1.4080001,1.332513,1.3883078,1.3489232,1.5885129,1.463795,1.0601027,0.6662565,0.78769237,0.827077,1.086359,1.273436,1.2176411,0.85005134,0.6892308,0.6301539,0.6170257,0.58092314,0.4660513,0.27897438,0.19692309,0.15097436,0.13456412,0.21333335,0.5218462,0.8730257,1.4605129,2.225231,2.8849232,3.5938463,4.5817437,5.687795,7.0104623,8.933744,12.022155,14.480412,15.527386,15.625848,16.469334,19.751387,21.881437,21.769848,20.027079,18.980104,19.659489,18.041437,15.540514,14.017642,15.770258,19.43959,24.746668,30.388515,35.862976,41.452312,42.033234,39.364925,35.0359,29.735388,23.250053,16.79754,11.625027,7.7718983,5.07077,3.1638978,2.6945643,2.537026,2.3794873,2.231795,2.412308,2.281026,3.0194874,3.8367183,4.342154,4.519385,4.7917953,3.5971284,2.162872,1.2012309,0.88943595,1.7591796,2.8389745,3.6135387,4.2174363,5.4416413,6.3573337,8.946873,13.512206,18.04472,18.231796,19.410053,20.41108,20.97231,21.11672,21.159386,20.30277,20.118977,21.464617,23.975386,26.082464,29.656618,33.194668,34.73067,34.47467,34.829132,34.747078,33.670567,31.48472,29.213541,29.003489,30.34913,31.11713,32.466053,34.179283,34.68472,35.718567,36.10585,34.97354,32.66626,30.756105,30.992413,30.25395,28.649029,26.919386,26.433643,27.798977,27.690668,27.316515,26.788105,25.120823,23.995079,23.745644,25.376822,28.432413,30.962873,28.777027,26.902977,26.315489,26.555079,25.737848,23.952412,22.816822,22.009438,20.453745,16.321642,13.938873,12.760616,12.563693,13.292309,15.064616,17.427694,20.562054,24.119797,27.204926,28.376617,25.426054,24.25108,22.459078,19.77436,18.051283,19.045746,17.24718,15.304206,14.634667,15.42236,18.100513,21.848618,24.513643,25.737848,26.948925,24.595694,23.19754,22.386873,22.370462,23.955694,26.020105,25.69518,23.5159,20.502975,18.15631,14.523078,12.868924,12.248616,11.444513,8.979693,7.250052,7.0400004,7.525744,9.386667,14.795488,16.328207,14.772514,12.652308,11.024411,9.4916935,9.416205,9.705027,9.662359,8.73354,6.5083084,6.091488,11.753027,13.22995,9.042052,6.47877,4.2830772,6.747898,6.7150774,3.7743592,4.266667,5.9634876,7.315693,8.979693,9.780514,6.7117953,12.356924,15.104001,16.416822,16.889437,16.272411,23.827694,16.676104,9.360411,6.8529234,4.568616,2.9997952,2.8750772,3.564308,4.1714873,3.5183592,2.412308,2.1891284,2.4746668,2.8455386,2.8389745,2.1989746,1.7920002,1.6180514,1.7526156,2.3630772,2.5961027,2.4155898,2.3663592,2.9965131,4.857436,7.3091288,5.172513,2.6551797,1.8281027,2.6289232,3.1343591,3.4756925,3.3772311,2.9636924,2.7470772,2.284308,2.5928206,3.6824617,5.0642056,5.7632823,6.055385,4.854154,2.8422565,0.98133343,0.512,0.47917953,0.34789747,0.24943592,0.2855385,0.54482055,1.8806155,1.2209232,0.8336411,1.3029745,1.522872,1.0404103,0.636718,0.45292312,0.44307697,0.36102566,0.2855385,0.14441027,0.11158975,0.17066668,0.1148718,0.055794876,0.016410258,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.01969231,0.026256412,0.04266667,0.09189744,0.2231795,0.36102566,0.7515898,1.2307693,1.6705642,1.972513,1.529436,1.5622566,2.422154,4.0402055,5.9503593,6.3277955,6.0291286,5.72718,5.7534366,6.0816417,3.5413337,1.7132308,0.574359,0.059076928,0.068923086,0.1148718,0.21333335,0.28882053,0.32820517,0.4135385,0.30194873,0.32164106,0.3708718,0.40697438,0.4266667,0.4004103,0.2986667,0.24615386,0.28882053,0.41025645,0.39056414,0.39056414,0.38728207,0.3708718,0.30851284,0.40697438,0.58092314,0.6498462,0.65641034,0.892718,0.8172308,0.8467693,0.98461545,1.1552821,1.2242053,1.2209232,1.5031796,1.8806155,2.176,2.228513,2.7044106,3.4658465,4.450462,5.6352825,7.0531287,8.257642,8.507077,8.15918,7.765334,8.073847,7.39118,6.5411286,6.0225644,5.986462,6.232616,5.802667,6.5345645,7.4797955,8.093539,8.234667,7.827693,7.765334,7.683283,7.3649235,6.7249236,6.485334,6.121026,5.8190775,5.6451287,5.5597954,5.5958977,5.3792825,4.9394875,4.3290257,3.623385,2.556718,2.5271797,2.7667694,2.8717952,2.802872,2.1924105,2.044718,2.1497438,2.3696413,2.6387694,2.2219489,2.176,2.28759,2.3663592,2.2482052,1.6935385,1.7132308,1.719795,1.657436,2.0020514,2.5337439,3.5249233,5.041231,7.0826674,9.6,9.682052,8.681026,7.824411,7.197539,5.7665644,2.865231,2.2580514,2.7634873,3.383795,3.308308,7.9458466,7.069539,4.713026,3.4724104,4.493129,3.948308,3.692308,3.4231799,2.934154,2.103795,2.1989746,2.7142565,2.425436,1.5195899,1.5819489,1.2209232,1.3292309,1.4375386,1.3292309,1.0404103,1.4309745,1.6016412,1.5622566,1.463795,1.6246156,1.1684103,1.1848207,1.2012309,1.1027694,1.1191796,1.2964103,1.5491283,1.6640002,1.6344616,1.6410258,1.7920002,1.7657437,1.6672822,1.6278975,1.8051283,1.9364104,2.1366155,2.3860514,2.7241027,3.2656412,3.2229745,3.2361028,3.0687182,2.6683078,2.169436,2.284308,2.3105643,2.2482052,2.2547693,2.6157951,2.865231,2.7634873,2.806154,3.058872,3.1540515,3.1606157,3.4297438,3.8104618,4.2502565,4.8049235,6.0717955,7.4174366,8.723693,10.000411,11.378873,13.853539,14.92677,15.258258,15.428925,15.970463,16.62031,17.64759,19.275488,21.287386,23.010464,24.159182,24.438156,25.120823,26.207182,26.420515,27.290258,27.890875,27.90072,27.700516,28.386463,29.443285,29.38749,28.898464,27.979488,25.977438,25.577028,25.813335,25.606565,24.917336,24.759796,23.968822,23.91631,24.795898,26.000412,26.115284,24.628515,24.22154,24.736822,25.403078,24.84513,23.522463,22.94154,23.09908,23.624207,23.7719,22.800411,22.258873,22.646156,23.801437,24.914053,24.116514,22.35077,19.702156,16.899282,15.287796,15.028514,14.037334,12.435693,10.601027,9.173334,8.362667,8.119796,7.9524107,7.7981544,8.03118,7.906462,7.3780518,7.197539,7.4699492,7.6701546,8.214975,8.39877,8.507077,8.421744,7.6176414,8.326565,9.6295395,10.912822,11.949949,12.918155,13.092104,12.928001,12.934566,13.3251295,14.03077,14.362258,14.168616,13.528616,12.694975,12.068104,12.232206,13.029744,13.269335,12.744206,12.248616,11.605334,10.758565,10.138257,9.957745,10.243283,9.944616,9.271795,8.5661545,8.018052,7.686565,7.322257,6.4557953,5.2381544,4.013949,3.3214362,3.2164104,3.255795,3.114667,2.865231,2.9669745,3.0523078,3.2787695,3.5610259,3.8564105,4.1747694,2.6683078,2.678154,2.7044106,2.7536411,2.7634873,2.5928206,2.3991797,2.3401027,2.300718,2.228513,2.1366155,2.2383592,2.4155898,2.481231,2.422154,2.3762052,2.5961027,2.8160002,3.190154,3.8432825,4.8607183,5.668103,6.426257,7.200821,7.9491286,8.503796,9.577026,10.194052,10.105436,9.458873,8.802463,7.7357955,8.772923,11.323078,13.147899,10.354873,5.47118,3.4100516,2.7733335,2.6518977,2.609231,2.7667694,2.6617439,2.422154,2.2908719,2.6157951,2.5993848,2.4943593,2.156308,1.7099489,1.5589745,1.6082052,1.8609232,1.9495386,1.8051283,1.6836925,1.7558975,1.6311796,1.5622566,1.5392822,1.3062565,1.2504616,1.214359,1.394872,1.6377437,1.4342566,1.4080001,1.339077,1.3226668,1.3456411,1.3095386,1.3686155,1.1323078,0.88943595,0.90256417,1.404718,1.8707694,2.03159,1.8018463,1.2504616,0.6268718,0.44964105,0.40697438,0.380718,0.3446154,0.34133336,0.26256412,0.19364104,0.13456412,0.11158975,0.16410258,0.32820517,0.58092314,1.0404103,1.6705642,2.28759,3.2065644,4.2962055,5.4482055,6.7117953,8.323282,10.397539,12.665437,14.411489,15.809642,17.929848,21.520412,22.33436,21.40554,19.46913,16.948515,16.160822,14.385232,13.344822,14.391796,18.487797,24.753233,31.054771,37.06749,42.04308,44.84267,44.022156,39.758774,33.81826,27.575796,22.029129,16.833643,12.314258,9.147078,6.997334,4.5128207,4.2141542,4.2272825,4.076308,3.7120004,3.5183592,2.5206156,2.8127182,3.5249233,4.201026,4.7983594,5.684513,5.4580517,4.8147697,3.692308,1.2603078,1.3226668,1.8379488,2.609231,3.3608208,3.7185643,5.2053337,7.529026,10.916103,14.519796,16.390566,18.796309,20.824617,20.181335,18.159592,19.639797,20.94277,20.785233,21.218464,22.721643,24.201847,25.872412,29.400618,32.833645,35.091694,35.981133,34.95713,34.704414,33.12903,30.683899,30.355694,31.504414,31.789951,31.701336,31.760412,32.512,32.800823,32.735184,32.01313,30.851284,30.004515,30.211285,29.850258,29.144617,28.146873,26.7159,26.479591,27.401848,28.73108,29.331694,27.67426,26.417233,25.846155,26.794668,29.075695,31.46831,28.970669,26.584618,25.98072,26.965336,27.490463,27.493746,26.558361,24.704002,21.786259,17.483488,15.202463,13.495796,12.58995,12.711386,14.086565,16.111591,18.678156,22.442669,26.971899,30.756105,29.892925,28.406157,25.265232,21.00513,17.723078,17.394873,16.052513,14.9398985,14.726565,15.471591,18.14318,21.297232,23.112207,23.985233,26.535387,26.738874,24.81231,23.315695,23.427284,24.95672,25.93477,24.51036,21.737028,18.582975,15.944206,12.422565,9.714872,8.966565,9.140513,7.000616,5.907693,5.5171285,5.7665644,7.6012316,12.987078,14.208001,11.923694,10.246565,10.095591,9.202872,9.120821,8.490667,8.55959,8.868103,7.2369237,6.170257,10.712616,10.886565,6.308103,6.166975,7.0859494,11.280411,9.622975,3.2262566,3.4527183,4.125539,7.581539,10.827488,11.464206,7.6668725,13.249642,14.162052,12.609642,11.139283,12.642463,21.041233,13.617231,6.4065647,4.7524104,3.2886157,2.5271797,2.3794873,2.7142565,2.9636924,2.1169233,1.3554872,1.4342566,1.9167181,2.297436,1.9954873,1.5261539,1.3029745,1.2800001,1.4900514,2.0545642,2.0841026,1.7296412,1.5261539,2.044718,3.882667,5.3760004,5.868308,5.1889234,3.8564105,3.0851285,3.9056413,5.1298466,5.097026,3.754667,2.6584618,3.1540515,2.9440002,3.5446157,4.9099493,5.428513,5.156103,4.07959,2.8127182,1.7657437,1.148718,0.8041026,0.64000005,0.55794877,0.8008206,1.9429746,1.8838975,1.3128207,1.4309745,2.3991797,3.3312824,1.5491283,0.702359,0.46933338,0.51856416,0.508718,0.34789747,0.14769232,0.036102567,0.026256412,0.006564103,0.009846155,0.016410258,0.009846155,0.0032820515,0.009846155,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.0,0.01969231,0.032820515,0.052512825,0.098461546,0.21333335,0.2297436,0.64000005,1.4408206,2.4057438,3.0851285,2.5271797,1.975795,1.9462565,2.5698464,3.5807183,5.717334,5.986462,5.9667697,6.2687182,6.547693,5.3234878,4.562052,2.8521028,0.60389745,0.055794876,0.06235898,0.14112821,0.22646156,0.2986667,0.37743592,0.32820517,0.3511795,0.42994875,0.49230772,0.39384618,0.36102566,0.33805132,0.33476925,0.36758977,0.4397949,0.40697438,0.36758977,0.39712822,0.45292312,0.34133336,0.34789747,0.574359,0.7318975,0.76800007,0.84348726,1.1191796,1.0272821,0.98133343,1.0765129,1.0929232,1.2307693,1.6508719,2.097231,2.3696413,2.3269746,2.2777438,3.0424619,4.2929235,5.7468724,7.1876926,7.860513,8.474257,8.392206,7.7423596,7.427283,6.7577443,6.1407185,5.8912826,5.989744,6.1013336,5.910975,6.951385,7.857231,7.9458466,7.200821,7.0465646,7.076103,7.069539,6.9120007,6.564103,6.1341543,5.720616,5.61559,5.6976414,5.4547696,5.540103,5.0642056,4.3060517,3.5446157,3.0490258,2.3958976,2.5271797,2.681436,2.5764105,2.422154,1.975795,1.9889232,1.9659488,1.8904617,2.2055387,2.2416413,1.9364104,1.7624617,1.847795,2.0184617,1.591795,1.6278975,1.6311796,1.5655385,1.8609232,2.6453335,3.748103,5.024821,6.6002054,8.891078,8.786052,7.7259493,7.3353853,7.2894363,5.3103595,2.5042052,1.3489232,1.0896411,1.2635899,1.7099489,4.020513,4.4307694,4.1189747,3.8465643,3.945026,3.3805132,3.062154,2.934154,2.7864618,2.231795,1.6705642,1.5064616,1.4834872,1.4473847,1.3587693,1.2012309,1.270154,1.2406155,1.0765129,1.0305642,1.3095386,1.3587693,1.273436,1.1782565,1.2012309,1.1060513,1.1684103,1.1979488,1.1257436,1.0305642,1.0404103,1.3423591,1.7723079,2.0118976,1.5753847,1.657436,1.7329233,1.8642052,2.0184617,2.048,2.100513,2.3433847,2.6387694,2.878359,2.9604106,2.8914874,2.9013336,2.6486156,2.2186668,2.1267693,2.03159,2.0250258,2.0808206,2.1431797,2.1530259,2.6322052,2.9144619,3.2000003,3.3641028,2.9538465,2.550154,3.1934361,3.8728209,4.332308,5.080616,5.861744,6.738052,8.444718,10.801231,12.701539,15.169642,15.602873,15.698052,16.278976,17.28,17.30954,18.20554,19.610258,21.251284,22.92513,23.732515,24.1559,24.884514,26.164515,27.80226,28.137028,28.918156,29.078976,28.475079,27.881027,28.209232,28.78031,28.82954,27.96308,26.14154,25.38667,24.891079,24.329847,23.880207,24.241232,23.768618,23.558565,24.310156,25.51795,25.472002,23.752207,23.542156,24.106668,24.795898,25.074873,24.169027,23.289438,23.017027,23.35836,23.745644,23.555285,23.095797,23.27631,24.270771,25.521233,24.425028,22.442669,19.744822,17.122463,15.986873,15.842463,14.729847,13.154463,11.355898,9.31118,8.92718,9.107693,8.973129,8.55959,8.789334,8.2215395,7.4863596,7.213949,7.529026,8.0377445,8.448001,8.576,8.569437,8.326565,7.4765134,8.251078,9.734565,10.994873,11.795693,12.596514,12.747488,12.599796,12.596514,12.941129,13.59754,14.191591,13.860104,13.154463,12.504617,12.212514,12.475078,12.960821,13.098668,12.740924,12.173129,11.618463,10.614155,9.741129,9.363693,9.622975,9.419488,8.687591,8.103385,7.906462,7.893334,7.328821,6.294975,5.0674877,4.0041027,3.5314875,3.5905645,3.748103,3.692308,3.4921029,3.5872824,3.4231799,3.4822567,3.6562054,3.7743592,3.6430771,2.5435898,2.6683078,2.537026,2.5337439,2.681436,2.6354873,2.4057438,2.3302567,2.2646155,2.1891284,2.1956925,2.1234872,2.3762052,2.5600002,2.5238976,2.3762052,2.6715899,2.7273848,3.0260515,3.7251284,4.6539493,5.536821,6.442667,7.1515903,7.7718983,8.753231,9.396514,9.829744,9.915077,9.396514,7.9228725,7.0367184,7.680001,9.458873,11.021129,10.049642,6.2884107,4.204308,3.3411283,3.1671798,3.062154,2.5764105,2.1136413,1.9035898,2.0118976,2.3696413,2.4943593,2.5206156,2.3302567,2.0217438,1.913436,1.9429746,2.1333334,2.100513,1.8149745,1.6114873,1.529436,1.3718976,1.3915899,1.4966155,1.2504616,1.1749744,1.2438976,1.4506668,1.595077,1.2996924,1.2537436,1.1585642,1.083077,1.083077,1.211077,1.2012309,1.0929232,1.0929232,1.3193847,1.782154,2.176,2.0709746,1.6246156,1.024,0.49887183,0.3314872,0.27569234,0.24287182,0.21989745,0.26256412,0.21989745,0.190359,0.17066668,0.14441027,0.1148718,0.14769232,0.3446154,0.6432821,1.0338463,1.5753847,2.556718,3.6627696,4.890257,6.2687182,7.8637953,9.366975,11.099898,12.901745,14.769232,16.843489,18.868515,18.62236,17.979078,17.273438,15.320617,14.293334,13.426873,13.308719,14.697027,18.517334,23.91631,28.806566,33.076515,35.974567,36.12226,34.94072,31.872002,27.700516,23.3879,20.082872,16.400412,12.983796,10.811078,9.357129,6.5936418,5.756718,5.2414365,4.962462,4.6900516,4.066462,3.1803079,3.186872,3.239385,3.2656412,3.9680004,4.886975,5.139693,5.5204105,5.2315903,1.8838975,1.2832822,1.1651284,1.5491283,2.2219489,2.740513,4.1682053,6.5837955,10.020103,13.994668,17.513027,20.118977,21.080618,19.859694,17.99549,19.114668,22.193232,21.983181,21.17908,21.248001,22.42954,23.824411,26.906258,30.759386,34.264618,36.115696,34.802876,34.304,33.16185,31.783386,32.466053,32.81067,32.915695,31.72431,30.116104,30.90708,30.500105,29.518772,28.678566,28.324104,28.419285,28.836105,28.616207,28.471798,28.182976,26.5879,26.22359,27.46749,29.200413,30.309746,29.69272,28.288002,27.047386,26.788105,27.736618,29.541746,28.022156,25.99713,25.330873,26.345028,27.815386,28.57026,27.96308,26.09231,23.138464,19.328001,17.007591,14.431181,12.790154,12.445539,12.944411,14.536206,16.827078,20.558771,25.465437,30.25067,31.780106,30.129232,26.151386,21.392412,18.074257,16.968206,15.261539,14.421334,14.788924,15.563488,17.893745,20.483284,21.563078,21.622156,23.410873,24.270771,22.79713,22.229336,23.571693,25.580309,25.829746,23.80472,20.850874,17.447386,13.190565,10.029949,7.026872,6.5017443,7.39118,5.2480006,4.854154,4.6572313,4.663795,6.12759,11.54954,14.04718,11.785847,10.036513,10.089026,9.278359,8.057437,7.8834877,8.726975,9.580308,8.487385,8.746667,11.254155,9.7673855,5.668103,7.9491286,13.735386,17.083078,12.406155,3.6430771,4.269949,4.0402055,7.79159,11.122872,11.355898,7.532308,12.86236,13.906053,10.8537445,6.7774363,7.6077952,16.705643,10.761847,5.110154,4.397949,2.5928206,2.3171284,2.097231,2.156308,2.231795,1.5688206,1.0962052,1.3686155,1.9692309,2.3236926,1.719795,1.1684103,0.92553854,0.90256417,1.142154,1.8051283,3.2131286,2.8521028,1.8806155,1.6475899,3.6627696,3.8728209,6.514872,7.3485136,5.7698464,4.818052,7.4830775,8.897642,8.3364105,6.380308,4.923077,4.919795,3.9384618,3.7054362,4.637539,5.8453336,6.409847,4.8607183,3.1343591,2.1300514,1.7033848,1.4769232,1.2570257,1.8248206,3.0162053,3.7185643,4.1846156,4.384821,4.135385,3.6758976,3.6627696,1.4145643,0.6268718,0.636718,0.8992821,0.9911796,0.44964105,0.15097436,0.026256412,0.0032820515,0.0,0.0,0.009846155,0.009846155,0.0032820515,0.009846155,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.006564103,0.026256412,0.032820515,0.04594872,0.08205129,0.15753847,0.108307704,0.4594872,1.1552821,2.0841026,3.0916924,3.2295387,2.3368206,1.6508719,1.5458462,1.5097437,4.578462,5.0609236,5.100308,5.425231,5.35959,5.428513,5.113436,4.013949,2.1891284,0.16410258,0.07876924,0.10502565,0.17066668,0.24615386,0.36102566,0.36430773,0.36102566,0.4397949,0.51856416,0.3446154,0.30194873,0.34133336,0.38400003,0.39712822,0.4135385,0.40369233,0.3511795,0.3708718,0.4201026,0.3117949,0.25928208,0.4266667,0.6170257,0.7384616,0.8041026,1.1158975,1.0568206,0.9682052,0.9944616,1.0732309,1.3587693,1.8576412,2.2383592,2.4188719,2.5435898,2.2219489,2.9538465,4.519385,6.377026,7.6570263,7.7981544,8.139488,8.192,7.719385,6.7249236,6.2851286,5.858462,5.737026,5.910975,6.0750775,6.2916927,7.0137444,7.5913854,7.565129,6.633026,6.62318,6.51159,6.422975,6.3967185,6.3934364,6.042257,5.756718,5.7632823,5.924103,5.7534366,5.6254363,4.906667,3.8695388,2.8914874,2.4615386,2.15959,2.4549747,2.605949,2.4385643,2.3368206,1.9364104,1.782154,1.5458462,1.3456411,1.7493335,2.1136413,1.8871796,1.6344616,1.6607181,2.0118976,1.8412309,1.719795,1.6246156,1.6311796,1.910154,2.7864618,4.017231,5.290667,6.3901544,7.1876926,7.0793853,6.5805135,7.197539,8.086975,6.048821,2.9833848,1.7165129,1.2373334,1.1848207,1.8674873,2.4451284,3.4002054,4.1222568,4.342154,4.135385,3.1507695,2.7076926,2.986667,3.3444104,2.297436,1.6344616,1.6049232,1.6902566,1.5688206,1.1257436,1.1618463,1.1749744,1.1093334,1.0305642,1.142154,1.214359,1.2340513,1.1684103,1.0338463,0.8960001,1.1027694,1.2242053,1.2668719,1.214359,1.0436924,0.9911796,1.1552821,1.6082052,1.9954873,1.5130258,1.6935385,1.9692309,2.2711797,2.412308,2.097231,2.2088206,2.5140514,2.806154,2.8849232,2.5895386,2.5731285,2.5698464,2.3302567,1.9922053,2.0611284,1.9561027,1.8838975,2.0020514,2.162872,1.9331284,2.4713848,2.9472823,3.2754874,3.2984617,2.7634873,2.2580514,3.0523078,3.9942567,4.644103,5.284103,6.0160003,7.1187696,8.910769,11.16554,13.111795,14.992412,15.527386,16.075489,17.106052,18.20554,18.54031,19.226257,20.28636,21.59918,22.905437,24.192001,24.65149,24.969849,25.777233,27.654566,28.054977,28.931284,29.462976,29.134771,27.72349,27.503592,28.21908,28.271591,26.981745,24.579285,23.745644,23.348515,22.869335,22.560822,23.446976,23.460104,23.296001,23.712822,24.4119,24.04431,22.596926,22.724924,23.496206,24.31672,24.90749,24.297028,23.273027,22.81354,23.158155,23.817848,24.388926,24.195284,24.297028,25.078156,26.246567,24.87795,22.6199,19.846565,17.444103,16.807386,16.754873,15.323898,13.686155,12.074668,9.780514,9.321027,9.793642,9.826463,9.347282,9.577026,8.480822,7.683283,7.50277,7.965539,8.832001,8.79918,8.546462,8.195283,7.8802056,7.75877,8.585847,9.609847,10.59118,11.47077,12.3766165,12.419283,12.12718,12.150155,12.675283,13.4400015,13.748514,13.144616,12.425847,12.048411,12.114052,12.278154,12.553847,12.612924,12.3076935,11.667693,11.273847,10.217027,9.360411,9.042052,9.068309,8.874667,8.342975,8.011488,7.958975,7.8080006,6.9677954,5.9602056,4.9099493,4.0369234,3.6726158,3.6726158,3.7021542,3.6135387,3.4921029,3.639795,3.5840003,3.5610259,3.629949,3.6562054,3.2886157,2.2744617,2.3433847,2.228513,2.231795,2.4057438,2.556718,2.3893335,2.428718,2.3991797,2.281026,2.3105643,2.0939488,2.2022567,2.3236926,2.3466668,2.3466668,2.5993848,2.6453335,2.9768207,3.6791797,4.4274874,5.3792825,6.426257,7.24677,8.001641,9.350565,9.452309,9.6984625,9.7673855,9.216001,7.460103,7.3452315,8.034462,9.114257,10.102155,10.469745,7.90318,5.1954875,3.5380516,3.0982566,2.986667,2.0053334,1.6377437,1.9659488,2.5731285,2.5271797,2.300718,2.1792822,2.0841026,2.0086155,2.0053334,2.103795,2.172718,1.9528207,1.5195899,1.2865642,1.2471796,1.1979488,1.1913847,1.1848207,1.0535386,1.0108719,1.1881026,1.2931283,1.204513,0.9944616,1.1027694,0.86317956,0.65641034,0.7056411,1.0601027,1.2242053,1.4244103,1.5786668,1.6672822,1.7165129,1.5622566,1.204513,0.85005134,0.5973334,0.45620516,0.34133336,0.27569234,0.24287182,0.2231795,0.17723078,0.13784617,0.15097436,0.18051283,0.190359,0.1148718,0.20348719,0.42994875,0.61374366,0.81066674,1.3128207,2.172718,3.058872,4.141949,5.4482055,6.8496413,8.080411,9.32759,10.794667,12.343796,13.482668,13.545027,13.351386,13.728822,14.503386,14.477129,14.063591,13.879796,14.076719,15.14995,17.946259,20.617847,23.115488,24.49395,24.576002,23.945848,23.289438,22.882463,21.861746,20.266668,19.029335,16.521847,14.332719,13.144616,12.258463,9.573745,7.397744,5.6320004,4.821334,4.604718,3.692308,3.7382567,3.8301542,3.2722054,2.5895386,3.5249233,3.8367183,3.6496413,4.5095387,5.609026,3.757949,2.2088206,1.5589745,1.4408206,1.8642052,3.2295387,3.5380516,6.4000006,10.8537445,15.547078,18.747078,21.26113,19.843283,18.78318,19.186872,18.976822,22.170258,22.235899,21.257847,20.67036,21.270975,23.686565,26.374567,29.341541,32.298668,34.668312,34.1399,32.84677,32.042667,32.531696,34.68472,34.195694,33.857643,32.039387,29.604105,29.909336,29.2759,28.058258,27.073643,26.656822,26.66995,27.208208,27.017849,26.916105,26.87672,26.029951,26.95877,27.582361,28.20267,28.954258,29.797747,28.45867,26.738874,25.491693,25.288208,26.384413,26.41067,25.521233,24.976412,25.380104,26.673233,26.886566,27.014566,26.50913,24.91077,21.871592,18.999796,15.409232,13.121642,12.491488,12.242052,13.400617,15.465027,18.881643,23.348515,27.831797,30.191591,28.99036,25.521233,21.494156,19.049026,17.624617,14.920206,13.846975,14.818462,15.783386,17.893745,19.889233,20.299488,19.34113,18.901335,17.588514,17.660719,19.40677,22.311386,25.048616,25.892105,24.549746,21.7239,17.427694,11.004719,8.379078,5.8847184,5.5269747,6.160411,3.4789746,3.8367183,4.135385,4.066462,5.208616,11.0145645,14.897232,13.679591,12.051693,11.411694,9.875693,8.152616,8.493949,9.419488,9.905231,9.380103,12.301129,13.6697445,10.837335,7.27959,12.563693,21.280823,21.612309,14.562463,5.874872,6.012718,6.1472826,8.280616,9.964309,9.531077,6.0947695,11.23118,13.4859495,10.561642,4.6211286,2.3138463,11.529847,9.212719,6.1472826,5.661539,3.620103,2.6322052,2.028308,1.8838975,1.9265642,1.5130258,1.4703591,1.7427694,2.2580514,2.550154,1.7788719,0.86646163,0.52512825,0.5021539,0.76800007,1.5392822,5.0576415,5.2315903,3.3411283,2.3072822,6.692103,5.0182567,7.0465646,7.7259493,6.616616,7.90318,13.026463,13.650052,12.314258,10.571488,8.992821,7.6931286,6.2523084,5.093744,4.9394875,6.7905645,8.487385,6.8660517,4.2272825,2.231795,1.9068719,1.9265642,2.8849232,5.037949,7.030154,5.874872,7.9950776,8.687591,7.273026,4.4996924,2.5337439,0.9321026,0.60389745,0.9419488,1.3620514,1.3161026,0.4135385,0.09189744,0.02297436,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.02297436,0.01969231,0.029538464,0.049230773,0.06564103,0.055794876,0.32164106,0.54482055,0.8533334,1.7887181,2.9472823,2.353231,1.7755898,1.6672822,1.1782565,3.3936412,3.5971284,3.4888208,3.5971284,3.2853336,3.889231,3.2164104,3.370667,3.6890259,0.74830776,0.2100513,0.07876924,0.101743594,0.18379489,0.37415388,0.42338464,0.39712822,0.4266667,0.47917953,0.36758977,0.2986667,0.32164106,0.35446155,0.35446155,0.3314872,0.35774362,0.3314872,0.30851284,0.29210258,0.23630771,0.20676924,0.23958977,0.35446155,0.5546667,0.8369231,0.761436,0.8369231,0.92553854,1.024,1.2438976,1.6082052,2.156308,2.4024618,2.3794873,2.6289232,2.6453335,3.4494362,5.1364107,7.1056414,8.083693,8.086975,7.6931286,7.6635904,7.752206,6.685539,6.23918,5.83877,5.7468724,5.989744,6.3573337,7.00718,7.1154876,7.250052,7.328821,6.6067696,6.6034875,6.2227697,5.979898,6.055385,6.2916927,6.170257,6.0225644,5.943795,5.937231,5.927385,5.4416413,4.644103,3.5938463,2.5632823,2.03159,1.8281027,2.1497438,2.3368206,2.2777438,2.428718,2.0184617,1.4867693,1.1093334,1.0699488,1.4539489,1.7624617,1.7723079,1.7624617,1.8707694,2.1070771,2.1924105,1.8543591,1.6672822,1.8182565,2.100513,2.8849232,4.2141542,5.799385,6.747898,5.5762057,5.5958977,5.874872,7.1844106,8.484103,6.8955903,3.6693337,2.4943593,2.15959,2.2547693,3.1737437,2.8816411,3.4822567,4.1124105,4.457026,4.772103,3.3608208,2.6945643,3.1442053,3.751385,2.2153847,1.9167181,2.097231,2.1792822,1.8576412,1.0994873,1.1323078,1.1060513,1.1126155,1.1782565,1.273436,1.1126155,1.1782565,1.1881026,1.0404103,0.8172308,1.1585642,1.2242053,1.1946667,1.1618463,1.142154,1.1979488,1.2603078,1.4408206,1.6377437,1.5392822,1.9364104,2.2678976,2.487795,2.4582565,1.9593848,2.3729234,2.5993848,2.681436,2.6354873,2.4418464,2.477949,2.412308,2.2088206,1.9429746,1.8018463,1.9035898,1.8543591,2.0151796,2.294154,2.1464617,2.6322052,3.0293336,3.0916924,2.8422565,2.5665643,2.3860514,3.18359,4.2962055,5.2512827,5.7698464,6.889026,8.621949,10.236719,11.513436,12.724514,13.590976,14.969437,16.423386,17.631182,18.422155,19.72513,20.17477,20.86072,21.979898,22.82995,25.163488,25.698463,25.577028,25.557335,26.020105,26.932514,27.907284,28.603079,28.553848,27.172104,26.66995,26.811079,26.450054,24.94031,22.137438,21.211899,21.471182,21.43836,21.13313,22.081642,22.65272,22.705233,22.961233,23.299284,22.774155,21.897848,22.226053,23.250053,24.356104,24.838566,24.001642,23.066257,22.836515,23.424002,24.234669,25.10113,25.216002,25.481848,26.180925,26.95877,25.409643,22.872618,20.04349,17.893745,17.673847,17.532719,15.78995,14.043899,12.570257,10.328616,9.488411,10.174359,10.584617,10.28595,10.236719,8.740103,7.8670774,7.8112826,8.490667,9.567181,8.979693,8.146052,7.4699492,7.381334,8.326565,8.992821,9.232411,9.921641,11.136001,12.156719,11.9860525,11.500309,11.605334,12.438975,13.364513,13.033027,12.301129,11.749744,11.602052,11.739899,11.776001,12.097642,12.114052,11.680821,11.109744,10.774975,9.701744,8.946873,8.763078,8.618668,8.4283085,8.251078,8.149334,7.962257,7.2992826,6.370462,5.504,4.667077,3.9680004,3.6627696,3.5347695,3.367385,3.190154,3.117949,3.314872,3.5807183,3.5872824,3.5971284,3.5938463,3.308308,2.2121027,2.1136413,2.1989746,2.4385643,2.6912823,2.7175386,2.7044106,2.737231,2.665026,2.4943593,2.3958976,2.1891284,2.2186668,2.1530259,2.041436,2.3335385,2.4320002,2.4746668,2.858667,3.5872824,4.2568207,5.2447186,6.1440005,6.99077,7.896616,9.032206,8.960001,9.344001,9.521232,9.084719,7.890052,8.779488,8.89436,8.41518,8.579283,11.641437,10.9226675,7.13518,3.889231,2.5009232,1.9987694,1.2898463,1.5163078,2.6518977,3.636513,2.3794873,1.6836925,1.4112822,1.3554872,1.3817437,1.4178462,1.332513,1.1191796,0.892718,0.7515898,0.761436,0.9944616,1.0896411,1.0043077,0.8336411,0.80738467,0.9911796,0.88287187,0.88287187,1.0568206,1.1290257,0.88615394,0.5874872,0.4397949,0.5218462,0.7778462,1.1191796,1.3686155,1.5360001,1.6049232,1.5556924,1.3259488,0.9911796,0.6071795,0.30851284,0.32164106,0.24615386,0.18379489,0.19692309,0.22646156,0.09189744,0.04266667,0.029538464,0.04266667,0.07876924,0.15097436,0.4955898,0.75487185,0.9682052,1.2504616,1.8018463,2.5928206,3.3509746,4.1813335,5.10359,6.042257,6.5444107,7.4732313,8.516924,9.429334,10.039796,10.834052,11.894155,12.983796,13.892924,14.404924,13.892924,13.590976,16.114874,21.146257,25.40636,29.67631,31.51426,29.958567,26.400822,24.582565,22.567387,22.41313,22.265438,21.582771,21.11672,19.275488,17.880617,17.220924,16.617027,14.418053,10.525539,7.427283,5.3103595,3.9975388,2.9604106,2.5928206,2.2908719,2.0709746,2.5731285,5.0510774,4.8049235,4.2502565,4.9788723,6.9087186,8.300308,4.5029745,2.5764105,1.9790771,2.1070771,2.28759,2.8127182,6.1768208,10.883283,14.841437,15.366566,18.369642,17.637745,16.384,16.118155,16.633438,16.682669,19.045746,21.815796,23.506054,23.04,23.735796,25.403078,27.904001,30.5559,32.105026,31.51754,29.633644,30.165335,33.539284,36.896824,36.785233,34.727386,32.180515,30.129232,29.06913,26.968618,26.755283,27.00472,26.755283,25.498259,24.825438,25.334156,26.14154,26.86031,27.618464,27.32636,26.820925,26.338463,26.22031,26.916105,25.941336,25.055182,24.769644,25.00595,25.11754,25.189745,25.38995,25.330873,24.77949,23.683285,24.20513,25.895386,26.729027,26.023386,24.398771,20.33231,16.800821,14.381949,13.266052,13.22995,13.899488,15.212309,17.690258,21.376001,25.816618,26.049643,26.666668,25.45231,22.54113,20.417643,17.339079,14.145642,13.380924,14.989129,16.295385,19.666052,20.854155,19.984411,17.99877,16.692514,13.154463,13.833847,16.213335,18.970259,21.973335,25.353848,27.158976,24.425028,17.545847,10.28595,8.979693,6.554257,6.3540516,7.00718,2.4418464,3.3444104,3.7448208,3.9942567,5.9963083,13.197129,15.090873,15.461744,15.638975,15.002257,10.985026,12.681848,9.737847,8.188719,9.15036,8.818872,11.211488,11.628308,9.344001,8.707283,19.11795,23.893335,21.769848,16.315079,10.857026,8.513641,11.493745,10.607591,9.258667,8.155898,5.32677,11.477334,13.298873,10.266257,4.71959,1.8609232,6.340924,8.41518,7.565129,5.7796926,7.5388722,4.3651285,2.4352822,1.8182565,1.9035898,1.404718,2.550154,2.5731285,2.6289232,2.9144619,2.6715899,0.9353847,0.38400003,0.36102566,0.46276927,0.5481026,4.322462,6.764308,5.179077,3.9942567,14.785643,6.803693,5.146257,5.07077,5.681231,9.91836,14.434463,14.263796,13.46954,12.996924,10.666668,12.179693,12.274873,10.686359,8.254359,6.9120007,4.604718,6.2162056,6.1078978,3.370667,1.847795,1.211077,7.276308,11.995898,12.173129,9.475283,8.109949,7.2992826,6.196513,4.522667,2.5928206,1.1782565,0.78769237,0.90912825,0.98461545,0.4135385,0.14441027,0.03938462,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01969231,0.029538464,0.029538464,0.029538464,0.029538464,0.15097436,0.2297436,0.27569234,0.4594872,1.276718,2.0020514,2.550154,2.6551797,1.8609232,1.7526156,2.540308,2.8553848,2.4549747,2.1989746,2.0512822,2.28759,2.4484105,2.4188719,2.4549747,0.5513847,0.059076928,0.052512825,0.108307704,0.28882053,0.47261542,0.49230772,0.44307697,0.4135385,0.48902568,0.34133336,0.29538465,0.30851284,0.32164106,0.25928208,0.28225642,0.28225642,0.26912823,0.25928208,0.25928208,0.25928208,0.21333335,0.27569234,0.50543594,0.88615394,0.5677949,0.50543594,0.65969235,0.96492314,1.3423591,1.7952822,2.3204105,2.5009232,2.4188719,2.6387694,3.3608208,4.1091285,5.2545643,6.633026,7.522462,7.7292314,7.525744,7.8014364,8.3593855,7.9195905,6.2227697,6.2555904,6.75118,6.954667,6.636308,7.785026,8.356103,8.470975,8.04759,6.7905645,7.02359,6.7774363,6.491898,6.340924,6.2555904,6.232616,5.786257,5.333334,4.890257,4.059898,3.9253337,3.5905645,3.2032824,2.8389745,2.4713848,2.2777438,2.1530259,1.9364104,1.6968206,1.7690258,1.9167181,1.4867693,1.1881026,1.2832822,1.5885129,1.9659488,1.719795,1.8871796,2.422154,2.228513,2.166154,1.8937438,1.847795,2.100513,2.3794873,3.0391798,4.3684106,6.1308722,7.125334,5.172513,5.7698464,6.3967185,6.701949,6.4065647,5.293949,3.18359,3.0851285,3.1409233,2.917744,3.4166157,3.9548721,4.023795,3.895795,3.8564105,4.210872,3.5511796,2.9111798,2.5764105,2.5698464,2.6551797,2.2383592,1.9364104,1.8543591,1.8806155,1.6475899,1.1848207,1.1126155,1.211077,1.3226668,1.3587693,1.1388719,1.0666667,1.1126155,1.1585642,0.97805136,1.3686155,1.2537436,0.97805136,0.85005134,1.1290257,1.5064616,1.8871796,2.0086155,1.9035898,1.8904617,2.0742567,1.9298463,1.8806155,2.0578463,2.28759,2.9472823,2.802872,2.3368206,2.0873847,2.6256413,2.6617439,2.5140514,2.2350771,1.8740515,1.4966155,1.5195899,1.8182565,2.1103592,2.3040001,2.487795,3.121231,3.436308,3.1606157,2.5173335,2.2121027,2.5796926,3.6594875,4.850872,5.9667697,7.24677,8.152616,9.557334,11.460924,13.056001,12.724514,12.800001,15.087591,17.096207,17.811693,17.716515,19.193438,20.036924,20.837746,21.842052,22.964514,24.612104,25.783796,26.548515,26.752003,26.029951,27.030977,27.749746,27.00472,24.98954,23.253336,22.20636,21.989746,22.06195,22.029129,21.638565,20.28308,19.941746,20.066463,20.115694,19.593847,20.630976,21.18236,21.700924,22.153849,22.019283,21.93395,22.452515,23.824411,25.32759,25.252104,23.361643,22.593643,23.089233,24.369232,25.344002,25.72472,25.892105,26.325335,26.90954,26.945642,25.055182,22.521437,19.951591,18.235079,18.54031,17.683693,16.07877,14.358975,12.635899,10.499283,9.67877,10.692924,11.657847,11.651283,10.712616,8.845129,7.762052,7.8441033,8.763078,9.504821,8.822155,7.6996927,7.24677,7.762052,8.726975,8.851693,9.019077,9.744411,10.896411,11.703795,11.546257,11.149129,11.08677,11.569232,12.435693,12.435693,12.1238985,11.904001,11.851488,11.703795,11.936821,12.304411,12.409437,12.1698475,11.841642,11.096616,9.856001,8.805744,8.3364105,8.546462,8.129642,7.8145647,7.5520005,7.250052,6.774154,6.1407185,5.330052,4.5062566,3.8695388,3.6627696,3.515077,3.4527183,3.383795,3.314872,3.3280003,3.6791797,3.9154875,3.9023592,3.6758976,3.4166157,2.1136413,2.162872,2.0512822,2.103795,2.3466668,2.5074873,2.612513,2.4943593,2.3663592,2.2777438,2.103795,2.1103592,2.2153847,2.281026,2.2482052,2.1398976,2.3433847,2.4713848,2.802872,3.3542566,3.879385,4.896821,5.737026,6.692103,7.8145647,8.910769,9.002667,9.7673855,9.796924,8.769642,7.4371285,7.509334,7.0498466,7.138462,8.766359,12.826258,12.790154,8.113232,3.7251284,1.7755898,1.6082052,1.8773335,2.294154,2.6387694,2.5600002,1.5885129,1.2340513,1.2635899,1.3456411,1.2635899,0.9189744,0.892718,0.955077,0.9747693,0.98133343,1.1782565,1.3423591,1.3226668,1.2077949,1.0732309,0.97805136,0.93866676,0.8008206,0.7811283,0.86974365,0.8369231,0.69907695,0.6170257,0.6071795,0.6826667,0.85005134,1.0568206,1.1913847,1.2800001,1.3161026,1.2865642,1.017436,0.7122052,0.51856416,0.47917953,0.5415385,0.52512825,0.571077,0.49887183,0.32164106,0.22646156,0.15753847,0.2297436,0.33805132,0.47261542,0.702359,0.88615394,1.014154,1.1224617,1.332513,1.8116925,2.5764105,3.3476925,4.1189747,4.8771286,5.602462,5.9963083,6.7249236,7.686565,8.736821,9.6984625,10.706052,12.609642,14.985847,16.994463,17.371899,16.17395,15.451899,16.758156,20.178053,24.320002,25.51467,25.347284,23.824411,21.737028,20.65067,21.097027,21.842052,21.559797,20.050053,18.248207,16.951796,16.31836,16.328207,16.15754,14.17518,10.535385,7.4863596,5.353026,4.0467696,3.058872,2.878359,3.4724104,3.383795,3.0916924,5.0018463,5.0215387,4.57518,4.0434875,6.0356927,15.40595,12.370052,9.314463,5.5893335,2.3729234,2.6551797,3.2886157,5.87159,9.4457445,12.324103,12.107488,14.611693,14.148924,14.339283,16.039387,17.352207,17.509745,19.70872,21.730463,22.478771,22.016,22.439386,23.719387,26.226873,29.029745,29.906054,29.193848,29.758362,31.849028,35.53149,40.704002,39.94913,36.804924,33.40144,31.366566,31.839182,27.93354,27.26072,27.930258,28.255182,26.742155,25.494976,24.352823,24.562874,26.10872,27.703796,27.0999,26.561644,26.049643,25.767387,26.161232,25.924925,25.760822,25.51795,25.048616,24.201847,25.153643,25.734566,25.360413,24.119797,22.777437,23.204103,24.618668,25.714874,25.770668,24.654772,21.392412,18.116924,15.563488,14.168616,14.083283,14.76595,15.954053,18.136618,21.195488,24.425028,25.429335,26.729027,26.522259,24.608822,22.406567,19.272207,15.908104,14.562463,15.563488,17.30954,20.923079,21.691078,20.476719,18.176,15.717745,13.328411,12.803283,13.689437,15.75713,18.993233,25.59672,29.302156,26.197336,17.952822,11.82195,7.6274877,4.926359,3.9384618,3.764513,2.3926156,2.993231,3.5380516,3.8564105,5.2545643,10.512411,15.960617,16.758156,15.714462,13.968411,10.985026,12.097642,8.828718,6.810257,7.8080006,9.7214365,10.962052,9.353847,6.3967185,4.7425647,8.182155,13.98154,17.946259,18.986668,17.650873,16.118155,11.382154,12.481642,12.189539,8.182155,3.006359,9.6065645,11.382154,9.196308,5.2611284,3.117949,4.4045134,11.017847,12.973949,9.321027,8.149334,4.57518,2.2678976,1.3522053,1.9396925,4.1124105,3.249231,2.6584618,2.3072822,2.2219489,2.487795,1.5753847,1.0010257,0.56451285,0.3314872,0.6235898,1.7493335,7.748924,7.640616,2.3794873,4.850872,3.4100516,2.737231,2.1497438,2.166154,4.4865646,7.4699492,10.056206,12.882052,15.258258,15.182771,14.78236,10.295795,10.86359,15.415796,12.685129,7.821129,5.297231,3.8695388,2.7700515,1.7132308,1.017436,5.796103,7.653744,5.87159,7.4141545,4.824616,3.9975388,4.4800005,4.585026,1.3981539,1.1913847,0.77456415,0.45292312,0.28882053,0.108307704,0.032820515,0.006564103,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.0032820515,0.009846155,0.032820515,0.049230773,0.029538464,0.068923086,0.13128206,0.19692309,0.2855385,0.46933338,1.0633847,1.6672822,1.8445129,1.8051283,2.3991797,2.044718,2.806154,2.8422565,1.8871796,1.270154,1.5524104,1.9790771,2.477949,2.6945643,1.9692309,0.48246157,0.06564103,0.03938462,0.06564103,0.13128206,0.3446154,0.3708718,0.3052308,0.27241027,0.40369233,0.33476925,0.27897438,0.29210258,0.33476925,0.28225642,0.21989745,0.24615386,0.26256412,0.24943592,0.25928208,0.33805132,0.3117949,0.2855385,0.32164106,0.446359,0.4397949,0.5152821,0.65312827,0.8467693,1.0994873,1.5491283,2.1333334,2.5173335,2.678154,2.9078977,3.4921029,4.33559,5.3136415,6.373744,7.5585647,8.185436,8.139488,7.9097443,7.719385,7.50277,6.51159,6.3310776,6.629744,6.9021544,6.4656415,7.000616,7.680001,8.195283,8.132924,6.9743595,6.4722056,6.308103,6.3442054,6.4065647,6.2916927,6.2194877,5.9536414,5.58277,5.0642056,4.204308,4.1189747,3.7809234,3.3345644,2.92759,2.7175386,2.2383592,1.913436,1.654154,1.463795,1.4276924,1.4572309,1.2471796,1.2504616,1.4441026,1.3292309,2.1300514,1.7558975,1.5064616,1.8149745,2.2646155,2.349949,2.2088206,2.0250258,2.1169233,2.9538465,3.5052311,4.6539493,6.3573337,7.50277,5.8912826,6.1505647,6.1538467,6.1997952,6.0356927,4.8672824,3.6430771,3.308308,3.367385,3.564308,3.8695388,4.3684106,3.9154875,3.1048207,2.540308,2.8455386,3.2984617,2.8914874,2.284308,1.8806155,1.847795,1.5622566,1.4933335,1.5786668,1.7394873,1.8674873,1.4900514,1.3554872,1.273436,1.1881026,1.1881026,1.2012309,1.1060513,0.99774367,0.9288206,0.892718,0.97805136,1.1552821,1.3259488,1.4309745,1.4572309,1.5360001,1.5655385,1.7132308,1.9331284,1.9889232,1.8904617,1.8707694,2.0906668,2.4320002,2.4976413,2.6486156,2.4681027,2.3171284,2.3860514,2.6978464,2.3729234,1.9692309,1.7591796,1.7591796,1.7033848,2.1267693,2.284308,2.3860514,2.5895386,2.986667,3.0752823,2.9965131,2.5895386,2.1234872,2.284308,3.5216413,4.6276927,5.661539,6.75118,8.090257,8.152616,9.357129,10.998155,12.527591,13.5548725,14.713437,16.072206,16.758156,16.955078,17.923283,19.242668,20.473438,20.992002,21.093744,22.01272,22.656002,24.270771,25.888823,26.624002,25.688618,25.626259,25.859283,25.3079,24.116514,23.634052,22.65272,21.894566,21.054361,20.164925,19.59713,19.738258,19.544617,19.666052,19.945026,19.419899,18.612514,19.209848,20.105848,20.575182,20.28636,20.932924,21.96349,23.96554,25.967592,25.422771,23.289438,22.452515,22.885746,24.1559,25.455591,25.403078,25.728003,26.194054,26.53867,26.4599,24.457848,22.199797,20.480001,19.74154,20.07631,17.572104,15.504412,13.636924,11.884309,10.315488,10.200616,10.929232,11.529847,11.303386,9.796924,8.231385,7.755488,8.12636,8.986258,9.849437,8.480822,7.3025646,7.1122055,7.9786673,9.265231,9.846154,9.980719,10.338462,10.8537445,10.752001,10.397539,10.010257,10.174359,10.834052,11.300103,11.339488,11.0605135,10.801231,10.827488,11.32636,11.625027,12.114052,12.373334,12.278154,11.9860525,10.459898,8.851693,7.9195905,7.716103,7.581539,7.3616414,7.1089234,6.8660517,6.5936418,6.1768208,5.346462,4.5554876,3.895795,3.5216413,3.626667,3.6069746,3.5807183,3.5052311,3.4133337,3.4231799,3.757949,4.017231,3.9286156,3.5610259,3.3444104,2.0644104,2.0841026,2.0086155,2.038154,2.2547693,2.6387694,2.8192823,2.6322052,2.540308,2.5665643,2.3040001,2.3663592,2.225231,2.1891284,2.2744617,2.2383592,2.4484105,2.5074873,2.7044106,3.1442053,3.757949,4.7294364,5.674667,6.7216415,7.824411,8.743385,9.252103,9.708308,9.45559,8.493949,7.4699492,6.7216415,5.9995904,6.163693,7.4929237,9.672206,9.7673855,7.4240007,4.7294364,2.8750772,2.15959,2.681436,2.4681027,2.0184617,1.5688206,1.1060513,1.0469744,1.1257436,1.0962052,0.92553854,0.79425645,0.8041026,0.90584624,0.9944616,1.083077,1.2832822,1.4276924,1.332513,1.2077949,1.1388719,1.086359,1.0633847,0.99774367,0.9911796,1.0404103,1.0469744,1.017436,0.9944616,0.9156924,0.82379496,0.8598975,0.9714873,1.020718,1.0338463,1.017436,0.955077,0.77128214,0.57764107,0.47261542,0.52512825,0.7515898,0.67610264,0.65641034,0.574359,0.446359,0.40697438,0.60389745,0.8467693,0.97805136,1.014154,1.1224617,1.1585642,1.1585642,1.2800001,1.6180514,2.1924105,3.0129232,3.7185643,4.4110775,5.1922054,6.1341543,7.1581545,7.968821,8.87795,10.056206,11.516719,12.960821,15.120412,17.122463,18.264616,18.021746,16.505438,14.769232,14.621539,16.521847,19.590565,20.975592,21.12,20.519386,19.51836,18.313848,18.110361,18.136618,17.34236,15.606155,13.74195,12.642463,11.881026,11.739899,11.703795,10.469745,8.182155,6.380308,5.1200004,4.2207184,3.2754874,2.9144619,3.5905645,3.6102567,3.3936412,5.4941545,5.2348723,4.8114877,3.9286156,4.397949,10.161232,9.481847,10.400822,8.333129,3.9745643,3.2787695,3.8038976,5.4514875,8.182155,11.021129,12.06154,14.578873,14.132514,14.217847,15.796514,17.302977,16.90913,17.634462,19.74154,21.953642,21.43836,21.205336,22.846361,25.042053,27.38872,30.38195,29.551592,30.244104,32.374157,35.731693,39.9918,40.51036,38.87262,37.54339,36.962463,35.51508,30.785643,30.040617,30.802053,31.0679,29.331694,28.242054,26.518976,25.298054,25.110977,25.875694,26.387693,26.318771,26.036514,25.85272,26.052925,26.633848,26.614157,26.427078,26.000412,24.766361,25.206156,25.662361,25.455591,24.356104,22.57067,21.441643,22.449232,23.430567,23.328823,22.193232,20.079592,17.59836,15.724309,14.752822,14.296617,15.186052,16.843489,18.806156,20.903387,23.253336,25.160208,26.978464,27.523285,26.518976,24.595694,20.81149,17.243898,15.832617,16.7319,18.330257,21.24472,21.638565,20.299488,17.844515,14.729847,12.3536415,11.769437,12.540719,14.5952835,18.22195,25.265232,29.377644,25.255386,15.642258,11.346052,6.1768208,5.6385646,4.6900516,2.7569232,3.7448208,3.4494362,3.7973337,3.9417439,4.4964104,7.53559,15.688207,18.067694,16.482462,12.980514,9.869129,12.416001,10.266257,7.4010262,6.1538467,7.210667,7.8047185,7.000616,5.5007186,4.2601027,4.4767184,8.195283,12.186257,15.346873,16.879591,16.282257,8.516924,8.979693,10.948924,9.616411,2.0611284,6.1013336,9.803488,11.109744,9.954462,8.267488,5.622154,11.139283,13.121642,9.8592825,9.645949,5.0642056,2.4024618,1.4506668,2.789744,7.8014364,4.1058464,2.7306669,2.2777438,2.1136413,2.349949,1.9856411,1.2274873,0.6268718,0.48574364,0.8795898,1.6213335,9.6295395,9.665642,2.3630772,4.240411,2.934154,1.9200002,1.1454359,0.86646163,1.6180514,4.0500517,6.0816417,9.370257,13.105232,13.994668,15.606155,11.592206,9.3768215,10.765129,11.959796,7.9261546,5.179077,5.72718,7.312411,3.3903592,3.1573336,5.156103,5.5269747,4.1025643,4.4242053,2.6387694,2.4648206,3.314872,3.879385,2.1333334,2.5961027,4.197744,3.5216413,0.83035904,0.059076928,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.009846155,0.01969231,0.032820515,0.04266667,0.03938462,0.052512825,0.14112821,0.20676924,0.26912823,0.48246157,0.65312827,0.8402052,1.0699488,1.3915899,1.8543591,1.6607181,2.4713848,2.5993848,1.8051283,1.2931283,1.1355898,1.5195899,2.3991797,3.1967182,2.806154,0.86317956,0.16410258,0.026256412,0.04266667,0.06564103,0.19692309,0.24943592,0.26912823,0.27569234,0.2986667,0.24943592,0.25271797,0.26584616,0.2855385,0.35446155,0.3117949,0.29538465,0.30194873,0.3117949,0.29538465,0.35774362,0.35446155,0.32820517,0.318359,0.3708718,0.41025645,0.5481026,0.7417436,0.9156924,0.9747693,1.394872,1.9823592,2.3072822,2.4188719,2.809436,3.3608208,4.201026,5.32677,6.6034875,7.788308,8.103385,8.214975,7.893334,7.4010262,7.4929237,6.747898,6.5444107,6.7544622,7.0137444,6.7249236,6.8693337,7.128616,7.433847,7.4699492,6.672411,6.521436,6.7216415,6.8233852,6.6494365,6.301539,6.2030773,6.117744,5.9930263,5.651693,4.8016415,4.2371287,3.8531284,3.308308,2.6978464,2.556718,1.9495386,1.5327181,1.3489232,1.3587693,1.4539489,1.3718976,1.2077949,1.2307693,1.3915899,1.3029745,1.7362052,1.6147693,1.3981539,1.4769232,2.1825643,2.3040001,2.3072822,2.2383592,2.356513,3.1442053,3.7940516,4.6178465,5.5171285,6.0619493,5.4974365,5.4908724,5.605744,5.7009234,5.5138464,4.6605134,4.5095387,3.8465643,3.5938463,3.895795,4.138667,4.2601027,3.4658465,2.7437952,2.5435898,2.7766156,3.318154,2.9243078,2.3302567,2.0086155,2.15959,2.1530259,1.9922053,1.7657437,1.6049232,1.6836925,1.5491283,1.4080001,1.3489232,1.394872,1.4998976,1.5392822,1.2570257,0.9747693,0.8336411,0.8041026,0.8992821,1.0633847,1.2537436,1.467077,1.7624617,1.9528207,1.8576412,1.7985642,1.8904617,2.0151796,1.7558975,1.7690258,2.0611284,2.422154,2.412308,2.5173335,2.481231,2.4484105,2.484513,2.5895386,2.100513,1.595077,1.332513,1.4145643,1.782154,2.2055387,2.3335385,2.6453335,3.2623591,3.9647183,2.9997952,2.4615386,2.2219489,2.2514873,2.6322052,4.2929235,5.605744,6.560821,7.282872,8.044309,8.372514,9.521232,10.952206,12.363488,13.673027,14.79877,14.976001,15.16636,16.026258,17.910154,19.383797,20.81149,21.48431,21.67795,22.662565,22.495182,23.2599,24.474258,25.432617,25.22913,24.782772,24.385643,23.94913,23.519182,23.2599,22.199797,20.814772,19.367386,18.185848,17.641027,18.770052,18.894772,18.274464,17.545847,17.729643,17.033848,17.339079,18.212105,19.029335,18.953848,20.266668,21.851898,23.811283,25.284925,24.441439,22.396719,21.99631,22.44595,23.440413,25.170053,24.996105,25.314463,25.714874,25.75426,24.917336,23.220514,21.62872,21.02154,21.080618,20.289642,16.902565,14.562463,12.859077,11.546257,10.535385,10.850462,11.017847,10.965334,10.427077,8.92718,7.860513,7.958975,8.664616,9.43918,9.760821,7.8047185,6.954667,7.259898,8.3823595,9.619693,10.102155,10.325335,10.545232,10.617436,10.010257,9.885539,10.148104,10.676514,11.050668,10.522257,10.35159,9.938052,9.69518,9.8592825,10.499283,10.7848215,11.264001,11.493745,11.32636,10.906258,9.685334,8.507077,7.634052,7.1581545,7.020308,6.7249236,6.6100516,6.308103,5.7731285,5.3136415,4.6178465,4.3585644,4.013949,3.6791797,4.073026,4.2929235,4.2568207,4.007385,3.7218463,3.7054362,4.027077,4.2469745,4.069744,3.6430771,3.5380516,2.0512822,1.9954873,1.9856411,2.0775387,2.2711797,2.5042052,2.858667,2.7963078,2.7044106,2.6387694,2.3335385,2.4943593,2.300718,2.2219489,2.3302567,2.3401027,2.477949,2.5009232,2.6551797,3.0523078,3.6824617,4.5029745,5.605744,6.747898,7.8014364,8.766359,9.682052,9.77395,9.485129,8.914052,7.8112826,6.885744,6.370462,6.314667,6.6067696,6.9809237,9.760821,10.988309,9.242257,5.398975,2.6354873,2.4057438,1.8412309,1.2898463,0.9353847,0.78769237,0.84348726,0.88615394,0.80738467,0.65969235,0.6662565,0.7450257,0.8795898,1.0305642,1.1684103,1.2832822,1.3850257,1.2373334,1.1257436,1.148718,1.2077949,1.3095386,1.3259488,1.2471796,1.1355898,1.1027694,1.1618463,1.1323078,1.020718,0.90256417,0.9353847,0.9878975,0.96492314,0.9288206,0.8960001,0.8402052,0.65312827,0.5481026,0.5415385,0.6432821,0.8533334,0.8008206,0.7089231,0.5907693,0.46933338,0.39384618,0.702359,1.0666667,1.3062565,1.3554872,1.2406155,1.1585642,1.1126155,1.273436,1.6968206,2.3204105,3.318154,4.1813335,4.962462,5.786257,6.8529234,8.425026,9.4916935,10.463181,11.523283,12.652308,13.899488,15.9573345,17.572104,17.867489,16.347898,14.6871805,13.141335,13.062565,14.785643,17.624617,18.924309,19.314873,19.091694,18.372925,17.079796,16.328207,15.665232,14.946463,14.066873,12.973949,11.9171295,10.515693,9.590155,9.235693,8.805744,7.0137444,5.917539,5.1922054,4.565334,3.82359,3.3247182,3.9056413,4.023795,3.892513,5.4580517,4.923077,4.519385,3.7284105,3.1737437,4.598154,4.9985647,8.116513,8.6580515,6.0192823,4.2830772,4.5029745,6.091488,8.1066675,10.082462,12.005745,14.185027,14.027489,14.362258,15.96718,17.595078,18.343386,19.90236,21.888002,23.236925,22.219488,21.13313,22.770874,24.42831,25.849438,29.243078,29.607388,30.280207,32.128002,35.150772,38.501747,40.310158,40.60226,41.16021,41.67549,39.732517,35.53477,33.94954,33.732925,33.572105,32.085335,30.454157,28.85908,27.313232,25.91508,24.832003,25.800207,26.04308,25.783796,25.823181,27.549541,28.711388,28.517746,28.035284,27.3559,25.586874,25.449028,25.59672,25.527798,24.644924,22.235899,20.696617,20.512821,20.352001,19.682463,18.793028,17.076513,15.760411,14.9628725,14.592001,14.372104,16.09518,18.06113,19.606976,20.722874,22.065233,24.838566,27.109745,28.09108,27.385439,25.00595,21.303797,18.481232,17.217642,17.621334,19.242668,21.014977,21.031385,19.459284,16.656412,13.161027,10.81436,10.587898,11.474052,13.364513,17.063385,23.640617,28.20267,24.01149,13.705847,9.3078985,7.003898,6.2884107,4.565334,2.609231,4.568616,3.4724104,4.06318,4.4865646,4.7556925,6.7544622,15.248411,18.087385,17.155283,13.709129,8.39877,12.642463,11.293539,7.5520005,4.4077954,4.634257,4.84759,5.661539,5.756718,4.850872,3.69559,5.0904617,7.2205133,9.616411,11.35918,11.08677,7.259898,7.6176414,11.474052,13.558155,4.023795,4.0434875,7.6570263,11.736616,14.17518,13.889642,11.313231,14.230975,13.364513,9.061745,11.283693,6.6034875,3.2525132,1.8937438,3.2098465,7.9261546,4.059898,2.7011285,2.3958976,2.4681027,3.0260515,3.1277952,1.8773335,0.9156924,0.8402052,1.214359,1.8445129,7.512616,7.3682055,2.1169233,4.010667,2.477949,1.467077,1.086359,1.8313848,4.588308,3.9253337,3.7743592,5.3136415,8.093539,10.029949,12.73436,13.472821,9.990565,5.2644105,7.506052,5.139693,4.2305646,6.294975,8.786052,5.100308,5.6254363,6.4557953,6.3310776,4.9952826,3.1967182,2.1530259,2.789744,3.5216413,3.3969233,2.0841026,2.6912823,4.2830772,3.5577438,0.85005134,0.118153855,0.029538464,0.006564103,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.013128206,0.01969231,0.02297436,0.026256412,0.03938462,0.052512825,0.20676924,0.2986667,0.33476925,0.53825647,0.44307697,0.3249231,0.58420515,1.0732309,1.0929232,0.9911796,1.6672822,1.972513,1.6410258,1.3128207,1.0010257,1.4080001,2.103795,2.6617439,2.6551797,1.1257436,0.33476925,0.049230773,0.029538464,0.052512825,0.11158975,0.17394873,0.2297436,0.25928208,0.21333335,0.19364104,0.24943592,0.256,0.24287182,0.35446155,0.36758977,0.318359,0.3117949,0.33805132,0.30194873,0.318359,0.34133336,0.3708718,0.4201026,0.50543594,0.446359,0.50543594,0.6629744,0.8336411,0.86317956,1.1881026,1.6804104,1.9495386,2.0578463,2.5042052,3.1474874,4.056616,5.297231,6.6625648,7.6668725,7.7718983,8.100103,7.8473854,7.2237954,7.4863596,7.131898,7.0531287,7.141744,7.1909747,6.872616,6.764308,6.698667,6.678975,6.616616,6.3277955,6.5706673,6.8627696,6.8529234,6.5411286,6.2884107,6.2916927,6.1374364,5.9602056,5.6976414,5.106872,4.0533338,3.5840003,3.1015387,2.5238976,2.2711797,1.7362052,1.3817437,1.214359,1.2012309,1.2438976,1.2242053,1.1881026,1.1979488,1.2603078,1.3161026,1.4080001,1.4572309,1.3620514,1.3456411,1.9626669,2.0545642,2.0873847,2.2219489,2.5928206,3.2951798,4.2141542,4.8672824,5.07077,4.886975,4.6539493,4.4964104,4.716308,4.962462,4.9329233,4.391385,4.6933336,4.013949,3.5905645,3.767795,3.9844105,4.0041027,3.1671798,2.7470772,3.0358977,3.3378465,3.249231,2.4976413,1.9396925,1.9200002,2.2514873,2.6026669,2.5107694,2.0841026,1.591795,1.4834872,1.5589745,1.4244103,1.4276924,1.6114873,1.719795,1.6902566,1.3751796,1.0666667,0.892718,0.82379496,1.020718,1.0732309,1.1585642,1.3915899,1.8149745,2.0118976,2.0184617,2.0086155,2.028308,2.0020514,1.7526156,1.6804104,1.9035898,2.2744617,2.3794873,2.4451284,2.297436,2.1431797,2.0873847,2.1103592,1.7066668,1.3522053,1.1552821,1.2307693,1.6672822,2.0020514,2.2514873,2.6978464,3.3214362,3.7874875,2.6223593,2.0611284,2.034872,2.4385643,3.114667,4.857436,6.2227697,7.062975,7.4830775,7.8506675,8.697436,10.059488,11.490462,12.829539,14.191591,14.611693,14.132514,14.381949,15.973744,18.507488,20.059898,20.975592,21.474463,22.01272,23.289438,22.71836,22.472206,23.026873,23.985233,24.057438,23.561848,22.800411,22.294975,22.09149,21.766565,21.638565,20.420925,18.763489,17.365335,16.978052,17.828104,17.8839,16.850052,15.589745,16.137848,16.38072,16.377438,16.777847,17.532719,17.893745,19.367386,21.35631,23.243488,24.290462,23.64718,21.59918,21.454771,21.920822,22.68554,24.408617,24.648207,24.891079,25.015797,24.687592,23.332104,21.78954,21.080618,21.251284,21.323488,19.268925,15.563488,13.354668,12.150155,11.483898,10.889847,11.21477,10.837335,10.171078,9.321027,8.070564,7.768616,8.402052,9.31118,9.8363085,9.32759,7.213949,6.813539,7.571693,8.858257,9.941334,10.151385,10.571488,10.765129,10.486155,9.6754875,9.954462,10.551796,11.142565,11.260718,10.30236,9.83959,9.380103,9.235693,9.432616,9.718155,9.993847,10.456616,10.394258,9.846154,9.577026,9.133949,8.349539,7.5191803,6.931693,6.8594875,6.422975,6.265436,5.8256416,5.093744,4.588308,3.9056413,3.948308,3.892513,3.7087183,4.1583595,4.4701543,4.4800005,4.2601027,4.0303593,4.1550775,4.394667,4.5029745,4.325744,4.0008206,3.9712822,2.1530259,1.9954873,1.9331284,2.0545642,2.231795,2.1070771,2.5829747,2.7634873,2.6584618,2.3663592,2.0709746,2.3401027,2.356513,2.3762052,2.4320002,2.3302567,2.4516926,2.605949,2.8553848,3.242667,3.7874875,4.348718,5.5105643,6.701949,7.781744,9.048616,10.177642,10.194052,10.075898,9.764103,8.162462,7.640616,7.6734366,7.53559,7.456821,8.628513,16.981335,20.132105,16.229744,7.9425645,2.4648206,1.2438976,0.8763078,0.8008206,0.7220513,0.61374366,0.60061544,0.61374366,0.6104616,0.574359,0.51856416,0.67938465,0.8402052,1.0305642,1.211077,1.2438976,1.2340513,1.079795,1.0305642,1.148718,1.3029745,1.4211283,1.4408206,1.270154,0.9878975,0.8172308,0.92225647,0.9156924,0.8960001,0.92553854,1.0305642,1.0338463,0.9517949,0.88287187,0.86317956,0.8795898,0.65641034,0.60061544,0.6695385,0.7778462,0.80738467,0.84348726,0.7778462,0.6170257,0.41682056,0.28225642,0.4955898,0.8598975,1.2077949,1.3587693,1.1126155,1.017436,1.024,1.2012309,1.5622566,2.0939488,3.1015387,4.201026,5.2053337,6.114462,7.1089234,8.723693,9.954462,11.139283,12.130463,12.3076935,12.885334,14.660924,16.111591,16.032822,13.528616,11.848206,11.739899,13.019898,15.458463,18.756924,18.91118,18.868515,18.376207,17.457232,16.426668,16.278976,15.872002,16.292105,17.444103,18.06113,16.777847,14.742975,12.822975,11.588924,11.296822,8.667898,7.1909747,6.3507695,5.7403083,5.074052,4.706462,5.737026,5.861744,5.0051284,5.3070774,4.5456414,3.9975388,3.2951798,2.6847181,3.0293336,2.8980515,4.6539493,6.38359,6.941539,5.9536414,5.920821,7.4108725,8.687591,9.4916935,11.047385,12.422565,12.937847,14.17518,16.459488,18.888206,22.308104,26.420515,27.687387,25.928207,24.329847,22.419695,23.2599,24.418463,25.127386,26.299078,28.310976,29.75508,31.671797,34.422157,37.687798,40.881233,42.384415,43.103184,43.362465,42.90626,40.956722,38.54113,36.72944,35.70544,34.7799,32.262566,30.697027,29.633644,28.314259,25.672207,25.829746,25.911797,25.583591,26.059488,30.119387,31.573336,31.058054,29.96185,28.583387,26.161232,26.095592,25.957747,25.593437,24.434874,21.507284,20.844309,19.222977,17.444103,16.065641,15.419078,13.627078,13.2562065,13.289026,13.46954,14.309745,17.030565,19.213129,20.608002,21.218464,21.27754,24.44472,26.978464,27.913849,26.735592,23.414156,20.60472,19.239386,18.149744,17.67713,19.666052,20.690052,20.54236,18.60595,15.235283,11.762873,9.642668,9.242257,9.8592825,11.477334,14.775796,21.428514,26.86031,23.706259,13.74195,7.890052,9.737847,6.11118,2.9735386,2.8422565,4.8016415,3.0490258,4.161641,5.0543594,5.3825645,7.5618467,13.955283,16.534975,17.083078,14.992412,7.2631803,12.0549755,10.768411,6.6625648,3.0654361,3.3903592,3.3312824,5.172513,6.058667,5.0477953,3.1113849,3.2984617,4.33559,5.152821,5.21518,4.5522056,7.4141545,8.999385,12.960821,15.82277,6.9743595,4.007385,5.3924108,9.911796,15.028514,16.899282,17.165129,18.031591,13.860104,7.9458466,12.504617,7.719385,4.276513,2.665026,2.9702566,4.896821,3.2918978,2.6551797,2.605949,3.0490258,4.164923,4.450462,2.733949,1.3784616,1.214359,1.5721027,1.8412309,3.7874875,3.7185643,1.7066668,1.5589745,1.1979488,0.85005134,1.2438976,3.7152824,10.233437,6.619898,4.5095387,3.2656412,3.170462,5.435077,7.13518,13.22995,12.06154,4.4734364,3.8071797,2.034872,3.5577438,5.533539,6.245744,5.113436,6.8660517,8.129642,7.7357955,5.7829747,3.629949,3.446154,4.2305646,4.381539,3.242667,1.1191796,2.228513,1.4539489,0.69907695,0.6268718,0.636718,0.3511795,0.26584616,0.18051283,0.059076928,0.02297436,0.006564103,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.013128206,0.016410258,0.01969231,0.029538464,0.06564103,0.23630771,0.3511795,0.40369233,0.5874872,0.4594872,0.29538465,0.4660513,0.8041026,0.60061544,0.45620516,0.7811283,1.1782565,1.3620514,1.1257436,1.1355898,1.6607181,1.7624617,1.401436,1.4342566,1.1848207,0.6465641,0.20348719,0.026256412,0.052512825,0.09189744,0.13456412,0.16082053,0.16738462,0.15425642,0.18051283,0.24287182,0.256,0.2297436,0.28882053,0.3314872,0.30194873,0.29210258,0.3117949,0.28225642,0.30194873,0.34789747,0.4266667,0.5284103,0.65312827,0.48246157,0.39712822,0.4397949,0.58092314,0.7220513,0.9321026,1.3062565,1.585231,1.7657437,2.097231,2.8521028,3.8596926,5.110154,6.3442054,7.072821,7.387898,8.090257,7.9819493,7.210667,7.2631803,7.325539,7.509334,7.6242056,7.4830775,6.9054365,6.616616,6.5247183,6.3343596,6.1078978,6.2720003,6.550975,6.5903597,6.413129,6.2129235,6.3277955,6.439385,5.986462,5.4908724,5.172513,4.9362054,3.7448208,3.1803079,2.8160002,2.4385643,2.0545642,1.7394873,1.5195899,1.273436,0.9911796,0.8008206,0.9682052,1.1224617,1.1782565,1.1782565,1.3062565,1.2931283,1.2832822,1.2373334,1.270154,1.6278975,1.6771283,1.7165129,2.0841026,2.7864618,3.515077,4.713026,5.2414365,5.10359,4.5489235,4.086154,3.9942567,3.9417439,4.2371287,4.6080003,4.20759,4.073026,3.7448208,3.5052311,3.4724104,3.623385,3.7842054,3.1376412,2.9768207,3.4855387,3.751385,2.7963078,1.6836925,1.1913847,1.4145643,1.7591796,2.2646155,2.4155898,2.1530259,1.6738462,1.4309745,1.6082052,1.5261539,1.5491283,1.7001027,1.6640002,1.5425643,1.3554872,1.1716924,1.0338463,0.9517949,1.1881026,1.2209232,1.2800001,1.467077,1.785436,1.7033848,1.8543591,2.0939488,2.2153847,1.9298463,1.8576412,1.6475899,1.7099489,2.0676925,2.3696413,2.2153847,1.7887181,1.4736412,1.3915899,1.4342566,1.2406155,1.1454359,1.1979488,1.3620514,1.522872,1.8116925,2.2088206,2.5107694,2.5993848,2.4681027,1.9954873,1.8346668,1.975795,2.4943593,3.5544617,5.1265645,6.2588725,6.948103,7.351795,7.785026,9.028924,10.84718,12.386462,13.538463,14.936617,14.7561035,14.299898,14.808617,16.610462,19.111385,20.388103,20.447182,20.41108,21.041233,22.728207,22.416412,21.904411,22.009438,22.505028,22.09477,21.520412,20.634258,20.096,19.968002,19.718565,21.146257,20.60472,19.003078,17.444103,17.243898,16.777847,16.528412,15.842463,15.018668,15.323898,16.374155,16.249437,16.02954,16.292105,17.112617,18.458258,20.558771,22.337643,23.27959,23.446976,21.251284,21.00513,21.343182,21.851898,23.072823,24.34954,24.500515,24.165745,23.499489,22.18995,20.581745,20.562054,20.867283,20.230566,17.394873,14.043899,12.3995905,11.85477,11.749744,11.378873,11.293539,10.427077,9.321027,8.297027,7.466667,7.965539,8.979693,9.878975,10.043077,8.841846,7.1023593,7.0826674,8.024616,9.242257,10.105436,10.203898,10.8537445,10.994873,10.390975,9.6065645,10.085744,10.597744,11.017847,11.07036,10.338462,9.6295395,9.265231,9.238976,9.370257,9.304616,9.557334,9.993847,9.626257,8.677744,8.582564,8.743385,8.1066675,7.4436927,7.1122055,7.069539,6.5050263,6.0356927,5.3891287,4.640821,4.2174363,3.4133337,3.3444104,3.4330258,3.4921029,3.7448208,3.9975388,4.1058464,4.164923,4.2994876,4.6572313,4.7983594,4.778667,4.6769233,4.5522056,4.457026,2.5337439,2.1300514,1.8379488,1.7952822,1.9462565,2.044718,2.1431797,2.422154,2.4582565,2.1956925,1.9364104,2.0611284,2.162872,2.3105643,2.4155898,2.2580514,2.6617439,3.2000003,3.623385,3.9581542,4.532513,4.8016415,5.691077,6.7840004,7.975385,9.475283,10.525539,10.824206,10.630565,9.8592825,8.103385,7.785026,8.300308,8.904206,10.889847,17.578669,31.944208,31.589746,21.27754,8.1066675,1.5261539,0.8795898,0.7089231,0.7515898,0.7975385,0.6859488,0.57764107,0.5481026,0.5546667,0.5907693,0.702359,0.8730257,0.7778462,0.81394875,1.024,1.0994873,0.892718,0.8205129,0.92553854,1.1191796,1.204513,0.92553854,0.79097444,0.75487185,0.7089231,0.48902568,0.574359,0.6859488,0.827077,0.94523084,0.94523084,0.8598975,0.7187693,0.5874872,0.53825647,0.67282057,0.6826667,0.7220513,0.69251287,0.61374366,0.6268718,0.60061544,0.65969235,0.6170257,0.48902568,0.48902568,0.7318975,0.9944616,1.1224617,1.1027694,1.0535386,1.1520001,1.2668719,1.4145643,1.6180514,1.9232821,2.1792822,2.9571285,4.0992823,5.349744,6.363898,7.509334,8.3823595,9.95118,11.720206,11.733335,12.320822,13.774771,14.129231,13.065847,11.9171295,10.453334,11.303386,13.000206,14.91036,17.243898,17.194668,17.207796,16.984617,16.452925,15.793232,16.269129,17.257027,19.889233,23.945848,27.877747,25.655796,23.663591,21.172514,18.438566,16.692514,12.872206,10.561642,9.554052,9.028924,7.5520005,7.6143594,10.496001,10.322052,7.1515903,6.941539,5.5269747,4.3027697,3.2361028,2.409026,2.028308,2.0053334,2.1169233,2.7109745,4.525949,8.713847,8.992821,7.506052,7.8539495,10.069334,10.620719,11.388719,12.635899,14.122667,16.518566,21.376001,26.322054,29.892925,30.14236,27.907284,26.811079,24.379078,23.847387,25.01908,26.4599,25.481848,26.555079,29.25949,31.763695,33.808414,36.713028,43.437954,45.32185,44.52759,42.95221,42.22031,44.58995,44.07467,41.67549,38.980927,38.16041,36.552208,33.667286,31.333746,29.833849,27.894156,26.83077,26.335182,26.518976,27.972925,31.770258,33.41785,32.518566,30.884106,29.141336,26.74872,27.480618,27.178669,25.767387,23.450258,20.690052,19.859694,18.271181,16.15754,13.942155,12.20595,11.54954,10.860309,10.637129,11.378873,13.627078,16.154257,19.301744,22.035694,23.289438,21.973335,24.329847,26.610874,26.758566,24.500515,21.362873,19.078566,18.464823,17.48677,16.649847,18.983387,20.775387,21.19877,19.035898,15.182771,12.619488,10.115283,7.834257,7.7357955,9.895386,12.481642,20.73272,26.706053,24.4119,15.849027,11.001437,11.257437,5.976616,2.7602053,3.8728209,6.23918,3.383795,4.20759,4.5390773,4.0467696,6.2555904,9.45559,14.135796,15.734155,12.816411,7.0793853,10.194052,9.16677,5.937231,2.9013336,2.9144619,2.6223593,4.1058464,5.0871797,4.322462,1.5885129,1.5392822,3.373949,4.4438977,3.882667,2.6256413,4.2371287,6.816821,7.8736415,6.925129,5.5072823,4.056616,4.8082056,7.5487185,11.346052,14.555899,13.190565,12.563693,9.5606165,6.8627696,12.954257,4.70318,3.9778464,3.945026,2.8717952,4.1058464,3.249231,2.8455386,2.9472823,3.495385,4.2863593,3.895795,2.5632823,1.5130258,1.3259488,1.9364104,2.5600002,8.146052,8.539898,3.0982566,0.65641034,0.31507695,0.2297436,1.1388719,3.7874875,8.92718,11.428103,9.6,5.9634876,2.6880002,1.6016412,2.678154,8.155898,10.541949,8.54318,7.0793853,3.5282054,6.987488,8.759795,6.0028725,1.7558975,5.796103,5.937231,4.33559,2.809436,2.8225644,6.0685134,5.2414365,3.636513,2.6322052,1.6935385,5.428513,3.3312824,1.7887181,2.4943593,2.4549747,1.5655385,1.270154,0.86646163,0.28882053,0.108307704,0.032820515,0.006564103,0.006564103,0.016410258,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.016410258,0.01969231,0.029538464,0.006564103,0.009846155,0.06564103,0.2100513,0.5021539,0.3446154,0.26912823,0.512,0.8336411,0.5021539,0.5152821,0.446359,0.83035904,1.4441026,1.2964103,1.2964103,1.8182565,1.8116925,1.2865642,1.3128207,1.4342566,1.2438976,0.67282057,0.026256412,0.016410258,0.06564103,0.0951795,0.08861539,0.068923086,0.108307704,0.13128206,0.16410258,0.20020515,0.23958977,0.28882053,0.30194873,0.3249231,0.3249231,0.30851284,0.32164106,0.45620516,0.52512825,0.54482055,0.54482055,0.58092314,0.41025645,0.33805132,0.35774362,0.44307697,0.56451285,0.77128214,1.1979488,1.4244103,1.4375386,1.6311796,2.281026,3.1737437,4.5095387,5.8912826,6.3179493,7.0498466,8.41518,8.63836,7.5913854,6.774154,6.445949,7.066257,7.837539,8.103385,7.3714876,6.941539,6.892308,6.7183595,6.4656415,6.698667,6.931693,6.75118,6.5312824,6.4623594,6.560821,6.426257,5.7435904,5.2053337,4.972308,4.6539493,3.8728209,3.2656412,2.6683078,2.1530259,2.028308,1.9200002,1.7099489,1.3423591,0.92225647,0.702359,0.95835906,1.0666667,1.148718,1.2438976,1.3423591,1.086359,0.93866676,0.9156924,1.017436,1.2373334,1.2964103,1.6311796,2.2908719,3.1015387,3.6627696,4.8705645,4.8147697,4.332308,4.086154,4.562052,4.9296412,4.2141542,4.276513,5.074052,4.6834874,3.4756925,3.6036925,3.8367183,3.7448208,3.7087183,3.5872824,3.1343591,3.2262566,3.6529233,3.1277952,1.723077,1.1355898,1.020718,1.1224617,1.2832822,1.270154,1.3686155,1.5458462,1.6640002,1.4802053,1.6869745,1.8051283,1.8149745,1.723077,1.5425643,1.332513,1.1520001,1.0929232,1.1224617,1.0994873,1.1946667,1.5031796,1.6935385,1.7985642,2.2121027,1.7624617,1.6836925,1.8116925,1.9167181,1.7099489,1.9396925,1.6968206,1.5622566,1.719795,1.9528207,1.4769232,1.2570257,1.1585642,1.1060513,1.0666667,0.92225647,0.85005134,1.1848207,1.7296412,1.7558975,1.975795,2.2678976,2.1825643,1.785436,1.6640002,1.4933335,1.6410258,1.9364104,2.4943593,3.7382567,4.95918,5.622154,6.232616,6.9677954,7.6767187,9.31118,11.605334,13.003489,13.459693,14.434463,14.91036,14.680616,15.202463,16.594053,17.670565,18.159592,18.290873,18.064411,18.225233,20.263386,21.192207,21.845335,21.625437,20.65395,19.77436,18.714258,17.476925,17.496616,18.520617,18.632206,20.30277,19.459284,17.841232,16.643284,16.508718,14.91036,14.959591,15.16636,15.028514,15.028514,15.9343605,15.983591,15.698052,15.707899,16.768002,18.576412,20.374975,21.349745,21.83549,23.299284,21.162668,20.785233,20.614565,20.374975,21.057642,23.926155,23.991796,23.168001,22.360617,21.4679,19.968002,19.830154,19.593847,18.261335,15.320617,13.4170265,12.635899,12.521027,12.576821,12.2847185,11.503591,9.977437,8.549745,7.712821,7.6143594,8.444718,9.465437,10.161232,10.072617,8.805744,7.827693,8.004924,8.67118,9.334154,9.688616,10.14154,10.912822,10.820924,9.888822,9.337437,9.288206,10.036513,10.673231,10.656821,9.826463,9.009232,8.713847,8.681026,8.864821,9.416205,9.501539,9.777231,9.649232,8.982975,8.116513,7.9950776,7.6996927,7.5520005,7.5946674,7.584821,6.8496413,5.907693,4.969026,4.3027697,4.240411,3.5938463,3.3969233,3.3903592,3.4133337,3.4034874,3.6824617,3.8367183,4.164923,4.6572313,4.97559,5.1954875,5.156103,5.110154,5.028103,4.637539,2.5435898,2.6387694,2.097231,1.7788719,1.8674873,1.8970258,1.9364104,2.0118976,2.1234872,2.1924105,2.0709746,2.1169233,2.1858463,2.3368206,2.5009232,2.477949,2.9013336,3.3509746,3.6791797,4.010667,4.7524104,4.8147697,5.5072823,6.5083084,7.637334,8.864821,9.816616,10.134975,9.941334,9.153642,7.4929237,7.857231,8.470975,10.023385,13.633642,20.86072,27.211489,22.54113,13.46954,5.211898,1.5622566,0.92553854,0.6170257,0.50543594,0.47589746,0.44307697,0.46933338,0.512,0.52512825,0.5546667,0.761436,0.8369231,0.95835906,1.1158975,1.2209232,1.0994873,1.0371283,1.083077,1.1388719,1.1651284,1.1946667,0.98133343,1.0535386,1.0994873,1.014154,0.892718,0.86974365,0.8172308,0.8402052,0.955077,1.0929232,1.086359,0.9288206,0.8336411,0.8172308,0.7089231,0.446359,0.48246157,0.6432821,0.761436,0.67282057,0.76800007,0.76800007,0.65641034,0.47261542,0.318359,0.62030774,0.8402052,0.9878975,1.0994873,1.2373334,1.3620514,1.3850257,1.4375386,1.5885129,1.8248206,2.0906668,2.733949,3.8104618,5.10359,6.1078978,7.39118,8.2904625,9.531077,10.925949,11.369026,13.495796,14.592001,14.897232,14.011078,10.893129,10.522257,11.119591,12.796719,15.271386,17.864206,18.556719,17.828104,16.449642,15.392821,15.816206,17.092924,21.18236,27.602053,34.550156,38.898876,40.136208,39.827694,35.826874,28.773746,22.088207,18.326975,16.81395,15.02195,12.57354,11.264001,8.884514,9.849437,9.757539,7.896616,7.259898,5.6976414,4.2994876,3.2065644,2.4418464,1.9068719,3.5413337,3.5446157,4.5456414,7.181129,10.079181,9.012513,7.958975,8.704,10.617436,10.66995,11.956513,14.450873,16.843489,18.809437,21.011694,24.208412,27.867899,30.319592,31.136824,31.143387,28.996925,27.250874,26.95549,28.498053,31.635695,30.454157,31.839182,33.621334,35.465847,38.85949,43.720207,45.446568,44.612926,42.932518,43.247593,44.452106,45.390774,43.976208,40.82216,39.21067,39.154873,38.173542,36.529232,34.747078,33.618053,29.879797,28.586668,28.642464,29.426874,30.792208,33.056824,33.828106,33.375183,32.019695,30.155489,29.784618,28.09108,25.301334,22.058668,19.446156,18.304,17.125746,15.320617,13.039591,11.168821,10.089026,9.386667,9.750975,11.533129,14.736411,17.703386,20.457027,22.649437,23.624207,22.422976,23.765335,24.605541,23.680002,21.083899,18.297438,17.558975,17.335796,16.935387,17.010874,19.554462,19.826874,20.306053,18.576412,15.0777445,13.11836,10.364718,7.4371285,7.0957956,8.914052,9.284924,18.139898,25.928207,24.999386,15.921232,7.463385,6.1078978,3.7316926,2.225231,2.281026,3.4100516,2.6617439,3.318154,3.6562054,3.7940516,5.671385,6.3474874,10.584617,14.532925,14.851283,8.704,10.624001,8.402052,5.142975,3.370667,5.0149746,4.3684106,4.8640003,4.71959,3.3936412,1.5885129,1.6443079,3.6036925,5.0051284,5.146257,5.0904617,8.467693,7.515898,5.3005133,3.620103,3.006359,2.3335385,2.353231,3.6890259,5.924103,7.6110773,7.017026,6.987488,8.021334,10.308924,13.722258,4.7983594,2.7241027,2.9472823,3.2032824,3.5183592,3.639795,3.56759,3.698872,4.20759,5.0215387,5.077334,3.892513,2.740513,2.176,2.034872,4.141949,7.4830775,8.779488,6.810257,2.425436,1.332513,0.61374366,0.52512825,1.8806155,6.0324106,11.388719,11.867898,11.9860525,11.457642,5.21518,2.6453335,3.9253337,5.720616,6.5706673,6.872616,7.890052,8.963283,9.16677,8.169026,6.245744,8.792616,11.1294365,9.540924,4.972308,3.0293336,3.0260515,2.5862565,2.1234872,1.7394873,1.2307693,1.7132308,2.297436,2.2908719,1.7887181,1.6738462,0.88287187,0.74830776,0.5481026,0.14769232,0.032820515,0.01969231,0.15097436,0.20676924,0.12143591,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.006564103,0.006564103,0.01969231,0.029538464,0.04594872,0.029538464,0.01969231,0.08205129,0.29538465,0.47917953,0.8336411,1.148718,1.2373334,0.90584624,0.4201026,0.2855385,0.44307697,0.81394875,1.273436,1.1355898,1.1618463,1.1126155,0.95835906,0.88615394,1.1716924,1.0699488,0.8369231,0.5415385,0.03938462,0.029538464,0.04594872,0.049230773,0.04266667,0.068923086,0.0951795,0.128,0.18379489,0.23958977,0.23958977,0.29210258,0.3314872,0.3117949,0.26256412,0.28225642,0.39712822,0.47917953,0.571077,0.6465641,0.60389745,0.4135385,0.36102566,0.3708718,0.38728207,0.380718,0.47261542,0.6498462,0.86974365,1.1191796,1.4145643,2.041436,3.0260515,4.1550775,5.146257,5.622154,6.4722056,8.434873,8.832001,7.381334,6.2129235,6.3245134,6.6592827,7.0432825,7.197539,6.747898,6.692103,6.6067696,6.5247183,6.452513,6.380308,6.4754877,6.314667,6.1440005,6.052103,5.9634876,5.661539,5.2676926,4.7556925,4.2305646,3.9220517,3.383795,2.6912823,2.1267693,1.8576412,1.9331284,1.6836925,1.3587693,1.0568206,0.8402052,0.7253334,0.86646163,0.90256417,1.014154,1.1979488,1.2570257,0.9911796,0.9288206,0.9878975,1.0272821,0.8566154,1.3686155,2.0512822,2.4516926,2.6256413,3.1376412,3.7021542,3.764513,3.4330258,3.1671798,3.7809234,4.4800005,3.8334363,3.7710772,4.5817437,4.903385,4.017231,3.5446157,3.498667,3.7087183,3.817026,3.0720003,2.5665643,2.7011285,3.2328207,3.2754874,2.359795,1.6869745,1.142154,0.81394875,1.0010257,1.2340513,1.3850257,1.6311796,1.8412309,1.5885129,1.5031796,1.6410258,1.8051283,1.8379488,1.6278975,1.467077,1.3718976,1.4769232,1.7165129,1.8182565,2.169436,1.9922053,1.7263591,1.6705642,1.9692309,2.034872,1.910154,1.7558975,1.6049232,1.3686155,1.3259488,1.3128207,1.4080001,1.5786668,1.6738462,1.6443079,1.6902566,1.4276924,0.9517949,0.8369231,0.827077,0.9419488,1.2242053,1.5885129,1.8281027,1.8510771,1.8904617,1.719795,1.3784616,1.1979488,1.1848207,1.4112822,1.9659488,2.802872,3.7251284,4.7327185,5.1856413,5.723898,6.5411286,7.394462,9.419488,11.828514,13.696001,14.9628725,16.436514,16.229744,15.740719,15.799796,16.213335,15.766975,17.483488,18.546873,18.842258,18.704412,18.898052,20.420925,21.083899,20.768822,19.99754,19.908924,19.689028,18.560001,17.686975,17.427694,17.312822,17.929848,17.956104,16.928822,15.566771,15.753847,14.749539,14.815181,14.651078,14.234258,14.808617,15.51754,14.811898,14.362258,14.710155,15.24513,18.074257,19.698874,19.872822,19.751387,21.858463,20.952618,20.306053,19.620104,19.288616,20.361847,23.007181,22.964514,22.308104,21.832207,21.077335,20.132105,19.820309,18.724104,16.518566,13.978257,13.46954,13.318565,13.157744,12.816411,12.3076935,11.224616,9.711591,8.474257,7.837539,7.748924,9.068309,10.079181,10.604308,10.512411,9.731283,8.989539,9.019077,9.337437,9.580308,9.504821,10.180923,10.541949,10.226872,9.416205,8.838565,8.759795,9.317744,9.90195,10.131693,9.83959,9.186462,9.173334,9.035488,8.861539,9.586872,9.396514,9.298052,9.156924,8.92718,8.65477,8.346257,8.267488,8.116513,7.834257,7.5946674,6.619898,5.799385,4.9526157,4.1189747,3.570872,3.5380516,3.436308,3.3312824,3.2853336,3.3411283,3.5347695,3.5347695,3.8104618,4.466872,5.2414365,5.9995904,6.1997952,6.052103,5.7698464,5.5532312,3.0162053,2.9801028,2.3335385,1.9462565,1.9561027,1.7690258,1.8674873,2.038154,2.1202054,2.1136413,2.1530259,2.038154,2.0742567,2.2580514,2.5304618,2.7700515,2.9571285,3.318154,3.7021542,4.07959,4.522667,4.667077,5.3924108,6.3868723,7.4765134,8.631796,9.45559,10.230155,9.829744,8.513641,7.9261546,8.674462,9.728001,12.235488,16.534975,22.15713,19.862976,13.932309,8.060719,4.0041027,1.5622566,0.88287187,0.79425645,0.7811283,0.6432821,0.49230772,0.49230772,0.508718,0.56451285,0.6859488,0.8960001,1.0699488,1.2800001,1.3620514,1.270154,1.0699488,1.024,1.0568206,1.1716924,1.2931283,1.2537436,1.2931283,1.3161026,1.3128207,1.2603078,1.148718,1.1060513,0.9747693,0.9288206,0.9944616,1.0469744,1.014154,0.9682052,0.88943595,0.8008206,0.761436,0.446359,0.47261542,0.5973334,0.7122052,0.81394875,0.86974365,0.8008206,0.6859488,0.56123084,0.39384618,0.5284103,0.67282057,0.7844103,0.88287187,1.0535386,1.1716924,1.204513,1.3161026,1.5425643,1.8018463,2.297436,3.2361028,4.417641,5.605744,6.5280004,7.837539,8.769642,9.632821,10.610872,11.753027,13.036308,13.495796,13.11836,11.963078,10.157949,10.699488,11.569232,13.51877,16.39713,19.14749,19.27877,17.988924,17.161848,17.769028,19.879387,24.228104,32.324924,42.830772,52.52595,56.32985,55.742363,53.66154,48.318363,40.457848,33.34236,27.59549,23.207386,19.862976,16.823795,12.924719,10.043077,9.40636,9.222565,8.65477,7.8047185,6.045539,4.821334,3.9811285,3.4067695,2.993231,3.6529233,4.2436924,5.668103,8.392206,12.461949,10.33518,9.472001,10.105436,11.234463,10.633847,12.081232,15.235283,19.633232,23.962257,26.066053,28.317541,29.810875,30.516516,30.37867,29.295591,28.20267,27.890875,28.077951,29.046156,31.625849,32.75159,34.898052,37.16267,39.48308,42.640415,43.91385,43.874466,42.86031,41.53108,40.87467,41.94462,43.49703,43.897438,42.912823,41.70831,41.96431,41.974155,41.137234,39.699696,38.757748,33.38503,31.3239,31.01867,31.186054,30.815182,32.226463,32.78113,33.106052,33.457233,33.716515,31.875284,29.879797,26.607592,22.478771,19.419899,17.51631,16.728617,15.563488,13.5548725,11.247591,9.6754875,9.199591,10.197334,12.566976,15.747283,19.035898,21.700924,23.250053,23.348515,21.796104,21.80595,22.393438,21.415386,18.91118,17.083078,16.971489,17.312822,17.85436,18.789745,20.752413,20.296207,20.184616,18.218668,15.087591,14.342566,11.319796,9.143796,8.333129,8.562873,8.667898,15.074463,24.44472,25.796925,17.152,5.543385,4.0992823,2.858667,1.9035898,1.5556924,2.3893335,2.556718,2.934154,3.3641028,3.9253337,4.9296412,4.6539493,8.369231,12.711386,14.677335,11.59877,12.294565,8.94359,5.2611284,4.010667,7.02359,8.326565,7.0498466,4.919795,2.9997952,1.6968206,1.6278975,3.0129232,5.395693,7.433847,6.925129,9.265231,6.1308722,3.0785644,2.225231,2.2350771,2.2482052,1.8609232,1.9396925,2.5107694,2.7634873,3.1343591,3.6463592,7.6110773,12.20595,8.487385,3.8465643,2.2514873,3.1934361,5.100308,5.3398976,3.9844105,3.7776413,4.1124105,4.709744,5.61559,5.970052,4.9985647,3.8990772,3.1507695,2.537026,3.4100516,5.85518,7.955693,7.9852314,4.397949,3.0129232,2.3236926,1.6016412,1.1782565,2.425436,4.8836927,7.072821,10.998155,13.449847,5.9995904,3.0030773,2.7864618,3.1606157,3.4198978,4.338872,5.5105643,5.398975,5.031385,5.0182567,5.5565133,7.312411,10.456616,10.515693,7.141744,4.135385,3.2820516,2.6617439,2.281026,1.9528207,1.2800001,2.1136413,2.4681027,2.3368206,1.972513,1.8740515,0.88615394,0.5907693,2.7076926,4.7491283,0.02297436,0.052512825,0.15753847,0.23630771,0.2100513,0.01969231,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.006564103,0.01969231,0.03938462,0.055794876,0.04594872,0.01969231,0.029538464,0.15097436,0.2231795,0.761436,1.1027694,1.0338463,0.7778462,0.40369233,0.30194873,0.34789747,0.512,0.8730257,1.1355898,1.148718,1.0371283,0.90256417,0.8336411,1.0896411,1.1684103,1.276718,1.2438976,0.5481026,0.128,0.026256412,0.026256412,0.026256412,0.04266667,0.06564103,0.0951795,0.15097436,0.21989745,0.2297436,0.28882053,0.3314872,0.3117949,0.256,0.26584616,0.30851284,0.38728207,0.5152821,0.63343596,0.6104616,0.51856416,0.446359,0.41682056,0.41682056,0.380718,0.38400003,0.43651286,0.58092314,0.8369231,1.1749744,1.6443079,2.6289232,3.623385,4.5554876,5.7764106,7.174565,8.914052,9.091283,7.7948723,7.1089234,6.8233852,6.9776416,6.994052,6.669129,6.180103,5.9536414,6.058667,6.23918,6.3540516,6.373744,6.2096415,5.937231,5.8289237,5.8453336,5.668103,5.149539,4.6572313,4.1124105,3.6069746,3.3903592,2.92759,2.3335385,1.9003079,1.719795,1.6968206,1.3193847,1.0535386,0.8992821,0.8172308,0.7318975,0.75487185,0.7778462,0.88615394,1.0469744,1.1158975,0.9156924,0.9419488,1.0272821,1.0436924,0.892718,1.1979488,1.9003079,2.349949,2.5337439,3.0687182,3.0260515,2.7766156,2.7798977,3.2295387,4.0434875,4.466872,4.076308,3.879385,4.1550775,4.46359,4.2535386,4.0369234,3.9187696,3.9844105,4.2830772,3.3509746,2.737231,2.6354873,2.9472823,3.2918978,2.6322052,1.8838975,1.2471796,0.9124103,1.0404103,1.1355898,1.3226668,1.6738462,2.0742567,2.2219489,1.8642052,1.910154,1.9954873,1.9298463,1.7033848,1.6213335,1.5819489,1.7132308,1.9528207,2.034872,2.048,1.9396925,1.8346668,1.8116925,1.8970258,1.7788719,1.5491283,1.4867693,1.5786668,1.4998976,1.142154,1.0699488,1.1224617,1.2438976,1.4998976,1.7329233,1.6475899,1.3587693,1.0469744,0.9353847,0.96492314,0.9747693,1.1158975,1.4112822,1.7624617,1.7624617,1.6049232,1.3489232,1.079795,0.9288206,0.9156924,1.2996924,2.103795,3.121231,3.895795,4.535795,4.8377438,5.402257,6.498462,8.04759,10.758565,12.560411,14.086565,15.586463,16.928822,16.475899,15.632411,15.419078,15.898257,16.167385,16.846771,17.739489,18.297438,18.399181,18.33354,18.871796,19.472412,19.728413,19.75795,20.227283,19.731693,18.169437,17.214361,17.115898,16.689232,16.20349,16.538258,16.141129,14.985847,14.565744,13.4859495,13.564719,13.6697445,13.620514,14.178463,14.887385,13.659899,13.213539,14.217847,15.264822,17.70995,19.035898,19.072002,18.707693,19.925335,19.561028,19.11795,18.504206,18.287592,19.692308,21.700924,22.137438,21.85518,21.30708,20.54236,19.538054,18.852104,17.411283,15.333745,13.915898,13.978257,13.978257,13.745232,13.141335,12.068104,10.840616,9.488411,8.5202055,8.113232,8.093539,9.488411,10.358154,10.738873,10.765129,10.640411,9.980719,9.895386,10.026668,10.036513,9.632821,10.322052,10.341744,9.852718,9.120821,8.5202055,8.868103,9.478565,10.006975,10.164514,9.741129,8.969847,9.019077,9.012513,8.861539,9.271795,9.360411,9.032206,8.864821,8.992821,9.117539,9.028924,8.94359,8.5891285,7.939283,7.213949,6.426257,5.8289237,5.097026,4.2305646,3.56759,3.6463592,3.4658465,3.3509746,3.3936412,3.4724104,3.636513,3.7087183,3.9942567,4.5817437,5.356308,5.904411,6.088206,6.0849237,6.0225644,5.976616,3.0818465,2.8258464,2.2777438,2.0053334,2.03159,1.8313848,1.8904617,2.1070771,2.1366155,1.9659488,1.9364104,1.8773335,1.972513,2.1300514,2.3794873,2.861949,2.930872,3.3280003,3.7940516,4.1485133,4.315898,4.519385,5.2709746,6.186667,7.13518,8.228104,9.07159,10.036513,9.547488,8.182155,8.6580515,10.075898,11.306667,13.715693,17.171694,20.073027,13.88636,8.533334,5.1889234,3.5347695,1.7526156,1.1749744,1.2373334,1.2603078,1.014154,0.7122052,0.5907693,0.61374366,0.7515898,0.9485129,1.1355898,1.3883078,1.5589745,1.5392822,1.3522053,1.1520001,0.9419488,0.93866676,1.1126155,1.332513,1.3587693,1.4080001,1.4276924,1.4342566,1.3981539,1.2274873,1.2865642,1.214359,1.1749744,1.2307693,1.339077,1.3161026,1.2668719,1.024,0.69251287,0.63343596,0.4266667,0.508718,0.6498462,0.78769237,0.99774367,0.9616411,0.8795898,0.764718,0.62030774,0.42338464,0.48574364,0.5513847,0.5973334,0.6629744,0.8467693,0.9878975,1.1126155,1.3062565,1.5688206,1.8051283,2.4155898,3.4921029,4.8114877,6.166975,7.3747697,8.986258,9.980719,10.541949,11.162257,12.632616,12.356924,12.058257,11.319796,10.469745,10.581334,12.107488,13.90277,16.082052,18.520617,20.854155,21.064207,21.707489,23.555285,26.479591,29.45313,34.45826,40.58585,47.382977,52.99857,54.193233,52.41108,50.100517,46.08,40.854977,36.578465,31.143387,25.737848,21.428514,17.78872,12.911591,10.79795,9.288206,8.848411,8.982975,8.251078,6.560821,5.5663595,5.35959,5.405539,4.5423594,4.1058464,5.924103,7.906462,9.488411,11.644719,11.093334,11.001437,11.638155,12.412719,11.874462,13.860104,17.188105,21.35631,25.219284,27.00472,28.813131,30.10954,30.162054,28.685131,25.842875,26.0759,28.22236,30.208002,31.251696,31.862156,34.550156,37.51713,40.66462,43.654568,45.90277,44.721233,42.837337,41.26195,40.359386,39.844105,39.9918,40.536617,41.62298,43.02113,44.114056,44.58995,44.973953,44.642464,43.651287,42.71262,37.36944,34.645336,33.473644,32.87631,31.944208,31.789951,31.458464,32.11159,33.870773,35.810463,34.12021,32.623592,29.105232,23.863796,19.718565,17.746052,17.220924,16.984617,15.858873,12.632616,10.906258,10.902975,12.2847185,14.6182575,17.401438,20.309336,22.629745,23.483078,22.665848,20.624413,19.734976,20.378258,19.843283,17.962667,17.138874,17.362053,17.913437,18.884924,20.276514,21.989746,21.497438,20.854155,18.983387,16.728617,16.856617,13.955283,11.67754,10.131693,9.393231,9.508103,13.984821,22.79713,25.504822,18.776617,6.413129,4.269949,2.8356924,1.7591796,1.1979488,1.8149745,2.3991797,2.789744,3.436308,4.1485133,4.092718,4.194462,7.6570263,11.21477,13.203693,13.551591,14.221129,10.919386,7.3747697,6.157129,8.687591,12.724514,9.990565,6.1472826,3.6102567,1.5458462,1.8674873,2.868513,6.121026,9.580308,7.5881033,8.681026,5.0215387,2.2219489,2.1497438,2.9046156,3.383795,2.4352822,1.404718,0.8598975,0.55794877,1.1552821,1.8707694,5.7140517,9.688616,4.775385,3.3805132,2.231795,2.8816411,4.965744,6.1997952,4.027077,3.6791797,4.125539,4.9099493,6.1538467,6.6822567,5.927385,5.2611284,4.844308,3.629949,3.3247182,4.2502565,6.4295387,8.260923,6.5083084,4.516103,3.2918978,2.2646155,1.3456411,0.9419488,1.0010257,2.861949,6.7577443,9.69518,5.4580517,2.8816411,2.3794873,2.3893335,2.428718,3.0818465,2.8914874,2.2449234,1.7066668,1.7887181,2.9571285,4.7622566,6.744616,7.2336416,5.8486156,3.501949,2.6715899,2.1891284,2.4352822,3.0982566,3.170462,3.9286156,4.0369234,3.5741541,2.8225644,2.300718,1.020718,0.67282057,2.9801028,5.2348723,0.3117949,0.8336411,1.3128207,1.0043077,0.16082053,0.04266667,0.055794876,0.07876924,0.06235898,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.01969231,0.032820515,0.049230773,0.052512825,0.04266667,0.04594872,0.108307704,0.04266667,0.51856416,0.90256417,0.9124103,0.6071795,0.71548724,0.56451285,0.5284103,0.65641034,0.6662565,1.214359,1.4309745,1.4572309,1.4178462,1.4178462,1.3915899,1.7132308,1.8871796,1.5786668,0.6104616,0.14769232,0.016410258,0.013128206,0.016410258,0.01969231,0.03938462,0.06564103,0.1148718,0.18379489,0.24615386,0.27897438,0.28882053,0.26912823,0.23630771,0.24615386,0.28225642,0.34133336,0.43651286,0.5284103,0.5481026,0.5284103,0.45620516,0.4266667,0.4397949,0.42338464,0.39384618,0.39712822,0.48902568,0.69251287,1.0043077,1.3554872,2.2219489,3.1638978,4.1550775,5.5926156,7.2172313,8.904206,9.554052,8.907488,7.522462,6.8332314,6.7150774,6.491898,5.973334,5.47118,5.074052,5.356308,5.6254363,5.7107697,5.979898,5.7731285,5.4843082,5.366154,5.35959,5.1232824,4.5522056,3.9089234,3.3575387,2.9735386,2.7569232,2.412308,2.0184617,1.7362052,1.5688206,1.3784616,1.0371283,0.88287187,0.8402052,0.81394875,0.6892308,0.69251287,0.72861546,0.81394875,0.9189744,0.9878975,0.9321026,0.9485129,1.0305642,1.086359,0.93866676,1.0338463,1.6278975,2.1267693,2.3991797,2.7963078,2.9078977,2.5173335,2.674872,3.6069746,4.6966157,4.6834874,4.420923,4.2371287,4.2371287,4.312616,4.4800005,4.417641,4.31918,4.2962055,4.381539,3.748103,3.245949,2.9210258,2.9078977,3.4034874,2.937436,2.162872,1.4867693,1.0896411,0.955077,0.9485129,1.270154,1.7132308,2.1169233,2.3696413,2.0841026,2.1530259,2.2416413,2.162872,1.8445129,1.7952822,1.7624617,1.8313848,1.9659488,2.0053334,1.8806155,2.0578463,2.1234872,1.9954873,1.910154,1.8248206,1.529436,1.4244103,1.5360001,1.5327181,1.086359,1.0108719,1.1093334,1.2865642,1.5491283,1.6213335,1.401436,1.2242053,1.148718,0.98133343,1.0535386,1.0338463,1.0896411,1.2996924,1.6410258,1.6049232,1.3062565,0.9714873,0.7450257,0.6662565,0.7811283,1.401436,2.3860514,3.4297438,4.056616,4.384821,4.775385,5.674667,7.207385,9.18318,11.67754,12.672001,13.636924,14.985847,16.06236,16.036104,15.291079,15.29436,16.308514,17.408,17.371899,17.772308,17.913437,17.706669,17.650873,17.509745,17.64759,18.228514,19.058874,19.616821,19.34113,17.923283,17.083078,17.063385,16.636719,15.635694,15.701335,15.353437,14.313026,13.522053,12.544001,12.445539,12.803283,13.321847,13.830565,14.224411,13.019898,12.721231,13.945437,15.442053,16.856617,18.011898,18.310566,17.969233,18.008617,17.824821,17.51631,17.178257,17.32595,18.888206,20.555489,21.382566,21.362873,20.640821,19.515078,18.386053,17.43754,16.075489,14.608412,14.227694,14.496821,14.345847,13.833847,12.944411,11.595488,10.522257,9.31118,8.65477,8.648206,8.812308,9.737847,10.453334,10.807796,10.893129,11.0375395,10.55836,10.686359,10.95877,10.889847,9.987283,10.568206,10.325335,9.655796,8.937026,8.52677,9.278359,9.895386,10.240001,10.187488,9.642668,8.871386,8.832001,8.825437,8.707283,8.89436,8.969847,8.5202055,8.444718,8.937026,9.485129,9.659078,9.6065645,9.101129,8.198565,7.2336416,6.413129,5.858462,5.2447186,4.5489235,4.0369234,4.066462,3.8695388,3.7874875,3.8596926,3.826872,3.7743592,3.9351797,4.2502565,4.706462,5.3366156,5.7435904,5.8223596,5.8847184,6.0291286,6.157129,2.681436,2.4385643,2.0939488,1.9462565,2.0053334,1.9922053,1.9331284,2.03159,2.0184617,1.8412309,1.6902566,1.7624617,1.975795,2.0775387,2.162872,2.6551797,2.8258464,3.31159,3.8038976,4.132103,4.276513,4.4734364,5.149539,5.927385,6.7117953,7.686565,8.562873,9.170052,8.858257,8.214975,9.061745,10.9226675,11.805539,12.937847,14.28677,14.565744,10.056206,6.298257,4.138667,3.2361028,2.03159,1.6902566,1.6180514,1.522872,1.2832822,0.9682052,0.7515898,0.78769237,0.9682052,1.1881026,1.3751796,1.654154,1.6935385,1.6114873,1.4769232,1.3292309,1.0043077,0.9944616,1.1585642,1.3653334,1.4998976,1.3423591,1.4178462,1.5327181,1.5163078,1.2209232,1.4244103,1.4802053,1.5622566,1.7723079,2.1530259,2.162872,1.910154,1.3554872,0.7122052,0.45620516,0.39712822,0.5907693,0.827077,1.0108719,1.148718,1.0371283,0.97805136,0.8467693,0.6170257,0.36430773,0.44964105,0.45620516,0.46276927,0.53825647,0.7581539,0.9419488,1.1520001,1.3686155,1.5622566,1.7263591,2.2416413,3.3017437,4.8016415,6.550975,8.280616,10.105436,11.657847,12.11077,12.064821,13.548308,12.156719,11.329642,10.965334,11.290257,12.872206,15.274668,18.146463,20.453745,21.983181,23.32554,24.927181,28.99036,33.654156,37.471184,39.41744,41.327595,40.48739,38.07508,35.30831,33.437542,32.68595,32.298668,31.471592,30.178463,29.200413,26.3319,22.692104,18.884924,15.24513,11.864616,11.011283,9.645949,8.999385,9.061745,8.585847,7.1647186,6.308103,6.7938466,7.8802056,7.2960005,5.6352825,8.43159,10.755282,10.44677,8.123077,10.000411,10.866873,12.012309,13.499078,14.178463,17.952822,20.453745,21.609028,21.979898,22.784002,24.244514,27.119593,28.547285,27.290258,23.742361,25.232412,28.603079,32.295387,34.665028,33.96595,36.15508,39.230362,43.00144,46.46072,47.776825,46.529644,43.907284,41.862568,41.199593,41.56062,39.844105,38.32123,38.593643,40.976414,44.48821,46.116108,46.71672,46.270363,45.25949,44.672005,41.458874,38.63959,36.36185,34.628925,33.312824,31.783386,30.71672,31.343592,33.53272,35.764515,36.158363,35.567593,31.845745,25.609848,20.256823,18.54031,18.422155,19.131079,18.930874,15.104001,13.341539,13.751796,15.169642,17.02072,19.311592,21.270975,22.951385,23.27631,21.96349,19.528206,18.41231,18.760206,18.802874,18.264616,18.353231,18.665028,18.970259,19.70872,21.280823,24.027899,23.578259,22.439386,21.03795,20.066463,20.49313,17.942976,15.113848,12.901745,11.746463,11.634872,14.916924,21.159386,23.7719,19.74154,9.6295395,5.546667,3.3378465,1.9167181,1.020718,1.2307693,2.1169233,2.802872,3.5938463,4.1780515,3.6102567,4.6802053,7.7456417,10.069334,11.441232,14.155488,14.8020525,12.3766165,9.977437,9.048616,9.38995,14.54277,11.759591,7.6209235,4.6867695,1.4933335,2.1989746,3.4034874,6.6100516,9.734565,7.1220517,8.155898,5.10359,2.7831798,2.9702566,4.4077954,4.916513,3.4067695,1.6213335,0.5349744,0.3708718,0.5349744,1.0338463,2.5140514,4.3651285,4.7261543,4.785231,3.2722054,2.1825643,2.6518977,4.965744,3.7054362,3.4560003,3.8596926,4.8147697,6.449231,7.13518,6.6625648,6.6133337,6.8004107,5.2512827,4.9362054,3.9778464,4.926359,7.1647186,6.9120007,4.630975,2.7700515,1.847795,1.7033848,1.4802053,1.7887181,2.048,2.8553848,3.9351797,4.141949,2.917744,2.231795,2.428718,3.1113849,3.1606157,2.169436,1.8281027,1.4506668,1.3522053,2.8389745,4.5456414,4.6276927,4.128821,3.4625645,2.4385643,0.94523084,0.86317956,2.2678976,4.312616,5.2315903,4.4800005,4.893539,4.5095387,3.1113849,2.2186668,0.98461545,0.8172308,1.3850257,1.8576412,0.8960001,1.7788719,2.9013336,2.1103592,0.03938462,0.118153855,0.12143591,0.15753847,0.13128206,0.04266667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0032820515,0.006564103,0.013128206,0.01969231,0.03938462,0.052512825,0.068923086,0.10502565,0.17066668,0.07876924,0.3052308,0.65312827,0.8336411,0.46933338,1.0469744,0.8172308,0.69579494,0.83035904,0.60389745,1.1815386,1.5491283,1.9035898,2.2022567,2.15959,1.7001027,2.359795,2.422154,1.4309745,0.17066668,0.055794876,0.009846155,0.0032820515,0.009846155,0.0,0.013128206,0.03938462,0.07876924,0.14112821,0.24943592,0.25271797,0.21989745,0.19692309,0.20020515,0.22646156,0.30851284,0.3511795,0.37743592,0.4135385,0.45620516,0.4266667,0.38728207,0.39712822,0.446359,0.4660513,0.45620516,0.446359,0.49887183,0.65312827,0.92553854,1.2832822,1.9200002,2.7602053,3.7415388,4.818052,6.304821,8.28718,9.96759,10.171078,7.3583593,6.4656415,6.0291286,5.737026,5.3891287,4.886975,4.381539,4.640821,4.7917953,4.7327185,5.139693,4.9985647,4.7491283,4.6112823,4.5489235,4.2568207,3.8367183,3.245949,2.740513,2.3893335,2.0676925,1.9167181,1.723077,1.5458462,1.3751796,1.1093334,0.9485129,0.86646163,0.8336411,0.79097444,0.6465641,0.69579494,0.7384616,0.78769237,0.8467693,0.90912825,1.0108719,0.9485129,1.0469744,1.2340513,1.0502565,1.0371283,1.4933335,1.9954873,2.3335385,2.5271797,3.2722054,3.0720003,3.0818465,3.8038976,5.0871797,4.900103,4.565334,4.532513,4.772103,4.772103,4.9362054,4.673641,4.5587697,4.630975,4.381539,4.1452312,3.876103,3.4756925,3.1770258,3.5741541,3.1474874,2.4681027,1.8149745,1.2898463,0.8041026,0.7778462,1.2438976,1.8215386,2.1989746,2.1169233,1.9889232,2.1464617,2.3630772,2.4057438,2.0250258,1.9692309,1.9068719,1.9429746,2.0217438,1.9593848,2.0250258,2.4418464,2.4648206,2.044718,1.8215386,2.028308,1.8379488,1.591795,1.4408206,1.3522053,1.0699488,1.1684103,1.4375386,1.6640002,1.6640002,1.3686155,1.1881026,1.1913847,1.2307693,0.9419488,1.0469744,1.142154,1.1749744,1.1979488,1.3817437,1.270154,0.9288206,0.5973334,0.4201026,0.44307697,0.9517949,1.8674873,2.9046156,3.7776413,4.204308,4.4340515,5.080616,6.38359,8.214975,10.052924,11.608616,12.225642,12.777026,13.574565,14.401642,15.051488,14.972719,15.507693,16.866463,18.116924,18.740515,19.006361,18.425438,17.332514,16.866463,16.935387,16.406975,16.649847,17.723078,18.376207,18.67159,18.176,17.32595,16.633438,16.679386,15.980309,15.488001,14.608412,13.433437,12.711386,12.07795,11.940104,12.389745,13.190565,13.745232,13.692719,13.036308,12.849232,13.607386,15.189335,15.573335,16.626873,17.332514,17.283283,16.679386,16.23631,15.80636,15.783386,16.459488,18.028309,19.813745,20.736002,20.74913,19.872822,18.179283,17.043694,16.072206,15.14995,14.480412,14.592001,14.884104,14.378668,13.371078,12.160001,11.034257,10.269539,9.186462,8.805744,9.252103,9.764103,10.006975,10.456616,10.778257,10.870154,10.8767185,10.7848215,11.365745,11.904001,11.785847,10.502565,10.955488,10.614155,9.8363085,9.078155,8.904206,9.724719,10.200616,10.289231,10.026668,9.531077,8.868103,8.674462,8.487385,8.277334,8.43159,8.2215395,7.768616,7.8703594,8.664616,9.626257,9.931488,10.072617,9.6295395,8.648206,7.634052,6.5083084,5.914257,5.47118,5.0674877,4.84759,4.7261543,4.4996924,4.3651285,4.2929235,4.0434875,3.7218463,3.879385,4.1813335,4.562052,5.2053337,5.832206,5.8814363,5.904411,6.117744,6.413129,2.546872,2.6453335,2.349949,2.0250258,1.8707694,1.9068719,1.9068719,1.8149745,1.785436,1.8970258,2.166154,1.8970258,2.1431797,2.3138463,2.2514873,2.228513,2.5435898,2.8980515,3.3509746,3.8498464,4.2272825,4.5817437,5.1265645,5.8912826,6.7840004,7.6143594,8.090257,7.9524107,8.050873,8.487385,8.621949,9.097847,9.170052,8.677744,7.778462,6.9743595,5.910975,4.345436,3.3509746,2.9243078,1.9823592,1.7887181,1.2898463,1.0535386,1.1388719,1.1126155,1.0043077,0.8566154,0.892718,1.1323078,1.3883078,1.8051283,1.6508719,1.4998976,1.5130258,1.463795,1.5392822,1.5556924,1.6180514,1.7066668,1.6935385,1.595077,1.5261539,1.6836925,1.8445129,1.3423591,1.5261539,1.6082052,1.9626669,2.6289232,3.3247182,3.2164104,2.6584618,1.8642052,1.1027694,0.6859488,0.6498462,0.90584624,1.0896411,1.1093334,1.1585642,1.0502565,0.9321026,0.7844103,0.6071795,0.4135385,0.31507695,0.318359,0.39056414,0.52512825,0.7318975,0.8795898,1.0436924,1.1585642,1.2406155,1.3718976,1.7526156,3.245949,5.1265645,6.9842057,8.743385,9.622975,13.128206,13.75836,11.897437,13.840411,12.3995905,11.85477,12.471796,14.385232,17.608206,20.148514,23.089233,25.652515,27.241028,27.451078,31.159798,35.83344,39.05641,39.72267,38.02585,35.13108,31.176207,26.735592,23.04,21.989746,21.733746,21.67795,21.779694,21.520412,19.899078,17.42113,14.647796,13.226667,12.731078,10.679795,10.706052,10.630565,10.276103,9.682052,9.110975,7.7292314,6.882462,7.381334,9.603283,13.472821,7.9425645,9.77395,11.385437,9.895386,7.1122055,6.340924,6.744616,9.07159,12.724514,15.776822,23.56513,23.122053,20.736002,19.80718,20.844309,21.553232,23.14831,24.815592,25.586874,24.352823,26.817642,27.26072,30.424618,35.222977,34.76021,37.054363,40.018055,43.618465,47.03508,48.64657,49.388313,47.983593,46.749542,46.017643,44.114056,41.09785,38.34749,37.51713,38.71508,40.497234,45.124928,46.408207,44.980515,42.88985,43.60862,44.878773,43.401848,40.549747,37.074055,33.079796,31.445335,30.20472,30.687181,32.564514,33.860924,36.90995,37.116722,33.539284,27.336206,21.760002,18.743795,19.830154,21.014977,20.36513,18.021746,15.51754,15.652103,16.8599,18.323694,19.958155,21.251284,22.482054,22.836515,21.812515,19.209848,18.271181,17.506462,18.116924,19.866259,21.087181,20.696617,20.627693,21.054361,23.125336,28.960823,27.53313,25.160208,23.722668,23.72595,24.336412,21.651693,20.86072,18.7799,15.786668,15.82277,15.530668,19.347694,21.205336,18.697847,13.108514,6.7610264,4.2568207,2.6584618,1.1552821,1.083077,2.2547693,3.062154,3.4756925,3.7316926,4.31918,5.7107697,7.0465646,8.395488,10.505847,14.815181,11.789129,9.275078,8.969847,9.842873,8.132924,9.475283,9.160206,7.318975,4.6900516,2.6387694,1.9331284,3.8137438,5.1889234,5.3760004,6.1341543,8.513641,5.8518977,3.8432825,4.4307694,5.799385,5.61559,4.342154,2.537026,0.9189744,0.380718,0.57764107,0.571077,0.98461545,2.3466668,5.080616,9.278359,6.9054365,3.239385,1.4736412,2.7306669,3.170462,3.2722054,3.620103,4.532513,6.058667,7.0465646,7.1122055,7.240206,7.509334,7.0957956,7.3747697,6.675693,4.5522056,2.103795,1.9692309,1.785436,1.3357949,1.1520001,1.2242053,0.9911796,2.2383592,2.5862565,2.7142565,2.6289232,1.6640002,5.2644105,3.7940516,1.785436,1.1355898,1.0994873,1.1093334,2.8521028,3.43959,4.204308,10.712616,10.06277,10.571488,10.095591,8.211693,6.2096415,1.7657437,1.3423591,2.8258464,4.0467696,2.7766156,1.1158975,0.60061544,0.5152821,0.571077,0.8992821,0.7417436,0.77456415,2.3433847,4.010667,1.5556924,1.0305642,2.1924105,1.8445129,0.0951795,0.3511795,0.068923086,0.0,0.029538464,0.06235898,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.016410258,0.016410258,0.009846155,0.006564103,0.029538464,0.029538464,0.03938462,0.08205129,0.17066668,0.3052308,0.13456412,0.06564103,0.04594872,0.04266667,0.029538464,0.51856416,0.4955898,0.28225642,0.09189744,0.029538464,0.71548724,0.93866676,1.5688206,2.3302567,1.8313848,1.0371283,2.2580514,2.484513,1.1355898,0.06235898,0.02297436,0.006564103,0.0,0.0,0.0,0.013128206,0.032820515,0.059076928,0.09189744,0.15097436,0.21333335,0.2100513,0.19364104,0.190359,0.21333335,0.2855385,0.3314872,0.380718,0.43323082,0.45620516,0.34789747,0.34789747,0.4135385,0.5021539,0.56451285,0.61374366,0.58092314,0.49887183,0.5218462,0.8992821,1.3751796,1.6968206,2.1366155,2.9013336,4.135385,5.796103,7.7948723,9.6754875,10.397539,8.346257,7.066257,6.5444107,6.3277955,5.9963083,5.142975,4.1911798,4.07959,4.1911798,4.273231,4.457026,3.892513,3.4527183,3.501949,3.7940516,3.4625645,3.2689233,3.1015387,2.6978464,2.1136413,1.723077,1.7132308,1.5819489,1.4112822,1.2406155,1.083077,1.0699488,0.92225647,0.7811283,0.7187693,0.7318975,0.7318975,0.7318975,0.7384616,0.77456415,0.88615394,0.9944616,0.95835906,1.1782565,1.5983591,1.7099489,1.3062565,1.5622566,2.2350771,2.9801028,3.3575387,3.9056413,3.9417439,3.6004105,3.4625645,4.562052,4.844308,4.4373336,4.516103,5.1987696,5.5532312,5.786257,5.421949,5.149539,5.2381544,5.5532312,5.0051284,4.630975,4.2272825,3.7940516,3.5249233,2.609231,2.2350771,2.0250258,1.719795,1.1585642,0.8795898,1.1946667,2.1103592,3.0096412,2.6551797,1.910154,1.9068719,2.1136413,2.2219489,2.1366155,2.0873847,2.028308,2.2482052,2.5206156,2.1070771,2.1431797,2.5731285,2.4943593,1.8346668,1.3587693,1.2603078,1.4933335,1.6311796,1.5360001,1.3259488,1.2307693,1.5885129,1.8215386,1.7132308,1.4178462,1.211077,1.1782565,1.3423591,1.4802053,1.1126155,1.1388719,1.2832822,1.1946667,0.892718,0.74830776,0.6268718,0.45620516,0.34133336,0.3446154,0.5021539,1.6738462,2.9111798,3.8038976,4.266667,4.5456414,4.962462,5.6976414,6.8266673,8.234667,9.613129,11.040821,12.47836,12.882052,12.507898,12.924719,13.436719,14.224411,14.982565,15.770258,17.027283,19.177027,20.263386,19.830154,18.294155,16.951796,17.391592,16.715488,16.026258,16.265848,18.218668,17.54913,18.002052,16.994463,15.094155,16.022976,16.229744,15.458463,14.12595,12.711386,11.733335,10.965334,11.74318,12.517745,12.806565,13.184001,13.453129,13.50236,13.078976,12.918155,14.723283,14.601848,15.287796,16.249437,16.899282,16.571077,14.936617,14.290052,14.660924,15.852309,17.440823,19.442873,20.41108,20.312616,19.203283,17.227488,16.042667,15.235283,15.064616,15.31077,15.274668,15.274668,14.247386,12.711386,11.2672825,10.620719,9.924924,9.091283,8.864821,9.449026,10.499283,10.679795,10.407386,10.35159,10.584617,10.55836,11.024411,11.825232,12.173129,11.835078,11.139283,11.542975,11.457642,10.860309,10.039796,9.613129,10.003693,10.28595,10.259693,9.885539,9.26195,8.3823595,8.100103,7.837539,7.4929237,7.430565,7.50277,7.240206,7.4043083,8.208411,9.3078985,9.626257,10.098872,10.006975,9.097847,7.584821,6.413129,6.193231,6.0816417,5.861744,5.933949,5.3136415,4.699898,4.194462,3.7874875,3.370667,3.2262566,3.318154,3.495385,3.8990772,4.97559,5.9503593,6.2129235,6.377026,6.705231,7.0957956,2.097231,2.359795,2.2744617,2.038154,1.847795,1.8838975,1.9626669,1.7952822,1.7099489,1.785436,1.847795,1.657436,1.847795,2.0545642,2.100513,2.0086155,2.4713848,2.8849232,3.3542566,3.8104618,3.9811285,4.1813335,4.6276927,5.464616,6.4065647,6.7610264,7.1680007,7.394462,7.2172313,6.7610264,6.485334,6.3474874,6.308103,6.1407185,5.917539,6.009436,5.172513,4.1517954,3.4658465,3.0884104,2.4582565,2.166154,1.7920002,1.4703591,1.3161026,1.4178462,1.211077,1.1355898,1.1782565,1.276718,1.3259488,1.9167181,1.8740515,1.6410258,1.4473847,1.3292309,1.4342566,1.5622566,1.7263591,1.8609232,1.8412309,2.0250258,2.100513,2.0906668,1.972513,1.6475899,1.5786668,1.8609232,2.2678976,2.6486156,2.937436,3.3641028,2.917744,1.9462565,0.95835906,0.60061544,0.54482055,0.5021539,0.5218462,0.5677949,0.53825647,0.4266667,0.37415388,0.35446155,0.34789747,0.33805132,0.34789747,0.42994875,0.5316923,0.6301539,0.7187693,0.827077,0.92553854,1.020718,1.148718,1.3620514,1.6016412,2.9407182,4.955898,6.9743595,8.04759,8.448001,10.400822,11.700514,12.100924,13.289026,14.280207,15.465027,16.8599,18.36308,19.767796,23.568413,27.264002,28.586668,27.608618,26.742155,26.880003,27.664412,28.245335,28.232206,27.687387,28.212515,26.151386,23.282873,21.057642,20.585028,19.780924,18.789745,18.100513,17.811693,17.650873,16.73518,14.9398985,13.83713,13.59754,13.000206,14.391796,14.355694,13.354668,11.943385,10.794667,9.7673855,9.7673855,9.783795,10.164514,12.619488,10.965334,12.698257,15.153232,15.983591,13.15118,9.990565,8.434873,9.846154,13.065847,14.39836,18.202257,19.328001,19.557745,20.017233,21.159386,23.089233,23.424002,23.80472,24.904207,26.417233,28.803284,32.07549,34.93416,36.66708,37.152824,36.450466,36.79508,38.340927,40.86154,43.762875,47.524105,49.867493,50.53375,49.775593,48.3479,45.35467,41.078156,38.324516,37.99631,39.105644,40.63508,41.30134,40.868107,39.92944,39.899902,41.862568,42.285954,41.06175,38.57395,35.70544,32.262566,29.374361,28.320822,29.646772,33.174976,37.848618,39.138466,35.35098,28.146873,22.54113,20.512821,20.739285,21.225027,20.814772,19.193438,16.515284,16.128002,17.45395,19.56759,21.202053,21.822361,22.298258,22.534565,22.245745,20.94277,19.662771,19.272207,20.516104,22.872618,24.54318,24.884514,24.454565,23.54872,22.505028,21.697643,19.840002,21.162668,23.282873,24.425028,23.433847,23.171284,21.234873,18.756924,17.161848,18.15631,17.51959,16.374155,18.405745,21.024822,15.366566,9.419488,5.98318,3.6036925,2.0250258,2.2055387,2.422154,3.7349746,4.4340515,4.4242053,5.2447186,4.273231,6.36718,8.254359,9.91836,14.608412,10.47959,6.2818465,4.263385,4.818052,6.498462,10.243283,9.238976,6.4295387,3.9154875,2.9702566,4.466872,6.813539,7.719385,6.931693,6.242462,6.9152827,5.149539,4.824616,7.125334,10.535385,9.580308,6.7872825,3.5938463,1.1552821,0.3446154,0.5021539,0.75487185,0.9419488,1.3554872,2.7634873,7.2336416,8.14277,5.658257,2.281026,2.8521028,2.6289232,2.7109745,3.062154,3.8990772,5.677949,7.653744,8.470975,8.379078,7.965539,8.146052,8.592411,9.288206,7.962257,5.2644105,4.788513,2.9243078,1.8740515,1.4080001,1.522872,2.4320002,2.4582565,3.7448208,3.876103,2.5961027,1.7985642,2.7044106,2.8422565,2.028308,0.8533334,0.7187693,0.49887183,0.85005134,1.0601027,1.332513,2.789744,3.8531284,5.85518,7.240206,6.806975,3.7316926,1.8379488,1.3915899,1.8149745,2.3040001,1.8248206,0.9156924,0.6268718,0.761436,1.1946667,1.8773335,1.1323078,0.8960001,1.2635899,1.972513,2.412308,2.7076926,2.3630772,1.8510771,1.2274873,0.15425642,0.18707694,0.098461546,0.03938462,0.032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.006564103,0.0032820515,0.016410258,0.026256412,0.01969231,0.009846155,0.009846155,0.04266667,0.04266667,0.059076928,0.08205129,0.128,0.23302566,0.21661541,0.16410258,0.11158975,0.072205134,0.029538464,0.13784617,0.15753847,0.108307704,0.03938462,0.006564103,0.15425642,0.20020515,0.3249231,0.47589746,0.36758977,0.29538465,0.6859488,0.7220513,0.2986667,0.02297436,0.006564103,0.0,0.0,0.0,0.0,0.0032820515,0.02297436,0.049230773,0.08205129,0.10502565,0.15425642,0.20020515,0.22646156,0.2297436,0.21333335,0.27569234,0.3052308,0.37743592,0.46933338,0.446359,0.2855385,0.27569234,0.32164106,0.3708718,0.39384618,0.48246157,0.54482055,0.5284103,0.52512825,0.7778462,1.3128207,1.6640002,1.9692309,2.3466668,2.878359,4.588308,6.1078978,7.50277,8.237949,7.174565,5.4843082,5.0182567,5.0642056,4.9821544,4.2141542,3.4297438,3.259077,3.5282054,3.9417439,4.066462,3.882667,3.3542566,3.0720003,3.1081028,3.0129232,2.5435898,2.3204105,2.1431797,1.9528207,1.8346668,1.9003079,1.5622566,1.273436,1.2274873,1.3522053,1.1355898,0.97805136,0.8960001,0.8960001,0.97805136,1.0338463,0.8730257,0.88615394,1.0404103,0.8960001,0.99774367,1.0404103,1.2537436,1.595077,1.7329233,1.847795,1.8543591,2.3630772,3.3312824,4.0533338,3.2820516,3.5610259,3.9089234,3.9581542,3.95159,4.8082056,4.9854364,5.1626673,5.609026,6.189949,7.3682055,7.0432825,6.452513,6.0291286,5.4186673,4.781949,4.1714873,3.82359,3.6824617,3.4034874,2.428718,2.228513,2.2219489,2.0873847,1.7690258,1.4703591,1.3981539,1.8838975,2.6322052,2.7273848,2.353231,2.0939488,2.041436,2.1398976,2.172718,2.4057438,2.5796926,2.6945643,2.5074873,1.5458462,1.522872,1.6246156,1.6672822,1.5786668,1.4080001,1.3587693,1.4572309,1.5195899,1.4966155,1.4736412,1.2603078,1.3128207,1.3784616,1.3587693,1.3095386,1.2471796,1.2209232,1.2898463,1.3686155,1.2471796,1.2340513,1.024,0.76800007,0.5546667,0.41682056,0.33476925,0.39712822,0.53825647,0.764718,1.1388719,2.1924105,3.0785644,3.698872,4.1156926,4.522667,5.024821,6.11118,7.3353853,8.717129,10.761847,11.260718,11.858052,12.140308,12.150155,12.3995905,12.461949,12.580104,13.548308,15.113848,15.980309,16.183796,16.712206,17.263592,17.368616,16.377438,16.406975,17.348925,16.971489,16.003283,18.133335,16.52513,16.613745,15.947489,14.608412,15.202463,14.972719,14.447591,13.791181,12.87877,11.306667,11.434668,12.373334,13.069129,13.292309,13.610668,13.840411,13.814155,13.377642,12.970668,13.627078,13.718975,14.017642,14.483693,14.995693,15.350155,15.051488,14.900514,15.356719,16.512001,18.087385,20.187899,20.923079,20.634258,19.561028,17.83795,16.321642,15.465027,15.392821,15.747283,15.701335,14.811898,13.558155,12.2387705,11.270565,11.168821,10.66995,9.862565,9.337437,9.32759,9.705027,10.180923,10.266257,10.512411,11.040821,11.523283,11.185231,11.621744,11.82195,11.59877,11.579078,11.864616,11.510155,10.794667,10.220308,10.515693,10.361437,10.322052,9.911796,9.229129,8.969847,8.041026,7.318975,6.931693,6.9152827,7.2369237,7.3386674,7.328821,7.460103,7.962257,9.051898,9.826463,9.96759,9.501539,8.54318,7.3025646,6.813539,6.744616,6.5017443,5.98318,5.5696416,5.474462,5.366154,4.9526157,4.273231,3.7021542,3.564308,3.9384618,4.348718,4.709744,5.3037953,6.0849237,6.6592827,6.885744,6.961231,7.4010262,1.9462565,2.0020514,2.176,2.1792822,2.0184617,1.9954873,1.9167181,1.8838975,1.9003079,1.9331284,1.9167181,1.8182565,1.9003079,2.0184617,2.0578463,1.9265642,2.294154,2.556718,2.9636924,3.4855387,3.8104618,3.9909747,4.598154,5.297231,5.901129,6.3442054,6.7938466,7.0104623,6.678975,5.9569235,5.474462,5.3202057,5.533539,5.651693,5.733744,6.3343596,6.2555904,5.179077,4.1682053,3.7021542,3.6594875,3.239385,2.7273848,2.1103592,1.5556924,1.404718,1.1355898,1.2373334,1.463795,1.6147693,1.5425643,1.8313848,1.8281027,1.7362052,1.654154,1.5721027,1.5130258,1.5491283,1.6705642,1.8116925,1.8674873,2.028308,2.0939488,1.8937438,1.5327181,1.3751796,1.3883078,1.7132308,1.9987694,2.156308,2.353231,2.3860514,2.0118976,1.3620514,0.72861546,0.56123084,0.6170257,0.49887183,0.4135385,0.41025645,0.35446155,0.29538465,0.28882053,0.3511795,0.46933338,0.5940513,0.7417436,0.7975385,0.8336411,0.90256417,1.0371283,0.9944616,1.0633847,1.1946667,1.3620514,1.5491283,1.8084104,2.8127182,4.397949,6.193231,7.6176414,9.494975,11.132719,12.901745,14.762668,16.246155,16.922258,18.002052,19.410053,20.890259,22.01272,24.923899,26.745438,26.824207,25.491693,24.047592,22.967796,22.166977,21.06749,19.80718,19.206566,20.62113,20.690052,20.168207,19.321438,17.942976,16.718771,16.144411,16.22318,16.787693,17.503181,17.900309,18.146463,17.828104,17.14872,16.938667,17.920002,17.152,15.415796,13.5318985,12.370052,12.540719,13.193847,13.371078,13.495796,15.353437,15.504412,16.183796,17.667284,18.819284,17.089642,14.690463,12.360206,11.716924,12.547283,12.800001,13.541744,14.614976,15.963899,17.637745,19.784206,21.513847,21.471182,21.733746,23.424002,26.722464,30.319592,34.92431,37.38257,36.998566,35.544617,33.257027,32.705643,33.119183,34.569847,37.98318,41.27508,45.4039,49.486774,53.044518,55.998363,51.564312,44.658875,39.043285,36.542362,37.034668,37.90441,37.428516,36.90339,36.90667,37.32349,38.948105,39.59795,38.95795,37.218464,35.062157,31.878567,29.61395,28.481644,29.101952,32.502155,37.753437,40.277336,37.284107,29.958567,23.450258,21.48431,20.867283,20.473438,19.866259,19.311592,17.621334,17.463797,18.582975,20.854155,24.270771,25.659079,25.685335,26.04308,26.932514,27.053951,23.88349,22.249027,22.974361,25.350567,27.126156,28.163284,28.15672,26.131695,22.550976,19.324718,16.305231,18.704412,21.028105,21.041233,19.767796,21.044514,19.777643,18.271181,18.176,20.476719,18.855387,14.096412,13.380924,16.278976,14.739694,11.090053,7.6898465,4.6933336,2.7011285,2.7700515,2.7470772,4.588308,5.654975,5.5171285,5.9634876,3.8728209,5.179077,7.1909747,9.498257,13.952001,10.601027,5.874872,3.7152824,5.5171285,10.125129,9.95118,7.515898,4.6867695,2.8160002,2.7306669,5.1265645,8.214975,9.133949,7.7259493,6.5378466,9.593436,7.7325134,6.1440005,7.3091288,11.0145645,9.990565,6.87918,3.8006158,1.8018463,0.8467693,0.58420515,0.81394875,3.7842054,6.6395903,1.4211283,4.2338467,6.8496413,6.7085133,4.2207184,2.802872,2.294154,2.1924105,2.5304618,3.2623591,4.2568207,5.7468724,6.948103,7.5421543,7.643898,7.77518,7.8834877,7.939283,6.948103,5.293949,4.7327185,3.249231,2.2580514,1.6672822,1.5425643,2.0873847,2.2088206,3.8596926,5.139693,5.041231,3.442872,2.231795,2.5304618,2.7700515,2.484513,2.3204105,2.1398976,1.5885129,1.2668719,1.4112822,1.8707694,3.2656412,4.7491283,4.7392826,3.2722054,2.0151796,1.7887181,1.3718976,1.3161026,1.4867693,1.0371283,0.8598975,0.86974365,1.2176411,1.6640002,1.5983591,1.148718,0.7975385,0.6432821,0.77128214,1.2865642,1.782154,1.5064616,1.3883078,1.3128207,0.14441027,0.2986667,0.19364104,0.06564103,0.013128206,0.009846155,0.009846155,0.009846155,0.009846155,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.026256412,0.02297436,0.029538464,0.026256412,0.013128206,0.006564103,0.036102567,0.059076928,0.072205134,0.08205129,0.12471796,0.24943592,0.3052308,0.23630771,0.15425642,0.10502565,0.049230773,0.032820515,0.049230773,0.049230773,0.026256412,0.009846155,0.118153855,0.072205134,0.02297436,0.02297436,0.01969231,0.049230773,0.118153855,0.11158975,0.036102567,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.029538464,0.06564103,0.09189744,0.118153855,0.16082053,0.21989745,0.26256412,0.23302566,0.24287182,0.24943592,0.3117949,0.4135385,0.45292312,0.39056414,0.3314872,0.2855385,0.26256412,0.25928208,0.2986667,0.41025645,0.51856416,0.58420515,0.62030774,0.97805136,1.3587693,1.7985642,2.2711797,2.681436,3.8990772,5.1889234,6.377026,7.1680007,7.1483083,5.907693,5.1331286,4.6802053,4.460308,4.4406157,3.9745643,3.5446157,3.5282054,3.8367183,3.892513,3.9187696,3.5741541,3.1671798,2.878359,2.7634873,2.0841026,1.723077,1.6180514,1.6672822,1.7165129,1.6607181,1.4441026,1.332513,1.3751796,1.4112822,1.0896411,0.88615394,0.8008206,0.7778462,0.69907695,0.78769237,0.78769237,0.86646163,0.96492314,0.80738467,0.97805136,1.2406155,1.4145643,1.4933335,1.6475899,1.9495386,1.9298463,2.3040001,3.0391798,3.3378465,3.0687182,3.5249233,4.023795,4.1911798,3.9909747,4.414359,5.1626673,5.8420515,6.265436,6.4754877,7.0334363,6.803693,6.3573337,5.858462,5.028103,4.194462,3.3444104,2.9636924,3.0884104,3.2886157,2.3827693,1.9889232,1.785436,1.6114873,1.463795,1.6278975,1.7427694,1.9232821,2.0578463,1.8116925,2.0086155,2.0709746,1.9823592,1.9167181,2.2186668,2.3269746,2.537026,2.5435898,2.2055387,1.522872,1.5163078,1.3423591,1.2964103,1.404718,1.4473847,1.5622566,1.585231,1.4998976,1.394872,1.463795,1.3587693,1.2931283,1.2603078,1.2471796,1.2373334,1.1815386,1.1684103,1.1716924,1.1520001,1.024,0.9124103,0.67938465,0.48246157,0.36430773,0.25271797,0.25928208,0.48246157,0.69251287,0.9747693,1.7165129,2.4155898,2.7831798,3.2722054,3.9417439,4.460308,5.35959,6.550975,7.50277,8.372514,9.993847,10.791386,11.227899,11.477334,11.684103,11.956513,11.835078,12.130463,13.29559,14.9398985,15.826053,15.875283,15.455181,15.852309,16.640001,15.684924,16.38072,17.188105,17.129026,16.57436,17.26031,16.026258,15.675078,15.00554,14.057027,14.093129,14.358975,14.050463,13.833847,13.46954,11.812103,11.21477,11.32636,11.585642,11.976206,13.049437,13.512206,13.558155,13.302155,13.10195,13.561437,13.489232,13.29559,13.53518,14.257232,15.0088215,15.37313,15.704617,16.456207,17.621334,18.73395,20.273232,20.693335,20.299488,19.331284,17.962667,16.66954,15.921232,15.812924,16.07877,16.072206,14.49354,13.239796,12.370052,11.900719,11.828514,11.1064625,10.187488,9.317744,8.730257,8.674462,9.596719,10.056206,10.722463,11.625027,12.150155,11.493745,11.592206,11.785847,11.766154,11.569232,11.657847,11.313231,10.84718,10.689642,11.401847,10.932513,10.262975,9.442462,8.628513,8.090257,7.128616,6.738052,6.741334,6.928411,7.059693,7.4108725,7.6570263,7.8112826,8.073847,8.832001,9.494975,9.051898,8.4512825,8.070564,7.719385,7.765334,7.532308,7.0104623,6.3376417,5.8157954,5.6418467,5.4416413,4.9526157,4.2141542,3.5840003,3.4625645,4.023795,4.7425647,5.32677,5.7074876,6.1308722,6.5903597,6.672411,6.5706673,7.072821,2.300718,2.0742567,2.28759,2.412308,2.294154,2.15959,1.9265642,2.0118976,2.169436,2.2350771,2.1300514,1.9692309,1.8970258,1.9298463,2.0250258,2.0775387,2.2646155,2.3958976,2.7634873,3.314872,3.6529233,3.9318976,4.5062566,4.9952826,5.398975,6.1078978,6.554257,6.7905645,6.5411286,5.87159,5.182359,5.0149746,5.2676926,5.4908724,5.7009234,6.373744,7.2205133,6.2916927,5.0871797,4.3618464,4.1222568,3.370667,2.6683078,2.0053334,1.4408206,1.0994873,0.9419488,1.2209232,1.5885129,1.8149745,1.785436,1.8116925,1.8642052,1.9167181,1.9626669,2.0118976,1.910154,1.7920002,1.8379488,1.9856411,1.9396925,1.8051283,1.6443079,1.4375386,1.2537436,1.2471796,1.3128207,1.5261539,1.723077,1.8412309,1.913436,1.5556924,1.2570257,0.9944616,0.8008206,0.7515898,0.7253334,0.61374366,0.5874872,0.62030774,0.4955898,0.33476925,0.2986667,0.38728207,0.56451285,0.7975385,1.0601027,1.1290257,1.1355898,1.1716924,1.276718,1.1815386,1.276718,1.4473847,1.6311796,1.8248206,2.231795,3.0358977,4.2207184,5.7731285,7.6898465,10.427077,12.347078,14.532925,17.237335,19.88595,19.48554,19.334566,20.230566,22.01272,23.538874,24.946875,25.124104,24.064001,22.28513,20.83118,19.889233,18.95713,17.450668,15.740719,15.133539,16.436514,18.12677,19.301744,19.088411,16.662975,15.58318,15.786668,17.017437,18.648617,19.698874,21.225027,22.311386,22.377028,21.474463,20.296207,19.958155,18.520617,16.78113,15.468308,15.248411,16.292105,16.820515,17.335796,17.972515,18.471386,18.320412,18.12349,18.340103,18.7799,18.57313,17.611488,15.356719,13.4170265,12.3306675,11.585642,11.008,11.37559,12.540719,14.332719,16.554668,17.834667,18.54359,19.551182,21.504002,24.854977,29.824003,34.356514,36.545643,35.741543,32.548103,29.850258,29.177439,29.167591,29.942156,33.112617,35.682465,39.000618,43.982773,51.101543,60.370056,60.609646,52.972313,43.109745,35.744823,34.674873,35.410053,34.592823,33.857643,33.86749,34.32041,35.62995,36.33231,36.115696,35.00308,33.345642,31.222157,30.102976,29.384207,29.558157,32.20677,37.3399,41.271797,39.83754,33.155285,25.639387,22.265438,20.516104,19.538054,18.980104,18.986668,17.920002,17.847795,19.232822,22.344208,27.280413,30.493542,31.360003,32.479183,34.070976,33.942978,28.150156,25.330873,25.560617,27.959797,30.723284,32.610462,32.262566,28.022156,21.605745,18.116924,15.179488,16.46277,18.274464,18.464823,16.452925,17.408,17.739489,18.06113,18.924309,20.808207,17.076513,11.460924,9.42277,11.474052,13.184001,13.568001,10.699488,6.439385,2.9505644,2.6847181,2.9440002,5.152821,6.5444107,6.449231,6.2818465,3.7940516,3.8498464,5.6385646,8.43159,11.602052,9.432616,5.3858466,4.1517954,6.889026,11.211488,8.441437,5.549949,3.2984617,2.3269746,3.1474874,5.0477953,8.484103,9.947898,8.487385,5.7140517,12.2617445,9.997129,6.7150774,6.1505647,7.968821,8.086975,6.0356927,3.9187696,2.5731285,1.5425643,0.7811283,0.77456415,5.07077,9.3078985,1.1946667,2.03159,4.1156926,5.4547696,5.080616,3.0654361,2.3663592,2.0808206,2.477949,3.3542566,4.020513,4.4406157,5.799385,6.8693337,7.0925136,6.5870776,6.416411,5.8518977,5.0543594,4.2502565,3.7316926,3.006359,2.294154,1.6836925,1.3029745,1.3292309,1.7165129,2.8750772,4.673641,6.166975,5.602462,3.501949,2.993231,3.0752823,3.3017437,3.7842054,3.7316926,2.6223593,1.910154,2.166154,3.0851285,5.2742567,5.3825645,3.692308,1.5491283,1.3686155,2.0217438,1.5885129,1.2865642,1.5458462,1.9954873,1.5261539,1.2832822,1.4473847,1.7165129,1.2996924,1.2438976,1.4244103,1.204513,0.6629744,0.5874872,0.9911796,0.79425645,0.7253334,0.8041026,0.3314872,0.3249231,0.19364104,0.072205134,0.016410258,0.009846155,0.02297436,0.026256412,0.029538464,0.029538464,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.006564103,0.0032820515,0.026256412,0.059076928,0.036102567,0.036102567,0.03938462,0.029538464,0.013128206,0.036102567,0.068923086,0.072205134,0.07548718,0.11158975,0.21989745,0.2986667,0.25271797,0.19692309,0.15425642,0.072205134,0.02297436,0.01969231,0.029538464,0.036102567,0.06564103,0.3314872,0.67282057,0.79097444,0.5874872,0.15753847,0.052512825,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.04266667,0.08533334,0.101743594,0.14112821,0.21333335,0.27569234,0.22646156,0.23630771,0.23302566,0.26584616,0.3314872,0.40369233,0.44307697,0.36758977,0.27241027,0.23630771,0.29538465,0.3052308,0.380718,0.48902568,0.5546667,0.48574364,0.7450257,1.1881026,1.7033848,2.2449234,2.8225644,3.7021542,4.7983594,5.7435904,6.314667,6.432821,6.186667,5.435077,4.768821,4.565334,4.9887185,4.8147697,4.2535386,3.9122055,3.8990772,3.826872,3.9253337,3.757949,3.308308,2.737231,2.3663592,1.8510771,1.4539489,1.3292309,1.4244103,1.4966155,1.4309745,1.4309745,1.4506668,1.4342566,1.3193847,1.0272821,0.827077,0.7450257,0.7089231,0.5284103,0.6498462,0.7581539,0.8172308,0.8205129,0.8041026,1.0075898,1.3751796,1.5064616,1.4572309,1.7394873,1.9692309,2.1103592,2.4516926,2.7798977,2.3696413,2.7470772,3.1803079,3.5478978,3.8498464,4.204308,4.1058464,4.8771286,5.717334,6.114462,5.865026,6.2916927,6.1440005,5.865026,5.4482055,4.457026,3.7120004,2.9669745,2.6157951,2.7634873,3.2295387,2.3204105,1.7755898,1.4408206,1.2537436,1.2406155,1.5064616,1.5556924,1.5360001,1.4933335,1.3981539,1.910154,2.100513,1.9889232,1.9331284,2.6289232,2.8324106,2.8816411,2.7109745,2.3138463,1.7296412,1.6311796,1.2668719,1.1651284,1.3620514,1.404718,1.5491283,1.4802053,1.3784616,1.3653334,1.4834872,1.3817437,1.270154,1.211077,1.204513,1.1684103,1.1093334,1.0535386,0.97805136,0.86317956,0.7089231,0.56123084,0.4266667,0.3249231,0.256,0.18707694,0.41682056,0.71548724,0.95835906,1.2603078,1.9429746,2.2186668,2.3040001,2.7569232,3.5741541,4.1813335,5.356308,6.449231,7.210667,7.788308,8.736821,9.875693,10.482873,10.9226675,11.411694,12.012309,11.644719,11.992617,12.947693,14.129231,14.874257,15.655386,15.225437,15.461744,16.393847,16.210052,16.853334,17.06995,16.971489,16.613745,15.996719,15.002257,14.309745,13.620514,12.987078,12.829539,13.883078,13.722258,13.581129,13.39077,11.782565,10.473026,10.115283,10.43036,11.260718,12.603078,13.197129,13.479385,13.499078,13.51877,14.01436,13.748514,13.380924,13.5548725,14.296617,14.995693,15.894976,16.420103,17.263592,18.356514,18.868515,19.570873,19.656206,19.334566,18.642054,17.424412,16.485744,16.06236,16.085335,16.226463,15.90154,14.329437,13.430155,12.931283,12.570257,12.114052,11.152411,10.272821,9.347282,8.55959,8.411898,9.465437,10.128411,10.916103,11.825232,12.363488,11.835078,11.595488,11.680821,11.782565,11.241027,11.244308,11.221334,11.21477,11.388719,12.035283,11.533129,10.44677,9.324308,8.379078,7.4797955,6.9809237,6.8266673,6.9677954,7.204103,7.181129,7.702975,8.100103,8.155898,8.001641,8.093539,8.612103,8.152616,7.8047185,7.939283,8.211693,8.513641,8.027898,7.204103,6.4623594,6.157129,5.7009234,5.159385,4.5456414,3.9942567,3.7415388,3.7940516,4.322462,5.0182567,5.612308,5.8912826,6.121026,6.449231,6.47877,6.409847,7.02359,2.6978464,2.4188719,2.5009232,2.5895386,2.5074873,2.2514873,2.048,2.1398976,2.3204105,2.409026,2.225231,1.913436,1.7362052,1.7558975,1.9528207,2.2383592,2.2711797,2.3893335,2.7733335,3.2853336,3.4691284,3.8859491,4.2207184,4.5554876,5.037949,5.8847184,6.2851286,6.678975,6.636308,6.048821,5.152821,4.854154,4.9099493,5.077334,5.290667,5.648411,7.076103,6.7282057,5.7435904,4.650667,3.3641028,2.2777438,1.5721027,1.1979488,1.0108719,0.761436,0.8566154,1.2077949,1.5655385,1.8018463,1.8970258,1.8806155,1.972513,2.0939488,2.2153847,2.3302567,2.3827693,2.1825643,2.176,2.3105643,2.0644104,1.5786668,1.1782565,1.1158975,1.3292309,1.4145643,1.3587693,1.4998976,1.6804104,1.7558975,1.5885129,1.2176411,1.0272821,1.0043077,1.0666667,1.0732309,0.7778462,0.67938465,0.761436,0.86974365,0.69251287,0.39712822,0.31507695,0.36430773,0.51856416,0.78769237,1.079795,1.2537436,1.3292309,1.3357949,1.2865642,1.3718976,1.591795,1.8510771,2.1169233,2.4024618,3.0720003,3.95159,5.041231,6.4754877,8.516924,10.850462,12.960821,15.537232,18.645334,21.733746,20.775387,19.61354,19.938463,21.891283,24.080412,24.146053,23.722668,21.753437,18.95713,17.824821,17.765745,17.401438,16.472616,15.356719,15.081027,16.459488,19.173744,21.142977,20.90995,17.654156,16.955078,17.368616,19.131079,21.395695,22.232616,23.995079,24.690874,24.618668,23.716105,21.559797,20.289642,19.111385,18.28431,18.087385,18.809437,19.810463,19.879387,20.5719,21.471182,20.207592,18.422155,17.660719,17.394873,17.58195,18.70113,18.225233,16.571077,14.749539,13.092104,11.264001,10.584617,10.456616,10.840616,11.700514,13.003489,14.296617,16.154257,17.985641,19.672617,21.563078,26.850464,30.585438,32.800823,33.024002,30.260515,28.074669,27.346054,27.19836,27.746464,30.083284,32.05908,33.332516,36.519386,43.96308,57.73785,68.164925,64.81067,52.56862,38.81026,33.362053,33.043694,32.42667,31.671797,31.090874,31.16308,32.137848,32.90585,33.201233,32.850056,31.760412,30.628105,30.296618,30.106258,30.46072,32.8238,36.837746,41.96431,43.01457,38.33108,29.794464,23.607798,20.397951,19.085129,18.753643,18.635489,17.578669,17.401438,19.419899,23.67672,28.947695,34.12349,36.995285,39.36821,40.772926,38.47549,30.998978,28.278156,28.78031,31.369848,35.29518,37.0839,34.46154,27.470772,19.30831,16.33477,14.884104,14.880821,17.066668,18.953848,14.831591,13.617231,15.258258,17.411283,18.645334,18.435284,12.504617,9.202872,8.093539,8.812308,11.076924,16.164104,14.700309,9.255385,3.5413337,2.3958976,2.989949,5.1298466,6.6133337,6.6822567,6.0061545,3.5807183,2.7667694,3.9548721,6.6002054,9.235693,7.3419495,4.263385,3.8728209,6.262154,7.7292314,6.0225644,4.069744,2.6420515,2.5074873,4.417641,5.2578464,8.283898,10.729027,10.174359,4.565334,11.805539,9.32759,5.8190775,4.634257,3.7842054,5.028103,4.8705645,4.2174363,3.4297438,2.3105643,1.1355898,0.8763078,3.69559,6.675693,1.8149745,1.4342566,1.6410258,3.0523078,4.601436,3.5380516,2.6354873,2.2777438,2.8521028,4.0041027,4.644103,4.844308,6.11118,7.0137444,6.7610264,5.208616,4.9132314,4.4767184,4.0303593,3.570872,2.9669745,2.5731285,2.097231,1.5130258,0.9747693,0.81066674,1.204513,1.4736412,2.6289232,4.6211286,6.3474874,5.0576415,3.5478978,2.5074873,2.428718,3.626667,3.7316926,2.7208207,2.5173335,3.4264617,4.138667,6.6527185,6.117744,4.138667,2.228513,1.8051283,2.300718,1.8379488,1.467077,1.8871796,3.43959,2.176,1.5195899,1.3554872,1.4145643,1.276718,1.3193847,2.100513,1.9823592,0.9714873,0.7220513,0.94523084,0.5349744,0.19692309,0.23302566,0.55794877,0.24943592,0.098461546,0.04594872,0.032820515,0.0,0.032820515,0.04266667,0.052512825,0.052512825,0.01969231,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.016410258,0.006564103,0.032820515,0.07548718,0.055794876,0.059076928,0.06564103,0.052512825,0.032820515,0.055794876,0.072205134,0.072205134,0.072205134,0.09189744,0.128,0.2100513,0.24287182,0.23958977,0.20020515,0.0951795,0.02297436,0.006564103,0.01969231,0.068923086,0.19692309,0.6662565,1.657436,2.2547693,1.9396925,0.6071795,0.18051283,0.03938462,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.02297436,0.072205134,0.0951795,0.14769232,0.21661541,0.25271797,0.190359,0.24943592,0.256,0.25928208,0.27569234,0.32164106,0.4004103,0.3511795,0.27241027,0.26584616,0.41682056,0.47261542,0.45620516,0.44964105,0.4594872,0.42994875,0.69907695,1.2340513,1.6771283,2.0578463,2.7864618,3.7054362,4.598154,5.228308,5.3694363,4.827898,5.661539,5.4153852,5.0674877,5.080616,5.3891287,5.362872,4.857436,4.345436,4.023795,3.8071797,3.8498464,3.7415388,3.2853336,2.556718,1.8937438,1.7427694,1.4276924,1.2406155,1.2406155,1.2504616,1.3554872,1.4933335,1.4834872,1.3161026,1.1323078,0.9714873,0.81394875,0.764718,0.79097444,0.72861546,0.84348726,0.88287187,0.8402052,0.79097444,0.892718,1.0502565,1.3456411,1.4834872,1.5425643,1.972513,2.0611284,2.3630772,2.6945643,2.7011285,1.8510771,2.4385643,2.793026,2.986667,3.314872,4.2863593,4.092718,4.46359,4.9887185,5.2053337,4.630975,5.605744,5.654975,5.398975,4.8607183,3.4691284,3.2754874,2.9801028,2.7766156,2.802872,3.131077,2.228513,1.7427694,1.5622566,1.5556924,1.5819489,1.3357949,1.0010257,0.90912825,1.1848207,1.7493335,2.2580514,2.2744617,2.1431797,2.3072822,3.3247182,3.7218463,3.446154,3.0851285,2.737231,2.0151796,1.6902566,1.273436,1.204513,1.4080001,1.2931283,1.2964103,1.148718,1.2438976,1.5524104,1.6180514,1.3095386,1.1585642,1.1323078,1.1520001,1.1126155,1.0371283,0.90256417,0.7384616,0.58420515,0.47261542,0.380718,0.3249231,0.27569234,0.23302566,0.24287182,0.69251287,0.93866676,1.2274873,1.5753847,1.785436,1.7788719,1.9232821,2.3958976,3.1573336,3.9581542,5.041231,5.805949,6.5280004,7.273026,7.90318,8.966565,9.714872,10.463181,11.362462,12.409437,11.69395,11.657847,12.041847,12.609642,13.124924,14.923489,15.271386,15.543797,16.341335,17.503181,17.11918,16.745028,16.331488,15.721026,14.65436,13.53518,12.796719,12.189539,11.795693,12.012309,13.272616,13.095386,12.672001,12.212514,10.955488,9.770667,9.639385,10.354873,11.477334,12.3306675,12.950975,13.466257,13.748514,13.899488,14.27036,13.945437,13.778052,13.98154,14.480412,14.907078,16.311796,16.89272,17.61477,18.477951,18.507488,18.41559,18.153027,17.962667,17.608206,16.374155,15.826053,15.885129,16.147694,16.134565,15.274668,14.332719,13.850258,13.436719,12.849232,11.976206,10.929232,10.243283,9.580308,9.012513,9.045334,9.819899,10.450052,11.0145645,11.588924,12.242052,12.07795,11.513436,11.395283,11.569232,10.902975,10.788103,11.191795,11.703795,12.117334,12.432411,11.995898,10.889847,9.714872,8.65477,7.456821,7.53559,7.3583593,7.3682055,7.6209235,7.781744,8.15918,8.329846,8.1066675,7.5487185,6.9842057,7.496206,7.5913854,7.716103,8.024616,8.395488,8.674462,7.9819493,6.997334,6.2818465,6.2687182,5.61559,4.841026,4.204308,3.945026,4.263385,4.535795,4.824616,5.146257,5.481026,5.7764106,6.1472826,6.514872,6.626462,6.6428723,7.13518,2.0151796,2.2350771,2.3893335,2.4615386,2.3991797,2.1070771,2.2646155,2.2777438,2.15959,1.9922053,1.9068719,1.6640002,1.585231,1.6804104,1.847795,1.847795,1.8215386,2.034872,2.4451284,2.9210258,3.249231,3.7152824,3.9942567,4.3716927,4.9427695,5.61559,6.0685134,6.5837955,6.5017443,5.7632823,4.896821,4.716308,4.844308,4.9788723,4.965744,4.8082056,5.796103,6.0619493,5.5302567,4.1452312,1.8609232,1.0305642,0.76800007,0.7318975,0.761436,0.86974365,1.1520001,1.394872,1.6082052,1.7624617,1.8018463,1.8116925,1.7788719,1.9790771,2.2711797,2.0742567,2.3302567,2.2482052,2.1825643,2.1956925,2.0742567,1.6114873,1.404718,1.3686155,1.4145643,1.463795,1.1848207,1.7001027,1.7985642,1.2832822,0.97805136,0.79425645,0.764718,0.81394875,0.9288206,1.1585642,0.7581539,0.636718,0.5874872,0.5349744,0.5349744,0.5218462,0.508718,0.49887183,0.51856416,0.64000005,0.78769237,1.1355898,1.3718976,1.3718976,1.1913847,1.7624617,2.228513,2.7766156,3.3903592,3.8301542,4.8804107,6.0750775,7.325539,8.687591,10.361437,12.314258,13.8075905,16.65313,19.866259,19.682463,19.232822,19.275488,19.64636,20.821335,23.909746,22.81354,21.586054,19.088411,16.042667,15.028514,16.384,16.640001,16.390566,16.022976,15.717745,18.218668,21.937233,24.697437,24.625233,20.155079,18.947283,18.113642,18.993233,20.841026,20.8279,20.46359,21.717335,21.625437,20.096,19.912207,19.8039,20.709745,21.270975,21.018257,20.371695,20.457027,21.18236,21.651693,21.369438,20.233849,17.060104,15.212309,15.849027,18.287592,20.020514,18.323694,17.440823,16.580925,15.048206,12.251899,10.811078,11.139283,11.372309,11.293539,12.343796,14.372104,16.059078,17.54913,18.635489,18.770052,22.002874,25.504822,28.14031,29.577848,30.273643,29.24636,28.048412,27.414976,27.716925,28.960823,27.9959,29.348104,31.704618,36.388103,47.35016,64.7319,73.87241,68.09272,50.7799,35.400208,32.0919,30.424618,29.45313,29.06585,29.968412,29.42031,29.144617,29.669746,30.575592,30.503387,29.817438,29.922464,30.58872,32.055798,35.03262,36.01067,41.3079,46.339287,46.286774,36.115696,26.423798,21.648413,19.659489,18.914463,18.46154,17.877335,18.159592,20.187899,23.955694,28.596516,34.392616,39.230362,42.624004,43.05395,37.96349,32.3118,31.69477,33.58195,36.273235,38.908722,37.251286,29.620516,21.766565,16.600616,14.221129,14.01436,16.15754,20.194464,22.130873,14.464001,10.253129,11.372309,14.155488,15.714462,13.932309,8.254359,9.856001,9.235693,5.671385,7.2336416,15.727591,17.752617,13.459693,6.2785645,2.8849232,3.1277952,4.378257,5.4547696,5.687795,4.9427695,3.0260515,2.3105643,2.4320002,4.571898,11.444513,7.7948723,4.069744,2.6551797,3.3608208,3.4330258,3.495385,2.9801028,2.2646155,2.5271797,5.737026,6.665847,8.454565,12.071385,13.952001,5.979898,6.298257,4.125539,3.0884104,3.5282054,2.5009232,1.8806155,3.190154,4.453744,4.5554876,3.249231,1.7723079,1.5688206,1.8674873,2.2449234,2.609231,2.3171284,1.7394873,2.740513,4.5029745,3.5249233,2.487795,2.228513,3.0884104,4.1550775,3.2656412,6.0717955,6.7840004,7.145026,7.003898,4.31918,3.6594875,3.4855387,3.8400004,4.076308,2.868513,2.4648206,2.0808206,1.5327181,0.88615394,0.45620516,0.90912825,1.0666667,1.1290257,1.5031796,2.809436,4.309334,2.678154,1.1355898,0.8533334,0.97805136,1.3686155,1.8773335,4.325744,7.128616,5.3103595,3.9680004,5.58277,5.0871797,2.5271797,3.0523078,1.7690258,1.394872,1.3686155,1.3653334,1.2668719,0.75487185,0.9353847,1.1684103,1.142154,0.88615394,0.71548724,0.52512825,0.2986667,0.11158975,0.13784617,0.12471796,0.17723078,0.190359,0.21661541,0.47261542,0.0951795,0.0,0.006564103,0.013128206,0.0,0.013128206,0.032820515,0.052512825,0.055794876,0.029538464,0.029538464,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.016410258,0.006564103,0.01969231,0.055794876,0.09189744,0.1148718,0.10502565,0.08533334,0.07876924,0.09189744,0.07876924,0.08533334,0.098461546,0.10502565,0.09189744,0.16410258,0.27569234,0.2855385,0.19364104,0.108307704,0.04594872,0.029538464,0.04266667,0.13456412,0.4266667,1.1224617,2.2219489,3.5413337,4.0008206,1.6311796,0.42338464,0.059076928,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.06235898,0.072205134,0.13128206,0.17394873,0.17723078,0.15097436,0.20020515,0.2231795,0.25271797,0.29538465,0.32164106,0.380718,0.3708718,0.29538465,0.23630771,0.32164106,0.5021539,0.42994875,0.38728207,0.45620516,0.5021539,0.6268718,1.270154,1.6344616,1.7132308,2.2744617,3.3476925,4.1550775,4.6145644,4.5587697,3.754667,5.182359,5.5007186,5.4547696,5.4383593,5.5236926,5.4383593,4.969026,4.4373336,4.0402055,3.8465643,3.6627696,3.570872,3.1737437,2.4681027,1.847795,1.6278975,1.3161026,1.083077,0.9944616,1.0075898,1.2865642,1.3587693,1.2668719,1.083077,0.8992821,0.8763078,0.6859488,0.65641034,0.8763078,1.204513,1.1454359,1.0732309,1.0075898,0.955077,0.9321026,0.97805136,1.1388719,1.3883078,1.6902566,1.9823592,2.1924105,2.3269746,2.4155898,2.3893335,2.0611284,2.8914874,3.5446157,3.7349746,3.6758976,4.1058464,4.348718,4.6834874,4.8804107,4.6900516,3.8596926,4.397949,5.0642056,4.8311796,3.4691284,1.5425643,2.2744617,2.428718,2.4976413,2.6551797,2.7766156,2.2153847,1.9200002,2.162872,2.6420515,2.4713848,1.4342566,1.0666667,1.1191796,1.4309745,1.9068719,2.3958976,2.5173335,2.5665643,2.8717952,3.8006158,3.5905645,2.917744,2.550154,2.5764105,2.3794873,1.8445129,1.5983591,1.4966155,1.404718,1.2209232,1.086359,1.0075898,1.463795,2.1300514,1.8609232,1.2504616,1.0633847,1.0666667,1.1126155,1.1126155,0.88287187,0.71548724,0.5546667,0.42338464,0.4135385,0.38728207,0.33476925,0.3249231,0.39056414,0.5481026,0.83035904,0.8467693,1.1126155,1.5524104,1.4802053,1.5425643,1.9331284,2.4385643,3.1638978,4.532513,5.0674877,5.1856413,5.733744,6.8430777,7.90318,8.720411,9.219283,10.049642,11.286975,12.419283,11.493745,10.978462,10.9226675,11.355898,12.2847185,15.067899,15.376411,15.153232,15.622565,17.319386,16.233027,14.907078,14.401642,14.447591,13.459693,12.849232,12.557129,12.064821,11.707078,12.694975,12.501334,11.976206,11.053949,10.174359,10.28595,10.066052,10.184206,10.496001,10.880001,11.244308,12.137027,12.560411,12.964104,13.377642,13.426873,13.121642,13.239796,13.525334,13.906053,14.480412,16.02954,17.08636,17.867489,18.336823,18.202257,17.591797,16.938667,16.594053,16.324924,15.274668,15.419078,15.8884115,16.108309,15.77354,14.8480015,14.54277,13.8075905,13.08554,12.488206,11.779283,10.742155,10.171078,9.77395,9.557334,9.826463,10.180923,10.59118,10.948924,11.339488,12.025436,12.071385,11.270565,11.08677,11.513436,11.063796,10.292514,10.79795,11.74318,12.544001,12.849232,12.176412,11.303386,10.466462,9.494975,7.7981544,7.322257,7.384616,7.752206,8.283898,8.940309,8.674462,7.827693,7.194257,6.889026,6.363898,6.813539,7.210667,7.53559,7.8080006,8.103385,8.224821,7.450257,6.6133337,6.1341543,6.012718,5.4383593,4.900103,4.5095387,4.3716927,4.59159,4.775385,4.7589746,4.7327185,4.9099493,5.5072823,6.3868723,6.918565,7.017026,6.7314878,6.2555904,2.1858463,2.930872,2.3401027,1.8904617,1.9954873,1.9954873,1.8609232,1.7362052,1.7558975,1.9035898,1.9922053,1.8642052,1.7001027,1.782154,1.9987694,1.8215386,1.8838975,2.0906668,2.349949,2.6584618,3.114667,3.892513,4.4406157,4.785231,5.0543594,5.481026,6.1472826,6.8627696,6.9842057,6.363898,5.362872,4.71959,4.97559,5.21518,5.024821,4.4767184,4.4406157,4.8804107,5.1265645,4.457026,2.1070771,1.0108719,0.6104616,0.5152821,0.5546667,0.77128214,0.88615394,1.0962052,1.3653334,1.6114873,1.7165129,1.657436,1.6738462,1.7690258,1.8281027,1.6246156,1.8510771,1.7033848,1.6213335,1.6180514,1.2832822,1.1290257,1.0305642,0.9878975,1.020718,1.148718,1.1191796,1.1520001,1.1716924,1.1388719,1.0371283,1.0601027,1.017436,0.90584624,0.75487185,0.63343596,0.43651286,0.5316923,0.6071795,0.56451285,0.48574364,0.5218462,0.6301539,0.6892308,0.6662565,0.65312827,0.7318975,0.8566154,0.9911796,1.1618463,1.4473847,2.1267693,2.8882053,3.7120004,4.6933336,6.052103,7.3747697,8.822155,10.059488,10.925949,11.434668,12.324103,13.656616,17.08636,20.312616,17.083078,16.584206,16.935387,17.490053,18.560001,21.431797,19.298464,18.471386,17.59836,16.341335,15.396104,16.905848,17.43754,17.542566,17.542566,17.509745,18.566566,20.929642,22.455797,22.088207,19.876104,19.049026,19.43959,20.322464,21.96677,25.626259,20.804924,20.171488,20.151796,19.272207,18.130053,18.392616,19.59713,20.348719,20.25354,19.91877,20.844309,20.969027,20.368412,19.39036,18.645334,15.051488,14.677335,15.701335,16.534975,15.809642,16.39713,16.758156,17.286566,17.14872,14.316309,12.658873,12.501334,12.586668,12.658873,13.456411,14.260514,14.976001,17.115898,19.43959,17.962667,18.074257,19.328001,22.78072,26.63713,26.26954,26.59118,27.283695,29.11836,31.104002,30.473848,29.686155,30.401644,31.616003,34.20554,40.94031,53.27426,66.67816,71.85395,64.748314,46.546055,33.83467,29.298874,27.634874,26.489437,26.466463,26.676516,26.446772,26.942362,28.271591,29.476105,29.282463,29.801027,31.369848,33.736206,36.0599,35.20985,39.663593,48.794262,56.352825,50.47139,35.984413,27.923695,23.561848,20.801643,18.182566,20.388103,20.07631,20.476719,22.839796,26.423798,32.610462,38.176823,41.96103,42.51898,38.12103,36.368412,38.262157,40.218258,39.821133,35.846565,31.382977,24.46113,18.707693,15.123693,12.048411,15.268104,18.865232,19.945026,17.867489,14.244103,10.729027,10.134975,10.404103,9.777231,6.813539,5.7665644,7.427283,7.39118,6.183385,9.258667,15.363283,17.870771,15.353437,9.442462,4.84759,3.9220517,4.3585644,4.7983594,4.8082056,4.893539,3.3214362,2.5140514,2.3663592,3.8367183,8.940309,7.000616,3.9384618,2.1924105,2.359795,3.2131286,3.1081028,3.501949,2.9833848,1.9200002,2.4549747,5.353026,8.493949,11.1064625,11.490462,7.00718,7.6767187,5.277539,3.0523078,2.0676925,1.2077949,0.95835906,1.8740515,3.0358977,3.8038976,3.8367183,2.8389745,2.3138463,2.0808206,2.1234872,2.5961027,2.5764105,2.4713848,3.7087183,5.5663595,5.1856413,5.3103595,4.5062566,5.668103,7.145026,2.7273848,5.0182567,4.670359,4.161641,4.263385,4.0369234,3.9942567,4.125539,4.164923,3.9089234,3.245949,2.9111798,2.3269746,1.6147693,0.97805136,0.67610264,0.9517949,1.4276924,1.5524104,1.4276924,1.8051283,1.8248206,1.404718,2.3204105,3.4231799,0.63343596,0.88943595,1.6804104,2.7602053,3.636513,3.564308,3.1967182,3.3509746,2.553436,1.1224617,1.1585642,0.78769237,0.67610264,0.8205129,1.0404103,0.9747693,0.8795898,0.92553854,1.1060513,1.3357949,1.4572309,1.2964103,0.76800007,0.36102566,0.2231795,0.15097436,0.108307704,0.101743594,0.14441027,0.20020515,0.19364104,0.049230773,0.013128206,0.009846155,0.0032820515,0.0,0.02297436,0.02297436,0.026256412,0.032820515,0.01969231,0.06564103,0.032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.02297436,0.032820515,0.068923086,0.1148718,0.10502565,0.098461546,0.072205134,0.059076928,0.06564103,0.07876924,0.07548718,0.072205134,0.059076928,0.049230773,0.06564103,0.11158975,0.16082053,0.20020515,0.20348719,0.16738462,0.07876924,0.14441027,0.24615386,0.41025645,0.7811283,1.2931283,2.5698464,3.6496413,3.4067695,0.571077,0.17394873,0.03938462,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.036102567,0.068923086,0.118153855,0.15097436,0.17394873,0.23958977,0.2297436,0.24287182,0.28225642,0.33476925,0.3708718,0.36102566,0.39712822,0.38400003,0.31507695,0.28225642,0.4955898,0.61374366,0.56123084,0.4266667,0.45620516,0.508718,0.90912825,1.3817437,1.8346668,2.3466668,3.3444104,4.1452312,4.598154,4.7228723,4.716308,5.7074876,6.1308722,6.0652313,5.7042055,5.3398976,4.9132314,4.7524104,4.667077,4.571898,4.5029745,4.164923,3.698872,3.1540515,2.5731285,1.9790771,1.4473847,1.1979488,0.9747693,0.7811283,0.8730257,1.0765129,1.148718,1.1651284,1.1454359,1.0601027,1.1126155,0.9419488,0.79425645,0.8369231,1.1552821,1.1355898,0.9944616,1.024,1.2012309,1.1881026,0.9517949,1.0338463,1.401436,1.8674873,2.0808206,2.2022567,1.9987694,2.0217438,2.300718,2.353231,2.6945643,2.9636924,3.1967182,3.4921029,4.007385,4.269949,4.5390773,4.4307694,3.817026,2.809436,3.3772311,4.1156926,4.3027697,3.751385,2.7995899,2.9735386,2.7995899,2.6518977,2.6322052,2.556718,2.103795,2.038154,2.1792822,2.297436,2.1070771,1.4211283,1.6278975,1.8543591,1.975795,2.6289232,2.6289232,2.3630772,2.7995899,3.6562054,3.4330258,2.989949,2.6256413,2.3466668,2.1366155,1.9396925,1.7066668,1.6836925,1.6640002,1.5458462,1.3423591,1.1585642,1.1716924,1.394872,1.5261539,0.94523084,1.0962052,1.1355898,1.142154,1.1027694,0.90584624,0.8205129,0.65312827,0.4955898,0.38728207,0.3249231,0.24287182,0.190359,0.190359,0.3249231,0.7581539,1.3095386,1.2176411,1.1618463,1.3029745,1.3095386,1.723077,2.2383592,2.7044106,3.2098465,4.066462,5.0642056,5.477744,5.924103,6.665847,7.6110773,8.448001,9.045334,9.586872,10.171078,10.79795,10.962052,10.985026,11.346052,12.117334,12.967385,14.588719,15.560206,16.052513,16.147694,15.842463,14.998976,13.751796,12.931283,12.504617,11.552821,12.058257,11.628308,11.434668,11.736616,11.864616,12.091078,12.842668,12.760616,11.58236,10.138257,10.31877,10.902975,11.16554,10.978462,10.807796,12.087796,12.960821,13.334975,13.443283,13.843694,13.000206,12.960821,13.236514,13.59754,14.053744,15.43877,16.377438,17.145437,17.46708,16.531694,15.783386,15.402668,15.392821,15.527386,15.346873,15.514257,15.803078,16.09518,16.003283,14.8709755,14.135796,13.11836,12.340514,11.861334,11.280411,10.515693,9.96759,9.878975,10.197334,10.584617,10.47959,10.581334,10.840616,11.35918,12.416001,12.668719,11.910565,11.437949,11.437949,10.978462,10.394258,10.9226675,11.634872,12.130463,12.544001,11.382154,10.453334,9.872411,9.409642,8.503796,7.834257,7.650462,7.7357955,7.939283,8.208411,8.369231,7.830975,7.1220517,6.7117953,6.997334,6.688821,6.701949,6.875898,7.0826674,7.24677,7.0957956,6.626462,6.3179493,6.301539,6.3540516,5.7501545,5.0904617,4.5554876,4.381539,4.824616,4.9493337,4.7491283,4.6145644,4.775385,5.277539,5.8223596,6.373744,6.5411286,6.262154,5.8157954,2.7142565,2.8389745,2.228513,1.7427694,1.6902566,1.8215386,2.0545642,2.1169233,2.0841026,2.0841026,2.3072822,1.9692309,1.6672822,1.5819489,1.6607181,1.6246156,1.7460514,1.9495386,2.1858463,2.4516926,2.7700515,3.5741541,4.332308,4.699898,4.8114877,5.2742567,5.796103,6.4754877,6.701949,6.1997952,5.0018463,4.5029745,4.4406157,4.460308,4.3552823,4.073026,3.7152824,4.1124105,4.647385,4.5489235,2.8914874,1.270154,0.76800007,0.67938465,0.6662565,0.7581539,1.014154,1.2438976,1.5360001,1.847795,2.0053334,1.910154,1.6672822,1.5130258,1.5163078,1.6016412,1.6968206,1.4966155,1.3751796,1.3456411,1.0568206,0.90912825,0.82379496,0.8172308,0.86974365,0.9124103,1.0502565,1.0075898,1.0272821,1.1060513,0.99774367,0.99774367,0.9878975,0.8533334,0.6170257,0.4397949,0.32820517,0.4201026,0.54482055,0.61374366,0.6104616,0.5940513,0.6826667,0.7122052,0.65641034,0.636718,0.7515898,0.892718,1.1388719,1.522872,2.0512822,2.7306669,3.6890259,4.670359,5.648411,6.8529234,7.975385,9.429334,10.673231,11.303386,11.053949,11.595488,13.380924,15.61272,17.046976,16.01313,15.376411,15.698052,16.347898,17.135592,18.323694,17.952822,18.235079,18.458258,18.527182,18.976822,21.083899,21.192207,20.906668,20.657232,19.72513,19.754667,20.151796,20.017233,19.163898,18.09395,18.842258,19.456001,20.348719,21.769848,23.814566,20.67036,20.706463,20.115694,17.893745,15.816206,15.540514,16.141129,16.790976,17.293129,18.084105,18.546873,18.730669,18.688002,18.38277,17.690258,15.163078,15.025232,15.566771,16.141129,17.161848,17.824821,17.831387,17.585232,16.843489,14.693745,13.328411,12.563693,11.828514,11.250873,11.654565,12.3076935,13.397334,14.516514,15.524104,16.544823,16.8599,16.981335,19.012924,22.478771,24.326567,24.743387,24.789335,26.098873,28.596516,30.513233,31.652105,32.99118,33.670567,34.888206,39.91303,47.52739,56.146057,63.612724,65.45067,54.859493,39.29272,30.47713,26.098873,24.448002,24.418463,24.264208,24.195284,24.838566,26.446772,28.918156,30.089848,30.854567,31.947489,33.552414,35.27221,34.97682,38.15385,48.436516,61.312004,64.105034,48.64657,36.873848,29.249643,25.097849,22.616617,22.327797,19.941746,19.446156,21.986464,25.833027,31.379694,36.52267,40.306873,41.196312,37.08062,37.56636,39.73908,39.11221,34.69785,28.973951,23.85395,22.038977,19.511797,15.386257,11.890873,15.468308,18.927591,19.968002,18.087385,14.601848,11.98277,10.732308,9.110975,6.5378466,3.6069746,7.312411,6.488616,4.7556925,4.8016415,8.36595,12.780309,15.780104,15.258258,11.424822,6.8233852,5.5893335,5.730462,5.5663595,4.7622566,4.352,3.0818465,2.5173335,2.5074873,3.5905645,6.9809237,6.8365135,4.519385,2.5796926,2.3401027,3.882667,4.007385,4.4045134,3.6824617,2.1202054,1.6771283,4.397949,6.987488,8.132924,7.3780518,5.113436,5.914257,4.6211286,2.8947694,1.5622566,0.6301539,0.6235898,1.2865642,2.281026,3.308308,4.092718,3.895795,3.5446157,3.2131286,3.121231,3.5183592,2.9801028,4.5390773,6.377026,6.928411,4.857436,6.2555904,6.3179493,8.444718,10.417232,4.4242053,13.11836,8.556309,3.6463592,3.0096412,3.006359,3.2984617,3.7874875,4.4340515,4.9985647,5.0182567,4.5390773,3.0982566,1.8740515,1.2307693,0.71548724,0.7778462,2.166154,3.045744,2.9013336,2.5271797,1.6443079,1.4802053,2.4484105,4.0008206,4.6244106,2.0808206,1.8904617,1.9626669,1.782154,2.4057438,1.9298463,1.7165129,1.6049232,1.5163078,1.4473847,0.83035904,0.5481026,0.574359,0.71548724,0.5874872,0.5349744,0.47589746,0.54482055,0.7450257,0.9419488,0.8205129,0.49887183,0.26584616,0.190359,0.108307704,0.06564103,0.04594872,0.06235898,0.098461546,0.11158975,0.108307704,0.06235898,0.02297436,0.009846155,0.009846155,0.013128206,0.01969231,0.01969231,0.013128206,0.016410258,0.098461546,0.16410258,0.1148718,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016410258,0.036102567,0.07876924,0.118153855,0.07876924,0.07548718,0.055794876,0.049230773,0.055794876,0.06564103,0.059076928,0.059076928,0.052512825,0.04266667,0.06235898,0.09189744,0.14112821,0.21333335,0.26912823,0.2297436,0.16738462,0.14769232,0.24287182,0.46276927,0.7515898,1.8313848,3.2032824,3.495385,2.3040001,0.2231795,0.18707694,0.08205129,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.029538464,0.06564103,0.09189744,0.12471796,0.18051283,0.24943592,0.2100513,0.24615386,0.28882053,0.3249231,0.39056414,0.32164106,0.36430773,0.40369233,0.380718,0.32164106,0.41682056,0.5940513,0.5907693,0.4594872,0.571077,0.56451285,0.80738467,1.2537436,1.8412309,2.5107694,3.5544617,4.493129,4.6867695,4.457026,5.106872,5.9634876,5.8880005,5.7009234,5.684513,5.5958977,4.827898,4.71959,4.644103,4.4340515,4.3749747,4.0336413,3.5380516,2.934154,2.300718,1.719795,1.2340513,1.1027694,0.9747693,0.7975385,0.81066674,0.9517949,1.0404103,1.0699488,1.0272821,0.90584624,1.0469744,1.1618463,1.1355898,1.024,1.0633847,1.0043077,0.92553854,1.0108719,1.214359,1.2340513,1.0535386,1.083077,1.3817437,1.7755898,1.8674873,1.9790771,1.9003079,1.8937438,2.166154,2.8488207,2.8980515,2.8488207,2.7503593,2.8947694,3.8367183,4.266667,3.9253337,3.4133337,2.9440002,2.3466668,3.0293336,3.501949,3.4166157,3.0654361,3.3608208,3.0654361,2.740513,2.5600002,2.4910772,2.284308,2.2055387,2.1366155,2.041436,1.8904617,1.6213335,1.3883078,1.6738462,1.9068719,1.9954873,2.3302567,2.4746668,2.2449234,2.3696413,2.861949,3.0293336,2.8816411,2.6289232,2.2055387,1.8674873,2.2055387,1.9889232,1.7001027,1.5195899,1.4834872,1.4736412,1.4112822,1.4112822,1.3817437,1.2307693,0.86317956,0.9944616,0.98461545,0.98133343,0.9714873,0.8008206,0.73517954,0.5874872,0.4266667,0.3052308,0.23302566,0.20020515,0.17066668,0.2297436,0.46933338,0.9911796,1.1881026,1.1782565,1.142154,1.1749744,1.2931283,1.7952822,2.3138463,2.7175386,3.1113849,3.8498464,4.903385,5.398975,5.7764106,6.2687182,6.8955903,7.4240007,8.3364105,9.088,9.616411,10.345026,10.81436,10.988309,11.346052,12.12718,13.338258,14.135796,15.012104,15.428925,15.320617,15.113848,14.027489,12.672001,11.969642,11.897437,11.47077,12.137027,11.526565,11.096616,11.254155,11.372309,11.35918,12.153437,12.448821,11.98277,11.52,11.191795,11.113027,10.8996935,10.673231,11.034257,11.608616,12.773745,13.722258,14.086565,13.938873,13.692719,13.6697445,13.8075905,14.03077,14.267078,15.419078,16.190361,16.827078,17.106052,16.361027,15.212309,14.565744,14.198155,14.063591,14.276924,14.716719,15.248411,15.783386,15.750566,14.089848,12.947693,12.051693,11.536411,11.270565,10.860309,10.59118,10.299078,10.299078,10.594462,10.893129,10.5780525,10.469745,10.70277,11.286975,12.117334,12.658873,11.864616,11.372309,11.457642,11.027693,10.70277,11.149129,11.546257,11.608616,11.579078,10.568206,9.888822,9.6065645,9.40636,8.618668,7.972103,7.6964107,7.506052,7.4010262,7.6603084,8.001641,7.5881033,7.020308,6.705231,6.872616,6.701949,6.5411286,6.4754877,6.4722056,6.36718,6.0816417,5.940513,5.940513,6.0160003,6.0258465,5.425231,4.706462,4.2896414,4.345436,4.8016415,4.850872,4.644103,4.5554876,4.7655387,5.2545643,5.661539,5.8945646,5.8289237,5.549949,5.3694363,2.9078977,2.5009232,2.0906668,1.8970258,1.9561027,2.1267693,2.3926156,2.3630772,2.1989746,2.0841026,2.2088206,1.8346668,1.6607181,1.5589745,1.4998976,1.5556924,1.6147693,1.7985642,2.048,2.3040001,2.4976413,3.0654361,3.882667,4.384821,4.571898,4.9920006,5.540103,6.2588725,6.4295387,5.792821,4.5817437,4.2207184,3.8728209,3.6890259,3.6562054,3.6036925,3.636513,4.020513,4.46359,4.453744,3.2754874,1.4473847,0.8467693,0.7220513,0.69579494,0.7515898,1.0896411,1.3161026,1.585231,1.910154,2.156308,2.03159,1.6771283,1.4408206,1.4211283,1.4736412,1.4408206,1.3029745,1.270154,1.2898463,1.0568206,0.85005134,0.79097444,0.7975385,0.8008206,0.7417436,0.79425645,0.77456415,0.8402052,0.955077,0.88943595,0.90912825,0.90256417,0.8008206,0.62030774,0.47589746,0.37743592,0.38400003,0.45620516,0.5481026,0.63343596,0.69907695,0.77456415,0.79097444,0.77456415,0.85005134,0.94523084,1.1881026,1.5622566,2.028308,2.5435898,3.1343591,4.0336413,4.900103,5.674667,6.5903597,7.686565,8.900924,9.980719,10.607591,10.407386,11.286975,13.99795,15.576616,15.629129,16.347898,16.603899,17.27672,17.818258,18.153027,18.694565,19.974566,21.106873,22.176823,23.292719,24.595694,25.918362,25.990566,25.619694,24.753233,22.485334,21.822361,20.978874,19.744822,18.346668,17.460514,18.36308,18.7799,19.67918,20.949335,21.395695,21.563078,21.3399,19.702156,16.8599,14.244103,13.732103,13.627078,13.994668,14.86113,16.229744,16.518566,17.030565,17.631182,17.99549,17.588514,15.835898,15.556924,15.770258,16.393847,18.25477,18.638771,18.46154,17.637745,16.256,14.592001,13.269335,12.163283,11.090053,10.33518,10.65354,11.132719,12.245335,12.754052,13.08554,15.346873,16.758156,16.83036,17.8839,20.617847,24.113234,24.54318,24.073849,24.398771,26.486156,30.58872,33.257027,35.43631,36.562054,37.49744,40.530056,44.02544,47.11385,52.48657,57.98072,56.576004,43.401848,32.961643,26.666668,24.244514,23.752207,23.46667,23.624207,24.021336,25.206156,28.498053,30.739695,31.520823,31.845745,32.44308,33.765747,34.92431,36.64739,45.98154,61.63693,74.0037,62.260517,48.390568,37.133133,30.450874,27.51672,24.198566,19.91549,19.012924,22.232616,26.725746,31.412516,35.764515,38.76103,39.14831,35.459286,36.775387,37.031387,33.089645,26.089027,21.454771,18.31713,21.287386,21.714052,17.952822,15.343591,19.347694,20.361847,20.420925,19.492104,15.481437,14.503386,12.78359,9.317744,4.9821544,2.5271797,6.4623594,4.7917953,3.751385,5.366154,7.456821,9.944616,12.360206,13.302155,12.087796,8.746667,7.02359,6.7774363,6.226052,4.9132314,3.6857438,2.8816411,2.6486156,2.8521028,3.6135387,5.3431797,7.4699492,5.940513,3.8400004,3.1376412,4.6867695,4.7425647,4.893539,3.9417439,2.2449234,1.719795,3.2754874,5.1626673,5.9569235,5.2414365,3.6168208,4.850872,4.7360005,3.7251284,2.2777438,0.8598975,0.7450257,1.2603078,2.1431797,3.2065644,4.3290257,4.7327185,4.598154,4.634257,5.179077,6.193231,3.5249233,5.3169236,7.5946674,7.680001,4.194462,5.4383593,5.677949,8.648206,11.533129,4.9427695,15.908104,9.974154,3.5347695,2.487795,2.225231,2.5961027,3.006359,4.1780515,5.786257,6.452513,5.6320004,3.5577438,1.9364104,1.2438976,0.7515898,0.65312827,1.7887181,3.0326157,3.636513,3.2525132,2.0676925,2.1070771,2.8225644,4.4242053,7.857231,4.1452312,2.6518977,2.0578463,1.8674873,2.4155898,1.3522053,1.4605129,1.7165129,1.6836925,1.4900514,0.9714873,0.67282057,0.56123084,0.52512825,0.37415388,0.32164106,0.20020515,0.16738462,0.256,0.3708718,0.3052308,0.2100513,0.14441027,0.11158975,0.052512825,0.026256412,0.016410258,0.013128206,0.03938462,0.16082053,0.14769232,0.098461546,0.072205134,0.06564103,0.02297436,0.0032820515,0.009846155,0.009846155,0.0032820515,0.02297436,0.128,0.26256412,0.2855385,0.17394873,0.013128206,0.108307704,0.2297436,0.27241027,0.21989745,0.14112821,0.08533334,0.14441027,0.15425642,0.08861539,0.055794876,0.128,0.08861539,0.055794876,0.059076928,0.06564103,0.049230773,0.059076928,0.06235898,0.052512825,0.06235898,0.08533334,0.14769232,0.23630771,0.3052308,0.27241027,0.29210258,0.22646156,0.26912823,0.4955898,0.8598975,1.7887181,2.6486156,2.3958976,1.1355898,0.14441027,0.24615386,0.12143591,0.013128206,0.0,0.006564103,0.006564103,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.029538464,0.072205134,0.108307704,0.14441027,0.18051283,0.20020515,0.18707694,0.24943592,0.30194873,0.3314872,0.40369233,0.36430773,0.34133336,0.34133336,0.34789747,0.3249231,0.318359,0.47261542,0.54482055,0.5284103,0.6301539,0.65969235,0.8205129,1.1913847,1.8116925,2.6945643,3.5905645,4.5128207,4.493129,4.059898,5.2447186,5.618872,5.3005133,5.146257,5.32677,5.330052,4.6276927,4.4274874,4.3060517,4.1813335,4.2962055,4.007385,3.5905645,2.9801028,2.2482052,1.5885129,1.1454359,1.0338463,0.955077,0.827077,0.78769237,0.8730257,0.96492314,0.9944616,0.9517949,0.8763078,0.96492314,1.2077949,1.2570257,1.083077,0.96492314,0.90256417,0.88615394,0.97805136,1.1585642,1.3193847,1.204513,1.2242053,1.4736412,1.8149745,1.8970258,2.172718,2.1267693,2.0611284,2.2055387,2.7306669,2.8127182,2.7503593,2.484513,2.4385643,3.5249233,3.9023592,3.4921029,2.9013336,2.4484105,2.1530259,2.878359,3.3476925,3.2131286,2.8750772,3.4592824,3.0490258,2.6978464,2.4582565,2.294154,2.100513,2.284308,2.176,2.422154,2.609231,1.2964103,1.3226668,1.6377437,1.9035898,2.0545642,2.294154,2.6551797,2.3171284,2.2383592,2.546872,2.537026,2.484513,2.3138463,2.041436,1.9035898,2.3335385,2.034872,1.6410258,1.394872,1.394872,1.5885129,1.5983591,1.5753847,1.4244103,1.1782565,0.9682052,0.90256417,0.8467693,0.83035904,0.8008206,0.65312827,0.5940513,0.47589746,0.32820517,0.20020515,0.15097436,0.16082053,0.17066668,0.3117949,0.6301539,1.0601027,1.1060513,1.1651284,1.1979488,1.2406155,1.4112822,1.8970258,2.4549747,2.878359,3.2164104,3.7973337,4.5456414,5.156103,5.602462,6.009436,6.6527185,7.204103,8.146052,8.897642,9.498257,10.5780525,10.522257,10.870154,11.408411,12.163283,13.3940525,13.8765135,14.7790785,14.972719,14.411489,14.139078,12.911591,11.749744,12.032001,13.266052,13.075693,12.62277,11.746463,11.250873,11.398565,11.904001,11.424822,11.477334,11.697231,11.920411,12.166565,11.851488,11.30995,10.893129,10.939077,11.772718,11.753027,12.977232,14.273643,14.880821,14.460719,14.857847,14.8250265,14.828309,14.946463,14.900514,15.645539,16.308514,16.853334,17.089642,16.682669,14.91036,13.676309,12.918155,12.662155,13.013334,13.472821,14.260514,14.916924,14.805334,13.095386,11.667693,10.971898,10.804514,10.866873,10.738873,10.7158985,10.676514,10.709334,10.840616,11.024411,10.893129,10.794667,10.955488,11.329642,11.605334,11.989334,11.369026,11.050668,11.244308,11.0605135,11.1294365,11.428103,11.513436,11.204924,10.584617,9.974154,9.714872,9.6,9.353847,8.648206,8.001641,7.653744,7.3583593,7.194257,7.5552826,7.9130263,7.568411,7.0498466,6.672411,6.554257,6.633026,6.518154,6.3507695,6.183385,5.9930263,5.5991797,5.549949,5.622154,5.671385,5.618872,4.9460516,4.3618464,4.1550775,4.352,4.6966157,4.841026,4.8607183,4.9329233,5.1232824,5.408821,5.612308,5.6418467,5.4416413,5.152821,5.106872,2.7175386,2.3401027,2.1989746,2.3794873,2.7273848,2.8455386,2.8127182,2.5600002,2.228513,1.9298463,1.7263591,1.5327181,1.585231,1.5885129,1.5163078,1.591795,1.5589745,1.7033848,1.9396925,2.1891284,2.3958976,2.6387694,3.2820516,3.882667,4.3027697,4.71959,5.5204105,6.3310776,6.2752824,5.3202057,4.2994876,3.8859491,3.5577438,3.3345644,3.2164104,3.1737437,3.7349746,4.096,4.3060517,4.135385,3.0785644,1.4506668,0.74830776,0.52512825,0.5218462,0.6498462,0.9419488,1.1782565,1.4178462,1.6869745,1.9987694,1.8806155,1.6443079,1.4933335,1.4244103,1.2176411,1.0896411,1.0338463,1.1191796,1.214359,1.0075898,0.8566154,0.86974365,0.8467693,0.7384616,0.6235898,0.45292312,0.43651286,0.53825647,0.67938465,0.72861546,0.82379496,0.8369231,0.7844103,0.6892308,0.58420515,0.47589746,0.42994875,0.39712822,0.39056414,0.47261542,0.761436,0.90584624,1.0010257,1.1290257,1.3489232,1.3357949,1.6180514,1.975795,2.3204105,2.6847181,3.2328207,3.9417439,4.568616,5.146257,5.979898,7.312411,8.388924,9.4916935,10.55836,11.18195,12.770463,16.23631,18.70113,19.541334,20.407797,21.451488,22.134155,22.065233,21.80595,22.89231,24.566156,25.93149,27.549541,29.348104,30.631388,30.28349,30.769234,30.759386,29.38749,26.246567,25.189745,24.152617,22.560822,20.535797,18.884924,18.28431,18.49436,19.446156,20.65395,21.221745,23.522463,22.088207,19.721848,17.493334,14.739694,14.404924,13.863386,13.833847,14.562463,15.786668,16.725334,17.59836,18.326975,18.697847,18.336823,16.59077,16.423386,16.708925,16.945232,17.240616,17.601643,17.59836,16.984617,15.786668,14.283488,12.777026,11.920411,11.339488,11.027693,11.352616,11.546257,12.274873,13.111795,14.01436,15.29436,17.132309,17.69354,18.747078,21.264412,25.429335,26.033234,25.537643,25.393232,26.843899,30.923489,33.7559,36.617847,38.79713,40.034466,40.516926,40.881233,41.70831,44.28144,48.3479,52.145233,43.953236,35.567593,29.371078,26.000412,24.33313,24.342976,24.720411,24.661335,24.960001,27.989336,30.641233,31.455181,31.389542,31.366566,32.262566,34.92103,35.600414,42.962055,58.95221,78.795494,73.94134,60.69498,46.240826,35.265644,29.912617,25.53436,20.726156,19.954874,23.808002,28.996925,32.879593,36.135387,37.70749,37.097027,34.386055,34.989952,31.471592,24.894361,18.103796,15.707899,15.816206,20.427488,22.744617,21.553232,21.225027,25.015797,22.79713,20.821335,19.994259,15.891693,17.03713,15.27795,10.571488,4.9329233,2.412308,2.7208207,2.359795,3.9253337,6.8365135,7.322257,7.8473854,8.779488,10.482873,11.907283,10.581334,7.8802056,6.5411286,5.58277,4.4274874,2.9013336,2.7241027,2.8258464,3.1606157,3.6463592,4.161641,7.9195905,7.1680007,5.287385,4.4340515,5.5138464,4.821334,4.4077954,3.370667,1.9922053,1.7165129,2.1956925,4.2305646,6.2096415,6.6461544,4.1878977,5.789539,6.931693,6.695385,4.9920006,2.5698464,1.3784616,1.6082052,2.3433847,3.2032824,4.348718,5.3136415,6.189949,7.0432825,8.237949,10.44677,4.6211286,4.857436,6.688821,7.0104623,4.066462,3.8137438,4.8771286,8.044309,10.098872,3.7973337,9.816616,6.4754877,2.802872,2.1169233,2.03159,3.239385,3.186872,3.8498464,5.435077,6.4065647,5.284103,3.314872,1.7624617,1.0568206,0.80738467,0.6629744,0.58420515,1.4441026,2.806154,2.934154,2.1300514,2.5698464,3.5610259,5.2381544,8.582564,6.449231,4.2863593,3.2065644,3.2131286,3.2065644,1.6508719,2.044718,2.0709746,1.2504616,0.9353847,1.3292309,1.0502565,0.7253334,0.574359,0.43323082,0.45620516,0.34789747,0.256,0.21333335,0.16410258,0.14112821,0.101743594,0.072205134,0.049230773,0.02297436,0.013128206,0.09189744,0.11158975,0.098461546,0.29210258,0.15753847,0.108307704,0.118153855,0.128,0.032820515,0.013128206,0.0032820515,0.006564103,0.016410258,0.04266667,0.17066668,0.29210258,0.4266667,0.47917953,0.25928208,0.48246157,0.7811283,0.81066674,0.56451285,0.3708718,0.20348719,0.35446155,0.36102566,0.16082053,0.1148718,0.31507695,0.26256412,0.17723078,0.14441027,0.11158975,0.08861539,0.09189744,0.08533334,0.068923086,0.068923086,0.09189744,0.15097436,0.23302566,0.30851284,0.3249231,0.4135385,0.40369233,0.48246157,0.76800007,1.332513,1.3226668,1.1782565,0.79097444,0.30194873,0.11158975,0.23630771,0.12471796,0.01969231,0.006564103,0.013128206,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.04266667,0.07876924,0.14112821,0.17394873,0.16410258,0.14769232,0.18379489,0.24943592,0.30194873,0.34133336,0.4135385,0.46276927,0.34789747,0.256,0.256,0.3117949,0.2855385,0.35446155,0.4594872,0.5415385,0.5546667,0.67938465,0.8336411,1.1651284,1.7952822,2.806154,3.370667,4.096,4.0500517,3.761231,5.208616,5.024821,5.0084105,5.0477953,5.0149746,4.772103,4.240411,3.8728209,3.8367183,4.1091285,4.450462,4.210872,3.8629746,3.2722054,2.4582565,1.595077,1.1158975,0.9616411,0.90912825,0.8533334,0.78769237,0.79097444,0.8598975,0.90584624,0.92553854,0.9747693,0.955077,1.083077,1.0962052,0.9714873,0.92553854,0.92553854,0.9288206,0.9714873,1.1060513,1.4080001,1.394872,1.4309745,1.6443079,1.9922053,2.2547693,2.7011285,2.5271797,2.4057438,2.4648206,2.2908719,2.4352822,2.5632823,2.477949,2.4484105,3.2098465,3.3903592,3.387077,2.9801028,2.353231,2.0939488,2.6945643,3.3411283,3.5216413,3.2918978,3.2853336,3.0687182,2.806154,2.5074873,2.2383592,2.1333334,2.1202054,1.9954873,2.7602053,3.4494362,1.142154,1.2668719,1.6836925,2.0545642,2.3663592,2.9210258,3.0490258,2.4549747,2.5173335,3.0030773,2.0939488,1.9528207,1.8806155,1.9790771,2.15959,2.1398976,1.782154,1.5688206,1.4276924,1.404718,1.6804104,1.6607181,1.5885129,1.4473847,1.2373334,0.9714873,0.8369231,0.79097444,0.7450257,0.65312827,0.5218462,0.4266667,0.32164106,0.21333335,0.12143591,0.101743594,0.108307704,0.17723078,0.39712822,0.7187693,0.9517949,1.1782565,1.2471796,1.3161026,1.4276924,1.5064616,2.0020514,2.6847181,3.2032824,3.515077,3.8728209,4.2305646,4.9362054,5.4383593,5.85518,6.9710774,7.896616,8.493949,8.923898,9.531077,10.8307705,10.148104,10.811078,11.670976,12.393026,13.4629755,13.974976,15.048206,15.051488,13.827283,12.724514,11.687386,11.099898,12.498053,14.79877,14.290052,12.678565,11.913847,11.848206,12.27159,12.911591,12.25518,11.497026,11.303386,11.562668,11.385437,11.926975,11.631591,11.362462,11.61518,12.511181,12.504617,13.584412,14.65436,15.16636,15.126975,15.845745,16.009848,16.128002,16.20677,15.730873,15.855591,16.28554,16.810667,17.14872,16.94195,14.674052,12.996924,12.1238985,11.949949,12.071385,12.22236,12.99036,13.50236,13.259488,12.133744,10.745437,10.240001,10.358154,10.71918,10.807796,10.692924,10.801231,10.929232,11.021129,11.155693,11.58236,11.661129,11.608616,11.503591,11.30995,11.158976,10.902975,10.781539,10.850462,10.965334,11.336206,11.477334,11.329642,10.811078,9.793642,9.593436,9.662359,9.527796,9.068309,8.503796,7.90318,7.571693,7.3714876,7.3550773,7.7718983,8.162462,7.8637953,7.250052,6.665847,6.416411,6.491898,6.5345645,6.3967185,6.1440005,6.058667,5.612308,5.4547696,5.428513,5.405539,5.3070774,4.568616,4.2568207,4.276513,4.4832826,4.6834874,5.031385,5.3037953,5.5204105,5.6352825,5.5565133,5.5072823,5.533539,5.4186673,5.182359,5.0871797,2.7306669,2.6453335,3.045744,3.3641028,3.3936412,3.2951798,3.626667,3.945026,3.370667,2.1300514,1.5556924,1.3128207,1.0962052,0.9747693,1.0305642,1.3718976,1.4966155,1.5983591,1.7690258,2.041436,2.3958976,2.5435898,2.7076926,3.0194874,3.6102567,4.6244106,5.4908724,6.0652313,5.7042055,4.604718,3.8006158,3.3476925,3.4166157,3.2820516,2.917744,2.989949,3.0654361,3.045744,3.2656412,3.4822567,2.8849232,1.4309745,0.65641034,0.3511795,0.30851284,0.32164106,0.6498462,1.0896411,1.3751796,1.4998976,1.6935385,1.6935385,1.529436,1.3161026,1.1946667,1.3259488,1.083077,0.83035904,0.7089231,0.71548724,0.702359,0.8369231,0.9353847,0.8730257,0.6826667,0.5481026,0.4397949,0.4660513,0.48574364,0.47261542,0.5349744,0.5218462,0.7187693,0.7450257,0.571077,0.5349744,0.48574364,0.48246157,0.4201026,0.30194873,0.2297436,0.6432821,0.95835906,1.2931283,1.6672822,1.9823592,1.8609232,1.9856411,2.0709746,2.1234872,2.4418464,3.2229745,4.0402055,4.7622566,5.395693,6.1046157,7.433847,9.176616,11.421539,13.817437,15.563488,17.650873,20.552206,25.081438,30.18831,32.958363,31.284515,29.466259,27.812105,26.886566,27.497028,28.92472,30.178463,31.67508,33.414566,34.986668,34.914463,35.344414,35.344414,34.28103,31.812925,30.66749,29.784618,27.98277,25.012514,21.546669,19.908924,20.178053,21.320208,22.478771,22.980925,25.104412,24.966566,23.611078,21.540104,18.707693,17.962667,17.161848,16.662975,16.873028,18.264616,20.118977,21.32677,22.002874,21.766565,19.728413,18.021746,18.609232,18.848822,17.801847,16.249437,16.20349,15.320617,14.582155,14.099693,13.121642,11.9860525,12.242052,12.5374365,12.317539,11.841642,12.57354,14.057027,15.14995,15.868719,17.394873,18.323694,18.855387,19.259079,21.290668,28.212515,28.445541,26.479591,25.783796,27.506874,30.470566,32.278976,35.987694,38.7118,39.443695,39.079388,37.81908,39.35508,41.46872,43.477337,46.25067,41.609848,36.92636,32.469337,28.639181,25.954464,25.72472,26.213745,26.440207,26.440207,27.283695,30.13908,31.530668,31.721027,31.287798,31.126976,35.09498,36.050053,41.750977,56.018055,78.73642,80.05252,70.34093,54.21293,37.67795,28.107489,24.90749,21.664822,21.93395,26.335182,32.561234,35.4199,36.617847,36.82462,36.42421,35.521645,33.362053,24.792618,17.207796,13.768207,13.413745,14.7790785,16.997746,19.941746,23.092514,25.557335,23.958977,21.50072,20.033642,18.697847,13.899488,16.610462,16.57436,12.898462,7.02359,2.7175386,1.5327181,1.4572309,1.9364104,3.2820516,6.636308,6.491898,6.491898,8.664616,11.972924,12.314258,8.579283,4.8344617,2.7536411,2.281026,1.6311796,2.0611284,2.5337439,2.9669745,3.3805132,3.9056413,6.042257,5.989744,5.5565133,5.7698464,6.882462,4.6834874,2.5961027,1.595077,1.6311796,1.6311796,2.1103592,5.3760004,9.337437,11.07036,6.8365135,7.4699492,11.234463,12.980514,10.9915905,6.987488,2.789744,2.1070771,2.3630772,2.5895386,3.4330258,5.7632823,10.410667,12.475078,12.228924,15.120412,7.0892315,5.8880005,5.5072823,4.2240005,4.578462,3.1737437,10.502565,12.921437,7.77518,3.4166157,2.172718,1.6508719,1.4506668,1.5064616,2.1070771,6.9152827,6.5805135,4.8344617,3.8662567,4.31918,3.3903592,2.4155898,1.6607181,1.1618463,0.74830776,0.69907695,0.6301539,0.75487185,1.0272821,1.1749744,1.6016412,2.2482052,3.5807183,5.7009234,8.362667,8.54318,7.2894363,5.5991797,4.1714873,3.4034874,2.0217438,1.6246156,1.5622566,1.522872,1.5097437,3.0851285,2.03159,1.0305642,0.92225647,0.702359,0.761436,0.8041026,0.702359,0.446359,0.15097436,0.07876924,0.08861539,0.07548718,0.032820515,0.04594872,0.04594872,0.42994875,0.5152821,0.3052308,0.48902568,0.24287182,0.108307704,0.072205134,0.08205129,0.04594872,0.032820515,0.02297436,0.026256412,0.055794876,0.09189744,0.23958977,0.32820517,0.43323082,0.6629744,1.1749744,1.3226668,1.6147693,1.3456411,0.64000005,0.45620516,0.24943592,0.54482055,0.7187693,0.58092314,0.39712822,0.6662565,0.7318975,0.6235898,0.41682056,0.25928208,0.23630771,0.20020515,0.14769232,0.0951795,0.108307704,0.118153855,0.16738462,0.23958977,0.33476925,0.45620516,0.46933338,0.53825647,0.93866676,1.6016412,2.0906668,1.6869745,0.80738467,0.23958977,0.16082053,0.13784617,0.16082053,0.08533334,0.029538464,0.02297436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.029538464,0.09189744,0.07876924,0.08533334,0.098461546,0.12143591,0.18379489,0.21989745,0.21989745,0.21333335,0.256,0.4266667,0.47589746,0.36102566,0.26256412,0.27569234,0.39712822,0.4201026,0.36430773,0.31507695,0.3249231,0.39712822,0.5316923,0.77456415,1.1913847,1.8313848,2.7470772,3.1245131,3.7152824,3.8071797,3.7185643,4.8049235,5.208616,5.786257,5.901129,5.5532312,5.3694363,4.076308,3.4888208,3.6824617,4.266667,4.3651285,4.1452312,3.8596926,3.2984617,2.4024618,1.2668719,0.86317956,0.80738467,0.9485129,1.0568206,0.82379496,0.65312827,0.6826667,0.7253334,0.72861546,0.7778462,0.88943595,0.9156924,0.9288206,0.9616411,1.020718,1.1191796,1.1257436,1.0699488,1.0404103,1.1749744,1.6508719,1.7165129,1.7099489,1.913436,2.546872,2.7798977,2.681436,2.6584618,2.806154,2.9144619,2.4615386,2.5140514,2.7700515,3.0391798,3.2361028,3.6004105,3.2623591,2.7175386,2.3138463,2.228513,2.4976413,2.7470772,2.9604106,3.0785644,3.006359,2.9440002,2.8750772,2.789744,2.6715899,2.487795,1.5360001,1.2800001,1.273436,1.2012309,0.88615394,1.3259488,1.7099489,2.1497438,2.7733335,3.7382567,2.665026,2.2416413,2.4484105,2.740513,2.044718,2.3630772,2.3696413,2.349949,2.3335385,2.0906668,1.7723079,1.6213335,1.5655385,1.595077,1.7558975,1.7066668,1.463795,1.2931283,1.2012309,0.94523084,0.8598975,0.702359,0.5907693,0.58420515,0.65641034,0.3249231,0.17066668,0.13456412,0.13784617,0.07548718,0.11158975,0.27897438,0.5284103,0.76800007,0.8533334,1.014154,1.1158975,1.3128207,1.4966155,1.3128207,1.9364104,2.7503593,3.318154,3.629949,4.1058464,4.4701543,4.900103,5.0477953,5.3727183,7.141744,8.155898,8.372514,8.621949,9.281642,10.269539,10.31877,11.283693,11.9171295,12.3766165,14.221129,14.575591,15.14995,14.690463,13.115078,11.490462,10.807796,10.8537445,11.625027,12.2617445,11.076924,11.090053,11.808822,12.576821,12.937847,12.619488,12.655591,11.995898,11.270565,10.689642,10.056206,11.533129,11.848206,11.552821,11.414975,12.389745,12.793437,13.617231,14.03077,14.066873,14.601848,15.701335,16.918976,17.765745,17.782156,16.52513,15.878566,15.442053,15.91795,16.932104,17.027283,15.051488,13.814155,13.059283,12.438975,11.536411,11.401847,11.723488,11.82195,11.510155,11.109744,10.374565,10.240001,10.512411,10.8307705,10.633847,10.354873,10.568206,10.9226675,11.204924,11.352616,12.547283,12.757335,12.268309,11.628308,11.628308,11.211488,11.191795,11.030975,10.709334,10.696206,10.745437,10.774975,10.561642,9.987283,9.048616,9.170052,9.101129,8.818872,8.297027,7.4929237,7.3583593,7.4075904,7.4075904,7.4174366,7.7981544,8.516924,8.185436,7.5388722,6.99077,6.636308,6.5280004,6.5739493,6.3901544,6.009436,5.874872,5.5926156,5.4875903,5.346462,5.110154,4.8672824,4.3060517,4.1846156,4.420923,4.7950773,4.9296412,5.293949,5.3694363,5.4908724,5.6320004,5.3858466,5.287385,5.2381544,5.2676926,5.3202057,5.2348723,1.8412309,2.858667,3.6594875,3.7218463,3.2656412,3.245949,3.4002054,3.3345644,2.789744,1.9823592,1.6049232,1.4309745,1.0994873,0.92553854,1.1520001,1.9232821,1.8674873,1.3883078,1.1027694,1.4539489,2.674872,2.8225644,2.7470772,2.9210258,3.5282054,4.453744,5.349744,5.408821,5.146257,4.821334,4.44718,3.564308,3.18359,3.1474874,3.3017437,3.501949,2.6486156,2.5074873,2.3827693,2.0841026,1.9429746,1.5064616,1.0666667,0.6629744,0.4266667,0.56451285,0.67938465,0.8730257,1.0404103,1.1552821,1.3029745,1.2537436,1.273436,1.270154,1.2209232,1.1684103,1.0404103,0.97805136,0.80738467,0.5513847,0.43323082,0.7450257,0.9517949,0.99774367,0.90256417,0.76800007,0.7089231,0.69579494,0.78769237,0.90912825,0.85005134,0.65312827,0.49887183,0.4135385,0.40369233,0.42338464,0.30851284,0.27897438,0.33476925,0.46933338,0.6695385,0.77128214,1.0075898,1.3915899,1.6672822,1.2996924,1.3456411,1.913436,2.097231,2.034872,2.917744,3.9811285,5.0182567,5.9963083,7.0104623,8.264206,9.760821,12.314258,15.300924,18.22195,20.690052,24.448002,29.144617,32.521847,35.45272,41.941338,42.262978,40.398773,38.85621,37.848618,35.285336,32.97149,32.242874,33.729645,36.644104,38.784004,40.421745,41.70831,43.739902,44.85908,40.66462,37.280823,33.81826,31.806362,30.995695,29.344822,28.763899,27.80226,26.57149,26.12513,28.45867,32.049232,32.298668,30.47713,27.559387,24.247797,21.75672,21.559797,22.967796,24.891079,25.846155,28.04185,31.43549,33.34236,32.57436,29.42031,25.905233,23.781746,21.99631,20.680206,21.13313,18.546873,16.889437,15.238565,13.3940525,11.890873,12.432411,11.881026,10.929232,10.108719,9.7903595,11.74318,13.705847,15.097437,16.006565,17.201233,16.866463,16.846771,17.385027,20.01395,27.542976,28.478361,27.142567,25.888823,26.43036,29.824003,33.749336,36.02708,36.73272,36.535797,36.696617,37.041233,37.300514,38.646156,40.805748,42.06277,41.445747,38.340927,34.6519,31.809643,30.765951,29.51549,29.35795,28.521029,27.30995,28.114054,30.237541,31.458464,31.606155,30.926771,30.116104,33.575386,35.859695,42.962055,56.92062,75.8318,80.37088,73.85929,58.56821,39.86708,26.213745,24.753233,23.96554,26.246567,31.625849,37.763287,36.0599,34.62236,34.832413,35.442875,32.6039,26.597746,18.481232,13.075693,12.015591,13.74195,17.227488,19.242668,20.168207,20.28308,19.761232,18.025026,17.700104,16.443079,14.194873,13.157744,17.526155,16.367592,13.252924,9.508103,4.194462,1.4769232,1.0601027,1.463795,2.3105643,4.3290257,5.435077,4.7360005,6.038975,8.828718,8.274052,5.2709746,3.2984617,2.231795,1.8609232,1.8904617,1.8871796,2.3269746,2.6617439,2.7667694,2.930872,3.1113849,3.6069746,4.857436,6.7117953,8.408616,3.6036925,1.4998976,0.9353847,1.0404103,1.2668719,1.3423591,3.9318976,6.75118,8.257642,7.653744,6.160411,8.697436,11.283693,12.704822,14.532925,9.317744,6.951385,5.024821,3.0293336,2.3466668,5.3924108,8.011488,9.947898,10.866873,10.361437,7.778462,7.506052,5.927385,2.9538465,2.038154,1.7099489,3.764513,4.896821,4.07959,2.5632823,1.8248206,1.5031796,2.0545642,3.4198978,5.034667,12.343796,12.780309,9.639385,5.8092313,3.7809234,2.2482052,2.7503593,3.1409233,2.477949,1.0272821,0.8730257,0.8960001,0.98461545,1.2274873,1.9200002,1.3029745,1.9593848,4.0467696,6.482052,6.944821,4.141949,3.8531284,4.417641,4.4438977,2.806154,2.3630772,2.225231,1.9364104,1.4112822,0.9485129,0.9321026,0.5940513,0.41025645,0.49230772,0.60389745,1.6902566,1.4998976,0.8205129,0.26584616,0.27569234,0.0951795,0.03938462,0.02297436,0.006564103,0.009846155,0.01969231,0.098461546,0.11158975,0.07548718,0.17066668,0.39712822,0.20348719,0.068923086,0.12471796,0.15425642,0.12471796,0.06235898,0.055794876,0.1148718,0.20020515,0.20020515,0.30851284,0.6465641,1.0666667,1.1388719,1.1388719,1.1618463,0.90256417,0.48574364,0.45620516,0.40697438,0.7778462,0.8763078,0.58420515,0.3708718,0.62030774,0.6629744,0.5874872,0.4397949,0.2231795,0.27569234,0.27569234,0.21661541,0.15425642,0.20348719,0.14769232,0.17394873,0.2297436,0.33476925,0.54482055,0.7122052,0.6629744,1.1257436,1.8084104,1.4080001,2.4681027,3.245949,2.7109745,1.273436,0.77128214,0.6892308,0.31507695,0.06564103,0.03938462,0.02297436,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.01969231,0.055794876,0.06564103,0.06564103,0.13128206,0.17394873,0.18379489,0.24287182,0.20348719,0.22646156,0.26912823,0.3117949,0.36758977,0.36758977,0.39056414,0.36102566,0.2855385,0.24943592,0.29538465,0.30851284,0.29210258,0.2855385,0.36102566,0.4266667,0.6662565,1.3128207,2.15959,2.5764105,3.892513,3.9023592,3.6824617,3.8104618,4.378257,4.391385,4.9526157,5.218462,5.0642056,5.0674877,3.8400004,3.5314875,3.9614363,4.5029745,4.082872,3.6890259,3.4264617,2.9472823,2.1497438,1.1815386,0.9156924,0.8369231,0.8336411,0.81066674,0.67610264,0.5152821,0.6071795,0.71548724,0.764718,0.85005134,1.1946667,1.148718,0.9911796,0.90912825,0.99774367,1.2209232,1.3259488,1.2603078,1.1323078,1.1881026,1.3029745,1.6869745,2.0053334,2.1858463,2.4024618,2.809436,2.930872,2.8882053,3.006359,3.817026,3.5511796,3.370667,3.1015387,2.8160002,2.8553848,3.3608208,3.0982566,2.4615386,1.9823592,2.3368206,2.6157951,2.9111798,2.930872,2.6322052,2.2383592,2.537026,2.6683078,2.9440002,3.2361028,2.9768207,1.6902566,1.3095386,1.2570257,1.3095386,1.5688206,1.8215386,2.3860514,2.9144619,3.0293336,2.3335385,1.7001027,1.8248206,2.2613335,2.5862565,2.3991797,2.4910772,2.550154,2.3958976,2.1070771,2.028308,1.585231,1.5327181,1.5163078,1.5031796,1.7788719,1.6311796,1.3751796,1.2931283,1.3226668,1.0568206,0.9616411,0.65969235,0.44307697,0.41025645,0.47261542,0.27897438,0.14441027,0.098461546,0.11158975,0.101743594,0.23630771,0.49887183,0.7384616,0.8763078,0.90256417,0.9353847,0.98461545,1.2012309,1.4572309,1.3718976,1.9954873,2.7306669,3.43959,4.066462,4.630975,4.391385,4.6178465,5.024821,5.5302567,6.2752824,7.0432825,7.6012316,8.697436,10.14154,10.817642,10.407386,11.017847,11.641437,12.310975,14.073437,13.774771,13.797745,13.817437,13.210258,11.050668,10.023385,10.463181,10.70277,10.171078,9.416205,11.139283,11.72677,11.835078,11.897437,12.107488,11.61518,11.204924,11.208206,11.346052,10.752001,10.587898,10.9915905,11.067078,10.948924,11.779283,12.212514,12.668719,13.000206,13.499078,14.897232,16.580925,17.864206,18.517334,18.34995,17.220924,16.282257,15.931078,16.219898,16.768002,16.79754,14.546052,13.380924,12.681848,11.940104,10.742155,10.489437,10.712616,11.2672825,11.792411,11.680821,10.774975,10.555078,10.732308,10.817642,10.134975,9.540924,9.596719,10.023385,10.722463,11.766154,12.816411,12.711386,12.173129,11.651283,11.30995,11.237744,11.388719,11.241027,10.880001,11.0145645,10.8767185,10.7158985,10.407386,9.9282055,9.32759,8.992821,8.73354,8.516924,8.073847,6.9054365,6.7216415,6.738052,6.76759,6.8299494,7.1515903,7.8408213,7.765334,7.2237954,6.6133337,6.4065647,6.432821,6.0816417,5.579488,5.225026,5.3727183,5.356308,5.146257,4.9985647,4.827898,4.2338467,4.197744,4.384821,4.7622566,5.179077,5.330052,5.677949,5.76,5.7501545,5.671385,5.398975,5.3202057,4.893539,4.6834874,4.906667,5.4153852,1.4703591,2.4582565,2.9505644,2.8389745,2.4024618,2.3368206,2.3072822,2.2449234,2.0086155,1.6246156,1.2865642,1.1224617,0.9419488,0.8960001,1.1093334,1.6672822,1.4375386,1.2964103,1.1520001,1.1454359,1.6475899,2.0873847,2.1431797,2.3466668,2.8947694,3.6496413,4.3027697,4.519385,4.781949,5.0116925,4.5817437,3.945026,3.3017437,2.9538465,2.986667,3.255795,2.6223593,2.3466668,2.0611284,1.785436,1.9298463,1.7526156,1.3029745,0.9189744,0.7384616,0.7253334,0.78769237,0.88287187,0.98461545,1.079795,1.1684103,1.2537436,1.270154,1.3620514,1.5163078,1.5589745,1.6738462,1.3883078,1.0436924,0.7811283,0.5415385,0.7253334,0.8566154,0.9485129,0.9911796,0.9517949,0.86646163,0.98461545,1.2898463,1.6114873,1.6443079,1.1881026,0.6432821,0.28882053,0.19692309,0.23302566,0.17723078,0.16410258,0.23302566,0.4594872,0.9616411,0.8467693,1.0272821,1.1618463,1.1027694,0.90912825,1.0601027,1.6049232,2.2153847,2.9046156,4.023795,5.2414365,6.439385,7.5421543,8.625232,9.921641,11.943385,15.225437,19.052309,23.61436,30.027489,31.215591,34.090668,36.26995,37.940517,41.892105,42.9719,43.093338,42.998158,42.706055,41.524517,36.959183,35.725132,37.159386,39.742363,41.078156,43.677544,45.22667,48.019695,50.924313,49.40472,46.29662,42.61744,40.68431,40.32985,38.8759,36.053337,32.580925,29.390772,27.969643,30.372105,34.13662,35.265644,34.609234,32.551388,29.013336,25.783796,23.584822,23.32554,24.658052,25.990566,28.018873,31.977028,35.41662,36.88698,35.94503,34.884926,34.12677,33.18154,32.08862,31.409233,26.646976,21.970053,17.716515,14.729847,14.345847,12.301129,10.463181,9.097847,8.687591,9.898667,11.352616,13.08554,14.408206,15.376411,16.804104,15.504412,14.674052,14.818462,17.345642,24.562874,24.95672,23.758772,23.131899,24.083694,26.469746,30.470566,32.958363,33.378464,33.21108,35.96472,38.350773,37.717335,38.032413,39.699696,39.568413,40.63508,38.803696,36.066463,34.067696,34.100517,33.00759,31.940926,30.434464,28.980515,28.996925,30.001232,31.0679,31.172926,30.431181,30.099695,32.068924,35.895798,43.861336,56.42175,72.20185,77.44,76.64575,64.47919,44.10421,27.204926,24.979694,26.555079,31.806362,38.47877,42.184208,36.864002,34.881645,35.045746,34.005337,26.256413,20.07631,14.208001,10.896411,10.880001,13.367796,17.851078,19.692308,20.266668,19.610258,16.416822,15.635694,18.038155,18.966976,18.474669,21.32677,24.149336,18.011898,12.33395,9.426052,4.4996924,3.43959,1.6607181,0.81394875,1.3292309,2.3893335,3.4625645,3.4625645,4.322462,5.933949,6.163693,3.7842054,2.989949,2.5764105,2.100513,1.9167181,2.356513,2.4385643,2.297436,2.0742567,1.9429746,1.6016412,2.0086155,2.9801028,4.1747694,5.080616,2.1956925,1.0338463,1.0010257,1.4276924,1.5688206,1.1782565,2.409026,3.623385,4.33559,5.2020516,3.7054362,5.5565133,7.4174366,9.563898,15.878566,12.005745,10.502565,9.366975,7.1187696,2.7995899,4.906667,7.9294367,10.850462,11.953232,8.832001,6.9743595,6.7150774,5.5630774,3.2164104,1.5589745,1.1848207,2.0118976,3.1376412,4.778667,8.274052,3.6135387,3.2295387,3.4560003,3.3411283,4.6605134,8.976411,11.398565,9.462154,4.7294364,2.7766156,1.7460514,2.156308,2.7536411,2.8192823,2.1792822,1.8412309,1.3883078,1.1224617,1.1716924,1.4736412,1.6705642,2.409026,3.4822567,4.4373336,4.5489235,2.930872,4.2469745,5.2644105,4.4734364,2.1070771,2.5796926,3.3444104,2.8553848,1.3718976,0.9353847,0.5513847,0.47589746,0.4955898,0.7187693,1.585231,1.719795,1.0929232,0.43651286,0.12143591,0.14112821,0.049230773,0.013128206,0.08205129,0.16082053,0.036102567,0.026256412,0.02297436,0.01969231,0.036102567,0.13784617,0.3708718,0.21661541,0.08861539,0.1148718,0.15425642,0.2231795,0.118153855,0.068923086,0.12471796,0.15425642,0.11158975,0.20348719,0.42994875,0.6892308,0.75487185,0.827077,1.0568206,1.0371283,0.7318975,0.45620516,0.65641034,0.90256417,0.9616411,0.7778462,0.47589746,0.54482055,0.6662565,0.636718,0.46276927,0.37743592,0.3708718,0.37743592,0.33805132,0.26912823,0.256,0.24287182,0.29538465,0.33805132,0.4266667,0.77456415,0.94523084,0.77128214,1.2209232,1.9889232,1.529436,2.0118976,2.7306669,2.7634873,1.9790771,1.0502565,0.9616411,0.5284103,0.21661541,0.18051283,0.2855385,0.1148718,0.029538464,0.0,0.0,0.0,0.0,0.009846155,0.036102567,0.06235898,0.06235898,0.07548718,0.14441027,0.18051283,0.17394873,0.21333335,0.26912823,0.29210258,0.30194873,0.31507695,0.3249231,0.318359,0.36430773,0.36102566,0.2986667,0.26912823,0.28225642,0.318359,0.36102566,0.39384618,0.4135385,0.37743592,0.57764107,1.2438976,2.1891284,2.8356924,3.879385,3.8728209,3.817026,4.0992823,4.46359,4.4734364,4.7524104,4.8147697,4.571898,4.322462,3.5971284,3.7087183,4.1846156,4.4701543,3.9581542,3.5774362,3.1934361,2.6617439,1.9692309,1.2242053,0.99774367,0.88943595,0.78769237,0.6859488,0.64000005,0.51856416,0.5349744,0.64000005,0.8041026,1.0338463,1.2176411,1.339077,1.3161026,1.1881026,1.148718,1.2996924,1.3423591,1.332513,1.3489232,1.5097437,1.5360001,1.8740515,2.3236926,2.6289232,2.4746668,2.8160002,3.121231,3.0260515,2.8291285,3.4658465,3.2032824,3.2065644,3.242667,3.0818465,2.4976413,2.9013336,3.045744,2.7536411,2.3171284,2.5107694,2.8356924,2.930872,2.6847181,2.3171284,2.3729234,2.5074873,2.2678976,2.5435898,3.0523078,2.3466668,1.5360001,1.4867693,1.6640002,1.8084104,1.9396925,2.2514873,2.7995899,3.0358977,2.737231,1.9922053,1.4080001,1.3489232,1.7788719,2.3794873,2.5600002,2.6912823,2.6945643,2.537026,2.2711797,2.0611284,1.6508719,1.5163078,1.5130258,1.5819489,1.7755898,1.5688206,1.3095386,1.204513,1.1848207,0.8992821,0.8598975,0.7220513,0.53825647,0.3708718,0.26256412,0.20676924,0.128,0.07876924,0.0951795,0.190359,0.43651286,0.6826667,0.8205129,0.83035904,0.8041026,0.8992821,0.9944616,1.1716924,1.4211283,1.654154,2.15959,2.8291285,3.3411283,3.6594875,4.020513,3.9647183,4.089436,4.44718,5.0149746,5.7009234,6.7314878,7.824411,9.16677,10.325335,10.249847,10.31877,10.843898,11.332924,11.851488,13.013334,13.4629755,13.495796,13.203693,12.58995,11.552821,10.8767185,11.9171295,12.675283,12.432411,11.749744,12.228924,12.058257,11.467488,10.955488,11.283693,11.188514,10.696206,10.712616,11.063796,10.522257,10.118565,10.528821,10.909539,11.109744,11.680821,11.98277,12.248616,12.629334,13.289026,14.401642,16.269129,17.67713,18.20554,17.801847,16.790976,16.121437,15.635694,15.399385,15.172924,14.395078,12.931283,11.926975,11.034257,10.197334,9.636104,9.93477,10.522257,11.408411,12.212514,12.1468725,11.434668,11.050668,11.044104,11.008,10.056206,9.258667,9.4916935,10.118565,10.84718,11.707078,12.228924,12.232206,12.120616,12.041847,11.907283,11.480617,11.116308,10.755282,10.564924,10.909539,10.873437,10.8307705,10.774975,10.561642,9.895386,9.110975,8.493949,7.975385,7.460103,6.8332314,6.7117953,6.6034875,6.488616,6.449231,6.669129,6.554257,6.5050263,6.363898,6.2030773,6.3474874,6.304821,6.0980515,5.7632823,5.402257,5.175795,5.113436,4.7261543,4.4406157,4.420923,4.5489235,4.6933336,4.7360005,4.7950773,5.0182567,5.579488,5.7731285,5.477744,5.2020516,5.1265645,5.080616,4.9493337,4.6769233,4.4701543,4.522667,5.0149746,1.1848207,1.8182565,1.9232821,1.7624617,1.5819489,1.6180514,1.5195899,1.4834872,1.4112822,1.2373334,0.9353847,0.83035904,0.7844103,0.8172308,0.93866676,1.1290257,1.0075898,1.1946667,1.2832822,1.1749744,1.0929232,1.4211283,1.4342566,1.6344616,2.1891284,2.930872,3.4658465,3.6168208,4.076308,4.6933336,4.4832826,4.0303593,3.4264617,3.0884104,3.1442053,3.4560003,3.0982566,2.4746668,1.9889232,1.8051283,1.8674873,1.7066668,1.3357949,1.0469744,0.9288206,0.84348726,0.8795898,0.8992821,0.955077,1.0404103,1.0765129,1.2603078,1.3587693,1.6246156,2.0676925,2.4516926,2.412308,1.6836925,1.0962052,0.92225647,0.8467693,1.017436,1.0010257,0.9911796,1.0535386,1.1355898,1.0601027,1.2012309,1.4769232,1.7526156,1.847795,1.4966155,0.9944616,0.54482055,0.256,0.14769232,0.14112821,0.18051283,0.27241027,0.45620516,0.80738467,0.8598975,0.99774367,0.9911796,0.88287187,1.0010257,1.273436,1.7263591,2.4976413,3.56759,4.7524104,6.048821,7.282872,8.598975,9.944616,11.080206,13.423591,16.466053,20.168207,25.183182,32.866463,35.57744,38.21621,39.909748,40.98298,42.945644,43.966362,43.35262,42.325336,41.98072,43.296825,40.224823,39.719387,40.786053,42.57477,44.35036,47.43549,50.093952,54.07836,58.522263,59.92698,57.780518,54.718365,52.52267,50.848824,47.245132,41.288208,35.83672,31.507694,29.367798,30.949745,32.76144,33.890465,34.546875,34.372925,32.449642,29.489233,26.098873,23.863796,23.233643,23.532309,24.923899,28.609644,32.41026,35.006363,35.94831,37.792824,40.041027,42.003696,43.090054,42.807796,35.925335,28.06154,21.313643,17.178257,16.538258,12.22236,9.688616,8.598975,8.94359,11.0605135,11.926975,13.078976,14.040616,14.739694,15.527386,14.316309,13.735386,14.424617,16.695797,20.535797,20.230566,19.488823,19.912207,21.553232,22.89231,25.419489,28.002464,29.010054,29.666464,34.067696,40.493954,40.76636,39.919594,39.683285,38.482056,39.489643,38.406567,36.26667,34.425438,34.569847,34.60267,33.276722,31.465029,30.024208,29.797747,29.574566,29.919182,29.83713,29.312002,29.305439,31.192617,36.775387,44.78031,54.69211,66.75037,72.47755,76.86893,68.6277,48.479183,29.161028,25.987284,29.732105,37.215183,44.061543,44.704823,37.408825,35.91221,35.981133,32.66626,20.315899,15.087591,10.9686165,8.812308,9.097847,11.907283,16.896002,18.819284,19.40677,18.710976,15.110565,14.8709755,17.51631,19.410053,20.936207,26.50913,25.856003,18.560001,11.858052,11.900719,23.745644,9.596719,2.605949,0.40369233,0.6662565,1.1093334,1.7657437,2.353231,3.242667,4.3027697,4.8836927,3.2098465,2.7700515,2.540308,2.1858463,2.0644104,2.3958976,2.3138463,1.9790771,1.5556924,1.1979488,0.8730257,0.98133343,1.3029745,1.6607181,1.9003079,2.1366155,1.7033848,1.4834872,1.6771283,1.8248206,1.6672822,2.1366155,2.2416413,2.1070771,2.9505644,1.9856411,3.6430771,4.6145644,6.012718,13.364513,11.201642,10.450052,9.711591,7.683283,3.1770258,5.149539,7.77518,10.151385,10.81436,7.7325134,6.3967185,6.265436,5.464616,3.6135387,1.8346668,1.6443079,2.176,3.636513,7.240206,15.205745,5.654975,5.1331286,6.741334,6.5050263,3.3969233,4.778667,8.119796,7.680001,3.9089234,3.4560003,4.1025643,3.0949745,2.3926156,2.9965131,4.955898,3.3312824,2.359795,2.048,1.9954873,1.401436,2.7864618,4.965744,5.661539,4.781949,4.4406157,3.7054362,4.6244106,4.965744,3.9778464,2.3794873,2.8356924,3.5052311,2.8882053,1.7723079,3.2623591,1.4408206,1.6147693,2.1136413,2.537026,3.7710772,1.6738462,0.77128214,0.41682056,0.29210258,0.38400003,0.53825647,0.77128214,0.6235898,0.29538465,0.65969235,0.18707694,0.10502565,0.09189744,0.052512825,0.101743594,0.2100513,0.18051283,0.12143591,0.098461546,0.15097436,0.22646156,0.15097436,0.098461546,0.108307704,0.108307704,0.13128206,0.2297436,0.30851284,0.35446155,0.43651286,0.6071795,1.0010257,1.3029745,1.4178462,1.4473847,1.5425643,1.339077,1.0633847,0.84348726,0.7089231,0.65312827,0.6498462,0.57764107,0.46276927,0.46276927,0.42338464,0.4955898,0.48246157,0.38728207,0.40369233,0.36758977,0.39384618,0.43651286,0.5513847,0.88615394,1.086359,0.9682052,1.1815386,1.6738462,1.6869745,1.8674873,2.172718,2.4582565,2.4057438,1.5392822,1.7394873,1.1782565,0.62030774,0.41025645,0.48246157,0.23958977,0.13784617,0.08861539,0.04594872,0.013128206,0.013128206,0.01969231,0.03938462,0.068923086,0.098461546,0.098461546,0.13128206,0.14769232,0.14769232,0.18379489,0.30194873,0.32820517,0.3446154,0.36102566,0.318359,0.30194873,0.3052308,0.29538465,0.27897438,0.2986667,0.25271797,0.29538465,0.4004103,0.51856416,0.5481026,0.43651286,0.5284103,1.1060513,2.048,2.8225644,3.3444104,3.5741541,3.8006158,4.056616,4.1058464,4.4406157,4.7392826,4.8344617,4.640821,4.125539,3.4592824,3.6430771,4.069744,4.2830772,3.9778464,3.7021542,3.31159,2.878359,2.3466668,1.5360001,1.0469744,0.892718,0.79425645,0.6629744,0.574359,0.5284103,0.5218462,0.62030774,0.8205129,1.0469744,1.0994873,1.3292309,1.4178462,1.3062565,1.214359,1.3259488,1.4802053,1.522872,1.5360001,1.8510771,1.9364104,2.0742567,2.4057438,2.740513,2.5665643,2.477949,2.7175386,2.7142565,2.537026,2.9111798,2.6322052,2.9702566,3.239385,3.0227695,2.166154,2.484513,2.7142565,2.678154,2.4713848,2.4615386,2.4320002,2.3335385,2.1202054,2.0086155,2.477949,2.5337439,2.2646155,2.4352822,2.7011285,1.6147693,1.394872,1.719795,2.1825643,2.4484105,2.2383592,2.7798977,2.7536411,2.4418464,2.0709746,1.8346668,1.7296412,1.3456411,1.3883078,1.9528207,2.5238976,2.9243078,2.858667,2.612513,2.297436,1.8707694,1.719795,1.6475899,1.7001027,1.8116925,1.8248206,1.4572309,1.2176411,1.1191796,1.0699488,0.86317956,0.69907695,0.6662565,0.6071795,0.44307697,0.17066668,0.13784617,0.09189744,0.068923086,0.128,0.35446155,0.5907693,0.8008206,0.86646163,0.7975385,0.7187693,0.90912825,1.0469744,1.1651284,1.3620514,1.7887181,2.2678976,2.9636924,3.383795,3.4658465,3.5872824,3.8137438,3.9942567,4.276513,4.7261543,5.32677,6.6133337,7.9819493,8.999385,9.412924,9.153642,9.826463,10.555078,10.975181,11.1983595,11.815386,13.072412,13.069129,12.491488,11.877745,11.579078,11.1294365,12.242052,13.3251295,13.643488,13.305437,13.266052,12.691693,11.690667,10.742155,10.70277,10.807796,10.581334,10.548513,10.614155,10.082462,9.849437,10.371283,10.9226675,11.247591,11.572514,11.9171295,12.219078,12.563693,13.121642,14.12595,15.707899,16.820515,16.840206,15.986873,15.314053,15.232001,14.8020525,14.201437,13.35795,11.946668,11.296822,10.541949,9.757539,9.229129,9.458873,10.04636,10.729027,11.487181,12.1468725,12.3536415,11.716924,11.293539,11.18195,11.0605135,10.171078,9.632821,10.131693,10.791386,11.234463,11.592206,11.664412,11.72677,11.956513,12.268309,12.33395,11.313231,10.5780525,10.220308,10.233437,10.538668,10.44677,10.729027,11.16554,11.352616,10.679795,9.435898,8.457847,7.709539,7.197539,6.954667,6.885744,6.7282057,6.445949,6.12759,5.98318,5.58277,5.6254363,5.8289237,6.038975,6.232616,6.0192823,6.0028725,5.920821,5.6451287,5.169231,4.955898,4.417641,4.141949,4.345436,4.8607183,4.886975,4.8016415,4.6834874,4.7524104,5.353026,5.4908724,5.110154,4.8016415,4.7556925,4.788513,4.7294364,4.6802053,4.5029745,4.2863593,4.342154,0.90584624,1.2800001,1.2931283,1.2209232,1.2307693,1.3915899,1.3095386,1.211077,1.1027694,0.9682052,0.761436,0.74830776,0.7220513,0.7253334,0.7384616,0.7056411,0.8369231,0.99774367,1.204513,1.4244103,1.5622566,1.3554872,1.1684103,1.204513,1.6016412,2.4418464,3.045744,2.8750772,3.1245131,3.9122055,4.279795,3.8465643,3.5052311,3.4494362,3.6496413,3.876103,3.495385,2.5829747,1.9823592,1.8576412,1.7001027,1.5360001,1.3456411,1.1552821,1.0075898,0.955077,0.9288206,0.8763078,0.892718,0.98461545,1.079795,1.2307693,1.5097437,1.9593848,2.5140514,2.989949,2.5796926,1.6475899,1.0075898,0.9485129,1.2406155,1.4572309,1.3259488,1.1716924,1.148718,1.2307693,1.1552821,1.1881026,1.2340513,1.273436,1.3718976,1.4244103,1.3981539,1.1881026,0.7844103,0.26584616,0.20676924,0.2855385,0.41025645,0.50543594,0.49887183,0.99774367,1.0962052,1.204513,1.4572309,1.723077,1.8970258,2.2547693,2.802872,3.6135387,4.818052,6.0849237,7.2927184,8.930462,10.755282,11.795693,14.322873,16.544823,19.580719,23.706259,28.366772,35.13108,39.473232,41.698463,43.582363,48.351185,49.887184,45.600822,41.16677,39.67672,41.629543,42.880005,44.058258,45.4958,47.478157,50.21867,53.63857,57.73785,62.880825,67.96472,70.42298,68.75242,66.50093,63.996723,60.563698,54.52144,46.72985,40.595695,35.82031,32.758156,32.449642,30.74626,30.500105,31.235285,32.324924,32.978054,31.363285,28.98708,26.36472,23.896618,21.858463,22.810259,25.62954,28.14031,29.495796,30.175182,33.158566,37.618874,42.725746,47.360004,50.13334,42.30236,33.29313,25.376822,19.895796,17.266872,12.662155,10.354873,9.888822,10.781539,12.524308,12.931283,13.161027,13.397334,13.6008215,13.525334,13.24636,13.906053,15.91795,17.923283,16.777847,15.96718,15.993437,17.414566,19.616821,20.804924,21.605745,23.995079,25.672207,27.083488,31.428925,43.664413,48.357746,46.739697,42.003696,39.312412,39.35836,37.78626,35.249233,32.98462,32.81067,34.166157,32.935387,30.9399,29.630362,30.076721,28.78031,28.294567,28.081232,27.910566,27.867899,31.573336,38.672413,46.063595,52.752415,59.86134,65.664,73.48185,69.805954,52.630978,31.461746,28.20267,33.184822,40.953438,46.53621,45.44985,37.684517,36.5719,36.43077,31.721027,17.079796,12.324103,8.648206,6.688821,6.9120007,9.632821,14.874257,17.214361,17.70995,16.935387,14.998976,14.034052,14.437745,15.648822,18.36636,24.556309,20.788515,16.866463,11.52,14.004514,44.07139,14.188309,3.1573336,0.7581539,0.702359,0.6268718,0.92225647,1.3981539,2.4451284,3.6430771,3.7710772,2.8849232,2.28759,1.9626669,1.9495386,2.349949,2.0578463,1.9823592,1.723077,1.2209232,0.76800007,0.49887183,0.43651286,0.5284103,0.69251287,0.8008206,3.1442053,2.993231,2.225231,1.8445129,1.972513,2.3827693,2.861949,2.6584618,1.9954873,2.1103592,1.4276924,3.1737437,3.9056413,4.6080003,10.692924,9.993847,8.812308,6.636308,4.125539,3.1409233,5.5171285,6.688821,7.4929237,7.837539,6.7183595,7.020308,7.13518,5.9569235,3.7809234,2.3040001,2.5600002,2.3991797,3.639795,7.8112826,16.17395,5.937231,6.0816417,9.524513,10.180923,2.9735386,3.4198978,6.308103,6.75118,4.8344617,5.6254363,7.5191803,5.1659493,2.8816411,3.3476925,7.6143594,5.0182567,3.8596926,3.817026,3.9187696,2.540308,3.9384618,8.185436,9.682052,7.9195905,7.463385,5.87159,4.663795,3.9778464,3.8301542,4.1058464,4.4767184,3.3476925,2.100513,2.3893335,6.1440005,2.7700515,4.073026,5.428513,5.5991797,6.7577443,2.6518977,1.7033848,1.2964103,0.6465641,0.7811283,1.4080001,2.3401027,1.8281027,0.48246157,1.2570257,0.3314872,0.17723078,0.16082053,0.052512825,0.009846155,0.07548718,0.13784617,0.128,0.07876924,0.14441027,0.17723078,0.18379489,0.15753847,0.128,0.15753847,0.2855385,0.380718,0.4004103,0.36102566,0.31507695,0.508718,0.96492314,1.6016412,2.300718,2.8947694,2.7306669,2.03159,1.3062565,0.8960001,0.9944616,0.9353847,0.6662565,0.48902568,0.46933338,0.43323082,0.4397949,0.6071795,0.61374366,0.49230772,0.6268718,0.49887183,0.44964105,0.50543594,0.65641034,0.84348726,1.1290257,1.2832822,1.1618463,1.0535386,1.657436,2.2088206,2.3893335,2.477949,2.4746668,2.1202054,2.6617439,2.1202054,1.4145643,0.9485129,0.6071795,0.4201026,0.47589746,0.44307697,0.25928208,0.108307704,0.118153855,0.098461546,0.08861539,0.11158975,0.18051283,0.14441027,0.12471796,0.118153855,0.13456412,0.17394873,0.26584616,0.318359,0.38728207,0.43323082,0.318359,0.2986667,0.28882053,0.27897438,0.28225642,0.32164106,0.2297436,0.24287182,0.3708718,0.5481026,0.64000005,0.5284103,0.5021539,0.9485129,1.7985642,2.5173335,2.878359,3.3805132,3.698872,3.7251284,3.564308,4.0041027,4.598154,5.037949,5.080616,4.5554876,3.4658465,3.3542566,3.6890259,4.0303593,4.010667,3.8990772,3.639795,3.436308,3.0851285,1.9692309,1.0666667,0.8566154,0.8172308,0.69579494,0.47917953,0.5021539,0.55794877,0.6826667,0.82379496,0.86317956,0.9517949,1.1520001,1.2406155,1.1913847,1.1848207,1.2996924,1.6902566,1.8084104,1.719795,2.103795,2.359795,2.3171284,2.353231,2.550154,2.6847181,2.0873847,2.0151796,2.103795,2.2153847,2.4516926,2.3105643,2.8947694,3.0391798,2.5173335,2.0250258,2.28759,2.2514873,2.1891284,2.2088206,2.2646155,1.6147693,1.4473847,1.5031796,1.7296412,2.2580514,2.4057438,2.425436,2.4516926,2.281026,1.3522053,1.6246156,2.1431797,2.7798977,3.0916924,2.3138463,2.9997952,2.556718,1.8609232,1.4572309,1.5622566,2.225231,1.7788719,1.339077,1.4802053,2.2580514,2.9013336,2.934154,2.6354873,2.1858463,1.6705642,1.7460514,1.8707694,1.9889232,2.0118976,1.8018463,1.2996924,1.1191796,1.0633847,1.024,0.9878975,0.61374366,0.5152821,0.5481026,0.52512825,0.20348719,0.0951795,0.04594872,0.07876924,0.22646156,0.54482055,0.6432821,0.8336411,0.90912825,0.8336411,0.7318975,0.9189744,1.0502565,1.1257436,1.2668719,1.7033848,2.231795,2.9702566,3.4822567,3.6594875,3.7152824,4.066462,4.391385,4.673641,4.9329233,5.21518,6.488616,7.5913854,7.9917955,7.8834877,8.149334,9.199591,10.213744,10.630565,10.587898,10.939077,12.452104,12.360206,11.861334,11.444513,10.909539,10.450052,11.099898,12.005745,12.678565,12.987078,13.75836,13.164309,12.035283,11.0145645,10.545232,10.571488,10.962052,11.004719,10.522257,9.875693,9.77395,10.31877,10.827488,11.093334,11.37559,12.097642,12.4685135,12.645744,13.00677,14.162052,15.0777445,15.55036,15.05477,14.020925,13.804309,14.080001,13.8765135,13.1872835,12.025436,10.41395,10.164514,9.77395,9.557334,9.754257,10.545232,10.8307705,11.113027,11.405129,11.772718,12.33395,11.628308,11.32636,11.21477,11.047385,10.538668,10.637129,11.395283,11.940104,12.002462,11.913847,11.795693,11.661129,11.841642,12.173129,11.98277,10.610872,9.974154,9.77395,9.826463,10.036513,9.849437,10.522257,11.460924,12.009027,11.460924,9.961026,8.749949,7.972103,7.5913854,7.3714876,7.125334,6.931693,6.485334,5.796103,5.156103,5.2348723,5.5204105,5.832206,6.0258465,5.9634876,5.6451287,5.654975,5.677949,5.5302567,5.152821,4.8804107,4.309334,4.197744,4.578462,4.772103,4.5554876,4.5095387,4.525949,4.604718,4.8377438,5.0182567,4.9460516,4.8311796,4.7556925,4.6966157,4.775385,4.7622566,4.5128207,4.069744,3.6562054,0.9321026,1.1388719,1.4834872,1.6049232,1.4408206,1.2209232,1.0633847,0.9485129,0.9189744,0.9321026,0.86974365,0.80738467,0.79425645,0.7515898,0.67938465,0.65641034,0.6301539,0.67938465,0.98461545,1.5885129,2.3794873,1.8806155,1.9298463,1.5688206,1.0371283,1.7690258,2.356513,2.428718,2.6486156,3.2295387,3.9351797,3.876103,3.761231,3.4724104,3.0818465,2.8389745,2.546872,2.1234872,1.972513,2.1267693,2.2744617,2.041436,1.7558975,1.5097437,1.3226668,1.1126155,0.97805136,0.9353847,0.9189744,1.020718,1.4966155,1.5195899,1.8084104,2.1333334,2.172718,1.5261539,1.3784616,1.2242053,1.1684103,1.2996924,1.6771283,1.5064616,1.3653334,1.3259488,1.3029745,1.020718,0.75487185,0.761436,0.8336411,0.92225647,1.1290257,1.2865642,1.719795,2.0644104,1.8642052,0.5940513,0.3511795,0.35446155,0.39712822,0.49887183,0.9156924,1.6475899,1.6935385,2.0611284,2.8356924,3.190154,2.4943593,2.4582565,2.7569232,3.3903592,4.6834874,5.648411,6.9710774,8.854975,10.916103,12.160001,15.419078,17.929848,21.658258,25.557335,25.557335,27.451078,30.953028,34.54359,40.40534,54.442673,59.483902,52.880413,46.070156,43.27713,41.517952,45.814156,49.316105,54.24903,59.264004,59.4478,63.4158,66.82257,70.44267,73.83959,75.378876,73.1799,72.18216,70.57724,67.64308,63.75057,57.40308,51.59385,46.408207,41.701748,37.123283,32.32821,29.709131,28.04185,27.16554,27.986053,28.947695,29.170874,28.274874,26.144823,22.934977,24.897642,25.957747,26.04308,25.183182,23.499489,25.232412,28.66872,34.271183,41.186466,47.241848,42.210464,36.42421,29.285746,22.111181,18.097233,13.922462,12.327386,12.340514,13.111795,13.915898,12.780309,11.418258,10.341744,10.203898,11.779283,12.097642,13.548308,15.875283,17.329231,14.680616,13.164309,13.446565,15.599591,18.766771,21.13313,22.071796,25.37354,27.083488,27.608618,31.72431,49.48349,64.15098,63.0679,49.650875,43.365746,42.62072,38.14072,33.490055,30.943182,31.478157,33.040413,30.739695,28.261745,27.608618,29.09867,27.109745,27.19836,27.470772,27.40513,27.831797,33.860924,41.330875,48.082054,52.47344,53.392414,56.136208,66.254776,68.91324,57.744415,34.819286,32.098465,35.977848,41.366978,45.072414,45.791183,38.114464,36.066463,35.46913,31.215591,17.286566,11.867898,8.041026,6.117744,6.055385,7.4469748,12.560411,15.589745,16.25272,15.366566,14.815181,11.641437,10.420513,11.641437,14.9398985,19.088411,15.8654375,13.594257,8.999385,4.772103,9.5835905,3.5413337,2.4976413,2.5206156,1.8576412,0.9321026,0.892718,0.92225647,1.4900514,2.3696413,2.6256413,2.3926156,1.9856411,1.7493335,1.8871796,2.4713848,2.5206156,2.0939488,1.4539489,0.8533334,0.5481026,0.28225642,0.4135385,0.6826667,0.8369231,0.64000005,2.9965131,3.367385,3.239385,3.131077,2.5928206,2.3991797,2.7437952,2.665026,2.0512822,1.6475899,1.014154,2.7503593,4.1156926,6.0061545,12.937847,14.221129,11.940104,6.9842057,2.4451284,3.6168208,3.9811285,5.346462,7.1581545,8.461129,7.890052,9.061745,8.5202055,6.6592827,4.391385,3.1573336,2.8291285,2.0217438,1.6278975,1.8281027,2.1234872,2.3171284,5.477744,5.917539,3.6562054,4.4242053,4.266667,6.9809237,8.214975,7.197539,6.7610264,6.173539,5.110154,3.9712822,3.7185643,5.904411,6.550975,5.733744,5.668103,6.23918,5.0215387,3.6529233,7.778462,9.970873,9.442462,12.0549755,9.465437,7.584821,6.380308,6.0849237,7.171283,10.052924,5.609026,2.0742567,2.3958976,4.2272825,3.383795,8.044309,9.947898,8.27077,9.613129,6.0356927,5.0510774,3.2918978,0.6465641,0.24287182,1.7690258,4.010667,3.6791797,1.0732309,0.06235898,0.02297436,0.02297436,0.02297436,0.02297436,0.04594872,0.2297436,0.14769232,0.04266667,0.02297436,0.04594872,0.26584616,0.3117949,0.28225642,0.26912823,0.36758977,0.46276927,0.43323082,0.446359,0.4594872,0.2297436,0.37415388,1.1979488,2.1891284,2.858667,2.7634873,3.006359,2.4615386,1.8576412,1.4834872,1.1913847,1.142154,0.9189744,0.7187693,0.5907693,0.45620516,0.54482055,0.65641034,0.6629744,0.61374366,0.74830776,0.60061544,0.58420515,0.6268718,0.7089231,0.8533334,1.1585642,1.6836925,1.5064616,0.98461545,1.7558975,1.8281027,2.103795,2.1202054,1.913436,1.9987694,2.2678976,2.6354873,2.7470772,2.281026,0.9616411,0.86317956,1.3062565,1.3423591,0.827077,0.4135385,0.47261542,0.4135385,0.3117949,0.23958977,0.28882053,0.25271797,0.190359,0.14769232,0.13784617,0.13784617,0.2100513,0.29210258,0.3708718,0.39056414,0.24287182,0.3052308,0.42994875,0.47917953,0.44307697,0.44307697,0.380718,0.29210258,0.29210258,0.38400003,0.45620516,0.43323082,0.43651286,0.7417436,1.467077,2.5796926,3.4100516,4.1025643,4.082872,3.7218463,4.332308,3.6004105,4.1517954,4.785231,4.95918,4.775385,3.56759,3.2656412,3.4592824,3.764513,3.8137438,3.948308,3.7251284,3.56759,3.2853336,2.0906668,1.1520001,0.86974365,0.80738467,0.7122052,0.5021539,0.4660513,0.5677949,0.7450257,0.86317956,0.7187693,0.86317956,1.020718,1.142154,1.2209232,1.2832822,1.2832822,1.585231,1.9003079,2.1267693,2.3335385,2.934154,2.8455386,2.612513,2.612513,3.0523078,2.550154,2.1234872,1.8806155,1.7788719,1.6311796,1.9626669,2.4943593,2.5107694,2.1497438,2.3794873,2.4155898,2.3269746,2.0808206,1.9232821,2.349949,1.5425643,1.3883078,1.4572309,1.6246156,2.0742567,2.038154,1.6804104,1.401436,1.401436,1.6935385,2.6223593,3.1277952,3.6758976,3.7054362,1.6180514,1.9232821,2.9965131,2.8389745,1.5753847,1.463795,2.0873847,2.0512822,1.719795,1.4769232,1.7099489,2.0873847,2.6486156,2.789744,2.4615386,2.1825643,1.8904617,1.9987694,2.0611284,1.847795,1.3718976,1.1651284,1.086359,0.97805136,0.86646163,0.97805136,0.76800007,0.5349744,0.42994875,0.4135385,0.2297436,0.068923086,0.03938462,0.15097436,0.3708718,0.64000005,0.60389745,0.7975385,0.9124103,0.8795898,0.8533334,0.86646163,0.9156924,0.97805136,1.142154,1.6180514,2.0217438,2.5796926,3.114667,3.5446157,3.8596926,4.3618464,4.706462,4.9920006,5.277539,5.5696416,6.5706673,6.738052,6.774154,7.1122055,7.90318,9.199591,10.134975,10.433641,10.315488,10.499283,11.864616,12.242052,12.012309,11.411694,10.545232,10.384411,10.765129,11.638155,12.694975,13.367796,13.8075905,12.642463,11.349334,10.66995,10.620719,11.23118,11.913847,11.884309,11.0605135,10.069334,10.144821,10.052924,10.210463,10.742155,11.474052,12.87877,12.898462,12.882052,13.285745,13.686155,13.820719,13.929027,14.099693,14.267078,14.204719,13.791181,13.4859495,12.754052,11.401847,9.5835905,9.521232,9.6525135,10.220308,11.204924,12.327386,11.9860525,11.680821,11.730052,12.07795,12.297847,11.848206,11.651283,11.536411,11.45436,11.490462,12.087796,13.154463,13.801026,13.732103,13.243078,13.08554,12.560411,12.248616,11.959796,10.725744,9.77395,9.4916935,9.081436,8.720411,9.537642,9.865847,10.837335,11.910565,12.475078,11.841642,10.778257,9.55077,8.746667,8.5202055,8.605539,7.6176414,7.141744,6.4590774,5.4613338,4.670359,5.2053337,5.7796926,5.937231,5.7074876,5.586052,5.4613338,5.395693,5.290667,5.106872,4.8377438,4.788513,4.391385,4.342154,4.6145644,4.457026,4.1517954,4.1485133,4.33559,4.5817437,4.716308,4.8377438,4.9493337,4.900103,4.7589746,4.8049235,4.7589746,4.5522056,4.089436,3.498667,3.1442053,1.4572309,1.2635899,1.2504616,1.2570257,1.2209232,1.1946667,1.0568206,1.0305642,1.0666667,1.0929232,1.0043077,0.892718,0.83035904,0.7975385,0.7581539,0.65641034,0.58420515,0.71548724,0.92553854,1.2537436,1.8937438,2.1431797,1.9626669,1.3423591,0.72861546,1.0010257,2.0939488,2.1202054,2.2514873,2.865231,3.5347695,3.754667,3.9220517,3.5872824,2.806154,2.1431797,2.356513,2.7733335,3.446154,4.325744,5.2512827,4.7556925,3.4822567,2.300718,1.5688206,1.1388719,1.3062565,1.4933335,1.4605129,1.2209232,1.0305642,1.4276924,2.1530259,2.359795,1.7788719,0.7318975,0.8205129,1.1913847,1.3718976,1.2242053,0.95835906,0.78769237,0.67282057,0.81394875,1.0502565,0.88943595,1.0404103,1.0272821,0.92225647,0.8402052,0.92225647,1.1585642,1.3981539,1.7263591,1.8871796,1.2898463,0.7450257,0.72861546,0.79097444,0.7778462,0.83035904,1.4539489,2.4910772,3.2918978,3.387077,2.481231,2.4681027,2.6912823,3.2623591,4.161641,5.221744,6.009436,7.250052,9.347282,12.100924,14.713437,17.864206,20.214155,22.78072,25.225847,25.85272,27.684105,31.01867,40.146053,53.1758,62.047184,61.1118,53.79939,46.053745,40.84185,38.12431,42.607594,49.778877,58.2958,65.67385,68.29621,78.24083,85.80267,90.11529,93.689445,102.41642,116.847595,116.713036,105.03878,88.933754,79.58318,68.42093,60.88862,55.676723,51.37067,46.46072,39.663593,36.053337,32.518566,28.74749,27.250874,24.848412,23.729233,23.535591,24.090258,25.399797,25.032207,24.992823,24.33313,22.918566,21.448206,21.90113,23.062977,26.312206,31.120413,35.0359,30.710155,25.842875,20.969027,16.676104,13.617231,12.058257,11.831796,12.219078,12.47836,11.828514,11.904001,11.546257,9.993847,8.096821,8.326565,6.8955903,7.194257,8.454565,9.449026,8.490667,7.748924,9.019077,13.610668,20.233849,25.002668,26.597746,32.800823,39.87036,44.26831,42.660107,59.103184,77.36452,76.79672,57.626263,40.960003,42.246567,38.150566,32.26913,27.789131,27.474054,29.817438,28.468515,26.151386,24.881233,25.947899,26.138258,27.3559,28.534157,29.909336,33.030567,40.1559,46.73313,50.852108,51.646362,49.28985,49.89703,58.58462,64.301956,58.876724,37.00513,34.448414,37.123283,41.16021,44.52103,46.998978,39.42072,35.44944,33.14544,28.983797,17.851078,10.272821,6.8365135,5.786257,5.9963083,6.957949,10.47959,13.065847,13.774771,12.452104,9.714872,8.805744,9.137232,10.729027,12.87877,14.158771,11.168821,7.748924,8.211693,12.448821,15.931078,5.425231,3.2656412,3.1474874,2.2580514,1.2603078,1.0765129,0.8566154,1.0436924,1.4998976,1.5130258,1.6935385,1.6443079,1.6804104,1.7526156,1.4572309,1.9462565,1.9528207,1.467077,0.76800007,0.40369233,0.41682056,0.5940513,0.7089231,0.7318975,0.8008206,1.2307693,1.595077,1.9856411,2.1825643,1.6672822,2.3204105,3.2361028,3.318154,2.5271797,1.8806155,0.84348726,1.3883078,2.4451284,4.962462,11.913847,13.751796,13.686155,10.86359,6.633026,4.5456414,5.543385,8.648206,10.614155,10.381129,9.084719,9.104411,7.64718,5.677949,3.9089234,2.793026,2.5993848,2.1792822,1.8740515,2.0906668,3.2918978,9.787078,9.366975,8.162462,7.213949,2.484513,2.4024618,4.2240005,5.5696416,5.481026,4.417641,5.2644105,10.056206,10.325335,6.2916927,6.8562055,8.940309,7.9228725,7.394462,7.8769236,6.8496413,7.0367184,6.314667,6.7314878,8.618668,10.564924,12.819694,13.482668,12.914873,12.409437,14.178463,11.588924,7.282872,6.11118,7.427283,5.0674877,14.001232,10.04636,5.421949,7.066257,16.630156,7.604513,4.073026,2.1103592,1.3489232,4.969026,2.0020514,1.2373334,0.92225647,0.39712822,0.098461546,0.06235898,0.032820515,0.02297436,0.03938462,0.08205129,0.22646156,0.17723078,0.08861539,0.04266667,0.059076928,0.20020515,0.32820517,0.44964105,0.55794877,0.63343596,0.5284103,0.29210258,0.2297436,0.33805132,0.30194873,0.23302566,0.6170257,1.0075898,1.2570257,1.4802053,1.8609232,2.0709746,2.0808206,1.9528207,1.8379488,2.4418464,2.2744617,1.5458462,0.76800007,0.7515898,0.4660513,0.43323082,0.44964105,0.5284103,0.90584624,0.7220513,0.7581539,0.88943595,0.9288206,0.63343596,0.9485129,1.1979488,1.148718,1.017436,1.4736412,1.595077,1.4441026,1.595077,2.2482052,3.2328207,4.2141542,3.7120004,3.2820516,3.3017437,2.9997952,2.0020514,1.847795,1.8707694,1.6246156,0.88943595,0.7056411,0.6071795,0.47917953,0.3249231,0.26584616,0.25928208,0.29538465,0.2986667,0.26584616,0.28225642,0.4266667,0.4660513,0.47261542,0.42994875,0.24287182,0.29538465,0.38728207,0.41682056,0.43323082,0.636718,0.47917953,0.27897438,0.16738462,0.17066668,0.22646156,0.28882053,0.39384618,0.60389745,1.020718,1.8084104,3.0884104,3.1409233,2.878359,3.0720003,4.345436,3.387077,3.692308,4.4274874,4.8836927,4.44718,3.4724104,3.3312824,3.6890259,4.07959,3.9253337,3.7842054,3.1573336,2.550154,2.0676925,1.4178462,0.93866676,0.80738467,0.80738467,0.7515898,0.5152821,0.39056414,0.41025645,0.58420515,0.77456415,0.7187693,0.7450257,0.8008206,0.9321026,1.1158975,1.2438976,1.0699488,1.2996924,1.8149745,2.409026,2.7733335,3.058872,3.1573336,3.0523078,2.8422565,2.733949,2.0775387,1.7723079,1.719795,1.7460514,1.6082052,2.1136413,2.7470772,2.7700515,2.3466668,2.540308,2.1464617,2.1891284,2.1431797,2.0020514,2.2514873,1.8084104,1.4867693,1.2406155,1.0994873,1.1716924,1.2340513,1.2603078,1.1946667,1.0371283,0.85005134,2.28759,2.9046156,3.190154,3.2886157,3.0096412,2.2383592,2.4320002,2.2088206,1.5524104,1.7952822,2.1431797,1.913436,1.7165129,1.8838975,2.4648206,2.7273848,2.9144619,2.8356924,2.5009232,2.1333334,1.975795,2.0775387,2.1333334,1.9528207,1.4572309,1.2603078,1.3161026,1.2996924,1.083077,0.7318975,0.7581539,0.56123084,0.35446155,0.2297436,0.14441027,0.052512825,0.08205129,0.25271797,0.5316923,0.8467693,0.8795898,0.86317956,0.827077,0.8336411,0.96492314,0.9485129,0.9517949,1.0994873,1.4145643,1.8116925,1.9035898,2.733949,3.4100516,3.5872824,3.495385,3.945026,4.138667,4.4767184,5.0609236,5.717334,6.422975,6.701949,7.069539,7.6143594,7.9885135,9.330873,10.568206,11.119591,11.050668,11.047385,12.199386,12.071385,11.526565,11.116308,11.067078,11.30995,12.547283,13.262771,13.400617,14.355694,13.203693,11.972924,11.323078,11.1983595,10.827488,11.290257,12.173129,12.018872,10.748719,9.632821,9.803488,10.203898,10.587898,10.794667,10.765129,12.179693,12.130463,11.88759,12.2387705,13.492514,13.636924,13.5318985,13.820719,14.388514,14.375385,14.332719,13.952001,12.918155,11.349334,9.813334,9.42277,9.80677,10.528821,11.336206,12.1468725,11.460924,11.424822,11.569232,11.638155,11.565949,11.493745,11.776001,11.684103,11.264001,11.319796,12.317539,13.233232,13.988104,14.424617,14.306462,13.689437,12.777026,11.933539,11.191795,10.249847,9.816616,9.40636,9.025641,9.055181,10.243283,10.466462,10.610872,11.329642,12.196103,11.707078,10.624001,9.911796,9.127385,8.4972315,8.923898,8.28718,7.3780518,6.5706673,5.920821,5.156103,5.546667,5.924103,5.9470773,5.7009234,5.7074876,5.586052,5.474462,5.3760004,5.290667,5.228308,4.44718,4.1878977,4.2371287,4.338872,4.197744,4.2371287,4.20759,4.348718,4.571898,4.4701543,4.2207184,4.2141542,4.1878977,4.138667,4.2929235,4.0992823,3.5282054,3.0260515,2.8882053,3.2787695,1.2668719,1.1355898,1.1520001,1.2176411,1.2504616,1.1716924,1.0535386,1.0601027,1.086359,1.0633847,0.96492314,0.9288206,0.95835906,0.97805136,0.92553854,0.72861546,0.6662565,0.69251287,0.79097444,1.0075898,1.467077,1.9954873,1.9987694,1.4145643,0.79097444,1.2931283,1.6804104,1.7690258,1.9889232,2.4746668,3.0752823,3.6627696,3.698872,3.4264617,2.9997952,2.481231,2.3991797,2.4451284,2.8127182,3.4888208,4.266667,3.8498464,2.8488207,2.038154,1.657436,1.4112822,1.4276924,1.4178462,1.2307693,0.8992821,0.6301539,1.3456411,2.0873847,2.1300514,1.463795,0.761436,0.85005134,1.0469744,1.0633847,0.8763078,0.7515898,0.50543594,0.40369233,0.508718,0.74830776,0.892718,1.1552821,1.1060513,1.0436924,1.1093334,1.2832822,1.522872,1.6016412,1.6869745,1.7591796,1.6016412,1.5064616,1.3554872,1.2274873,1.1782565,1.2570257,1.9298463,3.7874875,4.9821544,4.8114877,3.7218463,4.2174363,4.1124105,4.8016415,6.298257,7.240206,8.960001,9.67877,11.680821,15.635694,20.60472,22.688822,22.596926,23.341951,25.03877,24.917336,26.633848,31.868721,44.100925,56.963287,54.245747,53.536823,51.698875,47.520824,41.606567,36.397953,46.434464,61.206978,75.65457,86.20637,90.78811,99.48554,102.69539,104.53006,113.1717,140.85909,166.84637,152.17888,123.12288,98.85867,91.45108,86.974365,81.906876,75.204926,67.14093,59.30667,54.63631,49.19467,43.181953,37.2119,32.324924,28.593233,26.148104,25.193027,25.573746,26.74872,27.27713,27.56595,27.19508,25.412926,21.126566,20.184616,19.761232,21.221745,24.12308,26.213745,23.112207,18.996513,15.163078,12.212514,10.043077,9.4916935,9.905231,10.420513,11.168821,13.275898,22.787283,27.250874,22.186668,12.642463,13.22995,6.0291286,4.388103,5.0642056,5.9930263,6.2851286,7.030154,8.966565,13.328411,19.085129,22.94154,27.040823,41.869133,62.464005,75.648,60.04185,66.66503,78.99898,73.82647,51.734978,37.10031,39.699696,33.969234,26.82749,22.488617,22.44595,24.920618,27.057232,26.532104,24.425028,25.235695,26.942362,29.587694,32.036106,34.326977,37.69108,44.47508,49.618053,51.656208,50.149746,45.699287,46.07344,53.425236,60.66216,59.116314,38.55754,36.88698,38.964516,42.450054,46.2999,50.799595,41.38339,34.422157,30.10954,25.737848,15.721026,8.402052,5.504,4.95918,5.366154,5.9930263,7.076103,9.110975,9.984001,8.940309,6.5706673,6.088206,9.665642,12.156719,13.259488,17.473642,7.79159,10.348309,11.933539,9.301334,9.176616,4.0008206,2.9472823,4.594872,5.904411,2.2383592,1.522872,0.955077,0.84348726,1.014154,0.8041026,1.2537436,1.7526156,2.1530259,2.0939488,0.9944616,1.3883078,1.5327181,1.2635899,0.7089231,0.29210258,0.508718,0.69579494,0.7122052,0.69251287,1.0305642,1.1815386,1.5753847,2.0709746,2.3893335,2.1497438,2.356513,2.6223593,2.6847181,2.4681027,2.1103592,1.6278975,3.4330258,3.9318976,3.5774362,6.889026,15.228719,16.531694,14.55918,11.385437,7.4043083,7.860513,12.356924,13.528616,10.742155,10.069334,9.7214365,8.772923,7.0400004,4.9788723,3.6791797,3.3903592,4.0500517,4.3290257,4.7261543,7.568411,6.921847,6.124308,5.691077,4.896821,1.7887181,2.9505644,8.241231,8.234667,3.6463592,5.3398976,5.5893335,8.218257,8.841846,7.3058467,7.6898465,8.841846,7.27959,5.737026,5.1298466,4.571898,5.730462,6.370462,7.90318,9.642668,8.809027,12.694975,13.810873,14.444309,14.834873,13.164309,10.052924,7.9491286,7.893334,8.467693,5.802667,19.396925,12.2387705,7.640616,12.540719,17.499899,7.4240007,3.0096412,1.142154,1.1782565,4.9394875,1.6804104,1.6213335,1.3587693,0.18379489,0.108307704,0.1148718,0.06564103,0.04266667,0.07548718,0.14769232,2.484513,1.3161026,0.118153855,0.08205129,0.1148718,0.19364104,0.26584616,0.36758977,0.53825647,0.83035904,0.60389745,0.27569234,0.14112821,0.256,0.42994875,0.17066668,0.2297436,0.3446154,0.4397949,0.6301539,1.0075898,1.8346668,2.4976413,2.789744,2.9144619,2.3204105,1.8970258,1.3587693,0.764718,0.5218462,0.40697438,0.4004103,0.4201026,0.53825647,1.0010257,0.7844103,0.7515898,0.8008206,0.90584624,1.148718,1.2603078,1.1355898,1.4145643,1.9167181,1.6508719,1.5721027,1.1684103,1.3981539,2.1825643,2.3860514,2.9472823,2.9636924,2.9636924,3.2262566,3.7940516,3.0326157,2.3171284,2.0545642,1.9659488,1.0896411,1.3423591,0.9616411,0.7187693,0.77456415,0.6432821,0.92225647,0.7811283,0.57764107,0.48902568,0.5218462,0.61374366,0.58420515,0.5021539,0.4266667,0.4004103,0.4135385,0.4004103,0.380718,0.4004103,0.5316923,0.44964105,0.37743592,0.27897438,0.19364104,0.23958977,0.2986667,0.37743592,0.56123084,0.92225647,1.5360001,2.5173335,2.8324106,2.9997952,3.387077,4.2207184,2.6715899,3.1803079,4.325744,5.0149746,4.4996924,3.6890259,3.058872,3.0293336,3.4560003,3.6135387,3.318154,2.737231,2.3236926,2.0742567,1.5261539,1.0633847,0.8763078,0.8008206,0.7089231,0.49887183,0.44307697,0.4955898,0.67938465,0.8795898,0.86317956,0.81394875,0.86646163,0.9911796,1.1093334,1.0699488,0.955077,1.2274873,1.7690258,2.4155898,2.9571285,3.2229745,3.4297438,3.4888208,3.2951798,2.7273848,2.422154,2.15959,1.8379488,1.5261539,1.463795,2.1398976,2.6584618,2.9210258,2.92759,2.789744,2.487795,2.0151796,1.7493335,1.8248206,2.1366155,1.7296412,1.591795,1.4867693,1.401436,1.522872,1.3587693,1.5392822,1.5130258,1.2209232,1.0994873,2.1497438,2.9472823,2.9144619,2.2744617,2.0676925,1.9790771,1.9692309,1.7657437,1.719795,2.7831798,3.186872,2.9243078,2.6617439,2.7109745,3.0293336,2.9243078,2.9407182,2.7175386,2.300718,2.1300514,2.1530259,2.1136413,2.169436,2.176,1.6902566,1.3850257,1.4080001,1.404718,1.1782565,0.7089231,0.65312827,0.5021539,0.32164106,0.17394873,0.11158975,0.055794876,0.12471796,0.2986667,0.5284103,0.761436,0.92225647,0.86646163,0.7811283,0.7450257,0.761436,0.9517949,0.95835906,1.0633847,1.3784616,1.8510771,1.9462565,2.5140514,3.114667,3.4166157,3.1934361,3.3312824,3.511795,3.9548721,4.6867695,5.533539,6.2916927,6.678975,7.2205133,7.9130263,8.211693,9.419488,11.0605135,11.910565,11.785847,11.523283,12.189539,12.189539,11.638155,10.955488,10.850462,11.385437,12.685129,13.361232,13.285745,13.587693,13.6697445,13.262771,12.448821,11.510155,10.935796,10.9456415,11.096616,10.765129,9.898667,9.009232,9.488411,9.8592825,10.299078,10.725744,10.801231,11.45436,11.428103,11.293539,11.648001,13.111795,14.168616,14.234258,14.188309,14.39836,14.713437,14.240822,13.705847,12.6063595,11.178667,10.394258,10.650257,10.886565,11.050668,11.132719,11.175385,10.781539,10.857026,11.07036,11.208206,11.172104,11.431385,11.736616,11.588924,11.122872,11.113027,11.798975,12.324103,13.174155,14.257232,14.884104,13.896206,12.593232,11.316514,10.325335,9.810052,9.8592825,9.547488,9.380103,9.609847,10.240001,10.04636,9.941334,10.328616,11.116308,11.720206,10.57477,9.6754875,9.133949,8.802463,8.251078,8.155898,7.381334,6.4754877,5.730462,5.169231,5.5105643,5.687795,5.6943593,5.605744,5.5893335,5.8847184,5.7140517,5.2512827,4.827898,4.9394875,4.263385,3.9778464,3.9417439,4.023795,4.1091285,4.1058464,4.1058464,4.082872,4.069744,4.1550775,3.6069746,3.7185643,4.086154,4.378257,4.348718,3.9122055,3.4330258,3.2196925,3.255795,3.2295387,1.3522053,1.1027694,1.1552821,1.3095386,1.394872,1.2931283,1.2471796,1.2012309,1.1684103,1.1257436,1.0075898,1.0305642,1.1158975,1.079795,0.892718,0.6695385,0.6498462,0.67610264,0.7318975,0.8763078,1.2406155,1.8674873,1.8445129,1.2996924,0.8041026,1.3620514,1.3915899,1.5327181,1.7099489,1.9659488,2.4549747,3.1277952,3.1442053,2.92759,2.6847181,2.4155898,2.1497438,1.8740515,1.8707694,2.1464617,2.412308,2.231795,1.8707694,1.6672822,1.6475899,1.5425643,1.463795,1.4211283,1.2209232,0.9517949,0.9747693,1.5163078,1.972513,1.9200002,1.3784616,0.8041026,0.8402052,0.8336411,0.8008206,0.78769237,0.8598975,0.5513847,0.45292312,0.5349744,0.72861546,0.9156924,1.1191796,1.1881026,1.3226668,1.5425643,1.6738462,1.8937438,1.9167181,2.0545642,2.2711797,2.1825643,2.2908719,2.1333334,1.9265642,1.8412309,2.0217438,2.681436,4.7655387,6.514872,7.204103,7.141744,8.021334,8.352821,9.255385,10.315488,9.573745,10.253129,11.099898,12.875488,16.052513,20.818052,21.668104,21.27754,22.17354,24.448002,25.777233,27.733335,35.190155,46.45744,54.465645,46.785645,47.53395,49.78544,48.964928,44.455387,39.601234,58.53539,82.11693,100.033646,108.18298,108.6556,108.48821,104.34955,105.261955,118.68555,150.5313,167.16801,141.60083,107.79242,85.832214,81.89703,82.83242,84.70975,84.24698,80.3676,74.21703,70.02585,62.723286,55.059696,48.147697,41.47857,36.575184,32.39385,29.558157,28.885336,31.363285,33.447388,32.59077,30.683899,27.808823,22.255592,19.941746,20.164925,21.336617,21.881437,20.207592,17.024002,13.594257,10.755282,8.776206,7.3386674,7.4075904,8.605539,9.557334,11.30995,17.332514,37.812515,46.660927,36.755695,17.499899,14.828309,6.931693,4.2601027,4.2535386,5.1856413,6.173539,8.027898,9.990565,13.029744,17.178257,21.536821,30.762669,51.78421,76.56698,91.1557,75.67426,70.629745,73.22257,64.00001,43.940105,34.425438,34.756927,29.003489,22.767591,19.331284,19.633232,20.729437,23.45354,24.201847,23.506054,26.016823,28.639181,32.485744,36.128822,39.141747,42.085747,47.13026,50.425438,49.493336,45.528618,43.382156,44.058258,50.17272,57.10113,57.30462,40.359386,40.28718,41.668926,44.783592,49.266876,54.114464,41.908516,32.57108,27.073643,22.767591,13.364513,7.00718,4.594872,4.266667,4.640821,4.827898,4.9296412,6.4656415,7.719385,7.75877,6.4295387,5.7435904,10.594462,12.885334,12.130463,15.428925,5.796103,11.0145645,11.562668,4.535795,3.6332312,3.1376412,2.8422565,4.1485133,5.4875903,2.356513,1.5885129,1.142154,0.88287187,0.69907695,0.48902568,1.1027694,1.6968206,2.0841026,1.9692309,0.9288206,1.014154,1.2832822,1.3095386,0.99774367,0.574359,0.69907695,1.142154,1.5491283,1.719795,1.6311796,1.3357949,1.5885129,2.294154,3.3509746,4.650667,3.2918978,2.5304618,2.2055387,2.1497438,2.1858463,2.2908719,4.138667,5.0477953,4.706462,5.179077,14.808617,17.690258,16.8599,14.204719,10.443488,9.088,13.289026,14.808617,12.412719,11.851488,10.883283,10.512411,8.730257,5.6976414,3.7349746,3.2262566,4.466872,6.0160003,7.4075904,9.160206,4.9985647,4.6933336,4.1452312,2.665026,2.9669745,4.1124105,13.138052,12.501334,3.8334363,7.965539,6.2818465,5.979898,6.1341543,6.626462,8.15918,9.045334,7.509334,5.0674877,3.446154,4.571898,4.955898,6.4000006,8.231385,10.453334,13.771488,12.58995,11.401847,12.87877,15.658668,14.355694,9.856001,8.434873,8.572719,8.648206,6.948103,16.672821,11.772718,9.570462,13.584412,13.525334,5.9995904,2.1989746,1.1290257,1.9823592,4.128821,1.8674873,1.8510771,1.3784616,0.128,0.16082053,0.19692309,0.11158975,0.068923086,0.118153855,0.15753847,3.1081028,1.6836925,0.19692309,0.13784617,0.18379489,0.20348719,0.20676924,0.23630771,0.35446155,0.6301539,0.56123084,0.27569234,0.10502565,0.17066668,0.38728207,0.14112821,0.06564103,0.07548718,0.1148718,0.17723078,0.42994875,1.3029745,2.1497438,2.6683078,2.9078977,1.9922053,1.4244103,1.0666667,0.7515898,0.30851284,0.3708718,0.39056414,0.4004103,0.49887183,0.8730257,0.7253334,0.6826667,0.7187693,0.8730257,1.2438976,1.214359,1.0633847,1.5655385,2.3827693,2.048,1.7985642,1.339077,1.4998976,2.0742567,1.7952822,1.7427694,2.15959,2.4943593,2.789744,3.6758976,3.6890259,3.0982566,2.5928206,2.300718,1.7920002,1.8215386,1.4933335,1.2438976,1.1848207,1.1126155,1.339077,1.1158975,0.97805136,1.0371283,0.9616411,0.84348726,0.63343596,0.47261542,0.43323082,0.5021539,0.43323082,0.42338464,0.4397949,0.46276927,0.47589746,0.4397949,0.4266667,0.3314872,0.20676924,0.25928208,0.32164106,0.3511795,0.48246157,0.7844103,1.2668719,1.8281027,2.3926156,2.806154,3.1671798,3.8498464,2.5731285,2.7634873,3.7743592,4.71959,4.46359,3.7842054,3.0490258,2.8160002,3.0687182,3.1967182,2.858667,2.4713848,2.1924105,1.9823592,1.6049232,1.142154,0.90912825,0.7811283,0.6662565,0.51856416,0.48574364,0.56451285,0.77456415,1.0010257,0.9911796,0.92225647,0.9682052,1.0502565,1.0765129,0.9616411,0.9616411,1.214359,1.5983591,2.1169233,2.8849232,3.3509746,3.5971284,3.5905645,3.2918978,2.6683078,2.5173335,2.4188719,2.172718,1.9003079,2.038154,2.0545642,2.3433847,2.9144619,3.4034874,3.0654361,2.7503593,1.9396925,1.4736412,1.5425643,1.6672822,1.2964103,1.3620514,1.4276924,1.3817437,1.4572309,1.3029745,1.4309745,1.4211283,1.3062565,1.5688206,1.7887181,2.5435898,2.5731285,1.7755898,1.2176411,1.7132308,1.8576412,1.8871796,2.2022567,3.3509746,3.8629746,3.7448208,3.4330258,3.2098465,3.2000003,2.9144619,2.740513,2.484513,2.2153847,2.2383592,2.3269746,2.1234872,2.044718,2.097231,1.8806155,1.5688206,1.3784616,1.2570257,1.083077,0.6662565,0.508718,0.380718,0.24943592,0.128,0.08205129,0.059076928,0.190359,0.38728207,0.574359,0.702359,0.90584624,0.88287187,0.81066674,0.761436,0.71548724,1.0765129,1.0962052,1.1158975,1.332513,1.7985642,1.972513,2.2613335,2.6683078,2.9735386,2.7273848,2.917744,3.3969233,4.07959,4.844308,5.540103,6.235898,6.7117953,7.4043083,8.211693,8.480822,9.7903595,11.506873,12.432411,12.304411,11.785847,11.900719,11.992617,11.588924,10.81436,10.374565,11.185231,12.481642,13.561437,14.034052,13.83713,14.168616,13.53518,12.278154,10.978462,10.469745,10.036513,9.3078985,8.923898,8.960001,8.917334,9.691898,9.787078,10.033232,10.525539,10.617436,10.939077,10.840616,10.686359,10.9456415,12.1928215,14.39836,14.916924,14.710155,14.50995,14.808617,14.086565,13.354668,12.3076935,11.290257,11.303386,12.041847,11.904001,11.2672825,10.505847,9.941334,10.006975,10.269539,10.548513,10.722463,10.765129,11.188514,11.437949,11.191795,10.643693,10.525539,10.994873,11.408411,12.20595,13.3251295,14.204719,13.2562065,12.005745,10.748719,9.800206,9.468719,9.941334,9.938052,9.980719,10.134975,10.020103,9.616411,9.750975,10.213744,10.909539,11.828514,10.463181,9.540924,9.147078,8.822155,7.574975,7.7718983,7.204103,6.4000006,5.7042055,5.284103,5.6352825,5.474462,5.277539,5.2578464,5.333334,5.989744,5.8256416,5.0904617,4.2830772,4.135385,3.82359,3.639795,3.623385,3.7809234,4.076308,4.20759,4.197744,3.9811285,3.7284105,3.8301542,3.308308,3.4724104,4.017231,4.4701543,4.201026,3.751385,3.6135387,3.639795,3.5741541,3.0687182,1.8412309,1.270154,1.1979488,1.3489232,1.5031796,1.5130258,1.5983591,1.4933335,1.3751796,1.2865642,1.1158975,1.0962052,1.1257436,0.9714873,0.65969235,0.48902568,0.5316923,0.69579494,0.77128214,0.827077,1.1979488,1.7755898,1.4933335,0.9747693,0.7056411,1.0601027,1.4572309,1.5983591,1.585231,1.5983591,1.9003079,2.3663592,2.550154,2.425436,2.1136413,1.8937438,1.723077,1.5392822,1.4900514,1.5064616,1.3193847,1.3226668,1.3883078,1.4473847,1.4572309,1.3718976,1.4375386,1.5688206,1.5261539,1.401436,1.6410258,1.6836925,1.7526156,1.6968206,1.3981539,0.77128214,0.7581539,0.77456415,0.8795898,1.0075898,0.9682052,0.65969235,0.5973334,0.7318975,0.90584624,0.8467693,0.955077,1.2570257,1.5983591,1.8346668,1.8182565,2.100513,2.2416413,2.6354873,3.0916924,2.8488207,2.7634873,2.7437952,2.6453335,2.553436,2.7700515,3.7185643,5.835488,8.139488,9.997129,11.126155,12.048411,13.348104,14.683899,14.808617,11.552821,9.800206,10.965334,12.310975,13.318565,15.704617,15.38954,17.174976,20.128822,23.686565,27.670977,30.818464,40.004925,47.579903,49.91672,47.438774,47.780106,49.83795,50.369644,48.94195,47.9639,71.775185,98.98011,114.98668,116.24699,110.25067,101.26114,93.354675,95.72431,108.77375,124.1436,116.27324,91.723495,69.4679,58.39754,57.32103,58.660107,68.40124,79.5438,86.91857,87.21396,81.35221,72.914055,64.52513,57.08472,49.765747,43.887592,38.738052,36.637543,40.60226,54.31795,58.020107,48.452927,37.16267,29.433437,24.2839,22.291695,26.998156,30.930054,28.967386,18.353231,12.297847,9.045334,7.387898,6.432821,5.618872,6.1768208,8.316719,10.039796,12.596514,20.483284,43.986053,53.251286,41.360413,18.36308,11.280411,7.90318,5.3431797,4.5456414,5.3760004,6.633026,9.314463,10.788103,12.5374365,16.068924,22.895592,38.961235,57.508106,71.99837,79.05149,78.42462,68.38483,62.992416,52.608006,38.514874,32.90585,30.598566,25.951181,21.369438,18.563284,18.520617,18.084105,18.789745,19.859694,21.88472,26.83077,30.024208,34.336823,39.010464,43.05067,45.25621,47.4519,48.482464,44.550568,38.76103,41.110977,42.742157,48.321644,53.91098,54.242466,42.76185,44.576824,44.7639,47.202465,51.872826,54.85621,40.484104,30.096413,24.398771,20.506258,11.963078,6.166975,4.1091285,3.826872,3.95159,3.698872,4.5128207,5.796103,7.7423596,9.396514,8.664616,7.381334,10.496001,11.201642,8.562873,7.532308,5.5926156,9.143796,8.027898,2.7011285,4.2436924,3.501949,2.8553848,2.2449234,1.7427694,1.5786668,1.4375386,1.4998976,1.142154,0.4955898,0.45292312,1.0666667,1.4178462,1.5360001,1.4572309,1.214359,0.955077,1.3620514,1.7001027,1.6213335,1.1651284,1.0568206,1.7132308,2.6223593,3.0982566,2.2777438,1.1158975,1.1093334,1.9790771,3.698872,6.521436,4.637539,3.3805132,2.5665643,2.1070771,2.041436,2.678154,2.9505644,5.0543594,7.9097443,7.171283,13.820719,18.189129,18.005335,14.631386,13.046155,10.28595,11.940104,13.958565,14.39836,13.4400015,11.756309,11.542975,9.586872,5.835488,3.383795,2.3040001,3.1540515,5.5565133,7.8047185,6.8660517,6.7117953,6.7872825,5.175795,3.1376412,5.10359,4.8738465,17.250463,17.092924,5.651693,10.587898,7.6996927,7.748924,7.181129,6.1046157,8.293744,10.597744,9.668923,6.8397956,4.6834874,7.026872,6.518154,7.4699492,8.241231,10.771693,20.59159,12.550565,9.074872,10.404103,14.752822,18.294155,12.422565,10.210463,9.947898,10.085744,9.232411,10.407386,10.006975,9.731283,9.573745,7.8441033,3.9876926,1.5786668,2.793026,5.904411,5.284103,2.7175386,1.1749744,0.39384618,0.17394873,0.38728207,0.30851284,0.15753847,0.12471796,0.20020515,0.17066668,1.5524104,0.9944616,0.3249231,0.23302566,0.27241027,0.24287182,0.18051283,0.14112821,0.14769232,0.17394873,0.37743592,0.24943592,0.10502565,0.09189744,0.19364104,0.15425642,0.08533334,0.052512825,0.068923086,0.08205129,0.17394873,0.6498462,1.214359,1.6738462,1.9495386,1.975795,1.4834872,1.0765129,0.85005134,0.37415388,0.37415388,0.35446155,0.3446154,0.4004103,0.58420515,0.5546667,0.5874872,0.7220513,0.8763078,0.8467693,0.8336411,1.0896411,1.6049232,2.2153847,2.6157951,2.1530259,1.8149745,1.8313848,2.100513,2.2121027,1.6935385,1.9495386,2.281026,2.5271797,3.045744,3.564308,3.5741541,3.2229745,2.865231,3.0523078,2.2121027,2.2121027,2.0217438,1.5425643,1.6049232,1.3620514,1.3029745,1.4605129,1.6836925,1.6410258,1.4112822,0.92225647,0.6071795,0.55794877,0.52512825,0.36102566,0.46933338,0.6235898,0.6859488,0.5907693,0.47589746,0.38400003,0.27897438,0.19692309,0.21333335,0.3117949,0.3446154,0.40697438,0.58092314,0.92225647,1.211077,1.7493335,2.0644104,2.297436,3.2328207,2.9505644,2.5173335,3.0326157,4.1780515,4.20759,3.892513,3.5544617,3.2886157,3.0818465,2.8291285,2.5107694,2.3630772,2.038154,1.5688206,1.3686155,1.0436924,0.8467693,0.72861546,0.65312827,0.5874872,0.5152821,0.56451285,0.7778462,1.0371283,1.0601027,0.9878975,0.98461545,1.0108719,1.0502565,1.083077,1.1585642,1.276718,1.4276924,1.782154,2.6945643,3.2229745,3.4231799,3.242667,2.8160002,2.4713848,2.3335385,2.4352822,2.5698464,2.7273848,3.062154,2.0020514,2.1169233,2.8192823,3.4133337,3.0818465,2.6945643,1.9298463,1.467077,1.3686155,1.1093334,0.8566154,2.0053334,2.2121027,1.1946667,0.72861546,0.83035904,0.84348726,0.88615394,1.1060513,1.6738462,1.2209232,1.719795,2.034872,1.7755898,1.2996924,1.8313848,2.166154,2.484513,2.8914874,3.4231799,3.9548721,3.892513,3.501949,3.0818465,2.9636924,2.7076926,2.3433847,2.162872,2.225231,2.3696413,2.4024618,2.1464617,1.8707694,1.7558975,1.8904617,1.7001027,1.2898463,1.0075898,0.8730257,0.5481026,0.36758977,0.24287182,0.14441027,0.068923086,0.04266667,0.055794876,0.24287182,0.47261542,0.65641034,0.7384616,0.892718,0.90584624,0.8763078,0.8566154,0.8598975,1.2832822,1.3062565,1.2570257,1.3554872,1.7296412,1.9659488,2.1497438,2.3138463,2.4057438,2.3072822,2.865231,3.7316926,4.630975,5.349744,5.723898,6.2162056,6.73477,7.50277,8.346257,8.690872,10.348309,11.759591,12.448821,12.314258,11.621744,11.408411,11.392001,11.185231,10.755282,10.41395,11.250873,12.754052,14.224411,15.107284,14.992412,14.217847,12.383181,10.679795,9.685334,9.370257,8.789334,7.6931286,7.509334,8.402052,9.278359,10.092308,10.085744,10.131693,10.361437,10.157949,10.840616,10.748719,10.384411,10.28595,11.030975,13.906053,14.8939495,14.864411,14.54277,14.506668,13.974976,13.223386,12.3536415,11.766154,12.133744,12.619488,12.189539,11.175385,9.987283,9.114257,9.301334,9.800206,10.213744,10.407386,10.489437,10.886565,11.001437,10.617436,9.993847,9.842873,10.328616,10.896411,11.451077,11.96636,12.475078,11.913847,11.204924,10.410667,9.701744,9.363693,10.131693,10.505847,10.59118,10.400822,9.852718,9.734565,10.223591,10.8307705,11.323078,11.733335,10.174359,9.6065645,9.281642,8.661334,7.397744,7.5520005,7.020308,6.3868723,5.920821,5.5630774,5.865026,5.3005133,4.7917953,4.7228723,4.926359,5.622154,5.540103,4.821334,3.8334363,3.18359,3.1573336,3.2787695,3.4789746,3.7382567,4.092718,4.4832826,4.4701543,4.164923,3.7874875,3.6496413,3.3509746,3.2754874,3.5840003,3.9811285,3.7054362,3.4888208,3.620103,3.6430771,3.3444104,2.740513,1.9987694,1.4867693,1.1651284,1.1585642,1.3915899,1.5885129,1.8182565,1.8576412,1.6377437,1.2635899,1.0075898,0.8008206,0.7122052,0.62030774,0.49887183,0.4266667,0.5481026,0.75487185,0.7975385,0.7844103,1.1749744,1.3226668,1.1388719,0.85005134,0.79097444,1.3883078,2.0611284,2.1825643,2.0906668,1.9987694,1.9987694,2.2678976,2.4155898,2.6486156,2.7864618,2.2744617,1.8576412,1.6738462,1.5885129,1.463795,1.1585642,1.086359,1.0502565,0.94523084,0.8336411,0.9321026,1.2603078,1.270154,1.3128207,1.3850257,1.1290257,1.0929232,0.9353847,0.92553854,1.1027694,1.2964103,1.1749744,1.2898463,1.3259488,1.1126155,0.6268718,0.40697438,0.49887183,0.6859488,0.77128214,0.56451285,0.67282057,1.0765129,1.394872,1.5392822,1.7099489,2.294154,2.789744,2.9407182,2.7766156,2.5928206,2.5928206,2.6387694,2.6715899,2.733949,2.989949,5.431795,8.631796,10.971898,11.956513,12.2387705,12.347078,13.328411,15.304206,16.459488,13.029744,11.687386,11.316514,11.713642,12.872206,14.982565,13.262771,15.937642,20.073027,23.752207,26.04636,32.114876,42.646976,48.141132,49.08636,55.985233,52.847595,52.237133,53.202057,55.312416,58.669952,70.64616,86.21949,93.88637,92.353645,90.54852,88.52021,88.04103,91.15898,94.10954,87.312416,67.14749,53.06093,46.034054,45.236515,48.019695,50.021748,61.124928,75.3198,87.16473,91.76616,86.87262,78.72657,69.30052,59.470776,48.994465,44.320824,41.731285,50.143185,75.62503,121.40965,128.1477,92.993645,55.33539,33.828106,26.38113,29.604105,44.324104,56.195286,52.847595,23.893335,11.040821,6.4722056,5.4547696,5.2512827,5.142975,5.349744,7.781744,10.095591,12.268309,16.600616,22.92513,25.862566,21.48431,12.964104,10.55836,8.129642,5.5729237,4.4373336,5.044513,6.485334,11.0145645,12.0549755,13.239796,17.010874,24.628515,46.674053,49.74277,46.677338,46.467285,54.23262,56.231388,50.04144,40.385643,32.039387,29.830566,33.82154,26.801233,19.574156,16.374155,14.8480015,16.275694,18.399181,20.082872,21.812515,25.69518,29.551592,33.119183,38.89231,44.964108,45.013336,43.779285,42.036514,38.196514,34.23836,35.69231,40.52349,47.46503,52.56534,52.709747,45.59426,48.718773,47.12698,48.213337,52.158363,51.92534,38.170258,27.825233,22.065233,18.54359,11.414975,5.287385,3.4888208,3.249231,3.0884104,2.806154,4.1878977,5.684513,8.723693,11.897437,10.971898,7.9819493,7.9294367,6.7085133,4.6276927,6.409847,7.9458466,13.932309,11.792411,3.69559,6.5772314,2.5600002,1.5031796,2.4648206,3.446154,1.3587693,2.0184617,2.2744617,1.6082052,0.512,0.48902568,0.7811283,1.394872,1.7001027,1.6771283,1.9232821,1.3128207,1.6443079,2.1398976,2.228513,1.5556924,1.6049232,1.5524104,1.8937438,2.3860514,2.044718,0.88615394,0.8041026,0.93866676,1.1126155,1.847795,4.630975,4.4110775,3.6726158,3.1277952,1.723077,3.5446157,3.501949,6.0061545,9.465437,6.3179493,18.766771,22.87918,19.669334,14.230975,15.730873,15.402668,12.471796,11.080206,11.841642,11.841642,10.706052,10.604308,9.298052,6.8397956,5.5696416,2.993231,2.7175386,3.1573336,3.570872,4.059898,6.157129,6.892308,6.436103,5.579488,5.737026,4.9788723,23.138464,23.174566,6.180103,11.369026,11.428103,15.96718,15.323898,9.55077,8.392206,12.836103,12.1698475,9.563898,7.1220517,5.8912826,8.818872,13.269335,14.237539,12.09436,12.557129,9.176616,9.639385,9.504821,9.567181,15.855591,16.183796,15.396104,14.473847,13.883078,13.564719,12.649027,12.511181,12.199386,10.394258,5.402257,2.1924105,0.6826667,6.8299494,15.392821,9.947898,3.4527183,1.401436,0.8402052,0.5349744,0.9616411,0.42338464,0.21661541,0.27241027,0.4135385,0.36758977,0.63343596,0.53825647,0.41025645,0.39384618,0.44307697,0.39384618,0.18051283,0.03938462,0.03938462,0.07548718,0.17394873,0.21661541,0.17394873,0.0951795,0.108307704,0.25271797,0.18051283,0.118153855,0.16738462,0.28882053,0.36430773,0.6662565,0.9878975,1.3161026,1.8149745,2.097231,1.6738462,1.2996924,1.1323078,0.7187693,0.47261542,0.33805132,0.32164106,0.37415388,0.4135385,0.37415388,0.44964105,0.6071795,0.7975385,0.9321026,1.017436,1.8609232,2.2580514,2.3236926,3.495385,2.3466668,2.2416413,2.2678976,2.2613335,2.8225644,1.7001027,1.8412309,2.425436,2.7766156,2.349949,2.1070771,2.1103592,2.7011285,3.6627696,4.210872,3.2361028,3.0818465,2.7634873,2.2153847,2.28759,1.6049232,1.8838975,1.9364104,1.7624617,2.5337439,2.8389745,2.0808206,1.3423591,0.97805136,0.6104616,0.4266667,0.6104616,0.9288206,1.0929232,0.761436,0.48246157,0.33805132,0.33805132,0.3708718,0.21333335,0.3117949,0.446359,0.54482055,0.6301539,0.82379496,0.8960001,1.5392822,1.9528207,2.0611284,2.487795,2.4024618,2.4615386,3.3050258,4.378257,3.95159,4.71959,4.493129,3.5938463,2.6322052,2.487795,2.169436,2.412308,2.3204105,1.6968206,1.0371283,0.892718,0.7450257,0.64000005,0.6104616,0.67282057,0.65969235,0.6662565,0.7581539,0.9353847,1.1454359,0.98461545,0.8992821,0.9682052,1.204513,1.5721027,1.657436,1.6246156,1.6672822,1.9626669,2.6715899,2.487795,2.5238976,2.5665643,2.5074873,2.349949,2.8882053,2.8488207,2.7995899,2.9505644,3.1573336,2.2547693,2.4976413,2.8127182,2.7273848,2.349949,2.5074873,1.7788719,1.4309745,1.6114873,1.3423591,1.148718,6.2785645,6.921847,2.2678976,0.5349744,0.6071795,0.7089231,0.8008206,0.90584624,1.1126155,0.892718,1.2340513,1.3193847,1.1520001,1.5556924,2.5435898,2.793026,3.0194874,3.4724104,3.9351797,4.4012313,3.748103,2.9407182,2.5009232,2.487795,2.0841026,1.8084104,1.7624617,1.9396925,2.2580514,2.284308,2.2416413,1.9922053,1.657436,1.6311796,1.522872,1.2471796,0.9911796,0.7811283,0.48902568,0.256,0.14441027,0.0951795,0.06564103,0.029538464,0.04266667,0.20020515,0.37743592,0.5316923,0.702359,0.8369231,0.85005134,0.85005134,0.8598975,0.82379496,1.276718,1.3062565,1.2274873,1.3029745,1.7558975,2.048,2.166154,2.1070771,2.0873847,2.5632823,3.1113849,3.8071797,4.522667,5.139693,5.5532312,6.1046157,6.5805135,7.0990777,7.77518,8.726975,10.55836,11.648001,11.881026,11.424822,10.742155,10.804514,10.817642,10.811078,11.047385,12.025436,12.06154,13.817437,14.460719,13.748514,14.053744,13.883078,11.98277,9.856001,8.418462,7.965539,7.7948723,7.394462,7.748924,8.753231,9.216001,9.5835905,10.187488,10.59118,10.597744,10.269539,11.329642,11.861334,11.434668,10.545232,10.604308,12.86236,13.90277,14.099693,13.909334,13.88636,13.568001,13.351386,12.918155,12.340514,12.084514,11.585642,11.414975,11.247591,10.738873,9.504821,8.920616,9.42277,10.203898,10.781539,11.001437,11.234463,10.742155,10.174359,9.892103,9.964309,10.20718,10.627283,10.807796,10.755282,10.86359,10.594462,10.584617,10.295795,9.7903595,9.705027,10.522257,11.093334,10.909539,10.167795,9.764103,10.499283,10.817642,10.555078,10.197334,10.880001,9.622975,9.334154,9.403078,9.130668,7.752206,7.788308,7.1089234,6.2916927,5.7107697,5.540103,5.5269747,4.818052,4.33559,4.3027697,4.240411,4.594872,4.6112823,4.1156926,3.2918978,2.6715899,2.7306669,3.249231,3.7382567,4.020513,4.2272825,4.3716927,4.5456414,4.450462,4.1025643,3.8465643,3.4789746,2.7109745,2.546872,3.045744,3.3280003,3.314872,3.2196925,2.9768207,2.5698464,2.044718,1.8642052,1.6147693,1.3029745,1.1454359,1.2209232,1.463795,1.6869745,1.7165129,1.6344616,1.4769232,1.2504616,0.96492314,0.6892308,0.48902568,0.38728207,0.34133336,0.48246157,0.4955898,0.42994875,0.3708718,0.42994875,0.7811283,0.9124103,0.83035904,0.76800007,1.1815386,1.7066668,2.2088206,2.2744617,2.0151796,2.0709746,2.2416413,2.300718,2.3926156,2.3893335,1.9068719,1.5885129,1.4276924,1.339077,1.214359,0.9288206,1.0305642,1.2209232,1.014154,0.5546667,0.61374366,0.62030774,0.6235898,0.7778462,0.9911796,0.92225647,0.72861546,0.65969235,0.65641034,0.6629744,0.61374366,0.67610264,0.72861546,0.7450257,0.69579494,0.5415385,0.3511795,0.39712822,0.4397949,0.37743592,0.25928208,0.54482055,0.9419488,1.2865642,1.5425643,1.782154,2.3860514,2.7831798,2.7963078,2.6256413,2.861949,3.5249233,3.3345644,3.3509746,4.017231,5.1626673,9.344001,12.268309,13.492514,13.233232,12.373334,12.668719,13.604104,14.473847,14.913642,14.91036,15.209026,12.901745,12.018872,13.715693,16.278976,16.469334,17.536001,21.927387,27.992617,29.96513,31.872002,40.60554,45.78462,46.03734,48.978054,56.73026,60.350365,63.35344,64.72862,58.925953,63.136826,71.11549,78.0997,83.84985,92.65888,104.126366,108.888626,105.34073,93.167595,73.32431,61.748516,56.467697,53.73375,52.77867,55.794876,66.730675,81.29642,96.01314,107.47406,112.37088,108.186264,94.825035,78.85785,64.758156,54.879185,52.529236,50.85867,59.070362,89.5639,157.94545,182.4755,130.58955,68.89355,33.12903,28.163284,39.94913,60.373337,71.266464,60.596516,22.455797,10.410667,5.937231,4.8640003,4.8114877,5.1922054,5.5269747,7.000616,8.87795,10.748719,12.511181,13.88636,13.430155,11.362462,8.822155,7.860513,7.5913854,6.2162056,5.3366156,5.5565133,6.5083084,9.242257,11.188514,13.298873,16.242872,20.391386,31.22872,33.73949,35.524925,40.786053,50.336823,46.099697,36.84431,28.33067,24.34954,26.719181,30.34913,27.352617,21.80595,16.666258,13.771488,14.693745,16.039387,17.572104,19.590565,22.92513,27.858053,30.641233,34.15631,38.21621,39.59467,39.240208,36.850876,33.874054,31.442053,30.355694,31.215591,36.992004,45.380928,51.70872,48.93867,49.48349,45.991386,45.75508,48.830364,48.032825,36.023796,26.299078,20.680206,17.362053,10.939077,5.4153852,3.1474874,2.3893335,2.2153847,2.4910772,4.5029745,5.077334,6.5837955,8.687591,8.346257,5.6287184,4.9493337,4.089436,3.1081028,4.332308,12.081232,21.891283,18.504206,5.5630774,5.612308,2.484513,1.6771283,2.231795,2.7798977,1.5425643,2.0250258,1.5622566,1.0535386,0.82379496,0.63343596,0.5677949,1.0075898,1.3029745,1.467077,2.1792822,1.2274873,1.2898463,1.6475899,1.7624617,1.2865642,1.5031796,1.273436,1.086359,1.1585642,1.4211283,0.7811283,0.9616411,1.2077949,1.142154,0.761436,1.2373334,2.3762052,3.3214362,3.495385,2.5895386,3.1015387,4.71959,12.665437,20.79836,11.61518,14.907078,17.56882,15.350155,10.981745,14.181745,14.486976,13.722258,12.570257,12.425847,15.392821,14.276924,11.529847,9.353847,8.100103,6.2523084,5.228308,4.138667,3.9056413,4.522667,5.0609236,4.7294364,5.756718,6.0980515,5.723898,6.616616,6.9349747,15.881847,15.593027,7.7390776,13.551591,6.747898,14.096412,17.371899,12.3306675,8.710565,6.189949,7.8506675,10.233437,10.312206,5.474462,10.105436,17.109335,18.566566,13.673027,8.736821,20.598156,19.505232,14.8020525,14.408206,24.825438,17.158566,14.296617,11.536411,9.232411,12.819694,17.316103,16.712206,15.136822,13.354668,8.78277,2.681436,0.51856416,1.404718,3.1540515,2.2711797,1.3423591,0.96492314,0.60389745,0.24943592,0.42338464,0.3446154,0.3249231,0.33805132,0.44964105,0.83035904,1.2537436,1.5327181,1.2209232,0.5513847,0.44307697,0.42338464,0.3708718,0.2297436,0.101743594,0.23630771,0.29210258,0.25271797,0.20020515,0.16410258,0.118153855,0.17723078,0.17066668,0.16738462,0.256,0.5349744,0.77456415,1.1158975,1.214359,1.1454359,1.4145643,1.7624617,1.8740515,1.7329233,1.4244103,1.1552821,0.8041026,0.5415385,0.43651286,0.4397949,0.4004103,0.48902568,0.5218462,0.6235898,0.75487185,0.7220513,0.7778462,1.7066668,2.8192823,3.4855387,3.114667,2.2416413,2.2121027,2.2219489,2.0808206,2.2121027,1.657436,1.6804104,2.0676925,2.5107694,2.6322052,2.7273848,2.2678976,2.0644104,2.349949,2.7700515,3.1409233,3.2525132,3.0096412,2.6190772,2.5928206,2.5173335,2.3302567,2.2055387,2.1431797,1.9954873,3.3542566,3.2065644,2.5009232,1.9200002,1.8674873,1.0108719,1.2668719,1.3292309,0.9714873,1.0436924,0.69579494,0.57764107,0.62030774,0.6465641,0.3708718,0.39056414,0.50543594,0.5546667,0.571077,0.77456415,0.67282057,1.1585642,1.910154,2.4418464,2.1103592,2.4057438,3.0424619,3.7776413,4.4045134,4.768821,5.802667,5.149539,4.013949,3.131077,2.7798977,2.5304618,2.3433847,2.1825643,1.9298463,1.3784616,1.0469744,0.8041026,0.7089231,0.7253334,0.7089231,0.7253334,0.69579494,0.7975385,0.9878975,1.0108719,0.90912825,0.96492314,1.3226668,1.8806155,2.2547693,2.1464617,2.041436,2.038154,2.231795,2.7076926,2.5928206,2.5074873,2.5600002,2.6157951,2.300718,2.5173335,2.5271797,2.6289232,2.8750772,3.0720003,2.930872,2.8947694,2.5731285,2.048,1.8871796,1.7723079,1.2438976,1.2176411,1.5885129,1.2340513,1.3784616,11.769437,14.083283,5.920821,0.7778462,0.5677949,0.53825647,0.5349744,0.54482055,0.7220513,1.0108719,1.2800001,1.214359,0.93866676,1.020718,1.8313848,2.7306669,3.3903592,3.4691284,2.5928206,3.4494362,3.2525132,2.9013336,2.6486156,2.1103592,1.8806155,1.9298463,2.0020514,2.0250258,2.0873847,1.8576412,1.9889232,1.9232821,1.5753847,1.3259488,1.2373334,1.0568206,0.9321026,0.8336411,0.56123084,0.2231795,0.08861539,0.049230773,0.036102567,0.01969231,0.068923086,0.28882053,0.45620516,0.50543594,0.5316923,0.71548724,0.7122052,0.8041026,1.0043077,1.0568206,0.9714873,1.0502565,1.2570257,1.5327181,1.7788719,1.9364104,1.8970258,1.9068719,2.172718,2.8455386,3.4133337,4.348718,5.221744,5.8289237,6.163693,6.245744,6.744616,7.4043083,8.077128,8.717129,10.420513,11.113027,10.843898,10.072617,9.642668,9.705027,9.984001,10.374565,10.965334,12.06154,12.07795,12.576821,12.872206,12.918155,13.321847,12.389745,10.633847,8.792616,7.3485136,6.5247183,6.2752824,6.413129,7.39118,8.805744,9.386667,9.383386,9.915077,10.528821,10.7848215,10.269539,11.047385,11.477334,11.116308,10.358154,10.459898,11.670976,12.970668,13.541744,13.341539,13.092104,12.442257,12.3766165,12.150155,11.713642,11.730052,11.122872,10.8537445,10.584617,9.954462,8.553026,8.493949,9.481847,10.528821,11.168821,11.464206,11.158976,10.518975,10.210463,10.33518,10.427077,10.994873,11.172104,11.113027,10.988309,10.962052,10.545232,10.292514,9.7673855,9.265231,9.813334,10.44677,10.568206,10.144821,9.6984625,10.289231,10.778257,10.466462,10.092308,10.026668,10.282667,9.580308,9.777231,10.079181,9.688616,7.8112826,7.450257,6.948103,6.482052,6.0652313,5.5630774,5.435077,4.923077,4.44718,4.164923,3.9975388,3.9122055,3.6857438,3.308308,2.809436,2.2547693,2.4713848,3.18359,3.6496413,3.7185643,3.8498464,3.9745643,4.092718,4.128821,4.017231,3.7218463,3.5216413,3.117949,2.8127182,2.8160002,3.2525132,3.0260515,2.6420515,2.3401027,2.2416413,2.349949,1.3259488,1.2537436,1.0699488,0.9288206,0.93866676,1.1585642,1.3062565,1.3259488,1.2603078,1.1323078,0.955077,0.7318975,0.49887183,0.3511795,0.32164106,0.40369233,0.49230772,0.39056414,0.26584616,0.21661541,0.27241027,0.7122052,0.827077,0.7089231,0.5907693,0.8533334,1.1520001,1.5097437,1.6738462,1.6410258,1.6705642,1.7657437,1.8871796,1.8904617,1.7263591,1.4506668,1.2898463,1.1618463,1.0896411,1.0371283,0.88943595,1.1158975,1.3226668,1.1684103,0.80738467,0.8992821,0.76800007,0.63343596,0.69251287,0.8763078,0.8598975,0.98133343,0.9485129,0.86646163,0.80738467,0.8008206,0.7844103,0.61374366,0.4266667,0.30851284,0.30851284,0.21333335,0.25928208,0.37415388,0.44307697,0.33805132,0.56451285,0.8960001,1.2012309,1.4605129,1.7558975,2.1530259,2.5009232,2.7634873,3.121231,3.9548721,4.821334,5.024821,5.7698464,7.02359,7.5191803,12.038565,14.50995,15.730873,16.082052,15.527386,14.792206,14.378668,14.073437,13.912617,14.171899,15.589745,13.128206,12.3306675,14.578873,17.076513,16.328207,18.468103,22.216208,26.059488,28.291285,31.668516,37.536823,39.67016,40.02462,48.735184,56.28062,61.364517,65.47693,67.4757,63.596313,63.330467,68.74257,79.53067,96.22975,120.23796,140.07468,138.86032,119.450264,91.65785,72.241234,64.85334,60.032005,55.2238,51.75139,54.784004,69.19878,83.41006,93.531906,98.38606,99.51508,96.54483,92.13703,87.55201,81.69682,71.125336,61.65334,54.656006,54.101337,68.71303,111.9836,138.70605,102.495186,55.000618,26.28267,24.756516,36.516106,50.868515,56.385647,46.483696,19.429745,10.006975,6.678975,5.8912826,5.5663595,5.1200004,5.5893335,6.445949,7.8047185,9.133949,9.245539,8.254359,7.381334,7.0104623,7.276308,8.083693,7.4075904,6.445949,5.7501545,5.8880005,7.450257,9.6065645,11.588924,13.696001,16.02954,18.500925,23.860516,28.5079,35.96472,44.17313,45.508926,34.166157,26.056208,20.791796,19.049026,22.57067,27.408413,25.984001,21.3399,16.502155,14.473847,13.328411,13.019898,14.424617,17.424412,20.923079,23.003899,25.977438,29.535181,33.05354,35.620106,34.271183,32.36431,29.039593,25.767387,26.368002,27.06708,31.455181,40.917336,50.85867,50.73395,45.453133,41.636105,41.70831,44.07139,43.093338,32.74503,24.198566,19.495386,17.158566,12.182976,6.0356927,3.2032824,2.1234872,1.8576412,2.0808206,3.879385,4.056616,5.2545643,7.0531287,5.986462,4.2535386,4.516103,4.125539,4.164923,9.416205,25.531078,33.457233,24.234669,6.294975,5.4547696,4.1583595,2.4648206,1.8346668,2.1431797,1.6968206,2.2088206,1.9003079,1.3259488,0.90584624,0.8992821,0.5218462,0.7187693,0.90584624,1.014154,1.4998976,1.079795,1.1027694,1.276718,1.3883078,1.3128207,1.2242053,1.5491283,1.4375386,1.0666667,1.6508719,1.2570257,1.1257436,1.0469744,0.9288206,0.79097444,0.4004103,0.92553854,1.785436,2.4320002,2.3401027,2.868513,8.139488,18.615797,26.857027,17.526155,16.777847,17.27672,15.40595,12.081232,12.777026,12.882052,12.383181,11.474052,11.539693,15.156514,13.180719,11.001437,9.67877,8.818872,6.550975,6.245744,4.7556925,3.564308,3.636513,5.402257,7.8145647,6.7085133,5.0084105,4.460308,5.5991797,10.505847,15.268104,12.097642,5.6976414,13.2562065,4.8672824,6.7774363,10.873437,11.979488,7.8473854,3.8498464,7.2205133,11.286975,11.451077,5.1889234,9.275078,19.094976,21.858463,17.716515,19.764515,23.16472,20.59159,16.528412,14.36554,16.367592,11.575796,10.059488,8.349539,7.1056414,11.113027,14.720001,13.164309,11.556104,10.476309,5.9569235,2.7076926,1.2340513,0.5349744,0.190359,0.3511795,1.5556924,1.4309745,0.7778462,0.318359,0.6826667,0.8533334,1.5327181,1.7460514,1.2898463,0.7450257,1.148718,2.5337439,2.6354873,1.270154,0.3314872,0.35774362,0.4266667,0.34133336,0.20676924,0.4397949,0.37743592,0.256,0.2297436,0.30851284,0.3511795,0.30851284,0.2231795,0.16082053,0.18707694,0.40369233,0.84348726,1.4802053,1.6311796,1.3653334,1.522872,1.4408206,1.522872,1.5655385,1.5524104,1.6410258,1.1520001,0.78769237,0.5907693,0.5284103,0.45292312,0.5513847,0.574359,0.6235898,0.69251287,0.67282057,0.90912825,1.6640002,2.8127182,3.7218463,3.2131286,2.1792822,2.097231,1.975795,1.7066668,2.0676925,1.8379488,1.6869745,1.8281027,2.0742567,1.8313848,2.7241027,2.5435898,2.4648206,2.7634873,2.8324106,3.3280003,3.1934361,2.8127182,2.4943593,2.4681027,2.740513,2.2350771,2.0086155,2.3138463,2.5928206,3.8662567,3.5183592,3.006359,3.0227695,3.508513,2.353231,1.7263591,1.6475899,2.097231,2.9997952,1.020718,0.69579494,1.0732309,1.2996924,0.61374366,0.571077,0.52512825,0.46276927,0.4397949,0.5874872,0.5677949,0.7384616,1.276718,1.9200002,1.9954873,2.1956925,3.239385,4.069744,4.352,4.4898467,4.650667,4.7491283,4.417641,3.7218463,3.1638978,3.0194874,2.487795,2.0086155,1.7066668,1.4112822,1.0765129,0.8336411,0.7253334,0.69251287,0.5973334,0.61374366,0.6892308,0.77456415,0.8533334,0.93866676,0.9124103,1.3357949,1.9626669,2.5042052,2.6190772,2.3072822,2.1234872,2.0644104,2.162872,2.5042052,2.6354873,2.5632823,2.5632823,2.6420515,2.537026,2.4352822,2.3958976,2.5206156,2.740513,2.806154,3.190154,3.1606157,2.665026,1.9889232,1.7690258,1.5589745,1.273436,1.3817437,1.6344616,1.0601027,1.5983591,10.390975,14.998976,10.781539,0.88615394,0.7581539,0.6629744,0.60061544,0.60061544,0.7253334,0.9517949,1.1520001,1.3095386,1.3883078,1.3522053,1.4769232,2.03159,2.6847181,3.0260515,2.5796926,3.0096412,2.5796926,2.2646155,2.2547693,1.9495386,1.8543591,2.0545642,2.103795,1.9232821,1.7985642,1.5031796,1.8051283,1.9429746,1.6508719,1.1323078,1.1946667,1.0338463,0.8402052,0.6695385,0.45292312,0.20348719,0.072205134,0.026256412,0.02297436,0.032820515,0.12471796,0.2986667,0.50543594,0.6235898,0.48902568,0.7417436,0.7844103,0.8730257,1.0765129,1.2603078,1.0929232,1.0765129,1.2176411,1.4933335,1.8576412,1.9068719,1.8313848,1.9823592,2.4320002,2.9702566,3.7185643,4.775385,5.5762057,5.9569235,6.1341543,6.2720003,6.665847,7.312411,8.073847,8.684308,9.990565,10.243283,9.691898,8.881231,8.644924,9.130668,10.262975,10.985026,11.306667,12.297847,11.864616,11.956513,12.2617445,12.570257,12.763899,12.3995905,10.889847,9.16677,7.6898465,6.4295387,5.8092313,6.0980515,7.174565,8.631796,9.777231,9.219283,9.31118,10.089026,11.080206,11.303386,11.490462,11.414975,11.113027,10.807796,10.925949,11.152411,12.06154,12.662155,12.619488,12.235488,11.654565,11.572514,11.631591,11.661129,11.67754,10.561642,10.089026,9.852718,9.42277,8.372514,8.533334,9.386667,10.20718,10.555078,10.272821,9.760821,9.655796,9.796924,10.052924,10.331899,11.142565,11.533129,11.585642,11.447796,11.34277,10.745437,10.20718,9.6754875,9.475283,10.299078,10.607591,10.55836,10.072617,9.485129,9.55077,9.993847,10.000411,9.905231,9.980719,10.443488,9.580308,9.4457445,9.501539,9.245539,8.201847,7.6668725,7.000616,6.2523084,5.504,4.8836927,4.7392826,4.450462,4.128821,3.8071797,3.4527183,3.1671798,2.9965131,2.861949,2.678154,2.3630772,2.537026,3.1113849,3.515077,3.626667,3.7809234,4.086154,4.2240005,4.279795,4.2371287,3.9680004,3.7120004,3.511795,3.3345644,3.2131286,3.2361028,2.7864618,2.4418464,2.041436,1.6771283,1.7132308,0.955077,0.98461545,0.92553854,0.88615394,0.9517949,1.1651284,1.083077,1.0338463,0.9485129,0.8369231,0.8041026,0.73517954,0.50543594,0.33476925,0.3117949,0.3708718,0.4660513,0.39056414,0.3249231,0.33476925,0.37415388,0.69251287,0.8008206,0.6826667,0.52512825,0.69579494,0.7844103,0.9419488,1.1158975,1.2504616,1.3095386,1.3653334,1.5261539,1.5786668,1.4572309,1.2406155,1.1093334,0.98133343,0.92225647,0.9353847,0.9747693,1.204513,1.4342566,1.3522053,1.0601027,1.0666667,0.9288206,0.79097444,0.81066674,0.9353847,0.90256417,1.148718,1.3587693,1.339077,1.1158975,0.9353847,1.0075898,0.6826667,0.318359,0.128,0.18707694,0.2855385,0.3249231,0.38400003,0.4660513,0.47917953,0.61374366,0.83035904,1.0962052,1.4244103,1.8904617,2.3072822,3.0194874,4.0041027,5.044513,5.723898,6.8365135,7.6767187,8.736821,9.80677,9.96759,13.768207,16.90913,19.541334,20.565334,17.634462,16.167385,15.409232,14.956308,14.660924,14.65436,15.43877,13.764924,12.911591,13.718975,14.598565,13.791181,15.986873,19.213129,22.498463,25.88554,30.920208,35.413338,36.854156,39.27631,53.251286,56.44144,60.950977,64.39713,65.404724,63.63898,59.96308,62.641235,74.555084,96.108315,125.25622,149.15283,143.31406,114.75037,80.426674,67.24924,64.06564,60.452106,55.54544,51.826878,55.122055,69.691086,79.30093,82.50093,80.4037,76.668724,74.089035,77.26606,84.96247,91.703804,87.801445,70.04226,56.274055,47.323902,46.74626,60.8197,76.176414,58.962055,34.816,19.958155,21.185642,30.313028,37.044518,38.275284,32.502155,19.833437,12.612924,8.753231,7.138462,6.5017443,5.4153852,5.4383593,5.9963083,6.774154,7.1614366,6.242462,5.0609236,5.431795,6.698667,8.077128,8.651488,6.872616,6.4656415,6.419693,6.747898,8.480822,10.59118,12.396309,14.260514,16.226463,17.99877,21.999592,30.756105,40.84841,45.771492,35.94503,22.764309,18.970259,17.765745,17.125746,19.767796,25.294771,25.701746,21.907694,16.640001,14.444309,11.98277,11.145847,12.100924,14.483693,17.401438,18.30072,22.088207,25.619694,28.087797,31.01867,29.029745,28.1239,25.419489,22.170258,23.791592,24.766361,27.864618,37.415386,48.804108,48.48903,41.649235,37.779694,37.933952,40.021336,38.820107,30.385233,22.898874,19.236105,17.920002,13.115078,6.2523084,3.2787695,2.3204105,2.1202054,2.0644104,3.6036925,3.9712822,5.024821,6.1538467,4.2962055,3.436308,4.069744,3.9581542,4.5390773,10.919386,35.186874,39.01703,26.25313,8.461129,4.923077,5.225026,4.8114877,4.768821,4.460308,1.5064616,2.3630772,2.100513,1.5031796,1.1027694,1.204513,0.56451285,0.6104616,0.6826667,0.67938465,1.0436924,1.1093334,1.1454359,1.273436,1.4736412,1.5885129,1.6705642,2.5961027,2.5764105,1.7526156,2.1891284,1.6410258,1.211077,0.95835906,0.9156924,1.0666667,0.636718,0.4397949,0.6629744,1.1848207,1.585231,2.0808206,8.103385,17.05354,23.502771,19.203283,17.841232,15.691488,13.915898,13.072412,13.088821,14.083283,12.711386,11.621744,12.032001,13.732103,13.013334,13.430155,13.397334,12.2157955,10.079181,8.651488,6.5247183,5.149539,5.0609236,5.8518977,9.957745,6.892308,4.7556925,5.2348723,3.5905645,8.753231,12.117334,9.216001,4.781949,12.744206,6.99077,5.3366156,6.7183595,8.329846,5.6418467,4.824616,8.438154,11.221334,11.07036,9.045334,10.666668,15.744001,20.102566,22.081642,22.550976,23.985233,21.526976,17.257027,13.348104,12.058257,10.269539,8.205129,7.13518,7.6242056,9.5146675,10.246565,8.004924,6.173539,5.2709746,2.9735386,2.550154,1.4572309,0.5677949,0.4397949,1.3161026,5.4449234,6.498462,4.4340515,1.5327181,2.3991797,2.6453335,3.6168208,4.056616,3.3444104,1.4966155,1.0994873,2.3729234,2.7273848,1.6049232,0.47261542,0.318359,0.39056414,0.36758977,0.26256412,0.446359,0.34133336,0.21333335,0.23630771,0.39712822,0.47261542,0.4594872,0.37743592,0.27897438,0.23302566,0.3052308,0.67282057,1.2504616,1.4900514,1.4276924,1.6869745,1.3718976,1.3128207,1.4080001,1.5622566,1.6968206,1.339077,1.079795,0.84348726,0.6301539,0.4955898,0.56451285,0.6170257,0.6662565,0.7187693,0.7581539,0.9616411,1.401436,2.3302567,3.3050258,3.190154,2.4188719,2.1366155,1.7624617,1.4539489,2.0939488,2.1398976,1.9003079,1.913436,2.0020514,1.2504616,2.0086155,2.297436,2.4713848,2.6026669,2.4713848,3.0162053,3.045744,2.6617439,2.2711797,2.5665643,2.789744,2.2416413,1.910154,2.166154,2.7831798,3.5282054,3.1277952,2.809436,3.1015387,3.8498464,2.993231,1.9528207,1.8740515,2.8225644,3.7940516,1.3456411,0.7384616,1.0666667,1.4605129,1.083077,1.723077,1.3522053,0.8041026,0.51856416,0.5415385,0.5218462,0.446359,0.6301539,1.0929232,1.5688206,1.8018463,2.7569232,3.446154,3.639795,3.8531284,3.6791797,3.9680004,3.9581542,3.5052311,3.0851285,2.986667,2.4976413,2.0906668,1.8313848,1.3915899,1.0732309,0.8992821,0.8041026,0.7220513,0.5973334,0.55794877,0.6170257,0.6826667,0.7581539,0.92225647,0.94523084,1.4506668,2.1234872,2.665026,2.789744,2.4516926,2.1333334,2.034872,2.176,2.3762052,2.7569232,2.6453335,2.5173335,2.537026,2.5862565,2.412308,2.356513,2.4352822,2.556718,2.546872,2.934154,2.8324106,2.3368206,1.7591796,1.6246156,1.401436,1.211077,1.3062565,1.4900514,1.1093334,2.097231,8.369231,12.914873,11.10318,0.65312827,0.94523084,0.9517949,0.827077,0.7318975,0.8533334,0.9321026,0.955077,1.1618463,1.5360001,1.8215386,1.5163078,1.7591796,2.0873847,2.2547693,2.2383592,2.733949,2.176,1.8609232,2.0611284,2.048,1.8642052,1.9035898,1.8970258,1.7526156,1.529436,1.2668719,1.6278975,1.8970258,1.7001027,1.020718,1.1913847,1.1191796,0.88943595,0.5874872,0.3117949,0.16410258,0.055794876,0.009846155,0.01969231,0.059076928,0.21661541,0.31507695,0.46276927,0.5973334,0.47589746,0.76800007,0.81066674,0.8763078,1.083077,1.3587693,1.2176411,1.1355898,1.1782565,1.394872,1.8281027,1.9593848,1.8838975,2.1234872,2.6387694,2.8225644,3.764513,4.8836927,5.579488,5.7435904,5.7501545,6.009436,6.416411,7.0334363,7.834257,8.720411,9.573745,9.573745,9.091283,8.615385,8.756514,9.353847,10.614155,11.444513,11.69395,12.140308,11.329642,11.1294365,11.631591,12.402873,12.461949,12.370052,11.2672825,9.764103,8.293744,7.1122055,6.196513,6.2523084,7.0432825,8.146052,8.946873,8.4283085,8.743385,9.636104,10.742155,11.592206,11.83836,11.638155,11.339488,11.126155,11.027693,10.489437,10.902975,11.224616,11.0605135,10.660104,10.246565,10.404103,11.008,11.595488,11.362462,10.410667,9.931488,9.685334,9.347282,8.530052,8.789334,9.238976,9.498257,9.3078985,8.533334,7.860513,7.975385,8.516924,9.258667,10.131693,11.044104,11.556104,11.61518,11.401847,11.329642,11.260718,10.65354,10.102155,9.957745,10.325335,10.236719,10.259693,10.000411,9.508103,9.29477,9.468719,9.288206,9.271795,9.616411,10.187488,9.494975,9.196308,8.914052,8.539898,8.234667,7.565129,6.6067696,5.58277,4.7228723,4.266667,4.089436,3.8104618,3.5511796,3.3017437,2.9440002,2.681436,2.5304618,2.4943593,2.5009232,2.3926156,2.5042052,2.9604106,3.4592824,3.8432825,4.1091285,4.332308,4.417641,4.3290257,4.1747694,4.194462,3.948308,3.8137438,3.7907696,3.6693337,2.9965131,2.3926156,2.1956925,1.8838975,1.4375386,1.3456411,0.9517949,1.0633847,1.1191796,1.148718,1.1979488,1.339077,1.0305642,0.90912825,0.86646163,0.8960001,1.0666667,1.0568206,0.7187693,0.45292312,0.37415388,0.30194873,0.45292312,0.4594872,0.4955898,0.56451285,0.49887183,0.61374366,0.78769237,0.761436,0.6071795,0.7220513,0.6892308,0.77456415,0.8960001,1.020718,1.1815386,1.2274873,1.3226668,1.467077,1.5327181,1.2668719,1.1191796,1.024,0.9878975,1.0469744,1.2471796,1.4178462,1.6705642,1.5556924,1.1191796,0.9189744,0.8336411,0.85005134,0.93866676,1.0108719,0.9124103,1.0305642,1.5458462,1.6705642,1.2570257,0.7811283,1.1946667,0.8402052,0.39384618,0.19364104,0.23302566,0.5546667,0.58092314,0.4955898,0.48246157,0.73517954,0.8566154,1.0666667,1.4867693,2.1300514,2.8980515,3.5446157,4.6539493,6.2129235,7.683283,8.01477,9.235693,10.440206,11.021129,11.162257,11.848206,14.628103,19.226257,23.496206,24.402054,17.988924,16.91241,17.188105,17.430975,17.129026,16.636719,15.182771,14.27036,13.082257,11.569232,10.450052,10.985026,12.2847185,16.134565,21.743591,25.74113,30.017643,34.353233,37.526978,42.371284,55.78503,55.59467,58.207184,59.172108,57.068314,53.507286,48.00657,47.524105,56.142773,73.435905,94.477135,116.26011,111.32719,86.28513,57.701748,52.096004,54.21949,55.332108,54.741337,54.738056,60.58667,76.5637,80.55467,76.62606,68.94277,61.774773,59.316517,62.237545,72.126366,85.195496,92.28801,74.893135,58.335182,45.2759,37.730465,37.057644,36.50626,28.521029,20.614565,17.316103,20.17477,26.774977,28.996925,28.432413,26.184208,22.856207,17.946259,12.681848,9.03877,7.250052,5.8157954,5.225026,5.723898,5.9667697,5.366154,4.066462,3.9056413,5.4547696,7.6603084,9.130668,8.119796,6.2752824,6.9021544,7.7325134,8.149334,9.196308,10.971898,12.547283,14.073437,15.586463,17.010874,22.065233,34.248207,42.55508,39.906464,23.168001,14.572309,15.881847,17.719797,17.316103,18.484514,23.991796,26.427078,23.381334,16.790976,12.901745,10.627283,10.515693,10.929232,11.54954,13.367796,15.382976,19.393642,21.799387,22.495182,24.881233,24.198566,24.237951,23.213951,21.704206,22.642874,22.823387,24.822155,34.002052,45.44985,43.956516,38.787285,35.170464,35.190155,37.133133,35.475697,28.816412,22.367182,19.656206,18.98995,13.443283,6.2785645,3.4002054,2.789744,2.9013336,2.6387694,3.8432825,4.4964104,5.2381544,5.474462,3.387077,2.917744,3.82359,3.8071797,3.7382567,7.6603084,35.99426,36.01395,24.33313,11.923694,4.1025643,4.7622566,7.256616,9.340718,8.356103,1.2438976,2.2678976,1.7788719,1.4276924,1.6311796,1.5688206,0.7089231,0.7844103,0.76800007,0.571077,1.0404103,1.3686155,1.401436,1.6344616,1.9790771,1.7690258,2.4516926,3.6660516,3.620103,2.5107694,2.5271797,1.7558975,1.3062565,1.1684103,1.2242053,1.2603078,1.0436924,0.77128214,0.56123084,0.5546667,0.92553854,1.0272821,4.378257,9.330873,13.968411,16.121437,15.960617,12.304411,10.752001,12.393026,13.820719,18.487797,15.058052,12.3766165,12.839386,12.419283,14.549335,17.795284,18.960411,17.503181,15.547078,12.343796,9.3768215,8.139488,8.0377445,6.3868723,9.028924,5.5204105,5.2676926,8.316719,5.3694363,4.020513,6.413129,7.75877,8.408616,13.824001,11.178667,10.515693,8.178872,4.4800005,3.7054362,7.315693,10.230155,11.716924,12.885334,16.70236,15.809642,11.451077,14.953027,22.265438,13.958565,22.442669,22.107899,17.513027,13.515489,15.284514,12.84595,8.854975,8.018052,9.888822,8.887795,6.9743595,4.348718,2.1956925,1.3620514,2.3335385,2.0906668,1.1454359,0.63343596,1.142154,2.7175386,9.176616,12.228924,9.281642,3.698872,4.778667,5.0149746,6.340924,7.02359,6.11118,3.446154,1.8543591,1.6475899,1.8806155,1.9003079,1.3423591,0.46276927,0.33805132,0.34789747,0.27897438,0.31507695,0.24615386,0.17723078,0.256,0.42994875,0.44964105,0.57764107,0.636718,0.60389745,0.49887183,0.3708718,0.47589746,0.65641034,0.8763078,1.148718,1.5360001,1.3554872,1.2832822,1.3522053,1.4605129,1.3751796,1.2668719,1.2307693,1.0469744,0.72861546,0.5316923,0.571077,0.6662565,0.7318975,0.75487185,0.77128214,0.7450257,0.92553854,1.6804104,2.6912823,2.986667,2.7864618,2.4057438,1.8904617,1.6082052,2.231795,2.412308,2.162872,2.1202054,2.1431797,1.3095386,1.1191796,1.6311796,1.8182565,1.4933335,1.332513,2.1267693,2.6847181,2.5042052,2.041436,2.7306669,2.6945643,2.3269746,1.9364104,1.8051283,2.1956925,2.5042052,2.3958976,2.1497438,2.1136413,2.7044106,2.487795,1.9298463,1.9593848,2.605949,2.993231,1.3784616,0.65641034,0.6662565,1.1454359,1.7165129,2.937436,2.3105643,1.3095386,0.7056411,0.57764107,0.4660513,0.32820517,0.29210258,0.446359,0.86317956,1.3259488,1.8281027,2.1924105,2.537026,3.2623591,3.626667,3.4297438,3.0424619,2.7109745,2.5600002,2.4320002,2.28759,2.2646155,2.156308,1.3883078,1.0633847,0.96492314,0.9156924,0.83035904,0.69907695,0.57764107,0.51856416,0.5973334,0.7778462,0.9321026,0.9517949,1.2012309,1.6902566,2.294154,2.7503593,2.5698464,2.1070771,1.9922053,2.2613335,2.359795,2.8553848,2.737231,2.4746668,2.3072822,2.2613335,2.1891284,2.2153847,2.284308,2.3466668,2.3794873,2.3696413,2.0841026,1.6410258,1.273436,1.3357949,1.2242053,1.0371283,1.1552821,1.5163078,1.6213335,3.1474874,8.700719,11.021129,7.515898,0.27897438,0.99774367,1.1520001,0.9747693,0.78769237,0.9714873,0.9911796,0.892718,0.9353847,1.273436,1.9561027,1.7001027,1.9954873,1.9659488,1.522872,1.394872,2.3040001,2.0086155,1.8806155,2.2186668,2.2383592,1.7887181,1.4736412,1.4276924,1.529436,1.404718,1.1684103,1.3981539,1.6475899,1.585231,1.0043077,1.1355898,1.1848207,1.020718,0.6465641,0.21989745,0.108307704,0.032820515,0.0,0.016410258,0.07548718,0.29210258,0.33476925,0.37415388,0.4660513,0.54482055,0.77128214,0.7450257,0.81066674,1.0601027,1.3259488,1.1716924,1.1257436,1.1749744,1.3292309,1.6278975,1.9331284,1.9265642,2.1792822,2.6289232,2.546872,3.4921029,4.578462,5.2020516,5.277539,5.2512827,5.5729237,6.12759,6.764308,7.509334,8.562873,9.176616,9.196308,9.07159,9.140513,9.649232,9.984001,10.505847,11.10318,11.52,11.346052,10.417232,9.993847,10.696206,11.999181,12.225642,11.874462,11.224616,10.052924,8.677744,7.9524107,7.0793853,6.8397956,7.1614366,7.6012316,7.3452315,7.2992826,8.434873,9.45559,10.049642,10.912822,11.746463,11.782565,11.392001,10.873437,10.443488,9.570462,9.645949,9.544206,9.005949,8.621949,8.421744,8.87795,9.938052,10.925949,10.555078,10.525539,10.269539,9.974154,9.603283,8.884514,9.114257,9.156924,8.838565,8.139488,7.204103,6.5280004,6.380308,6.9842057,8.254359,9.80677,10.916103,11.424822,11.339488,11.024411,11.195078,11.989334,11.684103,11.175385,10.729027,9.977437,9.511385,9.613129,9.590155,9.383386,9.554052,9.416205,8.631796,8.444718,8.999385,9.344001,9.212719,9.255385,8.891078,8.185436,7.830975,6.9677954,5.7665644,4.7392826,4.132103,3.9417439,3.6660516,3.255795,2.92759,2.737231,2.5731285,2.4320002,2.297436,2.2416413,2.2613335,2.2547693,2.4582565,2.9078977,3.5511796,4.1846156,4.450462,4.4242053,4.4340515,4.164923,3.817026,4.1058464,4.066462,3.9548721,3.945026,3.7382567,2.556718,1.9462565,1.847795,1.7952822,1.6443079,1.5721027,1.1585642,1.4276924,1.7066668,1.6016412,1.1684103,0.8992821,0.7778462,0.72861546,0.9189744,1.2964103,1.6016412,1.2242053,0.79097444,0.56451285,0.55794877,0.5349744,0.65641034,0.5677949,0.52512825,0.56123084,0.48902568,0.67282057,0.77128214,0.7417436,0.6498462,0.6859488,0.6629744,0.69251287,0.7844103,0.9353847,1.1454359,1.1815386,1.1257436,1.1388719,1.204513,1.1454359,1.2898463,1.4276924,1.5195899,1.6278975,1.9068719,2.1136413,2.166154,1.782154,1.1257436,0.80738467,0.7220513,0.8205129,0.92553854,0.8992821,0.65641034,0.9124103,1.270154,1.2865642,0.97805136,0.79425645,1.5392822,1.1552821,0.636718,0.40369233,0.3052308,0.69579494,0.7844103,0.8402052,1.0535386,1.5425643,1.7591796,2.3466668,3.446154,4.841026,5.9503593,6.5378466,6.931693,7.6209235,8.854975,10.650257,10.9915905,11.654565,11.336206,10.614155,11.933539,14.555899,19.416616,22.882463,22.95795,19.272207,19.833437,20.94277,21.284103,20.027079,16.83036,13.082257,11.779283,11.237744,10.755282,10.620719,11.204924,14.500104,21.129848,28.133745,28.977234,30.33272,32.610462,34.980106,38.242466,44.84595,45.568005,45.636925,43.086773,37.7239,31.143387,28.691694,29.285746,33.870773,41.521233,49.457233,58.417236,55.72267,42.899696,29.09867,31.097439,37.38585,43.17539,47.872005,54.262157,68.5555,94.25067,98.49765,88.66462,74.32534,67.24596,67.049034,64.46606,61.535183,61.59754,69.27754,72.254364,62.926773,48.92554,36.10585,28.550566,23.545437,17.91672,15.786668,18.002052,22.14072,25.74113,25.662361,23.112207,20.588308,21.881437,22.662565,19.488823,13.843694,8.064001,5.3398976,5.366154,5.8847184,5.8420515,5.093744,4.4110775,4.972308,5.504,6.091488,6.498462,6.180103,6.9120007,8.805744,9.711591,9.403078,9.596719,9.842873,10.791386,11.437949,11.762873,12.727796,19.43959,29.797747,32.997746,26.095592,14.024206,12.6063595,16.098463,17.58195,16.105026,16.679386,23.171284,24.986258,21.782976,15.589745,10.804514,9.386667,9.527796,10.108719,11.011283,13.121642,14.221129,15.770258,16.239592,16.032822,17.47036,20.998566,21.385847,21.10031,21.507284,22.889027,21.5959,22.534565,30.693747,41.967594,43.152412,33.26359,31.589746,33.158566,34.146465,31.875284,25.72472,21.136412,19.524925,19.045746,14.601848,7.450257,3.9844105,3.2820516,3.8728209,3.7382567,3.6529233,3.639795,4.2929235,4.827898,3.0818465,2.5928206,6.738052,6.9710774,4.0467696,8.024616,30.949745,28.928001,20.74913,13.853539,4.332308,3.2951798,5.9667697,8.664616,8.178872,1.7690258,1.7099489,1.3357949,1.7263591,2.556718,2.1070771,1.079795,1.3653334,1.2307693,0.5513847,0.80738467,1.7132308,1.7723079,2.103795,2.4549747,1.2209232,1.8937438,3.0654361,3.1770258,2.3072822,2.1956925,1.9035898,1.6836925,1.6246156,1.6640002,1.6016412,1.2964103,1.2307693,1.1027694,0.9124103,0.9616411,1.0338463,2.1530259,4.95918,8.871386,12.071385,13.400617,12.442257,11.562668,11.392001,10.817642,23.40431,15.885129,8.644924,8.999385,11.185231,13.735386,17.61477,20.14195,19.905643,16.768002,14.50995,11.218052,8.477539,6.9120007,6.180103,6.2523084,3.882667,4.8082056,10.791386,19.590565,7.958975,7.3025646,12.849232,18.707693,17.851078,12.33395,12.458668,10.932513,6.7938466,5.402257,8.710565,11.907283,17.650873,23.80472,23.45354,23.440413,18.500925,13.74195,11.395283,10.834052,10.174359,13.269335,15.783386,15.284514,11.23118,7.680001,6.744616,9.02236,11.963078,9.888822,5.7009234,2.2646155,1.3423591,2.481231,3.006359,0.80738467,1.595077,2.6453335,2.8127182,2.5337439,3.7284105,7.0400004,7.6701546,5.5958977,5.586052,5.8289237,9.452309,10.59118,8.182155,5.933949,4.141949,2.7306669,2.793026,3.7842054,3.5413337,1.0010257,0.35774362,0.36430773,0.38728207,0.4135385,0.31507695,0.28225642,0.38400003,0.54482055,0.5349744,0.7417436,0.9944616,1.1060513,0.9419488,0.44307697,0.5874872,0.6629744,0.6859488,0.7056411,0.7778462,0.75487185,0.8041026,0.97805136,1.204513,1.2668719,0.9124103,0.85005134,0.8566154,0.8008206,0.64000005,0.65312827,0.7384616,0.7089231,0.5284103,0.32164106,0.3314872,0.58420515,1.3883078,2.5009232,3.0982566,2.6715899,2.8192823,2.7470772,2.4385643,2.6715899,2.4516926,2.1398976,1.8510771,1.6508719,1.5425643,1.2242053,1.4178462,1.394872,0.9911796,0.6268718,1.273436,1.7362052,1.7493335,1.5721027,1.9987694,2.0118976,1.7952822,1.5983591,1.5491283,1.6475899,1.9659488,1.9265642,1.5458462,1.1520001,1.3718976,1.4211283,1.654154,1.8248206,2.0053334,2.5796926,0.6629744,0.3117949,0.6301539,1.2274873,2.228513,1.5064616,1.2077949,0.90912825,0.5284103,0.32164106,0.30851284,0.3052308,0.3052308,0.3511795,0.5349744,0.9353847,1.211077,1.6016412,2.162872,2.7634873,3.5544617,3.7087183,3.3345644,2.6945643,2.1825643,2.034872,2.044718,1.910154,1.585231,1.2668719,1.0108719,0.892718,0.8730257,0.8467693,0.6268718,0.5021539,0.51856416,0.65969235,0.8467693,0.9321026,0.892718,0.92225647,1.1716924,1.6738462,2.3335385,2.3105643,1.8642052,1.7066668,1.9692309,2.2121027,2.5895386,2.878359,2.6322052,1.9922053,1.6640002,1.5031796,1.6836925,1.9396925,2.1366155,2.2580514,2.0020514,1.7362052,1.4244103,1.142154,1.0666667,1.3357949,1.339077,1.8510771,2.7076926,2.793026,5.0018463,11.175385,12.445539,7.0531287,0.3511795,0.8763078,0.86974365,0.75487185,0.78769237,1.0666667,0.98133343,1.273436,1.4145643,1.3587693,1.5425643,1.4802053,1.8412309,1.8510771,1.467077,1.3587693,1.467077,1.5425643,1.8773335,2.300718,2.166154,1.5195899,1.0469744,0.9419488,1.1848207,1.5261539,1.2209232,1.0535386,1.0765129,1.1881026,1.1126155,1.0404103,1.0305642,0.9353847,0.65969235,0.18379489,0.06235898,0.013128206,0.006564103,0.026256412,0.07548718,0.23630771,0.27569234,0.37743592,0.60389745,0.88615394,0.8598975,0.761436,0.8467693,1.0929232,1.1913847,1.020718,1.0765129,1.1946667,1.273436,1.2964103,1.5163078,1.8018463,2.0742567,2.3171284,2.546872,3.062154,3.8662567,4.3684106,4.519385,4.8377438,5.362872,6.0061545,6.701949,7.3058467,7.5979495,8.513641,8.779488,9.025641,9.416205,9.6754875,9.980719,9.938052,9.875693,9.931488,10.039796,9.110975,9.156924,9.862565,10.834052,11.565949,11.61518,11.158976,10.19077,9.015796,8.27077,7.9524107,7.9819493,7.9097443,7.6143594,7.3091288,7.076103,8.474257,9.764103,10.315488,10.620719,11.365745,11.16554,10.561642,9.931488,9.4916935,8.979693,8.858257,8.503796,7.827693,7.27959,7.5487185,7.5487185,8.080411,9.028924,9.383386,10.115283,10.069334,9.869129,9.750975,9.567181,9.4457445,9.278359,8.854975,8.109949,7.0957956,7.0826674,6.8496413,6.8397956,7.4141545,8.881231,10.811078,11.67754,11.638155,11.388719,12.1468725,12.658873,13.078976,13.072412,12.27159,10.269539,9.547488,9.29477,8.868103,8.372514,8.651488,8.933744,8.772923,8.644924,8.697436,8.759795,8.635077,9.199591,9.340718,8.674462,7.5388722,6.3901544,5.142975,4.269949,3.8564105,3.6004105,3.1967182,2.8947694,2.546872,2.2186668,2.1825643,2.0611284,2.3401027,2.4615386,2.3401027,2.3663592,2.986667,3.3805132,3.8137438,4.1682053,3.9351797,4.1550775,4.3290257,4.1517954,3.7152824,3.495385,3.8498464,3.892513,3.639795,3.0949745,2.228513,1.8609232,1.7066668,1.8084104,1.9856411,1.8149745,1.4900514,1.2603078,1.6246156,1.7788719,1.4769232,1.020718,1.0371283,1.3095386,1.4375386,1.4276924,1.6640002,1.4998976,1.273436,1.083077,0.892718,0.54482055,0.5218462,0.46276927,0.44964105,0.47589746,0.45292312,0.53825647,0.6071795,0.6892308,0.75487185,0.7220513,0.76800007,0.8598975,0.92225647,0.9616411,1.0699488,0.892718,0.892718,0.9353847,0.9616411,0.99774367,1.2504616,1.4244103,1.5064616,1.5688206,1.7624617,1.910154,1.6246156,1.1520001,0.75487185,0.7122052,0.9189744,1.1848207,1.204513,1.0043077,0.92553854,1.142154,1.1224617,0.92553854,0.69251287,0.6465641,0.98133343,0.9944616,0.764718,0.4660513,0.37743592,0.86646163,1.3456411,1.6804104,1.9003079,2.2121027,3.2525132,4.8640003,6.4754877,7.9097443,9.380103,9.38995,10.601027,11.270565,11.142565,11.431385,11.303386,10.883283,10.824206,11.638155,13.689437,16.177233,17.99877,19.74154,22.101336,25.875694,24.192001,23.913027,23.02031,20.519386,16.452925,13.945437,12.402873,11.185231,10.499283,11.401847,12.934566,15.205745,19.419899,24.31672,26.194054,27.264002,28.150156,30.0439,32.774567,34.786465,33.62462,31.977028,29.161028,26.272823,26.187489,25.314463,26.971899,28.905027,30.263798,31.609438,39.250053,40.61867,35.360825,28.455387,30.244104,32.92554,36.34544,41.347286,50.786465,69.53355,108.89847,124.48821,114.69129,89.908516,72.50708,63.36657,56.29703,48.640003,42.450054,44.48493,58.21375,62.027493,53.83549,38.308105,26.87672,20.788515,16.538258,14.989129,16.341335,20.138668,22.87918,22.052105,19.534771,17.483488,18.330257,20.371695,20.082872,16.351181,10.223591,4.9132314,5.0642056,5.622154,6.189949,6.3179493,5.4974365,5.0116925,5.074052,5.474462,5.927385,6.058667,6.75118,7.2664623,7.3780518,7.171283,7.0334363,7.062975,7.4240007,7.755488,8.329846,10.066052,15.392821,20.109129,19.433027,13.636924,8.03118,11.211488,13.984821,14.985847,15.238565,18.166155,23.158155,25.16677,21.051079,13.607386,11.585642,9.8363085,9.622975,9.852718,10.013539,10.194052,12.511181,14.158771,14.316309,13.771488,14.920206,18.710976,18.901335,18.94072,19.784206,19.872822,20.775387,22.442669,29.216824,38.245747,39.476517,30.526361,27.753027,29.239798,30.680618,25.393232,22.308104,20.33231,19.777643,18.386053,11.355898,5.920821,3.4789746,3.1015387,3.5446157,3.2623591,2.2088206,2.1169233,2.930872,3.7809234,2.9735386,3.5478978,6.7577443,7.4207187,6.7872825,12.540719,21.602463,19.810463,15.698052,12.035283,5.8223596,3.8367183,8.704,10.886565,7.6274877,2.917744,2.3860514,1.6640002,2.0644104,3.1376412,2.6683078,2.6584618,2.484513,1.8510771,1.0896411,1.1520001,2.1989746,2.3138463,2.5304618,2.7076926,1.5130258,2.3302567,3.5052311,3.4067695,2.2153847,1.9298463,1.5688206,1.7099489,1.9331284,1.9692309,1.723077,4.2502565,2.9735386,1.2570257,0.7975385,1.6082052,2.5895386,5.405539,6.816821,7.3452315,11.277129,10.722463,16.807386,17.188105,11.815386,12.931283,14.8709755,10.725744,8.195283,9.242257,10.098872,12.36677,15.734155,18.353231,18.563284,14.890668,11.644719,9.921641,8.100103,5.937231,4.568616,3.8400004,2.0611284,5.034667,9.91836,5.225026,6.6592827,8.234667,10.8307705,14.089848,16.436514,12.297847,9.363693,9.905231,12.074668,9.941334,8.444718,10.069334,15.07118,20.266668,19.032618,25.5639,19.59713,14.411489,15.232001,19.232822,15.878566,18.064411,16.262566,11.109744,13.403898,17.703386,14.299898,12.504617,13.587693,10.791386,4.279795,5.0674877,6.5378466,5.225026,0.80738467,0.5152821,0.95835906,1.4998976,2.1103592,3.3641028,4.4242053,8.1755905,9.468719,8.608821,11.369026,8.411898,9.636104,10.039796,8.356103,7.059693,7.2960005,5.5072823,4.4701543,4.414359,3.0260515,1.0535386,0.45620516,0.48246157,0.6662565,0.827077,0.74830776,0.6104616,0.5874872,0.67282057,0.67938465,1.2996924,1.4408206,1.394872,1.211077,0.7122052,0.702359,0.78769237,0.79097444,0.7187693,0.75487185,0.64000005,0.7253334,0.92225647,1.0699488,0.92553854,0.764718,0.702359,0.7089231,0.7187693,0.6301539,0.6498462,0.67282057,0.5940513,0.46276927,0.47917953,0.39384618,0.4594872,1.014154,2.0644104,3.2689233,3.2722054,3.367385,3.2295387,2.8521028,2.537026,2.4910772,2.3335385,2.0709746,1.7591796,1.4933335,1.2340513,1.4506668,1.5589745,1.2373334,0.44307697,0.9321026,1.2570257,1.4342566,1.7329233,2.6584618,2.034872,1.5589745,1.332513,1.3883078,1.6738462,1.529436,1.1716924,1.0272821,1.1815386,1.3620514,1.3128207,1.3226668,1.585231,2.034872,2.3335385,1.0043077,0.7187693,0.8205129,0.9878975,1.2274873,1.463795,1.4473847,1.0896411,0.65312827,0.74830776,0.3052308,0.2231795,0.28225642,0.35446155,0.4135385,0.64000005,0.8566154,1.1027694,1.4178462,1.8215386,2.166154,2.3302567,2.409026,2.4320002,2.3762052,2.3171284,2.231795,1.975795,1.5819489,1.2537436,0.9878975,0.84348726,0.827077,0.82379496,0.61374366,0.571077,0.53825647,0.65312827,0.85005134,0.8566154,1.0929232,1.2931283,1.3029745,1.2635899,1.5885129,1.847795,1.9068719,1.8806155,1.8674873,1.9429746,2.166154,2.2219489,1.9364104,1.4309745,1.1520001,1.2931283,1.6147693,1.7887181,1.785436,1.8674873,1.9528207,1.6836925,1.3587693,1.1815386,1.276718,1.8576412,1.8937438,4.4865646,7.9130263,5.6254363,11.943385,17.270155,15.563488,7.4830775,0.4004103,0.56451285,0.67938465,0.64000005,0.6301539,1.1060513,0.69579494,1.0075898,1.2373334,1.2996924,1.8346668,1.3817437,1.5425643,1.8149745,1.8740515,1.5885129,1.8576412,1.9692309,2.0841026,2.172718,2.0217438,1.8018463,1.3850257,1.0732309,1.0404103,1.3423591,1.4080001,1.2668719,1.1224617,1.0666667,1.0896411,1.1913847,1.0502565,0.7975385,0.49887183,0.17066668,0.03938462,0.0032820515,0.006564103,0.029538464,0.08861539,0.15097436,0.25271797,0.39712822,0.58092314,0.82379496,1.0338463,0.90584624,0.8960001,1.079795,1.1782565,1.017436,1.2012309,1.3161026,1.273436,1.3095386,1.5688206,1.6114873,1.8576412,2.422154,3.121231,3.3017437,3.6430771,3.945026,4.2338467,4.775385,5.7009234,6.3442054,6.7117953,7.0400004,7.781744,8.756514,8.546462,8.136206,8.067283,8.441437,9.068309,8.805744,8.461129,8.618668,9.636104,9.334154,9.107693,9.124104,9.590155,10.771693,11.542975,11.460924,10.587898,9.357129,8.562873,7.640616,7.3353853,7.525744,7.781744,7.3583593,7.653744,8.523488,9.216001,9.498257,9.655796,10.692924,10.774975,10.505847,9.987283,8.795898,8.625232,8.67118,8.388924,7.637334,6.669129,6.4590774,6.340924,6.6100516,7.171283,7.565129,8.073847,8.490667,9.065026,9.724719,10.069334,9.682052,8.992821,8.224821,7.509334,6.889026,6.885744,6.9349747,7.0892315,7.512616,8.490667,10.000411,10.791386,11.158976,11.651283,13.062565,13.955283,14.851283,14.834873,13.679591,11.844924,10.43036,9.485129,8.730257,8.352821,8.992821,9.488411,9.091283,8.720411,8.536616,7.9524107,8.661334,9.189744,9.176616,8.379078,6.7085133,5.540103,4.601436,3.9286156,3.511795,3.2951798,2.8455386,2.609231,2.4681027,2.3433847,2.2186668,2.0775387,2.4057438,2.5698464,2.5698464,3.0227695,3.3641028,3.3280003,3.498667,3.9614363,4.315898,4.164923,3.8432825,3.7087183,3.9811285,4.7261543,4.6112823,4.2601027,3.6430771,2.8882053,2.2777438,2.0086155,2.294154,2.553436,2.487795,2.0709746,1.3883078,1.2537436,1.3456411,1.3915899,1.3193847,1.2373334,1.2471796,1.3883078,1.4178462,1.3751796,1.5589745,1.3095386,1.1060513,0.96492314,0.8041026,0.45620516,0.4266667,0.42994875,0.44307697,0.45292312,0.46933338,0.58092314,0.58420515,0.636718,0.7318975,0.7056411,0.7450257,0.86646163,0.9485129,0.97805136,1.0633847,0.9189744,0.8172308,0.77128214,0.81066674,0.9878975,1.014154,1.086359,1.2242053,1.401436,1.5491283,1.463795,1.0666667,0.69907695,0.5349744,0.60389745,0.9156924,1.2668719,1.2438976,0.8795898,0.6892308,0.88943595,0.88615394,0.7089231,0.5349744,0.69251287,0.85005134,0.764718,0.6170257,0.5152821,0.48902568,0.60389745,0.9189744,1.401436,2.0118976,2.6912823,4.2502565,6.2096415,7.9852314,9.45559,10.94236,11.995898,13.551591,15.38954,17.030565,17.742771,15.527386,14.39836,14.549335,15.714462,17.142155,18.034874,18.596104,19.866259,22.304823,25.80677,24.592413,25.334156,24.096823,20.361847,17.043694,14.372104,12.84595,11.835078,11.654565,13.584412,13.367796,14.093129,17.234053,21.648413,23.555285,23.584822,23.768618,25.107695,26.857027,26.558361,25.993849,26.486156,27.421541,28.17313,28.114054,28.714668,30.375387,28.983797,25.232412,24.618668,34.917747,36.496414,34.68144,33.3719,35.045746,37.40554,38.63631,38.928413,42.13498,55.7719,96.141136,122.63714,123.60206,101.40883,72.47755,59.106464,53.43508,46.85457,38.95139,37.477745,55.397747,60.389748,54.37703,42.25313,31.878567,23.811283,19.577436,17.48677,16.626873,16.873028,18.36636,16.968206,15.189335,14.473847,15.169642,16.676104,17.667284,16.20677,11.972924,6.242462,5.1167183,5.865026,6.616616,6.633026,6.3343596,6.160411,5.6418467,5.474462,5.865026,6.547693,6.377026,6.173539,6.0685134,5.9503593,5.4580517,5.412103,5.3234878,5.684513,6.6625648,8.109949,11.565949,13.15118,11.71036,8.477539,7.0793853,9.567181,10.965334,12.2157955,13.860104,16.01313,20.83118,23.328823,19.86954,12.914873,11.021129,10.134975,10.660104,10.896411,10.417232,10.082462,11.395283,13.098668,14.089848,14.674052,16.561232,18.340103,17.046976,16.321642,16.981335,17.050259,18.58954,21.842052,28.114054,33.88718,30.841438,25.642668,23.54872,24.792618,25.859283,19.488823,17.54913,18.281027,19.495386,18.041437,9.783795,5.1889234,3.5183592,3.1671798,3.2065644,3.3805132,2.0217438,1.8379488,2.2711797,2.6978464,2.422154,3.3312824,4.824616,5.7468724,8.43159,18.697847,29.96513,34.28431,25.475285,9.540924,4.6834874,3.1803079,9.383386,12.461949,9.248821,4.240411,2.8225644,1.7920002,1.9495386,2.7831798,2.4582565,2.6683078,3.1081028,2.802872,2.0086155,2.1956925,2.537026,2.409026,2.4713848,2.4681027,1.2471796,3.2754874,4.9394875,4.7917953,3.121231,1.972513,1.3718976,1.4998976,1.8313848,2.4516926,4.0336413,4.2436924,3.2328207,2.0250258,1.2176411,0.9747693,1.654154,3.8301542,4.6145644,4.841026,9.065026,10.581334,16.44636,17.017437,13.528616,18.090668,12.097642,8.4053335,7.824411,8.845129,7.6570263,16.761436,26.095592,30.821747,28.78031,20.489847,11.579078,9.69518,7.4797955,3.9614363,4.5587697,3.6758976,2.0906668,2.7569232,4.325744,1.1552821,4.6769233,7.7718983,9.668923,11.211488,14.838155,10.433641,7.6012316,8.467693,11.510155,11.562668,11.670976,10.551796,11.936821,16.8599,23.670156,20.424206,18.01518,17.851078,19.580719,21.103592,16.31836,12.987078,11.250873,10.975181,11.766154,12.58995,12.041847,11.700514,10.699488,5.7435904,2.231795,3.3575387,4.0434875,2.6354873,0.8730257,1.4211283,1.1224617,1.0075898,1.9200002,4.5128207,4.0369234,6.636308,7.748924,8.602257,16.196924,9.997129,9.705027,9.984001,8.681026,6.8266673,6.9120007,5.402257,4.1452312,3.446154,2.0742567,3.3509746,3.18359,2.665026,2.2711797,1.8740515,1.4998976,0.98461545,0.67938465,0.67282057,0.8172308,1.6640002,1.9626669,2.0545642,1.9462565,1.3357949,1.1060513,0.99774367,0.86317956,0.69251287,0.636718,0.77456415,0.892718,1.1060513,1.2898463,1.086359,0.86646163,0.81394875,0.7975385,0.7450257,0.63343596,0.6235898,0.60389745,0.5152821,0.4594872,0.702359,0.58420515,0.5021539,0.79097444,1.6049232,2.9078977,3.383795,4.06318,4.089436,3.2886157,2.162872,1.8773335,2.0217438,2.0644104,1.8051283,1.3883078,1.2996924,1.339077,1.4703591,1.3718976,0.46933338,0.51856416,0.7253334,0.9747693,1.4998976,2.878359,2.0512822,1.4112822,1.1191796,1.1520001,1.2832822,1.0666667,0.86974365,0.84348726,0.9747693,1.1027694,1.0666667,1.1716924,1.4276924,1.7132308,1.7690258,1.2537436,0.79425645,0.6268718,0.73517954,0.8467693,1.2209232,1.6344616,1.5163078,0.99774367,0.9189744,0.37743592,0.3446154,1.1158975,2.1956925,2.294154,0.77128214,0.6170257,2.2908719,4.1747694,2.5665643,1.463795,1.2504616,1.6475899,2.1103592,1.8116925,1.8215386,1.6771283,1.4867693,1.3128207,1.1881026,1.0075898,0.86317956,0.78769237,0.78769237,0.8205129,0.761436,0.65969235,0.6268718,0.67282057,0.7122052,0.92225647,1.1454359,1.1881026,1.0732309,1.0469744,1.595077,1.9265642,1.9889232,1.8707694,1.8051283,1.9429746,1.8543591,1.6410258,1.4112822,1.2964103,1.2373334,1.5360001,1.7690258,1.8182565,1.8609232,1.8412309,1.6246156,1.4211283,1.4145643,1.7755898,2.1497438,4.9427695,9.032206,11.894155,9.590155,10.774975,16.098463,14.838155,6.550975,1.0699488,0.49230772,0.39384618,0.36758977,0.4266667,1.0043077,0.8172308,0.955077,1.1815386,1.4342566,1.8510771,1.5885129,1.4834872,1.6311796,1.8116925,1.5195899,1.7657437,1.8576412,1.9987694,2.103795,1.7920002,1.7558975,1.5721027,1.4703591,1.4736412,1.4145643,1.5392822,1.4506668,1.214359,1.0043077,1.1093334,1.2209232,0.99774367,0.6498462,0.3249231,0.10502565,0.01969231,0.0,0.013128206,0.059076928,0.15425642,0.17723078,0.3249231,0.47261542,0.6104616,0.86317956,1.1684103,1.0108719,0.9189744,1.0568206,1.2209232,1.1782565,1.276718,1.3062565,1.2537436,1.3128207,1.6114873,1.6475899,1.8215386,2.2744617,2.8717952,3.2689233,3.4592824,3.7087183,4.135385,4.7327185,5.4875903,6.298257,6.51159,6.4065647,7.197539,8.54318,8.441437,8.008205,7.9491286,8.562873,8.136206,7.578257,7.5520005,8.12636,8.786052,8.910769,8.4972315,8.608821,9.435898,10.328616,11.155693,11.385437,10.840616,9.757539,8.792616,7.4830775,7.0990777,7.3091288,7.634052,7.4141545,7.433847,7.6570263,8.024616,8.4512825,8.838565,9.93477,10.006975,9.544206,8.864821,8.136206,8.41518,9.035488,8.828718,7.6767187,6.5050263,6.052103,6.2194877,6.482052,6.5444107,6.370462,6.445949,6.695385,7.197539,7.860513,8.425026,8.041026,7.243488,6.6067696,6.373744,6.47877,6.377026,6.482052,6.8299494,7.387898,8.054154,9.019077,9.7903595,10.220308,10.742155,12.373334,13.709129,14.739694,14.723283,13.787898,12.914873,11.027693,9.344001,8.28718,8.093539,8.795898,8.789334,8.6580515,8.411898,8.021334,7.430565,8.441437,8.999385,8.726975,7.64718,6.160411,5.3398976,4.6834874,4.0369234,3.4264617,3.0720003,2.7470772,2.6322052,2.5632823,2.5271797,2.6584618,2.4320002,2.300718,2.2383592,2.4451284,3.3444104,3.570872,3.4034874,3.3805132,3.6004105,3.751385,3.6594875,3.4789746,3.8104618,4.535795,4.8049235,4.378257,3.6791797,3.0227695,2.5435898,2.2153847,2.3663592,2.5009232,2.5173335,2.3729234,2.0808206,2.3401027,1.7132308,1.3653334,1.0994873,0.94523084,1.1520001,1.2176411,1.2504616,1.204513,1.1093334,1.083077,0.8402052,0.702359,0.6826667,0.67610264,0.47589746,0.4201026,0.4135385,0.44307697,0.48574364,0.51856416,0.60061544,0.57764107,0.57764107,0.6170257,0.61374366,0.69251287,0.81394875,0.90256417,0.9682052,1.1158975,1.4276924,1.2406155,0.9747693,0.8992821,1.1158975,1.0469744,0.99774367,1.0338463,1.1323078,1.1848207,0.9878975,0.6498462,0.4955898,0.574359,0.65312827,0.8598975,1.1782565,1.1158975,0.6859488,0.39712822,0.62030774,0.702359,0.6071795,0.48902568,0.69907695,0.7975385,0.6071795,0.45292312,0.446359,0.46276927,0.33805132,0.56123084,1.1716924,2.1398976,3.3575387,5.3366156,7.515898,9.222565,10.390975,11.579078,13.659899,15.514257,18.372925,21.888002,24.132925,22.367182,21.03795,20.755693,21.293951,21.609028,21.907694,22.137438,22.816822,24.090258,25.721437,24.864822,25.330873,23.706259,20.289642,19.124514,15.07118,13.761642,13.387488,13.587693,15.458463,14.772514,14.490257,16.000002,18.84554,20.729437,21.343182,22.15713,23.240208,24.323284,24.769644,25.399797,26.607592,28.928001,31.474874,31.917952,31.855593,32.623592,31.560207,29.689438,31.721027,40.192,39.145027,36.657234,35.908924,35.186874,36.260105,37.572926,35.488823,32.41026,36.77867,65.237335,94.473854,107.733345,97.53601,65.69026,57.035492,54.86934,50.087387,42.404106,40.323284,53.868313,56.579285,52.864002,46.175182,39.01375,28.934566,23.046566,19.574156,17.06995,14.375385,13.824001,12.491488,11.867898,12.370052,13.344822,13.948719,14.943181,14.972719,12.950975,8.057437,6.2162056,6.518154,6.892308,6.701949,6.7183595,7.1581545,6.9842057,7.0793853,7.686565,8.434873,6.3376417,5.2480006,4.84759,4.644103,3.9778464,3.9581542,4.1189747,4.6605134,5.6976414,7.2664623,9.409642,9.222565,7.817847,6.5280004,6.8955903,7.972103,9.170052,10.886565,12.744206,13.61395,18.51077,20.969027,18.356514,12.599796,10.154668,10.371283,11.0375395,11.1983595,10.791386,10.663385,11.136001,12.888617,14.884104,17.001026,20.023796,18.182566,15.983591,15.222155,15.78995,15.658668,17.08636,20.676924,25.081438,27.720207,24.77949,22.928411,20.118977,19.465847,19.590565,14.598565,13.774771,16.01641,17.772308,16.128002,8.812308,4.5817437,3.767795,3.7743592,3.5544617,3.626667,2.3236926,2.2711797,2.4057438,2.2514873,1.9364104,5.98318,6.8365135,6.675693,9.475283,20.985437,32.518566,35.96472,25.1799,7.4469748,3.4625645,2.612513,8.625232,12.461949,10.581334,4.916513,3.383795,1.9889232,1.9364104,2.7208207,2.1300514,2.297436,4.017231,4.089436,2.5928206,2.8914874,2.674872,2.4024618,2.228513,1.9232821,0.86317956,3.4067695,5.933949,6.76759,5.5729237,3.3641028,1.9396925,1.5163078,1.719795,2.605949,4.6769233,3.7415388,3.4921029,3.05559,2.0578463,0.61374366,1.1027694,2.1858463,2.665026,3.239385,6.482052,8.461129,11.116308,12.182976,14.480412,25.895386,12.268309,7.0990777,7.752206,11.172104,13.8765135,20.112411,30.893951,35.70872,31.209028,21.19877,11.631591,7.890052,4.97559,2.349949,3.9187696,3.1409233,2.100513,1.2471796,0.78769237,0.7122052,2.7798977,5.874872,7.936001,9.235693,12.3766165,8.822155,10.873437,10.489437,7.325539,8.707283,12.304411,13.50236,14.024206,15.704617,20.483284,14.903796,15.540514,16.787693,16.57436,16.374155,13.397334,8.208411,6.8988724,9.170052,8.320001,5.9667697,6.7840004,7.2336416,5.5630774,1.8051283,0.88287187,2.3663592,2.9538465,2.0775387,1.8904617,2.7700515,1.7723079,1.1027694,1.9495386,4.4701543,3.895795,4.384821,6.4590774,10.59118,17.19795,11.208206,11.323078,11.1983595,8.838565,6.5903597,5.467898,4.5522056,3.498667,2.3827693,1.6771283,4.699898,5.113436,4.240411,3.0358977,2.0808206,1.6672822,1.1290257,0.955077,1.1585642,1.2931283,1.7723079,2.0512822,2.1530259,2.0151796,1.4834872,1.2307693,1.079795,0.88287187,0.64000005,0.49887183,0.7450257,0.9124103,1.1520001,1.394872,1.3423591,1.014154,0.97805136,0.9189744,0.7515898,0.6170257,0.63343596,0.67938465,0.6071795,0.4955898,0.6662565,0.6662565,0.60389745,0.6826667,1.079795,1.9626669,2.7208207,3.7743592,4.007385,3.2262566,2.162872,1.6443079,1.7427694,1.9003079,1.8018463,1.401436,1.2898463,1.2668719,1.3653334,1.3718976,0.81066674,0.6170257,0.52512825,0.5973334,1.0404103,2.2055387,1.7329233,1.2471796,0.9485129,0.8598975,0.8402052,0.7122052,0.7187693,0.77456415,0.8402052,0.8992821,0.9616411,1.0994873,1.2438976,1.3226668,1.2504616,1.0666667,0.7811283,0.6268718,0.6465641,0.7089231,0.9353847,1.4769232,1.522872,1.0699488,0.9124103,0.60389745,0.56123084,1.9692309,4.3290257,5.4613338,2.609231,1.2274873,3.2361028,6.672411,5.6976414,1.6672822,1.7591796,3.0391798,3.7382567,3.2656412,1.5885129,1.014154,1.0010257,1.142154,1.1618463,1.0404103,0.9485129,0.8566154,0.81394875,0.92553854,0.83035904,0.7253334,0.6465641,0.6071795,0.61374366,0.7122052,0.85005134,0.93866676,0.92553854,0.8205129,1.273436,1.6475899,1.8740515,1.9331284,1.8773335,1.8215386,1.7558975,1.6377437,1.5031796,1.4802053,1.3029745,1.4834872,1.6771283,1.7755898,1.8904617,1.9068719,1.719795,1.6508719,1.8116925,2.100513,2.2186668,6.235898,10.171078,11.451077,8.920616,9.360411,15.337027,14.188309,5.802667,2.6322052,1.1552821,0.5218462,0.256,0.27897438,0.892718,0.9878975,0.95835906,1.1158975,1.4473847,1.595077,1.7624617,1.585231,1.7329233,2.048,1.5556924,1.5491283,1.5261539,1.7001027,1.9200002,1.6508719,1.5983591,1.5688206,1.6672822,1.7657437,1.4998976,1.4736412,1.4211283,1.2406155,1.020718,1.0436924,1.0994873,0.8763078,0.51856416,0.18379489,0.036102567,0.006564103,0.0032820515,0.029538464,0.098461546,0.2297436,0.22646156,0.41025645,0.5973334,0.75487185,1.0108719,1.1848207,1.017436,0.92553854,1.0469744,1.2406155,1.1782565,1.2012309,1.2603078,1.3029745,1.2635899,1.5327181,1.5983591,1.7526156,2.0906668,2.487795,2.9768207,3.3280003,3.7809234,4.3684106,4.896821,5.228308,5.930667,6.1341543,6.038975,6.9152827,8.057437,8.001641,7.64718,7.5454364,7.9228725,6.8660517,6.3474874,6.8463597,7.958975,8.408616,8.726975,8.448001,8.805744,9.813334,10.253129,10.860309,11.034257,10.748719,9.997129,8.779488,7.5388722,7.2336416,7.0990777,6.9710774,7.282872,7.0400004,6.498462,6.5805135,7.433847,8.457847,9.488411,9.232411,8.484103,7.906462,8.064001,8.339693,8.960001,8.769642,7.7259493,6.9087186,6.3343596,6.5280004,6.6133337,6.2884107,5.8453336,6.1407185,6.311385,6.3967185,6.4656415,6.5903597,6.1341543,5.5171285,5.1167183,5.1265645,5.546667,5.408821,5.602462,6.23918,7.0859494,7.584821,8.03118,8.507077,8.851693,9.258667,10.282667,11.136001,12.320822,12.954257,12.914873,12.849232,11.474052,9.419488,8.162462,8.080411,8.448001,8.392206,8.562873,8.513641,8.119796,7.5946674,8.214975,8.3134365,7.722667,6.675693,5.802667,5.395693,4.857436,4.2371287,3.620103,3.1277952,2.8750772,2.7503593,2.7011285,2.7175386,2.8160002,2.681436,2.3794873,2.3302567,2.7602053,3.692308,3.8137438,3.5905645,3.4330258,3.4592824,3.5052311,3.69559,3.7185643,4.066462,4.5095387,4.086154,3.626667,2.9243078,2.5107694,2.5173335,2.6847181,2.8849232,2.6256413,2.3860514,2.284308,2.0644104,3.2623591,2.038154,1.529436,1.0994873,0.67938465,0.7778462,0.92225647,1.0469744,0.9878975,0.7450257,0.47261542,0.380718,0.37415388,0.47261542,0.5874872,0.508718,0.42994875,0.39712822,0.446359,0.5481026,0.6071795,0.5874872,0.56123084,0.52512825,0.4955898,0.49230772,0.6170257,0.69579494,0.7581539,0.8566154,1.0666667,1.8116925,1.6475899,1.2537436,1.0469744,1.214359,1.2242053,1.0929232,0.9419488,0.827077,0.761436,0.6432821,0.46933338,0.52512825,0.76800007,0.8205129,0.81066674,0.9616411,0.8598975,0.508718,0.318359,0.61374366,0.73517954,0.65312827,0.5021539,0.60061544,0.6826667,0.54482055,0.39712822,0.35446155,0.4004103,0.43323082,0.84348726,1.6114873,2.789744,4.519385,6.5444107,8.89436,10.463181,11.319796,12.704822,14.920206,17.184822,20.614565,25.028925,28.964106,30.112823,29.092104,28.025438,27.575796,26.945642,27.710361,27.585644,27.181952,27.00472,27.46749,25.655796,24.031181,22.032412,20.371695,21.051079,16.128002,14.621539,14.772514,15.602873,16.938667,17.857643,16.935387,16.06236,16.489027,18.802874,21.129848,22.806976,23.670156,24.421745,26.610874,28.580105,28.402874,28.639181,30.457438,33.631184,31.747284,31.140104,32.63672,36.47672,42.30236,46.57231,43.759594,39.683285,36.306053,31.744003,29.101952,31.215591,30.273643,25.16677,21.50072,33.046978,57.540928,77.177444,78.42462,52.017235,52.61785,52.9198,48.334774,41.38667,41.695183,48.003284,49.80185,49.14216,46.77252,42.09231,31.27795,23.378054,18.799591,16.292105,12.95754,10.689642,9.803488,9.964309,10.860309,12.209231,12.448821,13.318565,14.10954,13.449847,9.298052,7.574975,7.000616,6.875898,6.87918,7.059693,7.680001,8.480822,9.435898,10.266257,10.450052,6.5050263,4.450462,3.6430771,3.3280003,2.6683078,2.8225644,3.6036925,4.2830772,5.1265645,7.394462,8.845129,7.6767187,6.304821,5.865026,6.23918,7.1844106,9.271795,11.099898,12.130463,12.698257,16.823795,18.487797,16.390566,11.963078,9.380103,10.171078,10.427077,10.587898,10.765129,10.732308,11.670976,14.260514,16.987898,19.301744,21.632002,17.289848,15.468308,15.537232,16.144411,15.225437,16.278976,19.15077,21.008411,21.4679,22.610052,22.130873,17.703386,14.65436,13.755078,11.237744,11.664412,13.850258,14.831591,12.954257,7.8539495,3.9712822,3.9909747,4.6539493,4.59159,4.33559,2.934154,2.8521028,2.8553848,2.4451284,1.8642052,9.705027,12.048411,11.08677,11.398565,19.938463,24.697437,20.965746,14.329437,8.192,3.7710772,3.0851285,7.466667,10.9456415,10.305642,5.074052,4.3684106,2.4615386,2.2547693,3.3476925,2.03159,2.3204105,4.824616,4.900103,2.6354873,2.8750772,2.605949,2.4352822,2.0775387,1.4276924,0.57764107,2.3630772,5.2578464,7.27959,7.2369237,4.7458467,2.5632823,1.5130258,1.4539489,2.103795,3.0523078,3.626667,4.20759,5.287385,5.3694363,0.95835906,1.5097437,1.9856411,2.5665643,3.498667,5.1167183,4.630975,4.1714873,5.609026,12.435693,29.784618,13.745232,6.8693337,8.119796,15.143386,24.260925,21.589334,26.62072,27.585644,21.51713,14.260514,9.770667,4.5522056,1.910154,2.2088206,2.8488207,3.0096412,2.8127182,2.1202054,1.3883078,1.6804104,2.3630772,3.9253337,5.7632823,7.6996927,9.970873,8.595693,15.402668,13.755078,4.269949,4.84759,9.862565,15.172924,17.522873,15.560206,9.862565,11.434668,12.432411,10.870154,8.021334,8.448001,8.950154,6.875898,5.5171285,5.5565133,5.074052,3.2328207,2.553436,1.8609232,1.0404103,1.0568206,0.69579494,3.1737437,5.0674877,4.7917953,2.5895386,3.8301542,2.6486156,1.7493335,2.1497438,3.186872,4.06318,2.8356924,6.1013336,12.662155,13.522053,12.1928215,12.87877,11.664412,8.598975,7.686565,5.225026,4.2962055,3.3411283,2.2022567,2.1300514,4.2240005,4.8738465,4.0992823,2.5862565,1.6836925,1.467077,1.2471796,1.4408206,1.8576412,1.7033848,1.5819489,1.654154,1.5753847,1.276718,0.98133343,0.94523084,0.96492314,0.892718,0.69251287,0.44307697,0.5316923,0.7581539,1.0305642,1.2800001,1.4375386,1.1520001,1.1126155,0.9878975,0.7417436,0.6235898,0.7515898,0.9288206,0.8763078,0.60389745,0.42338464,0.574359,0.63343596,0.6071795,0.61374366,0.86317956,1.5195899,2.4155898,2.8488207,2.6912823,2.3926156,1.9790771,1.8543591,1.8609232,1.8018463,1.4539489,1.2307693,1.3062565,1.3915899,1.3751796,1.3259488,1.204513,0.73517954,0.44964105,0.571077,1.0010257,1.083077,1.024,0.8533334,0.65641034,0.5874872,0.60061544,0.64000005,0.7122052,0.79425645,0.8041026,0.9682052,1.024,1.0535386,1.0896411,1.083077,0.7253334,0.82379496,0.8598975,0.7122052,0.63343596,0.7056411,1.0338463,1.079795,0.827077,0.77456415,0.81066674,0.75487185,2.2449234,5.074052,7.200821,5.10359,2.7208207,3.623385,7.2664623,9.015796,2.9144619,3.9154875,6.0160003,6.550975,6.196513,2.8258464,1.5360001,1.3128207,1.3620514,1.0896411,0.97805136,0.99774367,0.9616411,0.8533334,0.827077,0.73517954,0.7187693,0.7187693,0.69907695,0.61374366,0.6301539,0.65641034,0.702359,0.764718,0.8336411,0.88287187,1.1388719,1.5360001,1.9003079,1.9364104,1.6672822,1.7723079,1.7526156,1.529436,1.4572309,1.394872,1.4539489,1.529436,1.6016412,1.7460514,2.03159,1.8576412,1.8510771,2.0939488,2.1202054,2.5665643,5.648411,8.402052,8.953437,6.518154,10.975181,15.8654375,13.748514,6.370462,4.6539493,2.809436,1.4375386,0.5316923,0.21333335,0.7187693,0.97805136,0.88943595,1.0272821,1.3718976,1.2800001,1.7591796,1.7165129,1.9954873,2.4024618,1.7165129,1.4506668,1.2898463,1.3686155,1.5885129,1.6278975,1.654154,1.5819489,1.6147693,1.6935385,1.4900514,1.2570257,1.2406155,1.214359,1.0929232,0.92553854,0.90912825,0.7089231,0.39712822,0.101743594,0.0,0.0,0.009846155,0.049230773,0.13128206,0.27241027,0.28882053,0.5021539,0.7384616,0.94523084,1.1946667,1.1257436,0.9747693,0.94523084,1.0666667,1.2077949,1.024,1.1027694,1.3095386,1.4408206,1.2274873,1.3850257,1.4342566,1.5885129,1.8937438,2.225231,2.6354873,3.2229745,3.9154875,4.565334,4.95918,4.9920006,5.3398976,5.602462,5.910975,6.954667,7.394462,7.1680007,6.738052,6.4065647,6.2916927,5.61559,5.5302567,6.363898,7.706257,8.411898,8.861539,9.055181,9.537642,10.180923,10.174359,10.55836,10.610872,10.469745,9.954462,8.549745,7.6635904,7.3714876,6.8594875,6.3376417,7.0367184,6.73477,5.661539,5.549949,6.7610264,8.28718,9.081436,8.487385,7.683283,7.4929237,8.3823595,8.306872,8.392206,8.172308,7.683283,7.4404106,6.9677954,6.885744,6.669129,6.2851286,6.189949,6.9710774,7.204103,6.961231,6.3967185,5.72718,4.969026,4.5587697,4.315898,4.210872,4.338872,4.414359,4.8344617,5.6943593,6.688821,7.1122055,7.0990777,7.2336416,7.6209235,8.077128,8.136206,7.890052,9.055181,10.325335,11.096616,11.480617,11.283693,9.478565,8.323282,8.349539,8.3823595,8.700719,8.930462,8.923898,8.621949,8.057437,7.8769236,7.2237954,6.3967185,5.7107697,5.477744,5.3169236,4.8607183,4.414359,4.027077,3.501949,3.186872,2.9965131,2.9604106,3.0030773,2.9243078,2.8816411,2.737231,2.937436,3.5052311,4.0369234,4.31918,4.1222568,3.7776413,3.5905645,3.826872,4.1058464,4.0992823,4.0041027,3.7710772,3.1015387,2.8225644,2.484513,2.4451284,2.809436,3.4133337,3.249231,2.681436,2.3696413,2.3729234,2.156308,0.5021539,0.7220513,1.024,1.1158975,0.9124103,0.5349744,0.5218462,0.77456415,0.8041026,0.55794877,0.4135385,0.33805132,0.32820517,0.34133336,0.31507695,0.16738462,0.26584616,0.4004103,0.49887183,0.58420515,0.7778462,0.72861546,0.6071795,0.5349744,0.5152821,0.44307697,0.42994875,0.41025645,0.4266667,0.4955898,0.58092314,0.67610264,0.6826667,0.6826667,0.7515898,0.94523084,0.8008206,0.6432821,0.5874872,0.61374366,0.56451285,0.56451285,0.574359,0.65969235,0.7975385,0.86974365,0.7220513,0.61374366,0.47261542,0.37743592,0.5481026,0.9517949,1.1520001,0.9353847,0.5021539,0.5021539,0.57764107,0.48574364,0.44307697,0.5218462,0.65641034,1.2176411,1.8609232,2.789744,4.2272825,6.422975,7.3649235,9.419488,11.021129,12.521027,16.219898,17.526155,20.233849,24.51036,29.72226,34.409027,36.630978,36.28636,35.305027,34.49108,33.539284,33.50318,31.954054,30.562464,29.630362,28.09108,24.441439,21.559797,20.25354,20.01395,19.012924,16.997746,13.7386675,13.653335,16.938667,19.561028,21.769848,19.157335,16.708925,17.02072,20.279797,22.06195,22.038977,21.769848,21.838772,21.851898,26.28267,26.555079,25.38995,25.64595,30.336002,29.469542,27.641438,26.755283,28.005745,31.875284,42.29908,44.950977,44.750774,42.962055,37.202053,29.741951,28.179695,26.90954,23.427284,18.326975,24.001642,45.38749,59.762875,55.620926,32.66954,34.0119,33.23077,27.670977,21.737028,26.886566,36.519386,39.906464,40.60226,39.187695,33.280003,24.759796,17.447386,13.938873,13.3251295,11.201642,10.210463,9.176616,8.487385,8.500513,9.537642,10.341744,12.905026,14.985847,14.424617,9.140513,6.918565,6.262154,6.5017443,7.240206,8.375795,8.352821,9.133949,9.852718,9.974154,9.278359,6.055385,3.9844105,3.259077,3.2656412,2.5928206,3.1671798,3.7415388,4.332308,5.3924108,7.7981544,8.260923,6.921847,6.2490263,6.741334,6.9120007,8.402052,10.456616,11.47077,11.71036,13.321847,14.713437,15.179488,13.574565,10.528821,8.454565,8.697436,9.77395,10.774975,11.0145645,10.026668,12.612924,18.376207,21.632002,20.397951,16.420103,15.465027,14.880821,15.051488,15.238565,13.564719,14.139078,17.742771,19.971283,19.767796,19.423182,18.386053,15.645539,13.505642,12.212514,9.980719,10.259693,11.346052,12.035283,11.004719,6.806975,3.7907696,4.0336413,4.9788723,5.654975,6.669129,4.240411,2.9636924,2.5665643,2.5961027,2.425436,6.8562055,13.072412,16.009848,16.66954,22.12431,20.903387,17.93641,16.8599,15.586463,6.2851286,5.1987696,7.3649235,8.94359,8.260923,5.7829747,6.0160003,3.3444104,2.802872,4.2174363,2.228513,3.0818465,3.9647183,3.623385,2.4484105,2.4713848,2.349949,2.4648206,2.2514873,1.5031796,0.380718,0.7122052,1.8740515,2.7766156,2.9144619,2.3663592,1.2176411,0.5021539,0.34789747,0.80738467,1.8313848,3.1967182,4.8049235,10.935796,15.360002,1.3128207,1.142154,1.5097437,3.18359,5.6418467,7.0957956,4.128821,2.5731285,2.0118976,4.9920006,17.030565,16.075489,9.67877,8.976411,15.228719,19.80718,26.312206,24.07713,17.447386,10.404103,6.547693,4.604718,2.4155898,2.5764105,4.4110775,3.9811285,7.4371285,7.5487185,5.346462,3.498667,6.3310776,5.4416413,4.706462,4.8705645,6.5280004,10.115283,9.93477,9.944616,9.941334,9.609847,8.4972315,9.43918,7.9261546,9.019077,11.815386,9.458873,7.9819493,7.430565,6.669129,5.408821,4.210872,4.772103,5.1232824,5.549949,5.5991797,4.073026,1.5458462,0.5940513,0.47261542,0.60389745,0.58092314,1.276718,2.7044106,4.900103,5.8978467,1.723077,3.9220517,3.564308,2.917744,2.6978464,2.0742567,3.3312824,2.858667,3.757949,5.979898,6.3343596,12.632616,9.472001,6.554257,7.821129,11.457642,8.224821,5.1987696,3.620103,3.373949,3.0227695,3.3378465,3.1245131,2.674872,2.356513,2.6256413,2.2219489,2.0217438,1.8871796,1.6049232,0.88615394,1.0568206,1.1815386,0.99774367,0.58092314,0.33476925,0.54482055,0.7417436,0.9911796,1.1027694,0.6268718,0.49230772,0.76800007,1.0633847,1.204513,1.2668719,1.3522053,1.2373334,1.0338463,0.8533334,0.79425645,1.0502565,1.2504616,1.2012309,0.8763078,0.4135385,0.42338464,0.4266667,0.45292312,0.49887183,0.5349744,0.54482055,0.9517949,1.6738462,2.2711797,1.9528207,2.2219489,2.5271797,2.4352822,1.8904617,1.2209232,1.2832822,1.4342566,1.591795,1.6804104,1.6311796,1.6443079,1.1454359,0.6071795,0.32820517,0.4266667,0.4397949,0.7450257,0.9156924,0.83035904,0.67282057,0.84348726,0.8041026,0.6629744,0.5481026,0.6104616,0.7450257,0.8795898,1.014154,1.1946667,1.5097437,1.1454359,0.9517949,0.82379496,0.7187693,0.67282057,0.5874872,0.7187693,0.7811283,0.67610264,0.51856416,0.54482055,0.78769237,1.5983591,2.6223593,2.793026,4.8672824,4.4438977,4.7655387,6.439385,7.4174366,5.290667,6.5444107,7.4732313,7.017026,6.7610264,6.892308,5.1954875,3.4560003,2.1989746,0.6859488,0.61374366,0.8041026,0.8730257,0.7417436,0.65641034,0.6432821,0.7318975,0.76800007,0.7220513,0.6859488,0.67282057,0.67282057,0.65312827,0.6629744,0.80738467,0.7122052,0.8041026,1.142154,1.5097437,1.4506668,1.3161026,1.6016412,1.7427694,1.5819489,1.3718976,1.3489232,1.4244103,1.5786668,1.6475899,1.3423591,1.7460514,1.6443079,1.5655385,1.7296412,2.0611284,4.197744,7.1647186,10.039796,12.327386,13.974976,14.293334,11.756309,9.888822,8.963283,5.9963083,5.47118,3.370667,1.3095386,0.19692309,0.24287182,0.65969235,0.6432821,1.0043077,1.595077,1.3259488,1.6311796,1.7001027,1.719795,1.7263591,1.6180514,1.6180514,1.4703591,1.270154,1.211077,1.6016412,2.3236926,2.0808206,1.7099489,1.5392822,1.404718,1.1224617,1.1913847,1.2570257,1.1684103,0.9616411,0.827077,0.54482055,0.26584616,0.072205134,0.0,0.0,0.01969231,0.06564103,0.15097436,0.25928208,0.44307697,0.6892308,0.84348726,0.9485129,1.2668719,1.1684103,1.0338463,1.0272821,1.1355898,1.1585642,1.0633847,1.339077,1.595077,1.6180514,1.3718976,1.3850257,1.3981539,1.4112822,1.5163078,1.9068719,2.6387694,3.0884104,3.4724104,3.8498464,4.1058464,4.4110775,4.6605134,4.9099493,5.3431797,6.2720003,6.564103,6.2720003,5.6418467,5.1200004,5.3398976,5.4153852,5.861744,6.449231,7.056411,7.6898465,8.582564,9.380103,9.938052,10.016821,9.3078985,9.613129,10.420513,10.532104,9.636104,8.329846,7.512616,6.806975,6.688821,7.02359,7.0498466,6.416411,5.733744,5.8880005,6.8233852,7.568411,7.77518,7.4797955,7.0531287,7.0400004,8.162462,8.1755905,8.214975,8.001641,7.5388722,7.1122055,7.282872,7.1876926,7.059693,7.1515903,7.752206,7.6668725,7.4896417,7.3550773,7.0957956,6.23918,4.9362054,4.378257,4.201026,4.069744,3.692308,4.4012313,5.1265645,5.792821,6.3310776,6.698667,6.186667,6.7183595,7.6274877,8.356103,8.454565,8.050873,8.260923,8.211693,8.086975,9.124104,9.357129,8.516924,8.077128,8.467693,9.078155,8.956718,8.907488,8.6580515,8.165744,7.6307697,6.9809237,6.226052,5.5105643,5.024821,4.9887185,4.71959,4.699898,4.6867695,4.5128207,4.073026,3.6332312,3.6529233,3.623385,3.5840003,4.1189747,3.570872,3.2032824,3.373949,3.879385,3.95159,5.3070774,5.481026,4.6933336,3.7284105,3.9351797,3.5216413,3.2164104,3.0654361,2.9407182,2.5632823,2.3926156,2.5435898,2.7667694,2.9735386,3.2032824,2.8750772,2.3991797,2.2022567,2.3269746,2.425436,0.2100513,0.44964105,0.78769237,0.9616411,0.88287187,0.6301539,0.46276927,0.4660513,0.508718,0.52512825,0.49887183,0.24943592,0.15097436,0.128,0.128,0.118153855,0.21661541,0.2986667,0.37415388,0.47261542,0.6695385,0.6695385,0.5513847,0.44964105,0.39712822,0.3446154,0.29210258,0.26912823,0.26912823,0.3052308,0.41025645,0.41025645,0.46276927,0.58092314,0.65641034,0.48246157,0.45292312,0.47917953,0.49887183,0.5021539,0.5513847,0.4660513,0.508718,0.5874872,0.6498462,0.7220513,0.5874872,0.56123084,0.6235898,0.73517954,0.8172308,1.3292309,1.2635899,0.892718,0.5415385,0.5874872,0.4955898,0.4955898,0.5513847,0.69579494,1.0338463,1.595077,2.7602053,3.9745643,5.182359,6.803693,8.621949,10.43036,12.461949,15.425642,20.49313,21.671387,24.54318,28.232206,32.74831,38.997337,42.243286,44.708107,45.09867,43.62831,42.023388,39.758774,37.398975,34.766773,32.177235,30.421335,27.477335,24.549746,21.746874,18.67159,14.447591,15.107284,16.384,20.128822,25.491693,28.934566,32.318363,29.673027,25.580309,23.072823,23.634052,25.311182,26.666668,27.214771,26.643694,24.82872,28.28472,31.954054,33.86749,33.729645,32.90913,29.525335,25.53436,24.44472,28.832823,40.359386,58.164516,66.88821,64.96493,54.672413,42.144825,36.637543,34.589542,31.711182,26.039797,17.959387,22.951385,39.486362,46.509953,36.97231,17.851078,17.378464,18.323694,17.58195,16.856617,22.662565,24.139488,23.72595,23.995079,23.96554,19.072002,15.189335,13.334975,13.472821,13.686155,10.174359,8.01477,6.941539,6.8004107,7.460103,8.828718,10.308924,11.503591,12.304411,11.841642,8.480822,6.816821,6.445949,6.5280004,6.6461544,6.813539,7.6307697,7.9261546,7.683283,7.2205133,7.1909747,6.75118,5.927385,5.5269747,5.330052,4.082872,3.436308,3.8662567,4.8147697,5.8912826,6.882462,7.3452315,8.421744,8.976411,8.4512825,6.875898,7.9852314,9.783795,10.420513,10.020103,10.683078,13.10195,13.459693,11.670976,8.802463,7.0498466,7.9097443,10.354873,11.96636,12.09436,11.85477,16.485744,20.086155,20.850874,18.960411,16.600616,14.555899,13.820719,14.007796,14.093129,12.42913,12.750771,15.66195,17.444103,17.345642,17.56882,16.971489,14.244103,12.140308,11.08677,9.186462,9.80677,10.072617,10.683078,10.512411,6.5870776,3.698872,4.57518,5.684513,6.298257,8.474257,6.114462,3.8596926,2.9801028,3.4330258,3.8662567,9.760821,12.698257,14.116103,16.20349,21.904411,18.710976,18.113642,23.210669,28.081232,17.785437,9.668923,9.252103,9.02236,6.8463597,5.979898,6.3573337,4.0533338,3.259077,3.945026,1.8379488,2.2022567,2.993231,3.1343591,2.6683078,2.7536411,2.6223593,2.609231,2.3269746,1.5819489,0.380718,0.25271797,0.47917953,0.6859488,1.4211283,4.1714873,9.399796,5.1364107,1.6443079,1.9462565,1.8182565,2.9111798,3.2918978,12.675283,22.278566,4.841026,7.384616,5.421949,4.388103,5.858462,7.5454364,6.954667,4.8640003,7.7390776,13.61395,12.097642,13.1872835,12.048411,11.513436,13.679591,19.928617,22.997335,19.482258,15.442053,13.02318,10.463181,8.533334,6.245744,4.571898,4.2436924,5.7403083,10.774975,7.6603084,6.701949,9.271795,7.7981544,6.8955903,7.381334,7.6110773,7.574975,8.907488,11.546257,11.697231,14.336001,18.051283,15.064616,11.444513,7.026872,7.171283,10.827488,10.522257,9.268514,9.147078,7.958975,5.602462,4.066462,2.9768207,2.6420515,2.7208207,2.9210258,3.0358977,3.6529233,3.4592824,3.0916924,2.5731285,1.2865642,1.4375386,2.2153847,3.7054362,4.6244106,2.3335385,3.0752823,2.553436,2.4352822,2.6486156,1.3915899,2.9407182,2.9538465,3.3017437,5.4449234,10.410667,8.887795,7.2303596,6.8955903,7.571693,7.1876926,6.99077,5.4843082,4.414359,4.023795,3.0949745,2.4746668,2.3040001,2.4549747,2.6683078,2.5764105,1.5885129,1.0043077,0.761436,0.69251287,0.51856416,0.62030774,0.69251287,0.60389745,0.42994875,0.45620516,0.6268718,0.9156924,1.1881026,1.2274873,0.77128214,0.5973334,0.65312827,0.81066674,1.0371283,1.401436,1.2504616,0.8205129,0.49887183,0.41025645,0.4266667,0.4397949,0.5152821,0.6268718,0.77456415,0.9747693,0.7318975,0.4955898,0.39712822,0.48574364,0.7187693,0.7384616,0.9714873,1.2832822,1.595077,1.8904617,2.0053334,2.540308,2.4352822,1.7591796,1.719795,2.0250258,1.7788719,1.5360001,1.4375386,1.1946667,1.3423591,1.2209232,0.9616411,0.69579494,0.5481026,0.43323082,0.6859488,1.0075898,1.204513,1.1848207,1.2176411,1.079795,0.8008206,0.53825647,0.56123084,0.5677949,0.65641034,0.761436,0.9353847,1.339077,1.3062565,1.1224617,0.955077,0.9353847,1.1585642,0.90912825,0.892718,0.9878975,1.0404103,0.8730257,0.4004103,0.48246157,0.892718,1.3784616,1.657436,2.609231,4.1452312,5.3924108,5.8223596,5.2545643,3.620103,6.262154,8.470975,7.6734366,3.4527183,6.875898,9.035488,9.051898,6.4689236,1.2373334,0.41025645,0.2986667,0.48574364,0.67938465,0.67938465,0.48246157,0.508718,0.6104616,0.67938465,0.6629744,0.6498462,0.69907695,0.69907695,0.64000005,0.60061544,0.60061544,0.6695385,0.9517949,1.2964103,1.2537436,1.1979488,1.1684103,1.142154,1.1355898,1.2012309,1.2471796,1.2307693,1.3686155,1.5721027,1.4539489,1.3587693,1.3522053,1.3423591,1.4703591,2.1333334,4.7294364,6.7872825,9.252103,11.762873,12.658873,11.559385,12.737642,13.682873,12.2847185,6.8397956,4.6244106,6.8397956,5.8092313,1.2209232,0.14769232,0.56123084,0.53825647,0.7318975,1.2471796,1.6311796,1.6640002,1.5753847,1.4802053,1.4441026,1.4703591,1.2964103,1.1191796,0.99774367,1.0108719,1.2832822,1.6344616,1.6016412,1.529436,1.5327181,1.4769232,1.204513,1.3357949,1.3883078,1.2209232,1.0338463,0.8598975,0.4594872,0.15097436,0.032820515,0.0,0.009846155,0.029538464,0.07548718,0.15097436,0.25928208,0.5021539,0.65312827,0.79097444,0.9714873,1.2307693,1.1618463,1.1158975,1.0929232,1.1027694,1.148718,1.214359,1.3883078,1.4998976,1.467077,1.3128207,1.2865642,1.3029745,1.401436,1.6114873,1.9429746,2.7142565,3.0654361,3.2787695,3.4789746,3.629949,4.07959,4.3749747,4.850872,5.477744,5.868308,5.720616,5.5236926,5.2512827,5.0477953,5.218462,5.1364107,5.2676926,5.668103,6.265436,6.8594875,8.201847,8.651488,8.73354,8.753231,8.809027,9.268514,9.199591,8.73354,8.136206,7.8080006,7.653744,7.131898,6.5378466,6.091488,5.937231,5.402257,5.4547696,5.8420515,6.363898,6.872616,6.5805135,6.6822567,7.076103,7.5520005,7.7981544,7.9163084,8.201847,8.0377445,7.4797955,7.256616,7.076103,6.5805135,6.3277955,6.5739493,7.250052,7.273026,6.7774363,6.2162056,5.8945646,5.9963083,5.648411,5.579488,5.1987696,4.598154,4.571898,5.024821,5.3431797,5.6320004,5.930667,6.1997952,6.183385,6.619898,7.1220517,7.4929237,7.6964107,7.509334,7.781744,7.762052,7.427283,7.4896417,8.01477,7.8473854,7.8637953,8.411898,9.334154,9.242257,8.907488,8.2904625,7.5881033,7.2270775,6.38359,5.4908724,4.9526157,4.9427695,5.405539,4.9394875,4.775385,4.667077,4.525949,4.4274874,4.309334,4.466872,4.493129,4.309334,4.1813335,3.757949,3.5774362,3.623385,3.8006158,3.95159,4.5456414,5.408821,5.3431797,4.3552823,3.6430771,3.318154,3.259077,3.190154,3.045744,2.989949,2.674872,2.477949,2.4352822,2.5632823,2.861949,2.5928206,2.4582565,2.5173335,2.6617439,2.6223593,0.108307704,0.24287182,0.67282057,1.083077,1.1881026,0.7187693,0.37415388,0.2297436,0.2100513,0.24287182,0.23630771,0.118153855,0.068923086,0.06235898,0.08205129,0.14441027,0.16082053,0.2100513,0.26256412,0.31507695,0.38400003,0.39056414,0.34789747,0.318359,0.30851284,0.26584616,0.23302566,0.22646156,0.2231795,0.2231795,0.27569234,0.37415388,0.4397949,0.508718,0.52512825,0.32820517,0.2986667,0.37743592,0.4135385,0.4004103,0.45620516,0.40697438,0.58092314,0.7056411,0.71548724,0.7515898,0.65312827,0.79425645,0.98133343,1.1454359,1.3161026,1.3259488,1.2373334,0.98133343,0.7089231,0.79425645,0.761436,0.69251287,0.761436,1.0404103,1.5031796,2.0217438,2.9768207,4.096,5.549949,7.9491286,10.65354,13.5778475,16.003283,18.425438,22.55754,24.930464,27.369028,30.608412,35.554462,43.29354,48.28554,50.58626,50.81272,50.107082,50.1399,45.72226,42.771694,40.52677,38.705235,37.504,30.720003,25.124104,21.238155,18.950565,17.526155,17.273438,18.553438,24.04431,32.902565,40.756516,46.093132,43.3559,37.254566,31.753849,30.066874,32.945232,34.304,33.870773,32.20677,30.680618,32.771286,35.94503,37.894566,37.32349,33.939693,30.201439,29.56472,34.36308,46.165337,65.78872,82.62237,84.55221,73.49498,54.77744,37.136414,32.551388,30.424618,28.064823,24.497232,20.466873,25.061745,33.57867,33.368618,22.505028,9.770667,9.741129,11.808822,14.27036,16.502155,18.934155,17.93313,16.73518,15.780104,14.690463,12.278154,11.497026,12.685129,13.551591,12.563693,8.946873,6.8955903,6.301539,7.177847,8.94359,10.417232,11.172104,10.978462,10.988309,10.758565,8.241231,5.9634876,5.3431797,5.428513,5.684513,5.9930263,6.961231,6.619898,6.2555904,6.439385,7.0334363,7.026872,6.3606157,5.930667,5.730462,4.8672824,3.9286156,4.194462,4.900103,5.5302567,5.8289237,6.738052,8.214975,8.848411,8.362667,7.6176414,8.562873,9.613129,9.754257,9.117539,8.973129,11.602052,11.861334,10.069334,7.4929237,6.3310776,7.4404106,10.384411,12.576821,13.512206,14.759386,15.750566,17.808413,18.274464,16.57436,14.204719,12.609642,12.107488,12.107488,12.032001,11.293539,12.189539,15.684924,16.485744,14.372104,14.204719,15.136822,12.642463,10.597744,10.085744,9.409642,9.019077,9.058462,9.734565,9.931488,7.2172313,4.1780515,4.7425647,5.8781543,6.5017443,7.4896417,5.6943593,4.1058464,3.6890259,4.2830772,4.6211286,10.932513,12.544001,13.843694,16.439796,19.167181,16.118155,19.072002,24.635078,27.250874,19.222977,13.3251295,11.720206,8.986258,5.0871797,5.3760004,5.405539,3.9614363,3.639795,4.0041027,1.6114873,1.8904617,2.612513,2.858667,2.737231,3.3542566,2.9997952,2.793026,2.3827693,1.6246156,0.56451285,0.23302566,0.20020515,0.18707694,0.49887183,2.0250258,4.650667,2.8553848,1.591795,2.103795,1.9068719,2.7798977,3.1606157,9.856001,16.922258,5.658257,9.130668,12.744206,12.737642,9.5606165,7.8802056,10.9686165,10.325335,14.667488,21.251284,15.852309,18.192411,17.578669,18.934155,21.192207,17.302977,16.216616,13.220103,10.706052,9.711591,9.924924,8.933744,12.895181,12.156719,6.7971287,6.629744,7.387898,4.969026,6.1407185,9.67877,6.3868723,7.4240007,10.827488,12.422565,10.94236,8.021334,11.175385,10.79795,12.514462,15.681643,13.384206,13.193847,11.365745,9.833026,10.226872,13.892924,9.334154,6.422975,4.5029745,3.367385,3.259077,2.0053334,1.654154,1.8871796,2.1891284,1.8346668,3.1277952,3.2525132,2.917744,2.359795,1.3456411,1.8707694,3.7907696,5.0018463,4.667077,3.2295387,2.3762052,1.7887181,2.3401027,3.1770258,1.7329233,2.2646155,2.3105643,3.639795,5.924103,6.7249236,5.477744,4.6769233,4.7294364,5.10359,4.332308,4.9920006,5.421949,4.886975,3.5183592,2.3269746,1.595077,1.6869745,2.048,2.2613335,2.041436,1.2209232,0.69251287,0.41682056,0.32820517,0.33476925,0.34133336,0.3511795,0.3052308,0.23958977,0.27897438,0.5316923,1.0732309,1.4473847,1.394872,0.86317956,0.75487185,0.7384616,0.7778462,0.9353847,1.3981539,1.0502565,0.65641034,0.446359,0.43323082,0.39056414,0.28225642,0.3052308,0.4397949,0.63343596,0.79425645,0.7089231,0.53825647,0.43323082,0.47589746,0.69907695,0.7318975,0.85005134,0.9485129,1.0765129,1.4572309,1.6607181,2.2121027,2.1300514,1.5885129,1.8904617,1.8116925,1.5983591,1.4080001,1.1946667,0.7253334,1.086359,0.90912825,0.67938465,0.571077,0.45292312,0.45292312,0.4955898,0.6465641,0.892718,1.1388719,1.3587693,1.3095386,1.1027694,0.86646163,0.7318975,0.57764107,0.64000005,0.77456415,0.94523084,1.2340513,1.404718,1.2504616,1.1126155,1.1684103,1.4572309,1.2635899,1.0994873,1.0272821,1.014154,0.92553854,0.4004103,0.35774362,0.58092314,0.8467693,0.9353847,1.6640002,3.117949,4.8640003,6.616616,8.2215395,5.366154,6.2490263,8.149334,8.3134365,3.9417439,4.7491283,7.020308,7.830975,6.0356927,2.281026,1.0601027,0.4266667,0.25928208,0.37743592,0.512,0.42338464,0.4004103,0.42994875,0.48574364,0.54482055,0.5481026,0.61374366,0.6465641,0.6071795,0.5218462,0.52512825,0.58420515,0.7811283,1.0502565,1.204513,1.1323078,1.1191796,1.0502565,0.9682052,1.0601027,1.0994873,1.0962052,1.1913847,1.3357949,1.3062565,1.2931283,1.3456411,1.3029745,1.2800001,1.6672822,3.5577438,5.5893335,7.6110773,10.217027,14.7561035,11.552821,10.679795,12.097642,12.832822,6.994052,4.532513,6.121026,5.4941545,1.9003079,0.11158975,0.30851284,0.36102566,0.48902568,0.827077,1.4342566,1.3456411,1.404718,1.394872,1.3062565,1.3259488,1.148718,0.94523084,0.83035904,0.8730257,1.086359,1.276718,1.404718,1.4145643,1.3259488,1.2406155,1.2406155,1.2438976,1.1651284,1.017436,0.90584624,0.7450257,0.37415388,0.101743594,0.016410258,0.0,0.0032820515,0.029538464,0.08861539,0.17394873,0.27897438,0.48902568,0.574359,0.6859488,0.86317956,1.020718,1.0404103,1.1126155,1.1060513,1.0272821,1.017436,1.1618463,1.270154,1.3718976,1.4309745,1.3259488,1.3095386,1.394872,1.5261539,1.6935385,1.9167181,2.3958976,2.8882053,3.1573336,3.2196925,3.3280003,3.6824617,4.3684106,5.0018463,5.408821,5.622154,5.349744,5.139693,4.850872,4.6539493,5.031385,5.0576415,5.1331286,5.47118,6.0291286,6.5444107,7.2205133,6.931693,6.6461544,6.9021544,7.821129,8.418462,8.372514,7.962257,7.450257,7.1154876,7.1647186,6.5870776,5.7796926,5.093744,4.8082056,4.896821,5.536821,5.868308,5.8125134,6.0947695,6.0980515,6.678975,7.1909747,7.3419495,7.2205133,7.6242056,8.080411,8.297027,8.123077,7.5487185,6.9087186,6.3606157,6.304821,6.6395903,6.741334,7.0465646,6.9776416,6.5017443,6.0849237,6.675693,6.5378466,6.3540516,5.8847184,5.2545643,4.965744,5.100308,5.1922054,5.4383593,5.917539,6.5870776,6.5706673,6.8627696,7.0990777,7.1876926,7.3321033,7.141744,7.2927184,7.506052,7.5520005,7.2369237,7.5913854,7.5454364,7.3747697,7.4404106,8.198565,8.408616,8.01477,7.4436927,6.8955903,6.3573337,5.284103,4.5456414,4.4340515,4.785231,4.969026,4.916513,4.650667,4.3716927,4.2896414,4.6080003,4.850872,5.1954875,5.211898,4.9099493,4.7261543,4.1911798,4.096,4.263385,4.532513,4.775385,4.4964104,4.59159,4.2929235,3.5872824,3.239385,3.4330258,3.387077,3.1606157,3.0030773,3.370667,3.0687182,2.7142565,2.7109745,3.0654361,3.3903592,3.0162053,2.7044106,2.5042052,2.3729234,2.176,0.07876924,0.12143591,0.5284103,0.9714873,1.1684103,0.892718,0.48574364,0.190359,0.052512825,0.03938462,0.026256412,0.04594872,0.03938462,0.036102567,0.055794876,0.11158975,0.0951795,0.15425642,0.190359,0.17394873,0.15097436,0.15097436,0.18707694,0.23958977,0.27897438,0.24615386,0.22646156,0.22646156,0.2100513,0.17723078,0.16410258,0.27897438,0.318359,0.32164106,0.2986667,0.22646156,0.21989745,0.27569234,0.29538465,0.28225642,0.33476925,0.32820517,0.5677949,0.7581539,0.81394875,0.8533334,1.1191796,1.3915899,1.8182565,2.1136413,1.5655385,1.3423591,1.2471796,1.086359,0.94523084,1.1848207,1.4211283,1.4933335,1.5360001,1.6968206,2.1267693,2.4385643,3.2918978,4.4438977,6.3967185,10.377847,13.748514,18.86195,22.849644,24.874668,26.154669,27.152412,29.4039,33.637745,40.277336,49.440823,53.03467,52.785236,52.450466,53.251286,53.868313,49.887184,46.742977,46.096413,46.831593,45.07898,37.041233,29.699284,24.98954,23.04,22.199797,21.290668,25.898668,39.78831,60.05826,77.16103,68.818054,54.659286,42.013542,35.19344,35.501953,36.59159,35.892517,34.6519,33.772312,33.808414,34.192413,34.48123,34.258053,32.935387,29.751797,29.32513,33.332516,41.48185,53.474464,68.98872,73.98401,69.29395,57.360416,41.94462,28.110771,25.819899,23.194258,22.209642,23.236925,25.03877,27.37231,33.00103,30.916925,20.073027,9.3768215,8.871386,11.175385,14.578873,17.769028,19.830154,18.816002,16.452925,13.377642,10.683078,9.9282055,9.642668,10.620719,10.732308,9.291488,7.0432825,7.276308,7.276308,8.224821,10.000411,11.18195,10.643693,9.682052,9.130668,8.825437,7.6143594,7.174565,5.6976414,5.159385,5.7435904,5.8486156,6.51159,6.4295387,6.9120007,7.972103,8.303591,7.4240007,6.5706673,6.117744,5.9634876,5.533539,4.8147697,4.7622566,5.169231,5.7829747,6.311385,7.79159,8.805744,8.802463,8.162462,8.198565,8.664616,9.16677,8.897642,7.9885135,7.512616,9.665642,9.849437,8.333129,6.2851286,5.7829747,7.3616414,10.860309,13.968411,15.67836,16.328207,13.522053,14.496821,15.067899,13.781334,11.907283,11.030975,10.725744,10.627283,10.640411,10.9226675,12.035283,15.081027,15.025232,12.041847,11.487181,12.921437,10.916103,9.140513,8.871386,8.999385,7.9097443,7.9491286,8.759795,9.324308,7.968821,4.644103,4.71959,5.874872,6.5378466,5.865026,4.57518,3.9680004,4.2174363,4.84759,4.7556925,8.644924,10.624001,12.507898,14.444309,14.913642,13.676309,17.98236,22.459078,23.151592,17.496616,13.764924,11.559385,7.8802056,3.8367183,4.6145644,3.892513,3.1540515,3.4560003,3.9318976,1.8116925,1.9035898,2.9111798,3.245949,2.9702566,3.82359,2.9965131,2.7864618,2.412308,1.6377437,0.7778462,0.40369233,0.31507695,0.25271797,0.7778462,3.255795,3.7874875,5.093744,5.986462,5.277539,1.785436,2.4910772,3.5347695,9.783795,17.283283,13.262771,10.240001,14.240822,16.787693,14.49354,9.074872,11.067078,10.305642,13.348104,19.14749,19.058874,20.86072,21.087181,23.026873,24.034464,15.540514,14.024206,11.72677,10.266257,10.243283,11.241027,10.689642,14.775796,14.119386,8.320001,5.943795,9.380103,5.3792825,4.204308,6.8988724,5.277539,8.185436,12.76718,17.77559,19.058874,9.563898,9.55077,8.12636,8.425026,10.029949,8.973129,12.859077,13.364513,10.666668,7.7390776,10.358154,6.1078978,3.0424619,1.5688206,1.5786668,2.477949,1.8642052,3.0916924,3.511795,2.9046156,3.4822567,3.2853336,2.3269746,1.6311796,1.4834872,1.4080001,2.097231,3.761231,4.3290257,3.5840003,3.186872,1.8806155,1.7920002,2.7831798,3.6693337,2.2022567,2.1891284,2.0118976,4.2601027,6.8463597,3.006359,4.1780515,3.6562054,3.1081028,3.1934361,3.5577438,3.508513,3.9942567,3.5938463,2.2580514,1.3062565,1.0535386,1.3456411,1.7362052,1.9265642,1.7788719,1.3784616,0.8041026,0.39056414,0.24287182,0.21989745,0.17066668,0.15097436,0.13784617,0.14112821,0.17394873,0.42338464,0.9419488,1.3522053,1.4244103,1.0535386,0.9616411,0.96492314,0.9878975,1.0633847,1.3292309,0.827077,0.56123084,0.5152821,0.57764107,0.54482055,0.41682056,0.44964105,0.508718,0.53825647,0.54482055,0.64000005,0.6170257,0.60389745,0.6465641,0.7220513,0.636718,0.67610264,0.73517954,0.8369231,1.1257436,1.4834872,1.9922053,2.0873847,1.8543591,2.0151796,1.6836925,1.463795,1.404718,1.2800001,0.5874872,0.827077,0.69907695,0.636718,0.6629744,0.40369233,0.39384618,0.29538465,0.2986667,0.47917953,0.8041026,1.0404103,1.1257436,1.148718,1.1158975,0.95835906,0.6662565,0.65969235,0.761436,0.90584624,1.1290257,1.3226668,1.2176411,1.1618463,1.2504616,1.3259488,1.2537436,0.9911796,0.7811283,0.7220513,0.77128214,0.39384618,0.3052308,0.40369233,0.55794877,0.5973334,1.4802053,2.162872,3.6529233,6.413129,10.35159,8.073847,6.3212314,6.4295387,7.145026,4.6276927,3.1409233,4.9985647,5.832206,4.4800005,2.9768207,2.0808206,1.1027694,0.39712822,0.12143591,0.256,0.3117949,0.2986667,0.28225642,0.30194873,0.35774362,0.4266667,0.47917953,0.5152821,0.52512825,0.508718,0.5021539,0.56123084,0.69251287,0.892718,1.1520001,1.1224617,1.2832822,1.2406155,1.0108719,0.99774367,0.94523084,0.98133343,1.1060513,1.2077949,1.079795,1.2274873,1.3128207,1.2438976,1.1684103,1.4769232,2.5173335,4.9985647,6.8955903,8.953437,14.6871805,12.865642,10.013539,10.643693,12.396309,6.042257,4.1583595,5.3760004,5.149539,2.5206156,0.118153855,0.128,0.256,0.3446154,0.48246157,1.0075898,1.0075898,1.1913847,1.2406155,1.1060513,1.0010257,1.0732309,0.9288206,0.79425645,0.7975385,0.93866676,1.1881026,1.3489232,1.2570257,1.0043077,0.9517949,1.1684103,1.0962052,0.98461545,0.90584624,0.77128214,0.5415385,0.26256412,0.072205134,0.006564103,0.0,0.0,0.02297436,0.108307704,0.2297436,0.30194873,0.48574364,0.5973334,0.7056411,0.81066674,0.8533334,0.9288206,1.086359,1.0962052,0.9517949,0.892718,1.083077,1.1651284,1.2570257,1.3620514,1.3850257,1.4342566,1.5195899,1.6246156,1.719795,1.7690258,2.0053334,2.5993848,2.9965131,3.0982566,3.2787695,3.4592824,4.132103,4.7228723,5.07077,5.4186673,5.1200004,4.844308,4.460308,4.1747694,4.5128207,4.529231,4.6834874,4.9821544,5.405539,5.901129,5.8945646,5.5171285,5.3924108,5.8880005,7.1122055,7.4863596,7.6734366,7.748924,7.653744,7.2205133,6.941539,6.2884107,5.661539,5.1659493,4.6080003,5.024821,5.7632823,5.9963083,5.7632823,5.979898,6.0750775,6.521436,6.678975,6.485334,6.4754877,7.1581545,7.7456417,8.2215395,8.3593855,7.7325134,7.056411,6.7840004,6.954667,7.2631803,7.076103,7.1876926,7.1909747,6.7577443,6.3179493,7.0793853,7.174565,6.8299494,6.3376417,5.865026,5.477744,5.425231,5.5236926,5.9634876,6.747898,7.683283,7.3714876,7.4174366,7.4929237,7.466667,7.394462,7.276308,7.256616,7.4929237,7.8112826,7.706257,7.5388722,7.433847,7.1187696,6.8529234,7.4075904,7.634052,7.322257,6.6560006,5.8256416,5.037949,4.4045134,4.010667,4.059898,4.3716927,4.394667,4.7589746,4.6605134,4.4734364,4.4012313,4.4734364,4.9394875,5.431795,5.6254363,5.4514875,5.0871797,4.4767184,4.4734364,4.9296412,5.431795,5.3202057,4.4734364,3.9712822,3.4822567,3.0293336,2.9604106,3.3247182,3.4592824,3.43959,3.4297438,3.7021542,3.4100516,2.8980515,2.7798977,3.121231,3.4527183,3.0391798,2.5600002,2.225231,2.041436,1.8149745,0.14441027,0.101743594,0.35774362,0.6104616,0.79097444,1.0732309,0.7581539,0.3249231,0.068923086,0.026256412,0.0032820515,0.04266667,0.029538464,0.016410258,0.016410258,0.026256412,0.036102567,0.14112821,0.16082053,0.08205129,0.06235898,0.08205129,0.14441027,0.26584616,0.4004103,0.4266667,0.41682056,0.37415388,0.2986667,0.20676924,0.13456412,0.13456412,0.14112821,0.12143591,0.098461546,0.14441027,0.19692309,0.2100513,0.190359,0.17723078,0.20676924,0.23302566,0.446359,0.67282057,0.8402052,0.9714873,1.6869745,2.1924105,2.92759,3.2918978,1.6246156,1.5392822,1.4211283,1.3161026,1.3522053,1.7394873,2.2121027,2.5238976,2.6256413,2.7109745,3.2098465,3.5774362,4.8607183,6.419693,8.835282,13.922462,17.670565,23.998362,29.029745,30.880823,29.663181,28.294567,31.360003,37.684517,46.004517,54.97436,55.70626,54.39016,55.83426,59.441235,59.20493,57.89539,55.41744,56.211697,58.752003,55.555286,48.873028,40.356106,34.021748,30.605131,27.569233,29.525335,42.847183,68.92308,99.551186,116.95262,83.74811,54.3278,36.17149,31.104002,35.285336,33.05354,30.106258,29.174156,30.565746,32.15426,31.678362,29.505644,26.98831,24.756516,22.734772,27.19836,33.61149,39.348515,42.87672,43.782566,35.5479,30.660925,27.848207,25.662361,22.482054,23.049849,20.43077,21.231592,25.882257,28.599796,28.484924,35.396927,34.69785,23.913027,12.724514,12.022155,14.057027,16.548103,18.921026,22.33108,21.408823,18.034874,13.840411,10.515693,9.813334,8.086975,6.882462,6.11118,5.664821,5.425231,8.320001,8.5891285,8.802463,9.714872,10.289231,8.809027,7.706257,6.6461544,5.976616,6.7249236,9.344001,7.2172313,5.9930263,6.8332314,6.413129,7.1876926,8.03118,9.268514,10.331899,9.750975,7.893334,7.0990777,6.9152827,6.8430777,6.36718,6.2523084,6.055385,6.6034875,7.8670774,8.979693,10.384411,10.561642,9.668923,8.43159,8.129642,8.0377445,8.375795,7.9852314,6.9152827,6.4065647,7.6077952,7.6996927,6.688821,5.421949,5.586052,7.906462,12.084514,16.022976,17.831387,15.812924,12.212514,12.150155,12.117334,11.08677,10.528821,10.089026,9.892103,9.931488,10.256411,10.9456415,11.792411,13.2562065,12.868924,10.860309,10.154668,10.617436,9.225847,8.054154,7.8539495,8.064001,6.7938466,6.8332314,7.722667,8.556309,7.9786673,4.8640003,4.7261543,5.786257,6.3967185,5.041231,3.820308,3.5478978,4.059898,4.6933336,4.2962055,4.5587697,7.177847,9.222565,9.90195,10.568206,11.175385,16.141129,19.876104,19.652925,15.629129,11.076924,8.598975,5.8453336,3.2328207,3.9351797,3.0851285,2.6190772,3.121231,3.8038976,2.4976413,2.0841026,3.4297438,4.0041027,3.5774362,4.197744,2.7700515,2.5698464,2.3368206,1.6475899,0.92553854,0.51856416,0.42338464,0.380718,1.6180514,6.8562055,8.001641,10.095591,11.296822,9.452309,2.100513,3.2722054,7.1483083,16.042667,25.491693,24.247797,13.387488,11.35918,14.424617,17.171694,12.527591,8.677744,5.549949,5.904411,10.230155,16.758156,22.04554,21.415386,19.790771,19.2,18.796309,16.292105,14.093129,14.391796,15.914668,13.912617,12.586668,11.096616,9.731283,8.067283,4.9526157,14.280207,8.195283,2.9997952,3.892513,4.955898,8.080411,11.884309,19.452719,24.730259,12.530872,7.4108725,4.906667,5.0642056,6.304821,5.428513,10.013539,11.073642,8.326565,3.7809234,1.7099489,1.3587693,1.2242053,1.2209232,1.4244103,2.0906668,2.3991797,5.0674877,5.287385,3.5741541,5.76,3.8662567,1.6246156,0.574359,0.94523084,1.657436,2.0250258,2.041436,1.7690258,1.5721027,2.1398976,1.7033848,2.6223593,3.6168208,3.8400004,2.8816411,2.8258464,2.4418464,4.578462,6.987488,2.3269746,4.1452312,3.6660516,2.8192823,2.7831798,3.9975388,2.9144619,1.9462565,1.3522053,1.0469744,0.5874872,0.90256417,1.1946667,1.4834872,1.7033848,1.7033848,1.6246156,0.9288206,0.38400003,0.2231795,0.118153855,0.108307704,0.118153855,0.13456412,0.17723078,0.27241027,0.508718,0.69251287,1.0108719,1.4080001,1.6016412,1.3489232,1.273436,1.2668719,1.2406155,1.148718,0.6432821,0.4660513,0.5021539,0.6235898,0.6859488,0.6104616,0.65641034,0.6268718,0.512,0.49887183,0.6498462,0.69907695,0.7844103,0.88943595,0.8467693,0.6301539,0.5874872,0.65641034,0.79097444,0.95835906,1.3751796,1.9528207,2.3893335,2.540308,2.4155898,2.0151796,1.6016412,1.5130258,1.529436,0.8730257,0.69251287,0.7515898,0.955077,1.017436,0.48574364,0.2986667,0.20676924,0.23302566,0.36430773,0.5677949,0.6235898,0.761436,0.9682052,1.1388719,1.0962052,0.7811283,0.69907695,0.6826667,0.7187693,0.94523084,1.0962052,1.1749744,1.2931283,1.3489232,1.017436,0.92225647,0.67282057,0.46276927,0.4135385,0.571077,0.34133336,0.27897438,0.2855385,0.33476925,0.47917953,1.3357949,1.4244103,2.1464617,4.4110775,8.648206,9.048616,6.0750775,4.46359,4.9493337,4.263385,2.6945643,4.4307694,5.0018463,3.636513,3.249231,3.0752823,2.0808206,0.88287187,0.032820515,0.04266667,0.14112821,0.16738462,0.17723078,0.18707694,0.18379489,0.33805132,0.4004103,0.4266667,0.46276927,0.52512825,0.51856416,0.55794877,0.65969235,0.8369231,1.0699488,1.1257436,1.3915899,1.4408206,1.2340513,1.1027694,0.92225647,0.9485129,1.1027694,1.2012309,0.955077,1.0929232,1.1651284,1.1355898,1.2012309,1.782154,2.3958976,5.037949,7.197539,8.562873,11.027693,12.822975,11.001437,11.07036,12.100924,6.741334,4.2240005,5.3431797,5.4514875,3.1442053,0.25271797,0.10502565,0.21989745,0.28882053,0.30851284,0.5940513,0.77456415,0.955077,1.014154,0.90584624,0.65641034,0.9747693,0.92553854,0.81066674,0.7844103,0.82379496,1.1323078,1.2307693,1.0436924,0.74830776,0.79425645,1.0305642,0.98461545,0.98133343,1.020718,0.77456415,0.380718,0.15425642,0.04266667,0.0032820515,0.0,0.0032820515,0.02297436,0.12471796,0.26912823,0.3052308,0.46276927,0.65641034,0.8041026,0.86646163,0.8566154,0.86646163,1.014154,1.024,0.8795898,0.8369231,1.0765129,1.1651284,1.1946667,1.2471796,1.4145643,1.5425643,1.591795,1.6475899,1.6836925,1.5721027,1.7558975,2.2613335,2.7076926,2.993231,3.2886157,3.2886157,3.56759,3.9844105,4.450462,4.906667,4.588308,4.2863593,3.9581542,3.6890259,3.7185643,3.7382567,3.9876926,4.210872,4.391385,4.7392826,4.59159,4.850872,5.221744,5.6943593,6.5378466,6.7872825,7.250052,7.857231,8.237949,7.7357955,6.931693,6.3474874,6.0291286,5.756718,5.0149746,5.2644105,5.668103,5.868308,5.861744,5.9995904,5.85518,5.8190775,5.622154,5.421949,5.792821,6.554257,7.24677,7.6603084,7.6964107,7.394462,7.1614366,7.4174366,7.7456417,7.9195905,7.9294367,7.5421543,7.1844106,6.701949,6.482052,7.456821,7.778462,7.4174366,6.99077,6.7314878,6.485334,6.048821,6.1768208,6.774154,7.6570263,8.546462,7.8506675,7.834257,8.054154,8.182155,8.004924,7.9786673,7.824411,7.837539,8.073847,8.329846,7.653744,7.3550773,7.0334363,6.76759,7.1581545,7.213949,7.059693,6.157129,4.775385,3.9942567,4.1485133,4.076308,3.9548721,3.9056413,3.9811285,4.460308,4.7392826,4.9099493,4.9132314,4.535795,4.8804107,5.3169236,5.7501545,5.8945646,5.2676926,4.716308,4.713026,5.2611284,5.792821,5.179077,4.3585644,3.9745643,3.5807183,3.0982566,2.8127182,2.878359,3.308308,3.7874875,4.027077,3.7940516,3.4330258,2.9144619,2.5829747,2.5665643,2.7667694,2.4648206,2.103795,1.9462565,1.9561027,1.7952822,0.47261542,0.21661541,0.318359,0.47589746,0.6465641,1.0371283,0.86646163,0.45620516,0.17066668,0.08861539,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.15097436,0.15097436,0.02297436,0.06235898,0.17066668,0.18051283,0.4004103,0.8041026,1.0371283,1.1355898,0.95835906,0.702359,0.47589746,0.3052308,0.256,0.27241027,0.24615386,0.20348719,0.28882053,0.31507695,0.3117949,0.24943592,0.14769232,0.06235898,0.18379489,0.3708718,0.55794877,0.761436,1.0666667,1.5819489,2.7798977,3.629949,3.4789746,2.0742567,1.8445129,1.847795,2.0151796,2.228513,2.349949,2.5698464,2.6322052,3.0720003,4.0402055,5.3103595,6.944821,9.222565,11.516719,14.020925,17.729643,21.67467,24.425028,25.38995,25.281643,26.12185,28.419285,33.98236,41.50154,48.797543,52.82462,56.43816,62.706875,72.61211,82.11693,82.16616,82.543594,82.32698,82.09724,81.250465,78.01765,68.24042,54.816826,44.10749,38.787285,37.871593,48.91898,72.608826,100.204315,115.64637,95.56678,51.649647,29.38749,22.088207,22.774155,24.201847,24.323284,23.35508,23.781746,25.780516,27.221336,29.052721,28.980515,27.369028,24.65149,21.333336,26.60431,30.34913,30.070156,25.176617,17.001026,15.619284,16.410257,20.516104,26.266258,29.157745,29.121643,29.689438,33.06995,35.21641,25.816618,28.563694,30.687181,25.212719,14.641232,10.939077,15.9343605,18.241642,19.433027,19.373951,16.249437,14.03077,14.290052,13.850258,11.999181,10.499283,7.77518,5.8223596,5.3037953,5.937231,6.5017443,7.9294367,7.6734366,8.044309,9.216001,9.216001,8.155898,6.8627696,5.2512827,4.417641,6.6527185,7.433847,6.5772314,6.5411286,7.5979495,7.8441033,10.637129,11.585642,11.204924,10.19077,9.383386,7.8080006,7.755488,8.316719,8.52677,7.3550773,8.4053335,9.032206,10.587898,12.740924,13.472821,12.924719,11.687386,10.161232,8.65477,7.384616,7.653744,7.8769236,7.8637953,7.456821,6.514872,6.626462,6.47877,6.009436,5.7074876,6.62318,9.4916935,13.659899,17.168411,18.011898,14.129231,13.5548725,11.818667,10.029949,8.953437,9.002667,8.904206,9.025641,9.478565,9.980719,9.872411,10.886565,11.753027,11.674257,10.656821,9.521232,8.753231,7.8014364,7.6242056,8.185436,8.454565,6.2555904,6.245744,6.9842057,7.2927184,6.2555904,4.9493337,5.044513,5.5072823,5.7731285,5.737026,3.9811285,2.789744,2.6847181,3.2722054,3.2361028,3.7120004,4.699898,4.9132314,5.0871797,7.9819493,7.637334,18.996513,21.920822,14.444309,12.770463,7.8408213,5.720616,4.1124105,2.7175386,3.2032824,4.7556925,4.2436924,3.95159,4.2305646,3.508513,2.3729234,3.1442053,4.1189747,4.6276927,5.0051284,3.1376412,2.3236926,2.0053334,1.6935385,0.9616411,0.3511795,0.446359,0.5677949,1.0962052,3.4625645,2.8291285,2.8914874,4.6802053,6.6034875,4.457026,7.88677,20.352001,28.517746,27.789131,22.308104,20.050053,16.226463,12.868924,12.882052,20.033642,11.769437,6.2063594,6.048821,9.104411,8.28718,33.70995,21.43836,9.4457445,14.427898,31.783386,14.729847,12.041847,16.564514,19.541334,10.604308,7.2861543,7.8834877,8.756514,8.283898,6.882462,5.028103,6.12759,6.189949,4.417641,3.2361028,3.761231,7.8080006,10.545232,11.139283,12.786873,5.5007186,2.6880002,4.4767184,7.4075904,4.4406157,5.6352825,8.169026,6.4590774,1.4769232,0.7318975,0.6826667,1.6246156,2.3302567,2.3827693,2.1530259,3.31159,2.858667,2.1530259,1.7066668,1.204513,1.024,0.69251287,0.7417436,1.2406155,1.8149745,1.9495386,2.1202054,1.9429746,1.467077,1.1749744,2.028308,3.8990772,4.4012313,3.761231,4.821334,3.5282054,3.2853336,3.9286156,4.46359,3.0982566,1.9265642,1.8806155,2.3794873,2.9604106,3.2656412,2.678154,1.7920002,1.2406155,1.0666667,0.6859488,0.892718,0.98133343,0.95835906,0.88615394,0.88615394,0.8369231,0.5481026,0.27569234,0.118153855,0.04594872,0.18051283,0.31507695,0.33805132,0.30851284,0.44307697,1.0404103,0.9419488,1.0404103,1.723077,2.8849232,2.1497438,1.6213335,1.2373334,0.93866676,0.67282057,0.5481026,0.41025645,0.39056414,0.49230772,0.56451285,0.57764107,0.54482055,0.512,0.512,0.5481026,0.7089231,0.6662565,0.67610264,0.81066674,0.94523084,0.92225647,0.761436,0.6695385,0.6662565,0.58092314,0.8598975,1.7920002,2.6289232,3.1113849,3.4789746,2.5009232,1.8904617,1.4966155,1.2996924,1.4342566,0.9714873,0.90912825,1.014154,1.0108719,0.5940513,0.3511795,0.35446155,0.52512825,0.761436,0.94523084,1.0305642,1.0535386,1.0535386,1.0469744,1.020718,0.9124103,0.9124103,0.761436,0.51856416,0.58092314,0.9353847,1.5622566,2.0151796,1.9692309,1.2373334,0.77128214,0.6826667,0.6104616,0.48574364,0.5349744,0.31507695,0.26912823,0.2986667,0.32164106,0.25928208,0.3446154,0.40369233,0.65969235,1.4211283,3.0818465,5.3760004,4.896821,4.6539493,5.0674877,3.9811285,2.0545642,2.3958976,3.1770258,3.5807183,3.8006158,3.751385,2.9505644,1.4933335,0.07876924,0.029538464,0.029538464,0.03938462,0.06564103,0.108307704,0.18379489,0.32820517,0.512,0.5973334,0.574359,0.5481026,0.52512825,0.49230772,0.571077,0.79097444,1.083077,1.0601027,1.0699488,1.3259488,1.6508719,1.4802053,1.2603078,1.1684103,1.1126155,1.0765129,1.1126155,1.0666667,1.024,1.1290257,1.4900514,2.1956925,2.917744,4.2962055,6.892308,8.966565,6.5017443,7.453539,9.714872,11.349334,12.42913,15.028514,7.2303596,3.3214362,2.937436,3.5971284,0.71548724,0.16738462,0.10502565,0.21989745,0.33805132,0.4135385,0.58420515,0.7187693,0.9124103,1.0469744,0.7778462,0.764718,0.65312827,0.67610264,0.81066674,0.761436,0.6892308,0.79097444,0.8467693,0.8172308,0.8533334,0.96492314,0.90912825,1.0371283,1.2504616,1.0075898,0.446359,0.15097436,0.032820515,0.013128206,0.0,0.013128206,0.032820515,0.108307704,0.20676924,0.24287182,0.29210258,0.46933338,0.7187693,0.955077,1.0535386,0.80738467,0.77456415,0.76800007,0.7515898,0.82379496,1.142154,1.2668719,1.2373334,1.1716924,1.2832822,1.4276924,1.585231,1.6640002,1.6311796,1.5097437,1.7427694,1.9364104,2.2482052,2.6420515,2.8980515,2.7044106,2.9768207,3.3608208,3.5905645,3.4789746,3.1967182,3.05559,3.062154,3.121231,3.0358977,3.7185643,3.9745643,4.0402055,3.945026,3.495385,3.7874875,4.519385,4.9099493,4.8771286,5.034667,6.5378466,7.6635904,8.274052,8.139488,6.941539,6.1505647,5.8518977,5.3431797,4.634257,4.4406157,4.46359,4.535795,4.713026,4.8049235,4.3651285,4.3749747,4.7360005,4.900103,4.9493337,5.586052,6.0258465,6.7840004,6.8627696,6.2588725,5.9667697,6.2096415,7.1220517,7.6603084,7.64718,7.781744,7.6110773,7.3583593,7.2369237,7.712821,9.504821,9.225847,8.805744,8.648206,8.631796,8.132924,6.2523084,5.9667697,6.242462,6.665847,7.4469748,6.5050263,7.243488,8.323282,9.055181,9.383386,9.055181,8.815591,8.723693,8.720411,8.635077,8.073847,7.194257,6.4722056,6.1341543,6.1341543,6.547693,6.5805135,5.8518977,4.8016415,4.6539493,4.59159,4.5029745,4.2896414,3.9581542,3.6168208,3.9089234,4.414359,4.900103,5.353026,5.9503593,5.5729237,5.5138464,5.7829747,6.11118,5.9503593,5.4875903,5.097026,4.906667,4.850872,4.6539493,4.604718,4.5456414,3.9680004,3.0326157,2.5928206,2.422154,2.737231,3.242667,3.5741541,3.2820516,2.806154,2.878359,2.806154,2.425436,2.1202054,2.0217438,2.0709746,2.1398976,2.1103592,1.8904617,0.28882053,0.16082053,0.17723078,0.21661541,0.2855385,0.5021539,0.4660513,0.33476925,0.20676924,0.12143591,0.026256412,0.016410258,0.016410258,0.009846155,0.006564103,0.026256412,0.006564103,0.14769232,0.3511795,0.5415385,0.6465641,0.7581539,0.98461545,0.9911796,0.8763078,1.1946667,0.8336411,0.9517949,0.88287187,0.53825647,0.4266667,0.45620516,0.46276927,0.52512825,0.6826667,0.92553854,0.95835906,0.827077,0.5546667,0.28225642,0.24287182,0.42338464,0.8467693,1.3423591,1.8346668,2.3236926,3.249231,5.297231,5.9536414,4.6802053,2.9046156,2.048,1.723077,1.7657437,1.9659488,2.0676925,2.7569232,3.4888208,4.7524104,6.5903597,8.592411,9.429334,11.211488,13.722258,16.66954,19.695591,21.67467,24.30359,25.606565,25.961027,28.100925,37.034668,45.4958,51.52821,55.12862,58.256416,70.912,85.98975,97.01416,100.535805,96.13129,90.12514,83.360825,78.332726,76.209236,76.82298,67.92206,59.46749,55.742363,56.8878,58.902977,68.39796,87.20411,104.4119,103.24349,61.046158,30.79877,17.72636,15.00554,16.800821,18.267899,18.369642,17.969233,18.182566,18.694565,17.762463,20.178053,21.159386,21.530258,21.26113,19.465847,17.345642,17.673847,16.613745,13.551591,11.116308,12.819694,16.439796,21.4679,26.308926,28.294567,27.221336,25.780516,26.689644,28.649029,26.318771,27.618464,23.83754,19.255796,17.880617,23.440413,19.321438,18.753643,21.185642,22.98749,17.47036,14.165335,13.413745,12.251899,10.535385,10.939077,12.422565,10.308924,7.643898,6.166975,6.2687182,6.1538467,6.1407185,7.1647186,8.766359,9.117539,7.9885135,8.3134365,7.5552826,6.0160003,6.8233852,6.921847,6.6395903,6.8529234,7.6734366,8.454565,11.628308,11.227899,10.594462,10.637129,9.810052,10.354873,11.52,12.002462,11.644719,11.418258,12.2847185,12.324103,12.859077,13.879796,14.034052,12.918155,12.025436,11.07036,9.878975,8.385642,9.025641,8.881231,8.339693,7.6734366,7.017026,6.921847,6.4590774,6.173539,6.518154,7.8539495,9.80677,12.580104,14.313026,14.375385,13.37436,12.721231,10.7158985,8.52677,7.1122055,7.2205133,8.198565,8.726975,9.344001,10.134975,10.725744,12.130463,13.820719,13.361232,11.172104,10.535385,9.481847,7.9327188,6.8332314,6.8397956,8.320001,7.2237954,7.000616,6.8365135,6.38359,5.756718,4.519385,4.6145644,4.8147697,4.6112823,4.2240005,3.0720003,2.0906668,2.0512822,2.7667694,3.1015387,3.879385,4.33559,4.2896414,5.110154,9.701744,8.812308,13.581129,16.180513,14.588719,12.612924,8.109949,5.651693,3.7973337,2.605949,3.629949,5.346462,4.5423594,3.751385,3.8695388,4.1550775,2.6880002,2.7733335,3.2787695,3.7907696,4.6276927,3.4625645,2.7044106,2.3991797,2.2514873,1.6443079,0.8795898,0.7417436,0.7975385,1.3029745,3.2328207,2.802872,3.5511796,6.4032826,8.89436,5.1626673,5.792821,7.194257,8.960001,10.14154,9.258667,12.117334,12.153437,8.979693,5.622154,8.487385,7.584821,7.5618467,6.6461544,5.481026,7.1122055,24.84513,20.916515,15.225437,19.570873,37.632004,18.048002,13.571283,13.239796,11.605334,8.713847,8.976411,8.493949,10.102155,11.388719,4.673641,3.2754874,4.2568207,4.7228723,5.2676926,9.961026,10.971898,9.813334,13.042872,17.027283,7.9524107,14.6182575,9.826463,5.2545643,5.028103,5.720616,7.778462,6.160411,3.186872,0.86646163,0.90256417,1.3718976,2.0250258,2.1366155,1.8281027,2.0644104,2.0742567,2.0086155,2.041436,2.0184617,1.4506668,0.8172308,1.401436,1.7263591,1.5721027,1.9495386,1.8313848,1.3751796,1.0371283,1.0272821,1.3095386,2.1825643,3.370667,3.6791797,3.2262566,3.4297438,3.1015387,3.5577438,4.4767184,5.0018463,3.7316926,2.8816411,2.537026,3.05559,3.820308,3.2164104,2.1825643,1.4605129,1.3161026,1.4408206,0.955077,0.7811283,0.7811283,0.8795898,0.98133343,0.98133343,1.0601027,0.9682052,0.955077,0.9189744,0.38728207,0.27897438,0.4397949,0.5218462,0.43651286,0.3446154,0.571077,0.56451285,0.6432821,1.0502565,1.9561027,2.0742567,1.595077,1.0732309,0.81066674,0.8533334,0.6826667,0.44307697,0.35774362,0.4266667,0.42994875,0.4135385,0.3708718,0.35774362,0.4135385,0.5973334,0.7581539,0.7056411,0.7778462,1.0896411,1.5556924,1.6377437,1.4736412,1.1191796,0.77456415,0.78769237,0.9419488,1.5688206,2.3368206,2.9407182,3.1113849,2.8882053,2.6256413,2.0873847,1.467077,1.3981539,1.1881026,0.9189744,0.90584624,0.9878975,0.5349744,0.25928208,0.3511795,0.53825647,0.6662565,0.702359,0.9353847,1.2274873,1.273436,1.1290257,1.1946667,0.96492314,0.892718,0.80738467,0.7450257,0.92225647,1.0305642,1.394872,1.7296412,1.7624617,1.2373334,0.636718,0.46276927,0.48246157,0.5481026,0.6071795,0.574359,0.38400003,0.23958977,0.19692309,0.18707694,0.21333335,0.256,0.32820517,0.512,0.9714873,1.8806155,2.540308,3.820308,5.4875903,6.229334,6.0685134,4.7261543,3.8564105,3.7349746,3.2623591,2.1989746,2.1924105,2.038154,1.273436,0.190359,0.12143591,0.04594872,0.026256412,0.06235898,0.08533334,0.1148718,0.26256412,0.44307697,0.571077,0.53825647,0.5021539,0.48902568,0.54482055,0.6629744,0.79097444,0.88287187,1.0994873,1.2832822,1.3522053,1.2964103,1.2340513,1.1881026,1.0732309,0.9517949,1.017436,1.211077,1.270154,1.3620514,1.8806155,3.4166157,3.318154,3.5905645,5.3070774,7.702975,8.185436,9.458873,10.006975,8.92718,7.8736415,11.050668,7.762052,4.84759,3.9548721,4.4996924,3.6594875,0.77456415,0.10502565,0.20676924,0.3446154,0.49887183,0.60061544,0.61374366,0.65969235,0.7778462,0.9485129,0.69251287,0.5415385,0.56123084,0.6826667,0.702359,0.6465641,0.81394875,0.9156924,0.8566154,0.7089231,0.69907695,0.7253334,0.8205129,0.88943595,0.71548724,0.34789747,0.12143591,0.026256412,0.013128206,0.013128206,0.0032820515,0.036102567,0.0951795,0.16738462,0.24287182,0.4397949,0.6104616,0.74830776,0.8566154,0.9419488,0.9124103,0.9714873,0.955077,0.8730257,0.8960001,1.1060513,1.2274873,1.3029745,1.3029745,1.1093334,1.1782565,1.3456411,1.3522053,1.211077,1.204513,1.339077,1.8412309,2.2088206,2.2580514,2.1070771,2.0873847,2.356513,2.7963078,3.0523078,2.550154,2.7602053,2.665026,2.556718,2.5928206,2.7798977,3.318154,3.5052311,3.6562054,3.8662567,4.0303593,3.945026,4.279795,4.7294364,5.149539,5.5729237,6.8299494,7.499488,7.9491286,8.254359,8.198565,6.9087186,5.605744,4.844308,4.5817437,4.1714873,3.7087183,3.6693337,3.8432825,3.9056413,3.436308,3.7218463,3.9154875,4.1550775,4.535795,5.1331286,6.0717955,6.954667,7.4732313,7.496206,7.076103,6.521436,6.419693,7.131898,8.392206,9.3078985,8.490667,8.3134365,8.828718,9.6754875,10.056206,9.324308,8.815591,8.736821,8.881231,8.644924,7.282872,6.882462,7.0859494,7.456821,7.506052,6.6067696,6.744616,7.5552826,8.576,9.238976,8.674462,8.326565,8.146052,8.178872,8.562873,7.9130263,7.1844106,6.5444107,6.232616,6.5739493,6.0028725,5.6320004,5.3398976,5.0904617,4.9362054,4.8738465,4.673641,4.44718,4.2305646,4.007385,4.086154,4.519385,4.8771286,5.07077,5.366154,5.2512827,5.0904617,5.221744,5.5302567,5.4514875,5.074052,4.640821,4.71959,5.0904617,4.7392826,4.086154,3.882667,3.8400004,3.754667,3.508513,3.4756925,3.3542566,3.3247182,3.3280003,3.0851285,2.8127182,2.7109745,2.6978464,2.7273848,2.802872,2.6289232,2.4615386,2.28759,2.097231,1.8674873,0.23630771,0.256,0.17394873,0.10502565,0.12143591,0.24615386,0.29210258,0.31507695,0.3511795,0.33476925,0.11158975,0.026256412,0.006564103,0.013128206,0.08861539,0.3314872,0.702359,1.0305642,1.2504616,1.339077,1.3062565,1.4736412,1.3226668,1.1027694,1.0010257,1.1454359,1.1093334,1.2996924,1.2603078,0.98133343,0.8960001,0.8566154,1.1848207,1.529436,1.6935385,1.6147693,1.3587693,0.99774367,0.6662565,0.48902568,0.6104616,1.0633847,1.8412309,2.7011285,3.43959,3.9023592,5.330052,6.803693,6.5903597,4.6605134,2.6912823,1.913436,1.7920002,1.9889232,2.2153847,2.2449234,3.0358977,5.159385,8.136206,10.994873,12.281437,11.690667,12.580104,14.818462,17.414566,18.520617,19.748104,22.452515,24.822155,27.247591,32.3479,42.436928,52.096004,60.05826,67.59057,78.50011,87.53888,88.940315,85.0478,78.47057,72.08698,65.48677,59.900723,60.333954,68.33231,81.99878,75.6677,70.52473,69.12985,69.46462,64.932106,77.17416,103.77847,111.44206,86.8956,36.92308,19.410053,12.888617,11.602052,12.251899,13.991385,14.112822,13.489232,12.816411,12.461949,12.465232,13.522053,14.053744,14.506668,14.447591,12.570257,9.849437,9.337437,9.088,8.828718,9.980719,12.563693,15.684924,20.325745,25.527798,28.406157,25.383387,25.193027,25.14708,24.211695,22.984207,24.74995,21.661541,20.46359,22.938257,25.898668,23.72595,23.70954,23.850668,21.707489,14.388514,10.315488,9.6295395,10.210463,10.7848215,10.939077,11.798975,10.374565,7.7390776,5.280821,4.71959,4.6933336,5.9667697,8.94359,11.82195,10.5780525,8.192,8.667898,8.201847,6.3245134,5.904411,6.8660517,8.083693,8.5661545,8.346257,8.487385,11.969642,11.16554,9.885539,9.619693,9.5146675,11.247591,12.668719,13.259488,13.275898,13.725539,14.04718,12.832822,12.452104,13.35795,14.073437,12.898462,11.841642,10.755282,9.882257,9.862565,9.189744,8.4283085,7.824411,7.4436927,7.197539,7.1220517,7.351795,7.781744,8.2445135,8.5202055,9.649232,10.955488,11.651283,11.779283,12.196103,10.463181,8.339693,6.6067696,5.799385,6.1997952,7.860513,8.73354,9.278359,9.862565,10.758565,12.425847,13.226667,12.373334,10.617436,10.266257,9.501539,7.243488,5.910975,6.0652313,6.416411,6.6625648,6.12759,5.4613338,5.0215387,4.8705645,3.5774362,3.4034874,3.495385,3.4330258,3.239385,2.3072822,1.6246156,1.9856411,3.3542566,4.8804107,4.9493337,5.0838976,5.333334,6.7577443,11.431385,9.908514,13.1872835,18.313848,21.746874,19.328001,16.200207,12.265027,8.89436,6.8430777,6.23918,6.0192823,5.1232824,4.1583595,3.7382567,4.46359,3.0982566,3.0949745,3.5314875,4.023795,4.7425647,4.2141542,3.3312824,2.7536411,2.5238976,2.0545642,1.5261539,1.0962052,0.8533334,1.2898463,3.2918978,3.1277952,7.8473854,9.826463,7.643898,6.0816417,9.488411,8.169026,6.7183595,6.373744,5.0084105,8.303591,10.036513,10.308924,8.772923,4.630975,6.806975,12.130463,14.073437,11.526565,8.805744,15.527386,13.948719,13.049437,16.922258,24.776207,15.113848,12.163283,11.690667,10.925949,8.54318,8.14277,8.690872,10.410667,11.802258,9.639385,5.464616,6.3245134,5.435077,3.446154,8.448001,11.963078,10.706052,9.442462,8.812308,5.32677,13.732103,13.124924,10.466462,8.615385,6.308103,9.941334,7.1154876,3.4264617,1.5819489,1.404718,1.6344616,1.7723079,1.9003079,2.0545642,2.2088206,2.300718,2.8258464,3.3280003,3.3608208,2.4910772,1.6508719,1.8379488,1.9364104,1.6738462,1.6344616,1.591795,2.3138463,2.540308,2.1956925,2.3958976,1.9626669,2.4910772,2.8750772,2.7241027,2.359795,2.7995899,3.1113849,3.6693337,4.1517954,3.5446157,2.7602053,2.484513,2.3827693,2.4681027,3.1048207,2.4615386,1.7690258,1.4572309,1.3587693,0.7187693,0.56123084,0.7450257,1.0962052,1.3292309,1.0436924,1.0010257,1.142154,1.1618463,0.9124103,0.39056414,0.30851284,0.43651286,0.46933338,0.34133336,0.24615386,0.4266667,0.7384616,0.7844103,0.72861546,1.2832822,1.6935385,1.4408206,1.1093334,0.9714873,0.98133343,0.84348726,0.5874872,0.4955898,0.5513847,0.45292312,0.44307697,0.39056414,0.35774362,0.39712822,0.56451285,0.7515898,0.7187693,0.7450257,0.94523084,1.2603078,1.723077,1.9035898,1.5491283,0.9878975,1.142154,1.2209232,1.3489232,1.8806155,2.6157951,2.809436,2.8192823,2.9669745,2.5796926,1.7920002,1.5524104,1.5688206,1.1946667,1.0371283,1.0994873,0.764718,0.4397949,0.4004103,0.5316923,0.67282057,0.61374366,0.764718,1.017436,1.2406155,1.3653334,1.401436,1.0633847,0.7975385,0.64000005,0.67938465,1.0699488,1.0699488,1.1651284,1.332513,1.394872,1.0436924,0.6498462,0.5218462,0.4955898,0.4955898,0.54482055,0.48902568,0.36102566,0.23302566,0.14441027,0.13128206,0.15753847,0.17394873,0.16410258,0.16082053,0.23302566,0.44307697,0.892718,1.9856411,4.3651285,8.914052,6.629744,4.4438977,3.7251284,4.2305646,4.07959,2.6945643,2.6518977,2.7963078,2.4713848,1.4998976,1.7165129,1.1520001,0.5021539,0.12471796,0.04266667,0.055794876,0.16410258,0.32164106,0.46933338,0.5349744,0.51856416,0.5481026,0.58420515,0.61374366,0.67282057,0.764718,0.9485129,1.020718,0.96492314,0.93866676,0.9682052,1.017436,0.98133343,0.90256417,0.98133343,1.1651284,1.2406155,1.467077,2.0151796,2.9538465,3.006359,2.858667,4.0303593,6.363898,8.001641,6.567385,7.9983597,7.276308,4.7589746,6.173539,7.2369237,5.691077,3.8728209,2.9243078,2.793026,0.7318975,0.14112821,0.18379489,0.380718,0.6104616,0.5349744,0.60061544,0.6662565,0.69251287,0.7450257,0.74830776,0.7778462,0.6892308,0.5284103,0.512,0.6104616,0.78769237,0.86317956,0.79425645,0.67282057,0.63343596,0.67610264,0.73517954,0.77128214,0.761436,0.34789747,0.1148718,0.01969231,0.006564103,0.006564103,0.0,0.036102567,0.08205129,0.13128206,0.21661541,0.39712822,0.5152821,0.6301539,0.761436,0.8598975,0.8402052,0.90256417,0.88287187,0.827077,1.0075898,1.1323078,1.148718,1.1979488,1.2274873,1.0043077,1.0371283,1.1191796,1.1027694,1.0404103,1.1651284,1.1716924,1.6902566,2.1333334,2.2121027,1.9364104,2.0118976,2.0578463,2.1103592,2.1333334,2.0184617,2.553436,2.537026,2.4188719,2.4615386,2.7602053,3.0358977,3.045744,3.0424619,3.1573336,3.387077,3.7842054,4.0500517,4.3749747,4.8147697,5.3037953,6.5805135,7.4075904,7.968821,8.329846,8.4512825,6.9677954,5.9470773,5.2315903,4.663795,4.1058464,3.3641028,3.0752823,3.2164104,3.4888208,3.314872,3.43959,3.5478978,3.7907696,4.2994876,5.1856413,5.805949,6.5903597,7.181129,7.384616,7.1909747,6.7840004,6.8988724,7.7981544,9.170052,10.128411,9.380103,9.380103,9.796924,10.118565,9.642668,8.595693,8.129642,8.444718,9.104411,9.02236,8.12636,8.280616,8.674462,8.704,7.9983597,7.128616,6.6822567,6.7872825,7.4075904,8.349539,8.050873,7.6898465,7.4896417,7.6898465,8.52677,8.01477,7.64718,6.8529234,5.8945646,5.868308,5.093744,4.972308,4.9985647,4.8738465,4.46359,4.397949,4.2896414,4.2272825,4.2371287,4.2962055,4.138667,4.457026,4.713026,4.8377438,5.218462,5.1922054,4.965744,5.0609236,5.398975,5.3070774,5.106872,4.8049235,4.8377438,5.0477953,4.6867695,4.2568207,3.9351797,3.7907696,3.7776413,3.7185643,3.8596926,3.6430771,3.43959,3.2361028,2.6518977,2.550154,2.609231,2.5895386,2.5173335,2.681436,2.9407182,2.858667,2.553436,2.1103592,1.5786668,0.24615386,0.256,0.15097436,0.06235898,0.052512825,0.12471796,0.19364104,0.34133336,0.46276927,0.45292312,0.21661541,0.06235898,0.016410258,0.1148718,0.36758977,0.74830776,1.8937438,2.359795,1.9823592,1.204513,1.079795,1.3554872,1.1191796,0.8763078,0.83035904,0.85005134,1.0043077,1.2274873,1.467077,1.8018463,2.4155898,1.9429746,1.9593848,2.1825643,2.2678976,1.8281027,1.3620514,1.0601027,0.92225647,0.95835906,1.1946667,2.359795,3.5052311,4.634257,5.7435904,6.806975,7.9195905,7.8670774,6.409847,4.135385,2.4582565,1.9823592,1.9429746,2.1858463,2.6453335,3.3575387,5.0215387,7.686565,10.561642,12.668719,12.836103,12.383181,13.029744,14.713437,16.745028,17.831387,19.88595,22.852924,25.928207,29.860106,36.942772,46.336002,60.402878,77.08883,93.6238,106.53539,99.74155,82.228516,64.84021,53.120003,47.323902,44.278156,42.61744,47.405952,59.62175,76.14688,79.03508,79.645546,76.00903,68.45703,59.6119,76.3438,102.19981,99.360825,62.94975,21.031385,13.866668,11.1294365,9.829744,9.196308,10.683078,11.418258,10.807796,9.317744,8.067283,8.822155,8.838565,8.776206,8.960001,8.960001,7.6143594,6.7905645,6.2752824,6.432821,7.6701546,10.459898,13.069129,15.048206,18.838976,24.329847,28.855797,28.09108,28.763899,26.807796,22.377028,19.840002,19.990976,19.6759,20.87713,22.994053,22.826668,24.664618,26.676516,24.405334,17.99877,12.179693,8.999385,8.093539,8.969847,10.341744,10.151385,10.8767185,9.741129,7.515898,5.2512827,4.2896414,4.57518,7.4863596,10.568206,11.746463,9.337437,7.0859494,7.131898,7.003898,6.2227697,6.2884107,6.8233852,8.812308,9.432616,8.54318,8.677744,11.739899,10.666668,9.18318,9.005949,9.833026,12.4685135,14.752822,15.353437,14.795488,15.471591,14.624822,12.566976,11.490462,12.028719,13.239796,12.553847,11.401847,10.105436,9.3078985,9.974154,8.756514,8.155898,7.781744,7.6307697,8.073847,8.300308,9.334154,10.04636,9.878975,8.851693,8.572719,8.999385,9.3768215,9.655796,10.47959,8.444718,6.7183595,5.737026,5.6352825,6.245744,7.9294367,8.94359,9.248821,9.278359,9.93477,11.749744,12.025436,11.001437,9.573745,9.288206,8.411898,6.5411286,5.723898,5.8223596,4.5062566,5.7632823,5.3792825,4.667077,4.3060517,4.345436,2.930872,2.3893335,2.356513,2.6256413,3.1507695,2.3762052,1.6771283,2.1956925,4.010667,6.1308722,5.4580517,6.439385,7.6570263,9.120821,12.2617445,10.988309,13.371078,20.17477,26.807796,23.345232,23.190975,18.648617,13.794462,10.489437,8.362667,6.4032826,5.8978467,5.3431797,4.5456414,4.630975,3.8498464,3.8498464,4.1682053,4.673641,5.5958977,5.8814363,4.59159,3.2623591,2.550154,2.231795,1.8838975,1.2931283,0.8041026,1.0699488,3.0358977,2.8258464,8.454565,11.250873,9.511385,8.51036,9.4457445,8.054154,8.132924,9.133949,6.1440005,6.5837955,9.291488,13.594257,15.031796,5.3694363,7.9130263,13.846975,20.926361,23.092514,10.486155,10.443488,8.766359,11.907283,17.539284,14.555899,13.147899,11.178667,11.090053,12.09436,10.164514,7.351795,7.5946674,8.720411,9.357129,8.933744,7.453539,12.895181,15.675078,12.448821,6.121026,12.635899,12.1468725,7.4896417,3.515077,7.062975,11.920411,17.434258,17.490053,12.196103,7.899898,7.955693,5.612308,3.1081028,1.8510771,2.412308,1.7099489,1.4966155,1.8018463,2.3171284,2.412308,2.2646155,2.7995899,3.5216413,3.7973337,2.868513,2.0775387,1.7296412,1.595077,1.4506668,1.0666667,1.6475899,3.7809234,4.7360005,4.0500517,3.5183592,1.9790771,2.2482052,2.6256413,2.425436,1.9987694,2.4320002,2.5173335,2.5961027,2.7044106,2.5862565,2.1333334,2.0644104,1.8543591,1.7887181,2.9440002,2.4582565,1.7952822,1.273436,0.92553854,0.4955898,0.41025645,0.6301539,1.0075898,1.3095386,1.2340513,0.82379496,0.8795898,0.8795898,0.65312827,0.39056414,0.40369233,0.42994875,0.36102566,0.23630771,0.23630771,0.5021539,1.3620514,1.5688206,1.0601027,0.9616411,1.3554872,1.2438976,1.1355898,1.1454359,1.0010257,0.892718,0.67938465,0.5973334,0.62030774,0.46933338,0.5284103,0.5021539,0.45620516,0.45292312,0.55794877,0.7089231,0.6498462,0.6235898,0.7220513,0.88287187,1.6278975,1.9561027,1.657436,1.1027694,1.2340513,1.3784616,1.211077,1.4342566,2.1234872,2.7241027,2.537026,2.7142565,2.6847181,2.2514873,1.595077,2.044718,1.7263591,1.3489232,1.2012309,1.1323078,0.78769237,0.65312827,0.81066674,1.0272821,0.7844103,0.7220513,0.78769237,0.9517949,1.1388719,1.2603078,1.270154,0.9485129,0.7122052,0.75487185,1.0601027,1.0601027,0.9747693,0.9747693,0.99774367,0.7384616,0.6465641,0.57764107,0.48246157,0.42338464,0.574359,0.5349744,0.5218462,0.39712822,0.20020515,0.13784617,0.1148718,0.10502565,0.11158975,0.12471796,0.1148718,0.07548718,0.13456412,0.571077,2.540308,8.054154,5.4580517,3.6857438,3.3903592,4.1124105,4.3060517,2.9702566,3.1540515,3.6890259,3.5610259,1.9232821,2.2153847,2.294154,1.7558975,0.79425645,0.19692309,0.08205129,0.108307704,0.20348719,0.3249231,0.4594872,0.47589746,0.508718,0.5349744,0.5677949,0.65312827,0.6662565,0.7581539,0.764718,0.6859488,0.6892308,0.73517954,0.79425645,0.82379496,0.84348726,0.9288206,1.1257436,1.2668719,1.6114873,2.1136413,2.422154,2.6715899,2.4484105,2.9833848,4.604718,6.7249236,4.650667,6.892308,6.9152827,4.096,3.7251284,6.5280004,5.5269747,3.367385,1.8182565,1.785436,0.5677949,0.13784617,0.13456412,0.3249231,0.6301539,0.52512825,0.5973334,0.7122052,0.764718,0.67282057,0.764718,0.8730257,0.77128214,0.5152821,0.446359,0.57764107,0.7089231,0.79097444,0.81394875,0.8041026,0.69251287,0.6629744,0.67610264,0.69907695,0.73517954,0.3314872,0.108307704,0.013128206,0.0,0.0,0.0032820515,0.036102567,0.072205134,0.118153855,0.20348719,0.36430773,0.5284103,0.67282057,0.77128214,0.78769237,0.77128214,0.86974365,0.86646163,0.82379496,1.086359,1.1520001,1.1060513,1.1224617,1.1520001,0.9353847,0.9321026,0.9517949,1.0043077,1.0929232,1.2340513,1.1520001,1.4703591,1.8281027,2.0184617,1.9593848,2.034872,1.8970258,1.7132308,1.6147693,1.6738462,2.2646155,2.3236926,2.3991797,2.6453335,2.8521028,2.9472823,2.865231,2.6617439,2.5304618,2.8389745,3.8728209,4.1747694,4.332308,4.71959,5.5105643,6.5969234,7.6242056,8.421744,8.802463,8.553026,7.2927184,6.5247183,5.664821,4.7294364,4.33559,3.3247182,2.7700515,2.8389745,3.2328207,3.2032824,3.131077,3.242667,3.3509746,3.636513,4.6539493,5.1364107,5.677949,6.262154,6.672411,6.5017443,6.675693,7.2992826,8.109949,8.956718,9.816616,9.517949,9.317744,9.163487,8.92718,8.39877,7.683283,7.5618467,8.395488,9.596719,9.655796,8.726975,9.07159,9.603283,9.616411,8.792616,7.7948723,7.204103,6.8627696,6.8594875,7.512616,7.9786673,7.5552826,7.1548724,7.3058467,8.149334,7.7948723,7.4469748,6.5411286,5.398975,5.21518,4.5817437,4.4865646,4.4045134,4.135385,3.8104618,4.0008206,3.9778464,4.0467696,4.263385,4.4373336,4.128821,4.3749747,4.637539,4.818052,5.2414365,5.2020516,4.8705645,4.818052,5.0543594,5.037949,4.893539,4.818052,4.896821,5.0116925,4.84759,4.5128207,4.135385,3.9122055,3.8531284,3.7940516,3.7874875,3.5249233,3.2000003,2.8455386,2.3401027,2.3860514,2.4418464,2.3368206,2.166154,2.3171284,2.7109745,2.7798977,2.5435898,2.1070771,1.6804104,0.34133336,0.17394873,0.08205129,0.036102567,0.02297436,0.059076928,0.101743594,0.29538465,0.41025645,0.37743592,0.28225642,0.118153855,0.052512825,0.21989745,0.57764107,0.9124103,2.8553848,3.2787695,2.2350771,0.6629744,0.37743592,0.7384616,0.71548724,0.6104616,0.57764107,0.62030774,0.77456415,1.0732309,1.6607181,2.5895386,3.820308,3.2196925,2.6715899,2.477949,2.3958976,1.6475899,1.1454359,1.1224617,1.3193847,1.6344616,2.1267693,4.2141542,5.654975,6.813539,8.077128,9.852718,9.944616,8.310155,5.8781543,3.6168208,2.5435898,2.3105643,2.2580514,2.802872,4.0369234,5.76,7.706257,9.344001,10.489437,10.975181,10.65354,11.992617,13.266052,14.621539,16.505438,19.6759,23.269745,26.551796,29.971695,34.756927,42.919388,53.24144,74.65026,103.57826,129.408,134.50504,105.73457,76.45867,55.46667,45.134773,41.4359,43.565952,46.41149,52.801643,62.35898,71.49621,82.52062,83.63324,72.96985,57.30462,52.03036,67.49211,78.34914,66.563286,35.987694,12.347078,11.437949,10.223591,8.687591,7.6209235,8.618668,9.734565,9.202872,7.4174366,5.5926156,5.786257,5.943795,5.7665644,5.98318,6.518154,6.5050263,7.456821,7.0334363,6.987488,8.267488,11.024411,14.55918,16.640001,19.498669,23.896618,29.121643,32.078773,30.972721,26.883284,22.042257,19.849848,15.750566,18.021746,20.066463,20.112411,21.195488,24.920618,26.469746,22.055386,14.401642,12.731078,11.542975,9.816616,8.868103,8.917334,9.107693,10.925949,9.547488,7.722667,6.449231,4.9788723,5.074052,8.562873,9.787078,7.6143594,5.431795,4.785231,4.706462,5.179077,6.121026,7.3550773,6.547693,8.172308,8.838565,8.231385,9.117539,11.011283,9.856001,8.87795,9.449026,11.1064625,14.395078,17.716515,18.048002,16.12472,16.420103,14.293334,12.356924,11.378873,11.628308,12.875488,13.075693,12.0549755,10.364718,8.891078,8.851693,8.553026,8.818872,8.740103,8.507077,9.412924,10.322052,11.592206,11.703795,10.541949,9.370257,7.79159,7.896616,8.123077,8.129642,8.792616,7.8769236,6.8529234,6.3376417,6.442667,6.764308,7.9425645,8.87795,9.042052,8.687591,8.848411,10.676514,11.323078,10.512411,9.042052,8.792616,7.0137444,6.2490263,6.2096415,5.835488,3.2951798,5.0149746,5.2578464,4.9427695,4.588308,4.322462,2.7470772,2.0184617,1.9528207,2.409026,3.3017437,2.9965131,2.5764105,3.2787695,5.5762057,9.173334,7.3452315,8.51036,9.826463,10.66995,12.652308,12.99036,13.551591,19.163898,25.91508,21.139694,22.79713,19.331284,14.953027,11.739899,9.636104,7.1680007,7.02359,6.8365135,5.858462,4.9427695,4.95918,4.8114877,4.7491283,5.1265645,6.422975,8.103385,6.6494365,4.338872,2.665026,2.349949,1.9265642,1.3193847,0.761436,0.79097444,2.2744617,2.412308,5.723898,11.264001,15.415796,11.910565,6.3868723,4.0402055,6.997334,11.657847,8.697436,5.6418467,8.080411,13.499078,16.118155,6.885744,9.051898,12.071385,22.478771,30.742977,11.273847,10.857026,8.805744,13.443283,20.54236,13.3251295,12.714667,10.384411,9.83959,11.319796,11.779283,9.980719,7.3583593,5.904411,5.142975,2.1300514,7.2894363,17.417847,26.656822,26.397541,5.280821,14.158771,14.907078,9.957745,5.3202057,10.594462,12.416001,19.889233,19.994259,12.356924,9.245539,3.0358977,1.7526156,1.7985642,2.0020514,3.629949,1.6902566,1.3981539,1.7985642,2.2416413,2.3991797,1.5392822,1.595077,2.3204105,2.986667,2.3762052,2.0053334,1.5064616,1.2570257,1.1618463,0.67282057,1.9167181,4.4110775,5.6385646,5.0182567,3.9056413,2.284308,2.5435898,2.789744,2.4484105,2.2613335,2.15959,2.162872,1.9265642,1.5195899,1.4178462,1.5556924,1.7723079,2.044718,2.3335385,2.5895386,1.9889232,1.7952822,1.3292309,0.65969235,0.58092314,0.37415388,0.45620516,0.67610264,0.96492314,1.3292309,0.6301539,0.42338464,0.47917953,0.5973334,0.6071795,0.6892308,0.53825647,0.36102566,0.2855385,0.36430773,0.69251287,2.0775387,2.6880002,2.0808206,1.1815386,1.2537436,1.0568206,1.0404103,1.1716924,0.92225647,0.8730257,0.7253334,0.65312827,0.63343596,0.45292312,0.55794877,0.5907693,0.5677949,0.5513847,0.6170257,0.64000005,0.51856416,0.48246157,0.5907693,0.7253334,1.4080001,1.7132308,1.6082052,1.2668719,1.0699488,1.2504616,1.1027694,1.1290257,1.657436,2.8356924,2.3105643,2.1497438,2.4418464,2.6847181,1.785436,2.540308,2.3302567,1.7788719,1.3751796,1.4736412,1.1388719,1.0404103,1.273436,1.529436,1.0929232,0.86317956,0.79425645,0.7122052,0.64000005,0.77456415,1.2865642,1.1355898,0.94523084,0.9353847,0.88615394,0.90256417,0.7581539,0.6826667,0.6662565,0.47589746,0.5349744,0.48246157,0.380718,0.3708718,0.6629744,0.7844103,0.8041026,0.6104616,0.30194873,0.19364104,0.0951795,0.055794876,0.098461546,0.16738462,0.14112821,0.0951795,0.052512825,0.072205134,0.90584624,4.013949,3.82359,3.4002054,3.1770258,3.190154,3.0818465,2.231795,3.3509746,4.420923,4.017231,1.3062565,1.591795,2.7044106,2.8324106,1.7394873,0.76800007,0.33805132,0.13784617,0.10502565,0.18707694,0.318359,0.36758977,0.3708718,0.38728207,0.46933338,0.63343596,0.5973334,0.64000005,0.6235898,0.56451285,0.60389745,0.6268718,0.60061544,0.6235898,0.7220513,0.8467693,1.142154,1.3686155,1.6836925,2.0676925,2.3368206,2.6518977,2.4681027,2.2744617,2.7306669,4.6802053,5.346462,6.9152827,6.8365135,5.074052,4.0992823,6.12759,5.097026,3.3214362,2.1070771,1.7296412,0.5218462,0.1148718,0.068923086,0.19364104,0.5349744,0.64000005,0.6235898,0.69251287,0.827077,0.7811283,0.6892308,0.7187693,0.7220513,0.6498462,0.55794877,0.56451285,0.6465641,0.7778462,0.8992821,0.92553854,0.73517954,0.6662565,0.67282057,0.67610264,0.5677949,0.27569234,0.08861539,0.006564103,0.0,0.0,0.013128206,0.036102567,0.07548718,0.13784617,0.23958977,0.42994875,0.65641034,0.7778462,0.7778462,0.7515898,0.80738467,0.92225647,0.9288206,0.8730257,1.0305642,1.0765129,1.079795,1.1224617,1.142154,0.8992821,0.8795898,0.8795898,1.017436,1.2307693,1.2537436,1.211077,1.2800001,1.4441026,1.6640002,1.8904617,1.8674873,1.7033848,1.6049232,1.5786668,1.4506668,1.8149745,1.9003079,2.2383592,2.802872,3.0227695,3.006359,2.8717952,2.5435898,2.2777438,2.6847181,3.9253337,4.2272825,4.315898,4.7556925,5.9569235,6.8693337,7.7948723,8.579283,8.914052,8.339693,7.7456417,6.99077,5.927385,4.8804107,4.644103,3.495385,2.793026,2.7044106,2.9636924,2.8882053,2.7470772,2.8422565,2.7536411,2.681436,3.436308,3.95159,4.31918,5.0084105,5.7731285,5.6287184,6.1538467,6.8266673,7.207385,7.4404106,8.260923,8.664616,8.267488,7.6635904,7.243488,7.200821,7.177847,7.496206,8.595693,9.96759,10.164514,9.019077,8.900924,9.199591,9.45559,9.353847,8.395488,7.9228725,7.5388722,7.204103,7.2303596,8.474257,7.8736415,7.0793853,6.889026,7.2664623,6.921847,6.262154,5.47118,4.8738465,4.9329233,4.562052,4.1550775,3.7185643,3.3772311,3.3805132,3.9253337,3.95159,4.073026,4.378257,4.420923,4.1452312,4.4767184,4.8836927,5.149539,5.349744,5.221744,4.7491283,4.46359,4.4964104,4.6145644,4.46359,4.644103,4.9329233,5.152821,5.175795,4.634257,4.3027697,4.2207184,4.2272825,3.9778464,3.5872824,3.2032824,2.7470772,2.3401027,2.2908719,2.4582565,2.3204105,2.103795,1.9954873,2.162872,2.2908719,2.4713848,2.4024618,2.1366155,2.1103592,0.6104616,0.256,0.07548718,0.016410258,0.02297436,0.04594872,0.02297436,0.006564103,0.06564103,0.18707694,0.25928208,0.16082053,0.09189744,0.049230773,0.08205129,0.28882053,2.3401027,2.4976413,2.2350771,1.9528207,0.97805136,1.270154,0.88615394,0.7515898,1.020718,1.083077,1.8510771,2.281026,2.5140514,2.5140514,2.0742567,3.2229745,3.564308,3.498667,3.0260515,1.7690258,1.2077949,1.1881026,1.5097437,2.225231,3.6168208,6.1440005,7.781744,8.569437,8.923898,9.642668,9.179898,7.2237954,5.044513,3.4133337,2.5928206,2.4484105,3.0326157,5.2315903,8.264206,9.705027,7.460103,6.6494365,7.4929237,9.212719,10.056206,12.849232,14.979283,17.060104,19.908924,24.536617,28.245335,31.67508,36.148514,43.139286,54.258877,70.468925,96.67611,131.4396,159.88185,153.7313,108.50462,82.14647,66.93088,58.587902,56.303593,61.83385,70.40985,83.68575,99.10811,109.9356,107.58237,84.45375,61.46298,50.95713,56.717133,52.676926,44.143593,31.783386,18.819284,11.017847,10.272821,9.435898,8.201847,7.4108725,9.032206,8.070564,6.3442054,4.9526157,4.2371287,3.7842054,4.713026,4.788513,5.110154,5.8223596,6.1046157,7.7259493,7.75877,8.500513,10.354873,11.795693,19.252514,23.781746,25.550772,26.194054,28.793438,26.328617,19.945026,17.434258,20.535797,24.917336,16.810667,21.451488,25.110977,25.238976,30.424618,34.54031,27.155695,18.225233,13.525334,14.647796,14.073437,11.661129,9.324308,8.3134365,9.216001,9.521232,8.388924,7.9327188,7.6274877,4.31918,3.7316926,4.565334,4.926359,4.2240005,3.1737437,3.2098465,4.1813335,5.333334,5.976616,5.4613338,5.976616,6.954667,7.8080006,8.448001,9.278359,9.852718,9.691898,9.632821,10.410667,12.678565,15.80636,17.867489,17.59836,15.714462,14.907078,12.662155,11.861334,12.806565,14.7790785,16.036104,17.135592,16.239592,13.131488,9.43918,8.621949,9.609847,10.315488,10.289231,9.777231,9.705027,11.864616,12.340514,11.027693,9.481847,10.909539,10.19077,9.800206,8.976411,8.034462,8.375795,9.511385,8.717129,7.781744,7.2172313,6.242462,6.948103,7.6931286,8.274052,8.602257,8.713847,10.397539,11.277129,11.122872,10.463181,10.57477,7.3025646,6.419693,6.36718,5.5663595,2.4418464,4.197744,5.024821,5.474462,5.481026,4.332308,2.5632823,2.2121027,2.5600002,2.802872,2.044718,2.9111798,4.70318,6.7282057,10.771693,21.087181,15.947489,12.018872,9.337437,9.258667,14.434463,17.742771,16.984617,18.267899,20.466873,15.24513,11.37559,10.305642,10.8996935,11.907283,11.992617,9.990565,8.89436,7.5520005,6.0685134,5.799385,6.2129235,5.786257,5.1265645,4.824616,5.4482055,9.69518,9.449026,6.629744,3.508513,2.7175386,2.0086155,1.3456411,0.86974365,0.761436,1.2373334,3.8859491,7.6767187,14.739694,20.54236,13.899488,11.286975,5.7632823,4.57518,7.75877,8.149334,4.8771286,3.2984617,2.6157951,2.809436,4.637539,8.057437,11.585642,16.66954,19.75795,12.297847,14.605129,12.711386,11.946668,13.105232,12.419283,7.709539,5.937231,5.5630774,6.419693,9.705027,20.201027,13.167591,4.673641,1.5195899,1.2504616,5.218462,6.23918,13.472821,20.050053,3.0818465,12.95754,18.87836,14.628103,5.5663595,8.605539,12.57354,9.875693,7.965539,8.257642,6.1341543,1.7887181,1.1782565,2.6978464,4.460308,4.3027697,1.5327181,1.2603078,1.6377437,1.7887181,1.8018463,1.020718,1.079795,1.6344616,2.1825643,2.0611284,2.681436,2.3269746,1.7755898,1.394872,1.1126155,1.8084104,2.6518977,2.9997952,2.868513,2.930872,2.3926156,2.2121027,2.4681027,2.8356924,2.5796926,2.5173335,2.228513,1.8740515,1.5163078,1.1126155,1.5524104,2.2383592,2.5764105,2.3433847,1.7099489,1.7460514,3.2098465,3.1376412,1.4703591,1.0666667,0.38400003,0.47917953,0.8205129,1.0010257,0.7318975,0.45292312,0.446359,0.7253334,1.0962052,1.1454359,1.2537436,0.86974365,0.5940513,0.6071795,0.65641034,0.88943595,2.2547693,3.4330258,3.5610259,2.2416413,1.4375386,0.88943595,0.81394875,1.0075898,0.82379496,1.020718,0.9124103,0.86317956,0.8533334,0.48902568,0.4397949,0.51856416,0.5874872,0.6170257,0.702359,0.5677949,0.4135385,0.4135385,0.54482055,0.58092314,0.71548724,1.4244103,1.9987694,1.9626669,1.083077,0.81394875,0.8402052,1.0469744,1.6016412,2.9440002,2.4188719,2.03159,2.228513,2.809436,2.9440002,2.9571285,2.6486156,2.2646155,1.9265642,1.6311796,1.2800001,1.2635899,1.4276924,1.5195899,1.1913847,1.1158975,1.1815386,1.1520001,0.88615394,0.33476925,0.45620516,0.6170257,0.7253334,0.71548724,0.51856416,0.36102566,0.27569234,0.32820517,0.46276927,0.48902568,0.29210258,0.23630771,0.24615386,0.32164106,0.5021539,0.9189744,0.79425645,0.50543594,0.28882053,0.2297436,0.18051283,0.10502565,0.06564103,0.07876924,0.09189744,0.10502565,0.068923086,0.06564103,0.37415388,1.5097437,2.5600002,3.3280003,3.1376412,2.0086155,0.64000005,1.1651284,3.7152824,4.5062566,2.9046156,1.404718,2.3926156,1.9068719,1.5458462,1.8051283,2.0742567,1.1946667,0.46276927,0.08533334,0.06235898,0.18379489,0.28225642,0.29538465,0.27241027,0.29210258,0.48902568,0.5973334,0.65312827,0.6104616,0.51856416,0.51856416,0.5316923,0.45292312,0.4266667,0.5415385,0.80738467,1.1257436,1.270154,1.2996924,1.4473847,2.1070771,2.9472823,2.802872,2.2153847,1.7033848,1.7394873,6.0356927,5.297231,4.4996924,5.037949,4.7458467,6.1505647,6.2063594,4.8344617,2.681436,1.1454359,0.5218462,0.16410258,0.04266667,0.13128206,0.4135385,0.88943595,0.7975385,0.6071795,0.56123084,0.67282057,0.5973334,0.5874872,0.67938465,0.79097444,0.7187693,0.5940513,0.74830776,0.86974365,0.81394875,0.5940513,0.58420515,0.7253334,0.90256417,0.92225647,0.51856416,0.22646156,0.06235898,0.0,0.0,0.0,0.013128206,0.04266667,0.09189744,0.17723078,0.33476925,0.5546667,0.5546667,0.46276927,0.46933338,0.82379496,0.95835906,0.88287187,0.80738467,0.78769237,0.702359,0.78769237,0.9353847,1.0896411,1.1323078,0.8992821,0.98461545,0.92553854,1.017436,1.204513,1.083077,1.3029745,1.3587693,1.467077,1.6213335,1.5721027,1.3653334,1.3292309,1.3686155,1.401436,1.3883078,1.3522053,1.3620514,1.654154,2.3269746,3.3411283,3.0490258,2.5895386,2.3105643,2.2711797,2.2580514,2.7963078,2.993231,3.2623591,3.8564105,4.8836927,6.554257,6.99077,6.889026,6.692103,6.6067696,7.1089234,7.003898,6.4000006,5.474462,4.4865646,3.8137438,3.190154,2.7864618,2.6551797,2.7175386,2.605949,2.4155898,2.2908719,2.300718,2.412308,2.1530259,2.7306669,3.7218463,4.772103,5.61559,5.4580517,5.1331286,4.9132314,5.024821,5.661539,7.0892315,7.748924,7.7292314,7.460103,7.6898465,7.6176414,7.8637953,8.4512825,9.127385,9.383386,8.933744,8.152616,7.522462,7.5454364,8.743385,8.779488,7.9195905,7.466667,7.6701546,7.706257,8.756514,7.899898,6.7544622,6.1078978,5.937231,5.3366156,4.59159,4.2272825,4.309334,4.457026,4.457026,4.0336413,3.7054362,3.5872824,3.4166157,3.7973337,3.9909747,4.210872,4.4110775,4.2863593,4.312616,5.0051284,5.687795,5.9470773,5.6320004,5.32677,4.781949,4.414359,4.3585644,4.457026,4.578462,4.97559,5.3694363,5.5302567,5.2480006,4.785231,4.650667,4.673641,4.6244106,4.197744,3.7087183,3.1474874,2.7306669,2.5238976,2.425436,2.6715899,2.5764105,2.3630772,2.2744617,2.5796926,2.6289232,2.9144619,2.8291285,2.353231,2.0611284,0.49887183,0.17723078,0.06235898,0.026256412,0.0032820515,0.009846155,0.0032820515,0.009846155,0.03938462,0.07548718,0.052512825,0.09189744,0.08533334,0.072205134,0.108307704,0.27897438,1.8215386,2.5731285,2.540308,2.1924105,2.4648206,3.1015387,2.048,1.3128207,1.4539489,1.585231,1.785436,2.097231,2.1825643,1.9987694,1.7952822,2.865231,3.370667,3.5741541,3.7218463,4.017231,3.501949,3.0194874,2.9505644,3.5347695,4.8377438,6.885744,7.312411,7.069539,6.9152827,7.4207187,6.997334,5.8486156,4.781949,4.1878977,4.0336413,4.161641,4.969026,5.8978467,6.738052,7.640616,7.6898465,8.664616,9.69518,10.581334,11.762873,13.35795,15.845745,19.236105,23.09908,26.574772,30.880823,35.649643,42.049644,53.14626,73.92493,100.60144,136.51694,181.6156,65535.0,195.4035,148.98544,127.300934,111.786674,97.72308,94.24083,99.29191,105.89211,112.01314,112.41026,98.599396,82.77991,66.77006,60.70154,70.19324,96.37416,76.22237,45.702568,23.61436,14.729847,9.770667,7.962257,6.941539,6.695385,7.39118,9.386667,9.127385,7.430565,5.284103,3.5544617,3.0162053,4.332308,4.7360005,5.605744,6.931693,7.2992826,7.6734366,8.444718,10.112,12.665437,15.589745,22.367182,22.81354,20.187899,19.186872,25.938053,26.880003,21.851898,18.546873,18.582975,17.496616,14.811898,19.140924,25.219284,30.129232,33.30626,28.836105,19.459284,13.226667,12.310975,13.013334,11.959796,10.348309,8.953437,8.152616,7.9228725,8.257642,8.4283085,7.716103,6.157129,4.5390773,4.2535386,3.882667,3.7251284,3.748103,3.5774362,3.31159,3.0982566,3.2098465,3.570872,3.7907696,4.585026,5.87159,7.273026,8.297027,8.3364105,9.360411,10.6469755,12.442257,14.431181,15.744001,16.485744,15.465027,13.423591,11.401847,10.732308,9.990565,12.527591,16.548103,19.377232,17.45395,18.074257,16.712206,13.850258,11.073642,11.08677,13.958565,14.381949,13.138052,11.510155,11.290257,12.796719,11.720206,11.441232,12.343796,11.789129,11.244308,10.075898,9.179898,8.937026,9.232411,10.581334,9.472001,7.962257,6.944821,6.1538467,6.6100516,7.128616,7.827693,8.54318,8.848411,10.561642,10.948924,11.008,10.998155,10.453334,7.6898465,7.525744,7.515898,6.242462,3.3312824,3.7316926,4.194462,4.778667,5.1232824,4.4438977,2.8192823,2.1464617,2.041436,2.2219489,2.5206156,4.9099493,5.5072823,6.885744,9.810052,13.239796,13.909334,14.677335,12.803283,10.049642,12.678565,12.859077,15.497848,18.271181,20.12554,21.248001,20.007385,23.77518,29.35795,32.52513,28.018873,22.71836,18.796309,16.042667,12.895181,6.445949,6.5280004,6.442667,6.242462,5.7534366,4.568616,7.430565,7.8769236,5.933949,3.0030773,1.8379488,2.7306669,2.169436,1.4572309,1.2077949,1.3226668,3.2853336,4.6244106,7.4240007,12.63918,20.089437,19.643078,13.351386,7.181129,4.4274874,5.7074876,3.9680004,3.8137438,4.073026,4.1222568,3.882667,5.874872,6.7085133,11.510155,18.070976,16.850052,9.734565,6.560821,5.408821,5.674667,8.073847,5.9602056,5.7731285,6.0028725,6.3310776,7.640616,10.581334,14.532925,14.372104,9.357129,3.1442053,3.4002054,5.1167183,8.795898,10.886565,3.8038976,6.5411286,11.533129,13.190565,10.079181,4.896821,16.272411,12.816411,8.736821,7.5585647,2.1070771,0.90584624,1.4309745,2.1956925,2.428718,2.0939488,2.4484105,2.1530259,1.8313848,1.6902566,1.5064616,1.6443079,1.9495386,2.1333334,1.9954873,1.4145643,1.9265642,1.9331284,1.8609232,1.8445129,1.7001027,2.1136413,2.100513,1.7394873,1.4900514,2.1858463,2.537026,2.1169233,2.172718,2.7995899,2.934154,4.46359,4.571898,3.7743592,2.5993848,1.5885129,1.2471796,1.276718,1.3587693,1.3686155,1.3784616,1.6114873,1.8740515,1.7066668,1.211077,1.0305642,0.5349744,0.5513847,0.6235898,0.7417436,1.3423591,1.7460514,1.7920002,1.7624617,1.6836925,1.3522053,1.6475899,1.3817437,1.211077,1.3095386,1.3751796,2.349949,2.9735386,3.1737437,3.1343591,3.2820516,1.8904617,0.9288206,0.636718,0.764718,0.5907693,0.62030774,0.54482055,0.5218462,0.5677949,0.56123084,0.44307697,0.43323082,0.43651286,0.43651286,0.48246157,0.43651286,0.42338464,0.49887183,0.58420515,0.446359,0.47261542,0.7187693,1.1290257,1.4605129,1.2537436,0.7515898,0.7187693,0.88943595,1.211077,1.8215386,1.8937438,1.6607181,1.5721027,1.7723079,2.103795,2.4681027,2.422154,2.4976413,2.806154,3.062154,2.228513,2.041436,1.9790771,1.654154,0.8369231,0.6662565,0.6695385,0.8533334,0.9944616,0.64000005,0.6071795,0.5152821,0.5021539,0.5349744,0.41025645,0.28882053,0.3314872,0.37743592,0.37743592,0.39056414,0.21333335,0.13128206,0.10502565,0.13128206,0.24615386,0.50543594,0.42994875,0.26584616,0.16082053,0.16738462,0.15753847,0.1148718,0.07548718,0.059076928,0.04266667,0.04594872,0.029538464,0.029538464,0.11158975,0.38728207,0.8336411,2.1070771,3.0490258,2.7109745,0.34789747,0.58092314,2.3958976,2.6518977,1.211077,0.93866676,1.0108719,1.079795,1.024,0.9189744,1.0633847,0.827077,0.48246157,0.19692309,0.055794876,0.06235898,0.128,0.16738462,0.17723078,0.18707694,0.256,0.36758977,0.42994875,0.44307697,0.4397949,0.45620516,0.51856416,0.4955898,0.446359,0.45292312,0.61374366,0.8336411,1.0929232,1.3062565,1.6082052,2.3269746,2.8947694,3.1409233,2.802872,2.0873847,1.654154,3.1770258,4.6605134,5.549949,5.474462,4.2338467,5.1298466,5.937231,5.35959,3.3444104,1.083077,0.29538465,0.049230773,0.01969231,0.07548718,0.27897438,0.83035904,0.86974365,0.7384616,0.64000005,0.6235898,0.67610264,0.65641034,0.6892308,0.77128214,0.764718,0.6432821,0.6662565,0.7122052,0.7384616,0.75487185,0.63343596,0.6268718,0.6629744,0.65969235,0.5316923,0.26584616,0.08861539,0.006564103,0.0,0.0,0.02297436,0.06235898,0.10502565,0.16410258,0.27569234,0.48574364,0.62030774,0.67282057,0.71548724,0.92225647,0.93866676,0.86317956,0.7844103,0.7384616,0.702359,0.7384616,0.73517954,0.8369231,0.9517949,0.7778462,0.9911796,1.1881026,1.3915899,1.5688206,1.6311796,1.4802053,1.2176411,1.2537436,1.529436,1.5097437,1.4211283,1.4834872,1.5031796,1.404718,1.2176411,1.2406155,1.4605129,1.7624617,2.1169233,2.5731285,2.484513,2.1530259,1.9889232,2.097231,2.2711797,2.8356924,3.3345644,3.876103,4.4832826,5.077334,6.1538467,6.6560006,6.5444107,6.052103,5.654975,5.3366156,5.0838976,4.919795,4.7228723,4.240411,3.308308,2.6584618,2.3105643,2.1924105,2.1530259,1.9856411,1.8674873,1.910154,2.1530259,2.5435898,2.4057438,2.4418464,2.917744,3.817026,4.8344617,4.9394875,5.179077,5.586052,5.976616,5.9667697,6.416411,6.5312824,6.6592827,6.99077,7.5552826,7.0826674,7.069539,7.5191803,8.103385,8.1755905,7.9097443,7.512616,7.181129,7.2336416,8.096821,7.830975,7.3616414,7.0925136,7.1844106,7.571693,7.6635904,7.3386674,6.675693,5.8157954,4.972308,4.3060517,3.9548721,3.9187696,4.082872,4.210872,4.269949,4.4274874,4.309334,3.9220517,3.6758976,3.9548721,4.1124105,4.1025643,4.0434875,4.2141542,4.562052,5.1364107,5.6352825,5.87159,5.789539,5.3858466,5.0084105,4.7556925,4.6933336,4.857436,5.0871797,5.861744,6.4557953,6.4656415,5.8223596,4.8705645,4.3290257,4.089436,3.9778464,3.7448208,3.3345644,2.8816411,2.3958976,2.0676925,2.2416413,2.556718,2.4713848,2.3991797,2.553436,2.9571285,2.868513,2.6912823,2.537026,2.4451284,2.3762052,0.22646156,0.1148718,0.06564103,0.036102567,0.006564103,0.0,0.006564103,0.006564103,0.016410258,0.026256412,0.0,0.036102567,0.059076928,0.07876924,0.118153855,0.21989745,0.9911796,2.0250258,2.8750772,3.3017437,3.259077,2.9768207,2.3893335,2.359795,2.7273848,2.3040001,2.3368206,2.1366155,1.7985642,1.5031796,1.5425643,2.349949,3.1048207,3.8432825,4.453744,4.670359,3.764513,3.0490258,2.802872,3.2229745,4.4110775,5.2480006,5.428513,5.3760004,5.405539,5.7403083,5.8814363,5.674667,5.421949,5.4153852,5.933949,6.3540516,7.141744,7.7259493,8.375795,10.230155,11.1064625,11.575796,11.828514,11.959796,11.953232,13.321847,16.361027,21.251284,27.16554,32.246155,36.240414,41.34072,48.295387,61.052723,86.78729,115.403496,146.67488,181.20863,203.56268,182.27202,145.22421,126.037346,111.83919,99.66277,96.452934,98.10052,95.69478,93.25949,88.75652,74.0956,65.253746,60.52431,66.08739,82.37293,104.05744,78.50011,46.94975,26.249847,19.065437,13.873232,11.805539,10.95877,10.233437,9.225847,8.231385,7.177847,5.832206,4.5029745,3.6791797,4.0041027,5.031385,6.088206,7.4010262,8.54318,8.41518,9.347282,9.8363085,10.469745,12.73436,19.012924,25.718155,24.346258,20.115694,17.532719,20.407797,23.571693,24.070566,23.476515,22.28513,19.93518,21.641848,27.59549,32.961643,34.93416,32.735184,26.463182,18.343386,13.328411,12.038565,10.755282,9.67877,8.996103,8.776206,8.438154,6.747898,5.989744,7.6734366,7.9458466,6.488616,6.514872,6.160411,4.7589746,3.446154,2.8258464,2.9538465,2.8389745,2.3991797,2.2547693,2.546872,2.9407182,3.4658465,4.59159,6.009436,7.3025646,7.965539,9.225847,12.481642,15.688207,17.42113,16.886156,15.488001,13.889642,11.71036,9.472001,8.582564,10.118565,14.683899,19.091694,21.205336,19.948309,20.558771,18.582975,15.619284,13.426873,13.909334,15.218873,14.368821,12.448821,11.08677,12.458668,13.938873,13.929027,14.01436,13.965129,11.74318,10.94236,10.295795,9.668923,9.3078985,9.865847,10.348309,9.078155,7.716103,6.8004107,5.7403083,6.0652313,6.9087186,7.6209235,8.169026,9.137232,10.843898,11.286975,11.080206,10.436924,9.156924,7.4075904,7.3550773,7.3025646,6.2916927,4.132103,3.9876926,4.4832826,4.706462,4.352,3.748103,3.062154,2.2416413,1.6968206,1.5885129,1.8445129,4.827898,5.156103,6.5378466,9.278359,10.305642,16.075489,17.972515,16.580925,13.833847,13.026463,11.319796,15.028514,16.512001,16.239592,22.787283,26.207182,32.259285,36.197746,36.128822,33.027283,24.65149,18.858667,15.78995,13.820719,9.544206,7.4863596,6.7216415,6.75118,6.3868723,3.7185643,4.9296412,5.3103595,4.197744,2.2350771,1.3784616,3.2229745,4.46359,3.8465643,2.034872,1.6278975,3.9614363,5.2381544,7.1614366,10.154668,13.351386,15.91795,14.486976,9.281642,3.8596926,5.1331286,3.5446157,3.1803079,3.5905645,4.092718,3.7743592,4.1878977,3.8400004,6.0291286,10.390975,12.901745,16.705643,19.659489,18.435284,12.918155,6.229334,4.4045134,4.9362054,10.79795,15.698052,4.086154,6.688821,10.505847,13.656616,14.785643,13.082257,4.604718,5.3169236,7.8441033,8.549745,7.5520005,5.07077,9.91836,13.568001,11.881026,5.110154,11.949949,12.865642,9.977437,5.4416413,1.4473847,0.6301539,0.82379496,1.1093334,1.2865642,1.8970258,3.0194874,2.5304618,1.8248206,1.5458462,1.6082052,1.8510771,1.9265642,2.0939488,2.3269746,2.3040001,2.0611284,1.7624617,1.7723079,2.166154,2.7536411,2.6683078,1.8707694,1.0765129,0.75487185,1.1093334,2.1300514,2.3302567,2.1497438,2.041436,2.4713848,4.9854364,5.7796926,4.7622566,2.858667,2.028308,1.529436,1.2898463,1.2603078,1.3062565,1.214359,1.1224617,1.086359,1.1158975,1.1257436,0.95835906,0.5940513,0.58092314,0.8566154,1.3981539,2.2088206,2.6354873,2.297436,1.9889232,1.972513,2.0086155,2.5928206,2.7963078,2.7142565,2.5862565,2.7831798,2.537026,2.172718,1.9003079,1.9462565,2.5337439,1.4769232,0.7417436,0.44964105,0.4660513,0.36102566,0.34789747,0.2855385,0.26584616,0.30194873,0.3511795,0.318359,0.33476925,0.36758977,0.4004103,0.4004103,0.4135385,0.4266667,0.50543594,0.574359,0.4201026,0.318359,0.4201026,0.7122052,1.1848207,1.8379488,1.2012309,0.9419488,0.8402052,0.8041026,0.8730257,1.1060513,1.1716924,1.1520001,1.1552821,1.3161026,1.7460514,1.8543591,2.0808206,2.4582565,2.6223593,2.3072822,2.353231,2.1497438,1.4736412,0.48246157,0.36758977,0.35446155,0.5021539,0.69907695,0.6432821,0.67938465,0.69907695,0.67282057,0.5907693,0.47261542,0.52512825,0.7581539,0.7975385,0.5973334,0.44964105,0.32164106,0.28225642,0.24287182,0.18051283,0.14769232,0.256,0.24615386,0.20676924,0.17066668,0.108307704,0.1148718,0.11158975,0.10502565,0.09189744,0.06564103,0.04594872,0.036102567,0.04594872,0.068923086,0.07876924,0.18051283,0.77128214,1.4309745,1.595077,0.55794877,0.37415388,1.0404103,1.1651284,0.6235898,0.5481026,0.40369233,0.47917953,0.47917953,0.41025645,0.571077,0.512,0.35774362,0.27241027,0.24943592,0.0951795,0.08205129,0.09189744,0.10502565,0.12471796,0.15097436,0.22646156,0.27569234,0.30194873,0.3249231,0.37743592,0.44307697,0.47261542,0.45292312,0.42994875,0.48246157,0.56123084,0.7581539,1.0502565,1.5031796,2.281026,2.7963078,3.2656412,3.2098465,2.6551797,2.1267693,2.028308,3.1474874,4.417641,5.1265645,4.900103,5.618872,6.2523084,5.658257,3.8695388,2.103795,0.7811283,0.19692309,0.016410258,0.032820515,0.14441027,0.6235898,0.7844103,0.77128214,0.702359,0.6826667,0.65969235,0.5907693,0.60061544,0.7450257,1.0075898,0.8205129,0.702359,0.6695385,0.69907695,0.72861546,0.65641034,0.98133343,1.3686155,1.4309745,0.7253334,0.36758977,0.13784617,0.026256412,0.0,0.0,0.02297436,0.08861539,0.14441027,0.18051283,0.23958977,0.4266667,0.6071795,0.7122052,0.7811283,0.9747693,0.81394875,0.7450257,0.764718,0.78769237,0.6465641,0.6498462,0.65969235,0.7581539,0.86317956,0.7187693,0.8336411,1.0994873,1.3522053,1.5819489,1.9626669,1.6443079,1.2996924,1.2176411,1.4211283,1.6410258,1.4769232,1.4998976,1.5360001,1.4998976,1.3751796,1.3259488,1.4309745,1.6508719,1.8904617,1.9856411,1.8773335,1.6508719,1.6147693,1.8838975,2.3827693,2.9505644,3.43959,3.8104618,4.092718,4.3684106,5.346462,5.98318,6.0061545,5.5696416,5.2611284,4.7655387,4.2601027,3.9023592,3.7021542,3.5413337,2.7667694,2.3335385,2.0906668,1.913436,1.719795,1.7493335,1.785436,1.9659488,2.2383592,2.349949,2.3204105,2.103795,2.3860514,3.18359,3.8498464,4.2568207,4.768821,5.3760004,5.8781543,5.868308,6.0258465,6.160411,6.121026,6.160411,6.944821,6.7314878,6.6822567,7.4075904,8.43159,8.185436,7.9786673,8.169026,8.267488,8.28718,8.740103,7.9524107,7.5191803,7.3452315,7.2927184,7.197539,6.340924,5.910975,5.6352825,5.2020516,4.2535386,3.9942567,3.9647183,3.9647183,3.9187696,3.8662567,4.128821,4.309334,4.1878977,3.8465643,3.6758976,3.7842054,3.8071797,3.7349746,3.7809234,4.3618464,4.7294364,5.031385,5.284103,5.402257,5.1889234,4.7983594,4.6900516,4.644103,4.634257,4.841026,5.3891287,6.3474874,7.059693,7.056411,6.0750775,4.8836927,3.9811285,3.5544617,3.4822567,3.3214362,2.9210258,2.4943593,2.162872,2.0020514,2.041436,2.349949,2.2678976,2.2449234,2.4746668,2.8947694,2.5993848,2.4713848,2.4418464,2.4418464,2.428718,0.055794876,0.068923086,0.06235898,0.04266667,0.016410258,0.0,0.013128206,0.006564103,0.0032820515,0.006564103,0.0,0.013128206,0.03938462,0.09189744,0.16410258,0.22646156,0.50543594,1.4276924,2.7536411,3.9056413,3.9778464,3.1409233,2.5731285,2.740513,3.2098465,2.6518977,2.6289232,2.5600002,2.2711797,1.8838975,1.8346668,2.428718,3.5216413,4.5522056,5.110154,4.926359,3.6332312,2.806154,2.3827693,2.4352822,3.1573336,3.4133337,3.6463592,3.95159,4.263385,4.3552823,5.3070774,5.858462,6.1013336,6.262154,6.701949,7.3714876,8.392206,9.110975,9.878975,12.048411,12.947693,13.243078,13.499078,13.4400015,11.936821,13.761642,18.7799,26.338463,34.192413,38.498463,39.781746,44.048412,50.691284,61.942158,82.85867,102.92513,118.40329,132.50955,139.47406,124.547295,103.68001,89.53436,79.54708,73.80678,75.067085,77.36452,72.3397,68.690056,67.01621,59.835083,57.235695,57.691902,65.68698,78.21129,84.76226,65.578674,45.052723,31.294361,24.822155,18.560001,16.137848,14.828309,14.04718,12.829539,9.849437,7.125334,5.3760004,4.4045134,4.522667,6.5378466,8.057437,9.301334,10.098872,10.358154,10.06277,10.6469755,10.57477,11.155693,14.36554,22.839796,26.568207,24.484104,20.457027,17.45395,17.54913,24.06072,29.417028,32.229748,32.036106,29.30872,30.67077,34.48123,35.83344,32.915695,26.98831,21.175797,16.039387,13.206975,11.989334,9.386667,8.297027,7.53559,7.4896417,7.5979495,6.373744,5.3727183,7.069539,8.119796,7.8145647,8.096821,8.743385,7.0334363,4.562052,2.6453335,2.3269746,2.2646155,2.100513,2.1136413,2.353231,2.6322052,2.8324106,3.7021542,4.903385,6.2851286,7.88677,10.331899,14.043899,16.853334,17.595078,16.134565,14.257232,12.553847,10.656821,9.140513,9.501539,13.942155,19.511797,22.656002,22.688822,21.822361,22.54113,19.990976,16.692514,14.516514,14.667488,14.139078,12.626052,11.280411,11.329642,14.063591,15.382976,15.560206,15.386257,14.5263605,11.500309,10.312206,9.609847,8.940309,8.549745,9.403078,9.3768215,8.310155,7.27959,6.5312824,5.464616,5.7468724,6.695385,7.394462,7.9097443,9.288206,10.843898,11.221334,10.71918,9.616411,8.169026,7.351795,7.13518,6.8332314,6.1538467,5.1889234,4.5423594,4.785231,4.4996924,3.5610259,3.1376412,3.0523078,2.4155898,1.6968206,1.2438976,1.2832822,3.4494362,4.644103,6.885744,9.67877,10.043077,18.432001,20.512821,19.442873,17.014154,13.666463,11.926975,15.133539,14.39836,11.195078,17.362053,25.4359,30.483694,31.540516,29.77149,28.478361,21.700924,16.400412,13.193847,11.923694,11.67754,8.310155,6.820103,6.560821,6.055385,2.9965131,3.3050258,5.979898,5.671385,2.349949,1.2996924,2.92759,5.435077,5.5926156,3.4002054,2.0841026,4.06318,5.868308,8.349539,10.289231,8.3823595,10.584617,14.408206,12.343796,5.799385,5.097026,4.5029745,3.9187696,3.9778464,4.33559,3.6529233,3.0358977,2.425436,2.740513,4.3684106,7.1876926,18.60595,25.363695,25.462156,20.608002,16.200207,6.180103,5.1200004,11.047385,15.222155,2.1398976,4.273231,5.602462,8.986258,13.312001,13.472821,4.8672824,5.602462,7.9163084,9.5835905,13.925745,7.466667,8.687591,13.656616,16.374155,8.772923,11.136001,12.153437,10.404103,6.432821,2.7470772,1.214359,0.8172308,0.7450257,1.0896411,2.8553848,3.2196925,3.117949,2.5764105,1.9003079,1.6869745,1.7723079,1.782154,1.972513,2.5009232,3.4264617,3.114667,2.412308,1.9922053,2.1530259,2.8389745,2.8422565,2.0808206,1.2373334,0.67610264,0.43323082,1.4408206,2.1431797,2.100513,1.7132308,2.2219489,3.764513,4.6244106,4.1747694,2.9013336,2.3893335,2.2121027,1.9593848,1.6344616,1.276718,0.9714873,0.7844103,0.81066674,0.92225647,0.9517949,0.71548724,0.5513847,0.7122052,1.273436,1.972513,2.1956925,2.356513,2.0709746,1.8740515,1.9626669,2.1956925,3.0851285,3.4658465,3.1934361,2.678154,2.9046156,1.9856411,1.2603078,0.9124103,1.0108719,1.5130258,0.9189744,0.54482055,0.38728207,0.36430773,0.29210258,0.318359,0.22646156,0.14769232,0.128,0.13784617,0.17066668,0.24287182,0.33476925,0.39384618,0.33805132,0.39056414,0.39712822,0.52512825,0.702359,0.5907693,0.30851284,0.38400003,0.6235898,1.0305642,1.8018463,1.2964103,0.92225647,0.636718,0.4266667,0.2986667,0.47917953,0.7187693,0.86974365,0.9189744,0.955077,1.6475899,1.6475899,1.5622566,1.591795,1.5163078,1.7132308,1.8674873,1.5983591,0.92553854,0.256,0.23958977,0.2231795,0.36102566,0.6235898,0.7975385,0.92553854,1.2668719,1.3489232,1.1224617,0.9353847,0.8566154,1.142154,1.3784616,1.2931283,0.761436,0.48574364,0.49887183,0.54482055,0.48246157,0.256,0.190359,0.2231795,0.28225642,0.27897438,0.08861539,0.13456412,0.15753847,0.14769232,0.118153855,0.10502565,0.06564103,0.059076928,0.06564103,0.07548718,0.06564103,0.052512825,0.08533334,0.25271797,0.4955898,0.62030774,0.41025645,0.5021539,0.6104616,0.5677949,0.34133336,0.19692309,0.15097436,0.15097436,0.21661541,0.44307697,0.38728207,0.23302566,0.20348719,0.26584616,0.118153855,0.052512825,0.03938462,0.055794876,0.07876924,0.098461546,0.14769232,0.19692309,0.21989745,0.2231795,0.26912823,0.318359,0.35774362,0.37743592,0.37743592,0.37743592,0.40369233,0.5677949,0.827077,1.2471796,1.9922053,2.605949,3.1967182,3.31159,2.9013336,2.3269746,1.6180514,1.8674873,2.8225644,4.07959,5.0904617,6.521436,6.009436,5.041231,4.2338467,3.3345644,2.3663592,1.0305642,0.18051283,0.009846155,0.052512825,0.40697438,0.6662565,0.74830776,0.7056411,0.7187693,0.6235898,0.58092314,0.5677949,0.6498462,0.9714873,0.8369231,0.69907695,0.64000005,0.6432821,0.5940513,0.574359,1.3587693,2.0873847,2.0545642,0.7187693,0.6629744,0.35446155,0.098461546,0.0032820515,0.0,0.013128206,0.08533334,0.14769232,0.18707694,0.2231795,0.36102566,0.5021539,0.57764107,0.636718,0.86317956,0.74830776,0.71548724,0.7811283,0.82379496,0.6104616,0.58420515,0.6071795,0.69579494,0.7778462,0.7089231,0.7187693,0.9682052,1.204513,1.4178462,1.847795,1.6213335,1.339077,1.214359,1.3259488,1.6049232,1.4703591,1.4834872,1.4998976,1.4539489,1.3686155,1.3718976,1.3883078,1.4769232,1.5721027,1.4736412,1.4408206,1.4506668,1.5556924,1.8313848,2.3893335,2.8225644,3.259077,3.570872,3.8104618,4.1780515,4.821334,5.277539,5.3136415,4.9887185,4.6769233,3.8432825,3.318154,3.0490258,2.930872,2.8192823,2.300718,2.097231,1.9922053,1.8904617,1.8248206,1.8642052,1.8379488,1.9790771,2.2121027,2.1431797,2.3171284,2.162872,2.3236926,2.8521028,3.2098465,3.767795,4.1747694,4.6178465,5.1364107,5.5991797,5.83877,6.1505647,6.009436,5.730462,6.4623594,6.4295387,6.442667,7.3025646,8.5202055,8.320001,8.054154,8.480822,8.822155,8.930462,9.271795,8.329846,7.830975,7.532308,7.253334,6.8988724,5.87159,5.077334,4.7261543,4.59159,4.017231,3.9614363,4.0041027,4.023795,3.9680004,3.8596926,4.1485133,4.1452312,4.007385,3.8301542,3.636513,3.4822567,3.4034874,3.4658465,3.7776413,4.4898467,4.716308,4.7950773,4.7327185,4.5554876,4.2896414,4.2240005,4.420923,4.6802053,4.903385,5.077334,5.8847184,6.636308,6.9677954,6.6560006,5.605744,4.8640003,4.027077,3.3542566,3.0162053,3.1113849,2.733949,2.4418464,2.3466668,2.3433847,2.1103592,2.2153847,2.100513,2.0545642,2.2088206,2.5435898,2.3368206,2.3663592,2.4484105,2.5074873,2.5928206,0.036102567,0.036102567,0.036102567,0.032820515,0.02297436,0.0,0.009846155,0.0032820515,0.0,0.0032820515,0.0,0.013128206,0.036102567,0.1148718,0.21989745,0.25928208,0.44964105,1.214359,2.6157951,4.1714873,4.844308,4.3290257,3.2361028,2.7142565,2.861949,2.7175386,2.681436,3.0227695,3.0654361,2.7241027,2.5140514,3.1540515,4.4800005,5.402257,5.5204105,5.113436,3.6594875,2.7569232,2.156308,1.8018463,1.847795,2.3762052,2.7241027,3.2032824,3.7251284,3.7874875,5.3136415,6.3376417,6.9152827,7.0367184,6.633026,7.5191803,8.769642,9.672206,10.325335,11.667693,12.297847,13.344822,14.201437,14.250668,12.859077,16.548103,24.365952,33.64103,40.84185,41.593437,39.93272,43.01457,48.518566,55.20739,62.93334,69.346466,67.81703,64.36759,61.026466,55.840824,49.847797,42.85703,38.866055,40.434875,48.689236,55.857235,55.46995,55.952415,58.597748,57.590157,53.809235,52.18462,55.325542,59.33621,53.8158,47.730877,40.533337,33.437542,27.086771,21.553232,19.416616,16.761436,15.415796,14.9398985,12.619488,9.048616,6.7085133,5.5269747,6.052103,9.45559,11.408411,12.360206,12.179693,11.565949,12.022155,11.424822,10.689642,12.484924,17.78872,25.911797,23.840822,21.48431,19.255796,18.176,19.872822,31.304207,38.344208,42.348312,42.932518,37.986465,34.868515,33.033848,29.426874,23.62749,17.860924,13.200411,11.280411,11.270565,11.385437,8.910769,7.716103,6.3212314,5.7074876,6.012718,6.514872,6.2720003,6.8660517,7.936001,8.87795,8.874667,11.286975,9.8363085,6.62318,3.515077,2.1366155,2.041436,2.228513,2.3827693,2.4451284,2.6289232,2.733949,3.4494362,4.4242053,5.7009234,7.755488,11.69395,14.145642,15.16636,14.949745,13.833847,12.777026,11.418258,10.381129,10.555078,13.10195,19.46913,24.851694,26.006977,23.588104,22.144001,22.4919,19.698874,16.518566,14.322873,13.08554,11.844924,10.866873,11.122872,12.875488,15.668514,16.482462,15.432206,14.588719,13.879796,11.080206,9.77395,8.513641,7.6635904,7.50277,8.237949,8.326565,7.64718,6.8004107,6.0717955,5.4186673,5.687795,6.4032826,7.138462,7.9327188,9.3078985,10.528821,10.617436,9.961026,8.982975,8.119796,7.8736415,7.2631803,6.5805135,6.117744,6.170257,4.893539,4.568616,4.135385,3.3936412,2.9768207,2.8127182,2.5042052,1.9593848,1.4244103,1.4736412,2.0676925,4.8738465,8.356103,10.883283,10.732308,19.328001,21.720617,20.926361,18.71754,15.602873,14.017642,15.698052,14.034052,9.504821,9.668923,17.69354,20.105848,20.171488,19.636515,18.73395,17.923283,14.7331295,11.398565,9.6984625,10.965334,8.018052,6.4032826,5.5729237,4.6539493,2.4582565,2.917744,8.477539,8.979693,3.7874875,1.8116925,2.3171284,4.9329233,6.3507695,5.5204105,3.636513,3.6627696,5.5630774,8.303591,10.240001,9.117539,8.621949,14.503386,15.0088215,8.841846,5.149539,6.380308,5.802667,5.4514875,5.733744,5.4482055,3.7743592,2.8192823,3.5774362,5.720616,7.6176414,12.987078,16.8599,18.031591,19.01949,26.056208,9.442462,6.557539,7.0990777,6.308103,4.9821544,3.9745643,3.4494362,5.280821,7.565129,4.6211286,3.5511796,4.972308,6.6494365,9.511385,17.660719,11.926975,7.962257,12.921437,20.709745,11.98277,14.454155,10.555078,9.186462,10.217027,4.453744,2.8127182,2.4910772,2.0775387,1.8576412,3.820308,3.058872,3.9056413,4.1878977,3.3411283,2.4418464,1.9167181,1.7985642,1.7427694,1.9954873,3.4002054,4.1682053,3.9253337,3.058872,2.172718,2.0742567,2.6256413,2.5600002,2.048,1.2996924,0.574359,0.9124103,1.4244103,1.657436,1.7001027,2.1792822,1.8543591,2.2022567,2.7273848,2.9702566,2.481231,2.6223593,2.5238976,1.9167181,1.0699488,0.78769237,0.9156924,0.955077,0.9124103,0.7515898,0.40697438,0.4266667,0.761436,1.3653334,1.8379488,1.394872,1.3161026,1.467077,1.6147693,1.6738462,1.7132308,2.6420515,2.7995899,2.297436,1.6443079,1.7591796,1.3489232,0.92553854,0.65312827,0.636718,0.955077,0.58420515,0.4594872,0.46933338,0.508718,0.46276927,0.574359,0.4004103,0.190359,0.08205129,0.08533334,0.098461546,0.18707694,0.29538465,0.3511795,0.28225642,0.38728207,0.40697438,0.6301539,0.9747693,0.9682052,0.46276927,0.4594872,0.636718,0.8336411,1.0535386,0.9321026,0.6498462,0.37415388,0.20676924,0.190359,0.30851284,0.51856416,0.7811283,1.0404103,1.2373334,2.3958976,2.156308,1.467077,0.8992821,0.6465641,0.9353847,0.90584624,0.6235898,0.2986667,0.27897438,0.32820517,0.27241027,0.46276927,0.892718,1.1716924,1.3850257,1.9167181,2.0841026,1.7723079,1.4276924,0.9714873,1.1257436,1.6377437,1.9528207,1.2274873,0.6859488,0.7056411,0.8172308,0.761436,0.46933338,0.25928208,0.25271797,0.34133336,0.36102566,0.108307704,0.19364104,0.21661541,0.18379489,0.13456412,0.13456412,0.101743594,0.08861539,0.072205134,0.059076928,0.072205134,0.10502565,0.118153855,0.108307704,0.14769232,0.37743592,0.48902568,0.6826667,0.7581539,0.6268718,0.32164106,0.16082053,0.08205129,0.08533334,0.18707694,0.4004103,0.3446154,0.15097436,0.06235898,0.098461546,0.072205134,0.013128206,0.006564103,0.026256412,0.049230773,0.055794876,0.10502565,0.16410258,0.18379489,0.16082053,0.15753847,0.19364104,0.20676924,0.23630771,0.27241027,0.27241027,0.3314872,0.5349744,0.7220513,0.95835906,1.529436,2.2383592,2.878359,3.0752823,2.7503593,2.1333334,1.4211283,1.3554872,1.847795,2.8291285,4.2272825,7.062975,5.865026,4.6539493,4.7392826,4.71959,4.647385,2.2383592,0.38728207,0.0032820515,0.013128206,0.24287182,0.5481026,0.6826667,0.63343596,0.6301539,0.5973334,0.65969235,0.61374366,0.512,0.6498462,0.72861546,0.6662565,0.6071795,0.571077,0.4594872,0.4266667,1.3193847,2.03159,1.8674873,0.5284103,0.90256417,0.56123084,0.16738462,0.013128206,0.0,0.0032820515,0.052512825,0.118153855,0.19364104,0.27897438,0.3446154,0.41682056,0.43651286,0.4660513,0.67610264,0.7581539,0.7844103,0.8041026,0.7975385,0.6695385,0.5973334,0.58420515,0.6301539,0.7056411,0.7253334,0.7450257,0.9878975,1.1848207,1.2668719,1.4080001,1.4178462,1.2537436,1.1815386,1.2635899,1.3751796,1.3850257,1.4605129,1.4342566,1.2898463,1.1782565,1.3620514,1.3850257,1.3357949,1.2537436,1.1355898,1.2800001,1.4703591,1.6246156,1.7920002,2.169436,2.4615386,2.8717952,3.2918978,3.757949,4.453744,4.634257,4.8311796,4.8049235,4.460308,3.8629746,2.612513,2.2482052,2.359795,2.5206156,2.284308,2.0939488,2.0151796,1.9954873,2.0512822,2.2744617,2.176,1.9298463,1.8674873,1.9987694,2.0217438,2.3204105,2.4188719,2.556718,2.7963078,3.0227695,3.4921029,3.6135387,3.8137438,4.3290257,5.1856413,5.533539,6.0258465,6.121026,5.927385,6.189949,6.012718,6.180103,6.918565,7.8506675,7.9852314,7.834257,8.0377445,8.352821,8.677744,9.074872,8.36595,7.8080006,7.3091288,6.921847,6.8562055,6.3376417,5.2020516,4.378257,4.1485133,4.1714873,3.9581542,3.8728209,3.9384618,4.06318,4.0303593,4.1222568,3.95159,3.820308,3.751385,3.5052311,3.1803079,3.131077,3.370667,3.8596926,4.4734364,4.585026,4.5554876,4.2272825,3.7743592,3.6857438,4.240411,4.562052,4.969026,5.4908724,5.8420515,6.422975,6.669129,6.416411,5.7042055,4.7622566,4.70318,4.20759,3.4133337,2.7667694,3.0227695,2.740513,2.7044106,2.8356924,2.878359,2.3958976,2.1956925,2.044718,1.9692309,2.0118976,2.2547693,2.2514873,2.3663592,2.5107694,2.6617439,2.878359,0.0,0.0,0.0,0.006564103,0.013128206,0.0,0.0,0.0,0.006564103,0.013128206,0.0,0.013128206,0.052512825,0.12471796,0.18707694,0.13784617,0.35774362,1.6475899,3.826872,5.8190775,5.661539,5.7829747,4.972308,3.95159,3.2656412,3.2656412,3.387077,2.674872,2.1989746,2.3302567,2.7470772,3.892513,4.9493337,5.536821,5.4580517,4.699898,3.3312824,2.3138463,1.719795,1.4473847,1.1913847,1.9232821,2.665026,3.4822567,4.384821,5.32677,6.5083084,7.821129,8.900924,9.18318,7.890052,9.048616,9.547488,10.243283,11.191795,11.641437,12.107488,13.384206,13.298873,12.750771,15.717745,24.395489,33.394875,38.229336,38.344208,37.126568,38.101337,41.439182,44.52103,44.560413,38.590363,38.980927,35.9319,32.200207,30.437746,33.158566,28.2519,24.937027,25.248823,30.720003,42.390976,52.00739,51.840004,49.043697,47.43549,47.471592,42.919388,39.84739,38.583797,38.275284,36.896824,39.43385,37.251286,30.431181,23.033438,23.056412,24.241232,19.849848,13.682873,9.104411,9.019077,8.211693,7.2861543,7.1647186,8.293744,10.650257,9.819899,10.758565,11.0145645,10.850462,13.22995,13.472821,11.592206,13.505642,19.6759,25.130669,18.136618,15.77354,17.476925,21.924105,27.03754,43.565952,48.951797,48.90257,44.783592,33.614773,26.817642,22.078362,17.414566,12.908309,10.696206,9.268514,9.314463,9.668923,9.399796,7.8112826,6.678975,6.1013336,5.9667697,6.0258465,5.904411,5.76,6.629744,7.3058467,7.972103,10.194052,13.072412,11.579078,8.264206,4.857436,2.2580514,2.612513,2.8488207,2.6322052,2.284308,2.7602053,3.0424619,3.754667,4.6080003,5.6320004,7.1548724,10.440206,11.536411,11.608616,11.283693,10.637129,9.55077,10.988309,12.931283,14.808617,17.532719,21.828924,25.202873,24.457848,20.985437,20.752413,19.423182,17.092924,15.750566,14.795488,11.047385,9.826463,10.171078,11.894155,14.165335,15.53395,15.852309,14.601848,13.02318,11.546257,9.810052,9.127385,8.848411,8.67118,8.418462,8.041026,7.955693,7.276308,6.340924,5.543385,5.3103595,5.5302567,6.189949,7.072821,8.136206,9.4916935,10.223591,10.269539,9.537642,8.621949,8.805744,8.792616,7.325539,6.377026,6.3540516,6.0717955,4.4734364,3.892513,4.325744,4.7458467,3.0982566,2.6322052,2.2613335,2.1530259,2.281026,2.425436,2.4615386,6.6461544,10.601027,12.1238985,11.185231,19.498669,21.832207,21.333336,20.791796,22.659285,17.47036,16.951796,18.235079,17.821539,11.595488,7.532308,9.7214365,11.533129,11.044104,11.034257,15.510976,13.124924,10.292514,9.061745,7.0957956,5.4482055,4.604718,3.69559,2.6289232,2.0906668,3.370667,5.7632823,7.0859494,6.2818465,3.387077,2.8750772,5.4547696,7.8670774,8.667898,8.237949,4.7491283,6.1013336,7.27959,7.200821,8.726975,9.508103,12.304411,13.062565,10.420513,5.720616,7.3321033,5.8880005,5.6418467,8.438154,13.686155,9.084719,6.2785645,9.892103,18.225233,23.253336,11.877745,7.210667,4.818052,2.9604106,2.5961027,7.3682055,8.021334,8.549745,11.08677,15.885129,11.329642,6.803693,5.901129,7.2927184,4.7294364,3.3378465,2.6880002,2.034872,2.8160002,8.651488,15.927796,13.3251295,12.383181,13.801026,7.4174366,11.628308,5.684513,5.937231,11.618463,4.8672824,5.4547696,6.5247183,5.7501545,3.6004105,3.3575387,2.5764105,4.164923,5.904411,6.518154,5.674667,3.1507695,1.7755898,0.90912825,0.43323082,0.764718,3.3378465,5.796103,5.5696416,3.1606157,2.1366155,2.6354873,2.8521028,2.934154,2.6978464,1.6475899,1.1946667,0.6170257,0.36758977,0.6301539,1.3128207,1.6902566,1.9495386,2.5107694,2.9440002,1.9692309,1.6016412,1.7493335,1.595077,1.142154,1.1913847,1.6410258,1.3883078,1.0962052,0.892718,0.380718,0.28225642,0.2231795,0.37415388,0.73517954,1.1126155,1.1126155,1.0765129,1.1093334,1.1618463,1.0535386,1.3095386,1.2537436,1.2537436,1.3686155,1.3423591,1.3915899,1.1290257,0.7089231,0.44307697,0.80738467,0.5152821,0.49887183,0.60061544,0.7318975,0.8533334,1.0633847,0.764718,0.380718,0.17066668,0.24287182,0.20676924,0.190359,0.21333335,0.27241027,0.32164106,0.5513847,0.636718,0.8566154,1.2242053,1.4802053,0.761436,0.50543594,0.4135385,0.3708718,0.44307697,0.761436,0.72861546,0.5218462,0.36102566,0.51856416,0.77456415,0.86646163,1.0666667,1.5195899,2.228513,3.570872,3.383795,2.284308,1.0502565,0.6104616,0.7318975,0.43323082,0.17066668,0.21661541,0.65641034,0.7187693,0.4955898,0.6235898,1.1355898,1.463795,1.8904617,1.9790771,1.8707694,1.5753847,0.97805136,0.45292312,0.4135385,0.8205129,1.3850257,1.5556924,1.0075898,0.9419488,0.77128214,0.45620516,0.51856416,0.34789747,0.16738462,0.13784617,0.20348719,0.108307704,0.14441027,0.16082053,0.17394873,0.18379489,0.18379489,0.17066668,0.13128206,0.07548718,0.036102567,0.06235898,0.21989745,0.24943592,0.22646156,0.19692309,0.18379489,0.34133336,0.51856416,0.60389745,0.5513847,0.380718,0.2231795,0.20020515,0.15097436,0.059076928,0.04594872,0.02297436,0.02297436,0.08533334,0.13456412,0.0,0.0,0.0,0.01969231,0.04266667,0.029538464,0.07876924,0.118153855,0.13784617,0.13456412,0.12143591,0.14769232,0.14441027,0.13784617,0.13784617,0.13784617,0.18707694,0.3708718,0.58092314,0.77128214,0.9911796,1.5524104,2.1431797,2.540308,2.5731285,2.1202054,1.3522053,1.5622566,1.9528207,2.2744617,2.8225644,6.7905645,8.247795,7.4436927,6.0160003,7.003898,6.442667,2.7667694,0.24615386,0.0,0.0,0.072205134,0.34789747,0.5316923,0.50543594,0.33476925,0.5677949,0.7253334,0.6465641,0.44307697,0.5021539,0.8467693,0.7844103,0.6301539,0.5349744,0.47261542,0.3511795,0.39384618,0.56451285,0.7122052,0.56451285,0.44307697,0.23958977,0.08533334,0.02297436,0.0,0.013128206,0.04266667,0.108307704,0.25271797,0.5349744,0.5218462,0.58420515,0.636718,0.6662565,0.702359,0.71548724,0.7811283,0.761436,0.7187693,0.8992821,0.7417436,0.6826667,0.702359,0.7515898,0.761436,0.8960001,1.2603078,1.4506668,1.3456411,1.1126155,1.211077,1.1454359,1.1454359,1.2406155,1.2668719,1.2668719,1.3751796,1.3817437,1.276718,1.2504616,1.4834872,1.394872,1.2406155,1.1848207,1.2832822,1.3686155,1.1782565,1.086359,1.2668719,1.6935385,2.1825643,2.487795,2.7306669,3.062154,3.6463592,4.20759,4.9362054,5.110154,4.535795,3.508513,2.7273848,2.231795,2.1267693,2.1989746,1.9068719,2.409026,2.349949,2.2022567,2.1891284,2.2744617,2.4188719,2.1924105,1.9232821,1.8051283,1.8773335,1.7558975,2.0184617,2.537026,3.0129232,2.9768207,3.121231,3.239385,3.636513,4.20759,4.4406157,4.525949,5.32677,6.1505647,6.419693,5.677949,5.284103,5.802667,6.491898,6.948103,7.0957956,7.79159,7.680001,7.834257,8.342975,8.329846,7.6603084,7.017026,6.692103,6.770872,7.125334,6.820103,5.5729237,4.3716927,3.8531284,4.31918,3.9384618,3.7809234,3.7448208,3.7251284,3.6168208,3.5314875,3.318154,3.0654361,2.8947694,2.9440002,2.934154,3.1113849,3.2722054,3.5216413,4.3027697,4.5587697,4.450462,4.161641,3.9417439,4.089436,5.346462,5.2480006,5.1200004,5.671385,6.987488,6.2916927,6.12759,6.091488,5.7501545,4.637539,4.161641,3.56759,3.3050258,3.242667,2.6715899,2.6223593,2.7831798,3.0752823,3.1770258,2.5173335,2.1989746,2.0939488,2.100513,2.231795,2.609231,2.156308,2.3663592,2.6387694,2.7667694,2.9144619,0.0,0.0,0.0,0.0,0.0032820515,0.0,0.0,0.0,0.0,0.0032820515,0.0,0.0032820515,0.026256412,0.08205129,0.20020515,0.40697438,1.2209232,2.9243078,5.3169236,7.6143594,8.43159,6.961231,6.1341543,6.436103,7.1056414,6.1078978,5.293949,4.919795,5.074052,4.9132314,2.674872,4.3585644,4.604718,4.588308,4.4045134,3.0523078,2.4746668,1.910154,1.5819489,1.5983591,1.9462565,2.356513,2.9801028,3.751385,4.7261543,6.0947695,7.3353853,8.493949,9.747693,10.748719,10.633847,10.358154,11.336206,12.475078,13.184001,13.364513,14.10954,15.665232,17.42113,19.672617,23.61436,29.138054,31.996721,33.618053,34.596104,34.68472,33.82482,32.213337,31.126976,30.516516,29.0199,28.278156,28.032001,25.892105,22.610052,22.111181,21.90113,20.850874,22.4919,28.01231,36.273235,42.886566,40.149338,37.632004,38.823387,41.133953,35.03918,30.595284,27.897438,27.300104,29.426874,38.908722,37.060925,28.734362,21.53354,25.813335,27.408413,24.146053,18.789745,14.201437,13.315283,15.507693,12.813129,9.399796,7.824411,9.03877,9.097847,9.472001,9.396514,9.176616,10.19077,11.96636,12.645744,15.048206,18.435284,18.491077,15.596309,17.174976,18.75036,19.754667,23.522463,26.870155,26.696207,28.199387,30.057028,24.425028,22.409847,22.104616,19.26236,14.129231,11.441232,9.701744,8.772923,7.433847,5.618872,4.4438977,4.2863593,5.110154,6.2194877,7.2270775,8.054154,8.356103,7.896616,7.4699492,7.6996927,9.032206,8.116513,6.695385,5.3727183,4.2994876,3.1737437,3.6824617,3.636513,3.0752823,2.5140514,2.934154,4.201026,4.7458467,5.3136415,6.226052,7.4010262,8.4972315,9.015796,9.143796,9.055181,8.92718,9.196308,9.915077,11.651283,14.985847,20.50954,24.44472,23.991796,20.102566,15.96718,17.004309,16.915693,15.350155,13.147899,10.807796,8.4972315,9.209436,10.417232,11.382154,12.442257,15.02195,15.356719,13.361232,11.1064625,9.734565,9.458873,10.41395,10.587898,9.947898,8.923898,8.418462,8.303591,7.450257,6.245744,5.1626673,4.7228723,4.6605134,5.228308,6.3606157,8.004924,10.102155,10.804514,10.499283,9.892103,9.554052,9.90195,10.164514,9.803488,9.488411,9.216001,8.320001,5.832206,5.284103,5.182359,4.854154,4.4274874,4.4045134,3.3280003,2.4943593,2.2908719,2.1956925,2.6912823,6.6527185,12.051693,16.193642,15.714462,18.566566,24.070566,29.210258,30.224413,22.610052,19.160616,13.965129,11.119591,11.45436,12.511181,7.830975,10.604308,12.78359,11.963078,11.385437,15.396104,15.75713,13.515489,10.282667,8.231385,6.669129,5.733744,5.037949,4.394667,3.8006158,3.7349746,4.8836927,5.799385,6.038975,6.183385,7.1548724,7.1548724,7.056411,7.315693,7.972103,4.821334,6.7282057,7.939283,6.629744,4.896821,5.7829747,16.472616,19.528206,12.740924,9.114257,11.506873,9.238976,6.058667,4.644103,6.5837955,8.700719,10.164514,9.196308,10.029949,22.898874,27.24431,18.34995,8.644924,3.754667,2.5206156,4.529231,5.113436,9.458873,15.399385,13.420309,18.41559,16.964924,11.467488,5.4482055,3.5577438,5.858462,11.667693,11.874462,6.409847,4.2568207,7.030154,8.891078,10.177642,9.800206,5.2315903,6.4065647,3.9811285,3.6660516,5.943795,6.0750775,4.788513,4.6145644,3.8564105,2.5009232,2.1989746,2.4320002,3.4560003,4.926359,6.038975,5.5302567,3.9778464,3.1737437,2.4582565,1.7165129,1.3718976,1.9659488,2.7634873,3.373949,3.8400004,4.650667,3.5971284,2.5337439,1.9232821,2.1825643,3.6627696,4.6080003,3.18359,1.4473847,0.60061544,0.9714873,1.9068719,2.6256413,3.3444104,3.8006158,3.2754874,2.2153847,2.1136413,1.913436,1.4736412,1.5819489,1.7887181,1.3784616,0.86646163,0.5021539,0.27241027,0.38728207,0.49230772,1.0633847,1.7329233,1.2603078,1.211077,1.404718,1.332513,1.086359,1.3587693,1.5064616,1.3817437,1.214359,1.1191796,1.0732309,1.083077,0.9156924,0.7220513,0.6826667,0.97805136,0.71548724,0.6826667,1.1585642,1.6804104,1.0502565,0.955077,0.7450257,0.5218462,0.36102566,0.318359,0.446359,0.55794877,0.67610264,0.7581539,0.69907695,0.7253334,0.88287187,1.2570257,1.6443079,1.5786668,0.8369231,0.5940513,0.43323082,0.2986667,0.47917953,0.6892308,0.65969235,0.7318975,1.0732309,1.6902566,1.4112822,1.4408206,1.4966155,1.591795,2.044718,2.3138463,1.9396925,1.4769232,1.2209232,1.2209232,0.8336411,0.4004103,0.17394873,0.20348719,0.3511795,0.5481026,0.5874872,0.75487185,0.9911796,0.892718,0.63343596,0.54482055,0.6268718,0.79425645,0.8795898,0.45292312,0.25928208,0.34133336,0.636718,0.98133343,1.1158975,1.083077,0.79097444,0.40697438,0.36102566,0.33476925,0.19364104,0.09189744,0.08861539,0.118153855,0.108307704,0.128,0.19364104,0.26256412,0.23302566,0.16082053,0.108307704,0.06564103,0.04266667,0.049230773,0.15753847,0.29538465,0.35774362,0.30851284,0.17066668,0.38728207,0.49230772,0.5152821,0.446359,0.23630771,0.702359,0.85005134,0.55794877,0.07548718,0.032820515,0.049230773,0.03938462,0.118153855,0.27569234,0.36758977,0.09189744,0.009846155,0.013128206,0.029538464,0.01969231,0.03938462,0.068923086,0.098461546,0.11158975,0.108307704,0.1148718,0.128,0.108307704,0.068923086,0.08861539,0.16738462,0.30851284,0.45620516,0.5973334,0.74830776,1.1618463,1.6705642,1.9987694,2.0217438,1.7657437,1.0371283,0.7089231,0.7778462,1.079795,1.2964103,3.8301542,5.405539,5.474462,4.585026,4.391385,2.7273848,1.214359,0.3052308,0.032820515,0.013128206,0.08533334,0.17723078,0.2855385,0.39056414,0.43323082,0.53825647,0.61374366,0.58420515,0.49230772,0.5021539,0.6301539,0.6695385,0.60061544,0.47917953,0.44964105,0.5415385,0.5284103,0.5218462,0.5415385,0.49230772,0.58420515,0.37415388,0.14441027,0.02297436,0.0,0.013128206,0.055794876,0.13784617,0.24943592,0.36430773,0.42994875,0.44964105,0.5021539,0.5513847,0.48246157,0.45620516,0.5481026,0.6432821,0.6662565,0.5940513,0.6695385,0.7089231,0.7253334,0.7318975,0.71548724,0.7417436,0.98133343,1.1257436,1.1224617,1.1618463,1.2406155,1.1257436,1.014154,1.0075898,1.1191796,1.1881026,1.2340513,1.3423591,1.4211283,1.2012309,1.463795,1.339077,1.2012309,1.1618463,1.0732309,1.1684103,1.0633847,1.024,1.1552821,1.3883078,1.8576412,2.0906668,2.3204105,2.6289232,2.9505644,3.5511796,4.1189747,4.4438977,4.394667,3.9253337,3.1048207,2.9111798,2.5337439,1.9626669,1.9922053,2.0841026,1.7755898,1.7624617,2.0841026,2.1530259,1.8281027,1.7263591,1.7723079,1.8510771,1.7657437,1.9462565,2.359795,2.8389745,3.1573336,3.0227695,2.917744,2.993231,3.2295387,3.4789746,3.4756925,3.4527183,3.8695388,4.4373336,4.8344617,4.6769233,4.7524104,5.1232824,5.671385,6.340924,7.131898,7.5946674,7.5487185,7.5421543,7.706257,7.781744,7.5191803,6.701949,5.7829747,5.21518,5.4416413,5.6254363,4.8147697,3.9417439,3.6069746,4.0500517,3.5938463,3.2918978,3.1474874,3.131077,3.1770258,3.131077,2.9768207,2.7470772,2.609231,2.8717952,2.8291285,2.937436,3.2328207,3.636513,3.948308,3.8728209,4.2436924,4.4701543,4.457026,4.6145644,5.412103,5.293949,5.113436,5.100308,4.8771286,4.640821,4.7655387,4.9493337,4.903385,4.3716927,3.308308,3.43959,3.8038976,3.8531284,3.4133337,3.3280003,3.4133337,3.5774362,3.6004105,3.1277952,2.359795,2.2153847,2.1956925,2.2219489,2.609231,2.7634873,2.609231,2.6551797,2.806154,2.3663592,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.16410258,0.78769237,1.5753847,1.6082052,1.8182565,3.4297438,6.3901544,9.672206,11.277129,9.6,8.598975,8.493949,8.618668,7.4240007,6.747898,6.73477,6.685539,5.914257,3.7251284,4.2994876,4.4110775,4.962462,5.5269747,4.332308,3.1770258,2.7241027,2.7700515,3.062154,3.2984617,3.3444104,3.9220517,4.854154,5.835488,6.432821,6.738052,7.39118,8.333129,9.416205,10.397539,12.143591,13.751796,14.857847,15.491283,16.055796,16.659693,18.868515,21.622156,24.598976,28.215797,30.57231,31.415798,31.051489,30.050465,29.210258,26.240002,23.5159,22.393438,22.738052,22.938257,23.433847,25.609848,24.530054,20.322464,18.166155,18.65518,18.993233,21.152822,26.0759,33.683697,38.560825,35.53149,33.795284,35.298466,34.707695,27.060514,22.54113,19.163898,17.604925,21.231592,33.473644,32.902565,27.073643,22.482054,24.562874,23.975386,22.839796,22.009438,21.316925,19.570873,27.382156,28.26831,22.419695,13.682873,9.580308,10.394258,10.056206,9.544206,9.577026,10.59118,12.688411,14.135796,15.668514,16.666258,15.172924,17.59836,20.470156,22.396719,23.61436,26.003695,23.739079,21.970053,23.568413,26.479591,23.719387,23.450258,22.245745,20.168207,17.398155,14.244103,14.096412,12.471796,9.691898,6.76759,5.3760004,4.6572313,5.5269747,7.4075904,9.133949,8.956718,8.809027,7.4174366,6.3967185,6.11118,5.684513,4.8147697,4.460308,4.604718,4.821334,4.263385,4.388103,4.013949,3.4330258,2.9801028,3.0293336,3.6660516,3.9975388,4.493129,5.543385,7.433847,8.277334,8.641642,8.789334,8.818872,8.674462,8.940309,9.852718,12.455385,17.56882,25.777233,29.653336,24.982977,17.490053,12.107488,12.973949,15.025232,14.585437,12.511181,10.125129,9.238976,9.193027,10.026668,10.617436,11.575796,15.232001,15.169642,12.186257,9.55077,8.818872,9.8363085,10.765129,10.699488,9.691898,8.352821,7.8473854,8.595693,7.9130263,6.436103,4.900103,4.1550775,4.44718,5.540103,6.9842057,8.608821,10.545232,10.627283,9.964309,9.921641,10.902975,12.347078,12.580104,13.243078,13.400617,12.790154,11.828514,8.759795,6.944821,5.805949,5.1954875,5.3727183,5.3431797,4.3749747,3.8662567,3.9384618,3.4264617,4.089436,8.2215395,13.331694,17.178257,17.769028,17.289848,23.394463,30.598566,33.217644,25.37354,24.07713,18.07754,14.79877,15.819489,16.869745,12.1468725,11.621744,12.721231,13.147899,10.896411,12.586668,12.708103,11.487181,10.006975,10.217027,8.664616,7.430565,6.76759,6.51159,6.0750775,5.2644105,5.398975,5.8289237,6.308103,6.99077,9.682052,8.835282,7.026872,6.38359,8.598975,5.865026,6.3901544,6.6527185,5.730462,5.2742567,11.477334,15.638975,16.853334,14.887385,10.174359,17.72636,18.241642,14.099693,8.602257,5.940513,5.4974365,5.756718,4.59159,4.0434875,10.299078,15.038361,11.044104,6.4722056,4.279795,2.228513,4.2141542,3.817026,7.716103,14.460719,14.477129,16.229744,17.650873,13.879796,6.560821,3.8432825,4.2240005,8.300308,11.697231,12.028719,8.917334,7.716103,8.146052,9.068309,8.753231,4.857436,3.5807183,3.1409233,3.8432825,4.9887185,4.857436,4.713026,4.6178465,3.5314875,1.9954873,2.1464617,2.5304618,3.0949745,4.1747694,5.172513,4.568616,3.6069746,3.43959,3.508513,3.3345644,2.5042052,1.6443079,1.3718976,1.847795,2.9801028,4.44718,3.43959,2.6978464,2.0709746,1.8609232,2.8389745,4.315898,5.1298466,4.388103,2.5764105,1.5819489,2.162872,3.0260515,3.9876926,4.637539,4.325744,4.1747694,3.9712822,3.748103,3.4166157,2.7766156,2.556718,1.6114873,0.86974365,0.5940513,0.35446155,0.34789747,0.5907693,1.2406155,1.8576412,1.4145643,1.4506668,1.7033848,1.6902566,1.4506668,1.5524104,1.9626669,1.8018463,1.4802053,1.3587693,1.7591796,1.9856411,1.5491283,1.1618463,1.1388719,1.3981539,1.3620514,1.2373334,1.4572309,1.8215386,1.4998976,1.1913847,1.083077,0.90584624,0.60389745,0.3249231,0.32820517,0.45292312,0.7318975,1.0568206,1.1782565,0.8763078,0.9944616,1.2077949,1.3095386,1.2077949,0.65312827,0.45620516,0.34789747,0.29210258,0.47917953,0.69907695,0.79097444,0.9485129,1.401436,2.4057438,1.8510771,1.5524104,1.339077,1.1716924,1.1388719,1.0732309,0.892718,0.9321026,1.2274873,1.529436,0.88287187,0.39056414,0.15425642,0.14112821,0.15425642,0.39384618,0.49887183,0.7778462,1.079795,0.8205129,0.4004103,0.190359,0.23958977,0.47917953,0.73517954,0.47261542,0.3708718,0.32820517,0.318359,0.41025645,0.7056411,0.88943595,0.7450257,0.39712822,0.30194873,0.2855385,0.21333335,0.12471796,0.059076928,0.07548718,0.118153855,0.118153855,0.14441027,0.19364104,0.17066668,0.1148718,0.07548718,0.055794876,0.06235898,0.09189744,0.12471796,0.25271797,0.33476925,0.30851284,0.19692309,0.3249231,0.4397949,0.47589746,0.40369233,0.23630771,0.49887183,0.61374366,0.4594872,0.17394873,0.13128206,0.20676924,0.16410258,0.15753847,0.23630771,0.33805132,0.48902568,0.3249231,0.12471796,0.01969231,0.006564103,0.009846155,0.02297436,0.04594872,0.07548718,0.08861539,0.0951795,0.128,0.118153855,0.068923086,0.059076928,0.108307704,0.19692309,0.318359,0.4594872,0.5940513,0.8205129,1.1257436,1.3981539,1.5163078,1.3686155,0.8008206,0.40697438,0.27897438,0.3708718,0.512,1.5589745,2.4910772,3.4527183,4.066462,3.4560003,2.665026,1.3423591,0.37743592,0.049230773,0.02297436,0.04594872,0.07876924,0.17723078,0.33805132,0.4955898,0.52512825,0.5349744,0.512,0.47261542,0.45620516,0.48574364,0.6498462,0.6629744,0.5021539,0.39712822,0.49887183,0.52512825,0.49887183,0.45620516,0.45620516,0.5940513,0.380718,0.14441027,0.032820515,0.009846155,0.013128206,0.03938462,0.10502565,0.2100513,0.3117949,0.43323082,0.574359,0.78769237,0.9124103,0.56451285,0.512,0.512,0.55794877,0.6071795,0.58420515,0.67938465,0.6662565,0.67282057,0.7417436,0.81066674,0.79097444,0.86974365,0.94523084,1.0075898,1.148718,1.3522053,1.1585642,0.9189744,0.8402052,0.9747693,1.2340513,1.270154,1.3489232,1.4473847,1.2438976,1.3095386,1.1684103,1.0404103,0.97805136,0.86646163,0.90584624,0.85005134,0.88615394,1.0601027,1.2570257,1.5392822,1.847795,2.1825643,2.477949,2.5928206,2.9538465,3.2853336,3.4034874,3.2689233,2.9833848,2.4188719,2.4516926,2.3269746,1.9889232,2.0775387,1.9429746,1.8773335,1.8379488,1.8313848,1.8937438,1.6508719,1.5885129,1.7263591,1.9462565,1.9790771,1.910154,2.1366155,2.5862565,3.0096412,2.9801028,3.2000003,3.6036925,3.7021542,3.4198978,3.114667,3.0654361,3.3345644,3.7907696,4.2962055,4.709744,4.8607183,5.0051284,5.3169236,5.940513,7.003898,7.39118,7.0465646,6.7840004,6.941539,7.397744,6.616616,5.865026,5.0674877,4.466872,4.6276927,4.5522056,3.95159,3.3247182,3.0162053,3.2229745,2.740513,2.4976413,2.4418464,2.5435898,2.8192823,2.665026,2.4484105,2.3335385,2.3663592,2.487795,2.3958976,2.5665643,2.9013336,3.2918978,3.6135387,3.4691284,3.7448208,4.073026,4.2994876,4.4800005,5.435077,5.6451287,5.3103595,4.6211286,3.761231,3.9548721,4.0336413,4.1550775,4.3716927,4.640821,4.31918,4.667077,4.8082056,4.4373336,3.7940516,3.8432825,3.95159,3.826872,3.4231799,2.9604106,2.5632823,2.28759,2.2088206,2.3335385,2.5895386,2.7208207,2.5862565,2.5074873,2.4648206,2.100513,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.029538464,0.10502565,0.86317956,2.4976413,4.06318,3.4756925,2.4320002,3.1573336,5.5072823,8.717129,11.405129,11.739899,11.631591,11.0145645,10.020103,8.956718,8.89436,8.55959,7.857231,6.875898,5.8486156,5.668103,5.32677,5.98318,7.0432825,6.1768208,4.8311796,5.3202057,6.058667,6.2162056,5.720616,4.768821,4.919795,5.622154,6.294975,6.340924,5.9634876,6.4000006,7.394462,8.756514,10.377847,13.236514,15.130258,16.082052,16.840206,18.888206,18.888206,20.25354,22.121027,24.034464,25.970873,26.65354,26.4599,25.337439,23.706259,22.468925,20.683489,18.83241,18.57313,19.669334,19.977848,20.539078,23.686565,23.650463,19.899078,17.155283,17.51631,18.356514,20.59159,24.86154,31.527388,34.287594,32.28554,30.680618,30.12267,26.774977,20.224,16.482462,13.574565,12.143591,15.458463,25.03549,26.440207,24.730259,22.869335,21.707489,20.929642,22.360617,24.080412,24.969849,24.697437,40.175594,44.914875,36.81149,21.940514,14.54277,15.556924,11.818667,8.982975,9.219283,11.1983595,12.609642,13.722258,14.972719,16.433231,17.814976,22.715078,25.639387,27.520002,28.33067,27.096617,22.25231,20.690052,22.452515,25.091284,23.657028,23.236925,21.254566,20.26995,20.608002,20.33559,19.72513,16.137848,11.588924,7.893334,6.6592827,5.832206,5.8486156,7.0957956,8.530052,7.680001,7.3550773,6.445949,5.6287184,4.9394875,3.7743592,3.9975388,4.164923,4.2929235,4.3651285,4.325744,4.194462,3.9975388,3.8006158,3.636513,3.4822567,3.4756925,3.9712822,4.5817437,5.4908724,7.453539,9.380103,9.363693,9.07159,9.120821,9.081436,9.977437,11.493745,15.176207,22.17354,33.23077,34.510773,24.740105,14.378668,9.330873,10.939077,13.4859495,13.705847,12.425847,10.889847,10.771693,10.256411,10.368001,10.794667,12.212514,16.305231,16.249437,12.668719,9.6525135,8.946873,9.980719,10.187488,9.750975,8.720411,7.5618467,7.174565,8.418462,7.8539495,6.4557953,5.1232824,4.699898,5.142975,6.5805135,8.231385,9.6754875,10.850462,10.489437,9.833026,10.617436,12.937847,15.24513,15.632411,16.54154,17.092924,16.853334,15.839181,12.048411,8.749949,7.0334363,6.8430777,6.99077,6.052103,5.609026,5.549949,5.395693,4.3060517,5.041231,7.752206,11.073642,13.991385,15.858873,18.176,25.248823,32.623592,35.324722,27.844925,25.61313,22.478771,22.340925,24.083694,21.569643,17.09949,13.824001,13.522053,14.841437,13.279181,13.013334,12.714667,11.697231,10.873437,12.737642,13.220103,11.779283,9.69518,8.132924,8.139488,7.574975,7.3091288,6.87918,6.2851286,5.9667697,8.690872,8.077128,6.2720003,5.5926156,8.533334,7.2861543,6.4032826,5.622154,5.5597954,7.6898465,14.9628725,13.285745,12.491488,13.574565,8.690872,17.417847,22.659285,22.22277,17.72636,14.572309,8.474257,4.972308,3.2131286,2.6617439,3.0818465,4.6178465,3.7448208,3.058872,2.9604106,1.6311796,3.6102567,2.8324106,5.0642056,10.932513,15.954053,12.937847,14.86113,13.312001,7.643898,4.9952826,3.062154,4.141949,8.214975,12.626052,12.07795,9.622975,8.832001,8.815591,8.2215395,5.225026,3.259077,3.117949,4.0402055,4.850872,3.9778464,4.4865646,4.8344617,4.092718,2.5993848,1.975795,2.5304618,2.7667694,3.3936412,4.023795,3.1573336,2.7273848,3.1048207,3.5905645,3.6594875,2.934154,1.7624617,1.3062565,1.404718,1.9790771,3.0129232,2.8389745,3.2131286,3.170462,2.605949,2.294154,3.1409233,5.1856413,5.7764106,4.670359,4.010667,3.6890259,3.879385,4.568616,5.152821,4.44718,5.024821,5.0510774,4.844308,4.394667,3.3641028,2.8356924,1.6311796,0.8992821,0.7975385,0.51856416,0.3052308,0.48902568,1.079795,1.7296412,1.7591796,1.723077,1.7952822,1.6278975,1.3128207,1.3817437,2.0775387,2.0184617,1.7460514,1.782154,2.6420515,3.0129232,2.540308,2.0118976,1.7952822,1.8543591,1.975795,1.6902566,1.5753847,1.7690258,2.0020514,1.9003079,1.7329233,1.3883078,0.90256417,0.44307697,0.33805132,0.35446155,0.6432821,1.1323078,1.5195899,1.1618463,1.404718,1.5688206,1.3718976,0.9288206,0.4660513,0.34133336,0.4135385,0.5677949,0.7122052,1.1979488,1.7788719,1.9954873,2.028308,2.7109745,1.7657437,1.2242053,0.9747693,0.81066674,0.42338464,0.32820517,0.30194873,0.5021539,0.8730257,1.1454359,0.6268718,0.28882053,0.15097436,0.14112821,0.101743594,0.26584616,0.36758977,0.60389745,0.83035904,0.571077,0.43323082,0.26584616,0.2297436,0.3708718,0.60061544,0.508718,0.5021539,0.41025645,0.23630771,0.14769232,0.28882053,0.49887183,0.512,0.3446154,0.28225642,0.2231795,0.20020515,0.15097436,0.08533334,0.08861539,0.14441027,0.11158975,0.08533334,0.10502565,0.14112821,0.128,0.09189744,0.07548718,0.08861539,0.128,0.11158975,0.19692309,0.24943592,0.2231795,0.190359,0.24615386,0.380718,0.4594872,0.42338464,0.30851284,0.34133336,0.36102566,0.33805132,0.31507695,0.4004103,0.44964105,0.41682056,0.3708718,0.34133336,0.30194873,0.6235898,0.512,0.30851284,0.16738462,0.08533334,0.032820515,0.006564103,0.016410258,0.04266667,0.059076928,0.059076928,0.101743594,0.1148718,0.08533334,0.06564103,0.07548718,0.10502565,0.17723078,0.29538465,0.45620516,0.6465641,0.7778462,0.9353847,1.0666667,1.0010257,0.61374366,0.34789747,0.16738462,0.08533334,0.15097436,0.3511795,0.6859488,1.6640002,2.8127182,2.6683078,2.9801028,2.1136413,1.024,0.27569234,0.055794876,0.052512825,0.052512825,0.12471796,0.27897438,0.4955898,0.45620516,0.43323082,0.44307697,0.47261542,0.48902568,0.45292312,0.57764107,0.61374366,0.50543594,0.4201026,0.446359,0.48574364,0.47261542,0.4266667,0.44964105,0.60389745,0.40697438,0.17394873,0.04594872,0.016410258,0.016410258,0.029538464,0.08205129,0.18051283,0.318359,0.42994875,0.6104616,0.827077,0.9156924,0.5874872,0.5481026,0.48574364,0.49230772,0.58092314,0.69907695,0.7384616,0.6662565,0.6662565,0.77456415,0.8795898,0.80738467,0.79097444,0.8172308,0.8960001,1.0436924,1.3226668,1.1093334,0.85005134,0.77456415,0.892718,1.1158975,1.1618463,1.2635899,1.4244103,1.3915899,1.2012309,1.0404103,0.92553854,0.85005134,0.7811283,0.7089231,0.69251287,0.764718,0.9321026,1.1848207,1.3029745,1.5360001,1.8445129,2.1366155,2.2514873,2.4582565,2.6683078,2.674872,2.4648206,2.2449234,2.1924105,2.3663592,2.2711797,1.9790771,2.1464617,2.0578463,2.0873847,1.9823592,1.8084104,1.9462565,1.7296412,1.5688206,1.595077,1.7723079,1.8674873,1.8018463,1.910154,2.2219489,2.612513,2.8160002,3.3280003,3.8695388,3.892513,3.3936412,2.9144619,2.986667,3.1737437,3.4264617,3.8629746,4.7327185,4.9788723,5.1659493,5.540103,6.1997952,7.1023593,7.6898465,6.8562055,6.058667,5.9503593,6.4032826,5.8223596,5.4514875,4.8640003,4.1747694,4.0402055,3.817026,3.3345644,2.793026,2.4057438,2.4057438,2.0545642,1.8445129,1.9003079,2.2186668,2.6551797,2.3171284,2.038154,1.9265642,1.9232821,1.8281027,1.7788719,2.0808206,2.537026,2.9735386,3.2295387,3.1967182,3.2196925,3.3280003,3.5413337,3.8629746,4.8804107,5.333334,5.024821,4.1714873,3.3969233,3.6824617,3.6758976,3.7776413,4.1583595,4.7392826,4.9788723,5.172513,5.146257,4.7655387,3.9384618,4.0369234,4.0402055,3.6594875,3.0260515,2.6978464,2.605949,2.3794873,2.349949,2.540308,2.6584618,2.6617439,2.4549747,2.228513,2.0775387,1.9889232,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.03938462,0.15097436,0.55794877,2.3433847,4.8082056,6.4295387,4.8836927,2.9472823,2.5632823,3.2689233,5.146257,8.79918,12.688411,14.332719,13.748514,12.07795,11.592206,12.2157955,11.250873,9.714872,8.569437,8.713847,8.710565,7.456821,7.4010262,8.464411,8.03118,7.456821,8.969847,10.368001,10.433641,8.923898,6.38359,5.7731285,5.8814363,6.1538467,6.701949,6.2588725,6.73477,8.034462,9.80677,11.441232,13.568001,15.43877,16.433231,17.322668,20.26995,19.659489,18.996513,18.638771,18.714258,19.127796,19.403488,17.929848,16.787693,16.534975,16.213335,18.44513,18.422155,18.70113,19.524925,18.835693,18.264616,20.982155,22.098053,20.374975,18.215385,18.258053,18.707693,20.404514,23.640617,28.166567,28.74749,27.48718,24.982977,21.779694,18.372925,14.828309,12.3306675,11.050668,11.250873,13.292309,17.352207,21.507284,24.297028,24.549746,21.38913,21.99631,25.583591,27.136002,26.59118,28.85908,47.665234,52.90667,43.03098,26.210464,20.338873,21.59918,14.336001,9.265231,9.764103,11.867898,11.195078,11.716924,14.342566,18.983387,24.579285,27.408413,28.786875,29.256207,28.084515,23.27631,18.070976,17.900309,20.506258,23.250053,23.138464,22.839796,21.559797,21.349745,22.980925,25.93477,22.278566,16.193642,10.466462,7.0104623,6.8660517,6.7577443,5.7829747,5.428513,5.691077,5.0576415,5.2381544,5.7140517,5.5302567,4.6769233,4.096,4.7458467,4.568616,3.7448208,2.9571285,3.383795,3.3608208,3.7710772,4.2436924,4.519385,4.466872,4.768821,5.4908724,6.0291286,6.416411,7.3386674,10.036513,9.705027,9.147078,9.488411,10.177642,12.724514,14.483693,19.10154,28.212515,41.46544,36.736004,22.35077,10.962052,7.7456417,10.368001,11.979488,12.544001,12.265027,11.759591,12.071385,12.3306675,11.890873,12.301129,14.460719,18.612514,18.789745,14.749539,11.264001,10.154668,10.308924,9.416205,8.467693,7.565129,6.928411,6.892308,7.77518,7.276308,6.363898,5.792821,6.11118,6.2752824,7.972103,9.91836,11.280411,11.680821,10.860309,10.28595,11.54954,14.50995,17.306257,18.392616,19.27877,20.529232,21.48431,20.246977,16.239592,11.979488,9.970873,10.240001,10.341744,8.267488,8.096821,7.7718983,6.554257,5.0215387,5.684513,5.792821,6.6100516,8.595693,11.428103,20.522669,29.029745,36.55549,40.280617,34.966976,29.83713,29.735388,32.439796,33.729645,27.362463,21.602463,17.94954,16.846771,17.529438,18.011898,17.7559,17.778873,16.33477,14.313026,15.235283,18.891489,17.64431,13.275898,8.999385,9.458873,9.429334,9.110975,7.8473854,5.83877,4.1517954,5.2381544,5.3103595,4.827898,4.8804107,7.197539,8.2215395,7.2172313,5.9503593,6.058667,9.028924,12.173129,10.650257,9.796924,9.990565,6.6461544,10.499283,18.65518,23.722668,23.890053,22.938257,15.881847,10.105436,6.7183595,5.5663595,5.2447186,5.674667,3.259077,1.2274873,0.76800007,1.0272821,2.1497438,1.782154,2.6584618,6.7249236,15.133539,10.827488,11.424822,10.57477,7.197539,5.4613338,3.5905645,3.7382567,5.47118,7.8014364,9.179898,8.155898,8.667898,9.232411,8.677744,6.1440005,4.201026,3.242667,3.4494362,4.3290257,4.716308,4.096,4.5390773,4.8771286,4.164923,1.6771283,2.3072822,2.5304618,2.9243078,3.249231,2.4582565,2.162872,2.7142565,3.058872,2.8356924,2.4155898,1.8543591,1.7526156,1.6672822,1.5491283,1.7329233,2.284308,3.5511796,4.240411,3.9975388,3.3936412,2.8553848,3.9122055,4.8738465,5.362872,6.3277955,5.290667,4.6867695,4.7655387,4.9427695,3.7907696,4.2174363,4.4734364,4.3027697,3.7021542,2.917744,2.4582565,1.3817437,0.81394875,0.86646163,0.636718,0.30194873,0.318359,0.7975385,1.5360001,1.9823592,1.9035898,1.7099489,1.2340513,0.77128214,1.086359,1.8182565,1.8642052,1.7723079,2.0545642,3.1934361,3.4625645,3.2164104,2.7766156,2.3991797,2.2547693,2.4057438,2.1136413,1.9659488,2.1792822,2.6026669,3.0424619,2.7175386,2.097231,1.4769232,0.9714873,0.79425645,0.5546667,0.571077,0.92553854,1.4572309,1.5031796,2.0906668,2.3138463,1.8248206,0.8598975,0.380718,0.39384618,0.7450257,1.1355898,1.1126155,1.8313848,2.917744,3.318154,2.9210258,2.5862565,1.2406155,0.764718,0.79097444,0.83035904,0.27569234,0.15097436,0.108307704,0.20348719,0.36430773,0.40369233,0.2231795,0.16082053,0.20348719,0.27569234,0.2297436,0.19364104,0.23958977,0.29210258,0.2855385,0.17066668,0.4004103,0.39712822,0.33805132,0.3511795,0.5021539,0.56123084,0.55794877,0.43651286,0.25928208,0.19364104,0.118153855,0.14769232,0.21989745,0.2855385,0.30851284,0.256,0.20020515,0.15097436,0.118153855,0.13784617,0.18379489,0.12143591,0.055794876,0.055794876,0.15753847,0.21989745,0.16082053,0.108307704,0.108307704,0.13128206,0.11158975,0.17066668,0.190359,0.16738462,0.19692309,0.23630771,0.36430773,0.4594872,0.4660513,0.4004103,0.4397949,0.45292312,0.43651286,0.48246157,0.74830776,0.6268718,0.65312827,0.7450257,0.7417436,0.38400003,0.42338464,0.43651286,0.4397949,0.40697438,0.23958977,0.108307704,0.059076928,0.03938462,0.026256412,0.02297436,0.013128206,0.049230773,0.072205134,0.07548718,0.07548718,0.06564103,0.055794876,0.059076928,0.1148718,0.28225642,0.55794877,0.62030774,0.65312827,0.7056411,0.69579494,0.49230772,0.36102566,0.2297436,0.08861539,0.02297436,0.08861539,0.19692309,0.45292312,0.88287187,1.4309745,2.1398976,2.3302567,1.8182565,0.85005134,0.09189744,0.10502565,0.07548718,0.0951795,0.21661541,0.46276927,0.37743592,0.34789747,0.39056414,0.47589746,0.54482055,0.47589746,0.45292312,0.4660513,0.5021539,0.5513847,0.46933338,0.4594872,0.44307697,0.4135385,0.4266667,0.60389745,0.49230772,0.26584616,0.068923086,0.016410258,0.016410258,0.029538464,0.07876924,0.17066668,0.32164106,0.38728207,0.4955898,0.5481026,0.52512825,0.47261542,0.48246157,0.46933338,0.5152821,0.6432821,0.79425645,0.7778462,0.6892308,0.69579494,0.80738467,0.8566154,0.7515898,0.7450257,0.75487185,0.77128214,0.88287187,1.0666667,0.9288206,0.78769237,0.7811283,0.8467693,0.85005134,0.9124103,1.0962052,1.3259488,1.3981539,1.1060513,0.9682052,0.8992821,0.8598975,0.8402052,0.65969235,0.6859488,0.75487185,0.8402052,1.0732309,1.1454359,1.1881026,1.3423591,1.6147693,1.8904617,2.044718,2.2383592,2.3138463,2.2383592,2.103795,2.5140514,2.7798977,2.4549747,1.8543591,2.03159,2.2022567,2.156308,2.0217438,1.9593848,2.1530259,1.8740515,1.6147693,1.5163078,1.5491283,1.4998976,1.654154,1.8445129,2.0545642,2.281026,2.540308,3.121231,3.4855387,3.5380516,3.2820516,2.809436,3.05559,3.1540515,3.2065644,3.4527183,4.279795,4.673641,5.3103595,6.0324106,6.7117953,7.2369237,7.9130263,6.764308,5.543385,5.031385,5.0215387,5.2414365,5.2742567,4.8377438,4.073026,3.5314875,3.3936412,3.0162053,2.487795,2.0118976,1.8970258,1.7066668,1.4900514,1.6311796,2.1202054,2.556718,2.103795,1.8116925,1.5885129,1.3784616,1.1585642,1.2340513,1.657436,2.231795,2.7109745,2.8192823,2.8980515,2.7602053,2.5698464,2.5731285,3.114667,3.889231,4.384821,4.2994876,3.757949,3.2820516,3.3312824,3.2787695,3.4888208,3.9712822,4.3716927,4.601436,4.5554876,4.6769233,4.7622566,3.9745643,3.95159,3.7710772,3.3247182,2.7831798,2.6157951,2.3991797,2.4516926,2.605949,2.737231,2.7602053,2.6912823,2.2908719,1.9396925,1.8215386,1.9495386,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01969231,0.128,0.45620516,1.8018463,4.663795,6.6527185,6.4590774,3.8465643,2.8553848,2.553436,2.409026,3.0358977,6.2096415,13.02318,15.658668,15.297642,14.132514,15.366566,16.52513,16.082052,13.682873,10.994873,11.703795,11.98277,10.039796,9.399796,10.594462,11.168821,11.707078,11.667693,12.78359,14.073437,11.841642,7.788308,6.636308,6.4656415,6.9349747,9.278359,8.874667,8.920616,9.731283,11.063796,12.100924,14.139078,16.249437,17.808413,18.402462,17.85436,17.585232,16.180513,14.411489,13.6237955,15.747283,14.916924,12.603078,11.244308,11.490462,12.22236,16.738462,19.324718,20.59159,20.28636,17.273438,17.8839,19.88595,22.029129,23.476515,23.817848,21.43836,20.594873,20.407797,20.978874,23.40759,24.067284,20.97231,16.968206,13.978257,13.000206,10.230155,9.124104,10.243283,12.658873,13.978257,16.065641,24.109951,31.661951,34.2679,29.495796,27.638157,31.8359,34.68472,34.53703,35.475697,41.08144,41.327595,31.40267,17.64431,17.532719,20.706463,17.444103,15.96718,17.362053,15.579899,10.404103,11.1064625,16.922258,24.74995,29.144617,26.006977,22.137438,18.763489,16.403694,14.87754,14.437745,17.78872,21.602463,24.65149,27.80226,31.097439,29.29231,26.82749,25.055182,22.249027,15.875283,9.741129,5.865026,5.097026,7.1122055,7.3058467,6.229334,5.100308,4.3618464,3.6758976,4.6769233,5.4416413,5.3005133,4.585026,4.6080003,4.4012313,3.892513,3.239385,2.7142565,2.7011285,2.934154,3.7152824,4.7950773,5.737026,5.920821,7.77518,7.7357955,7.315693,7.0826674,6.669129,7.1187696,7.765334,8.809027,10.433641,12.803283,16.794258,17.408,22.954668,34.888206,47.78995,34.68144,19.400208,9.885539,7.6701546,7.890052,10.134975,11.877745,12.189539,11.900719,13.610668,14.805334,14.116103,14.726565,17.85436,22.75118,22.226053,16.722052,12.806565,12.370052,12.603078,9.905231,7.722667,6.5017443,6.370462,7.125334,7.0892315,6.997334,6.7282057,6.491898,6.820103,6.6625648,9.5146675,12.3536415,13.843694,14.342566,11.900719,10.541949,10.86359,13.046155,16.83036,19.429745,21.720617,24.654772,27.060514,25.619694,23.640617,19.311592,16.003283,15.199181,16.49559,14.857847,13.781334,11.716924,8.989539,7.781744,7.9163084,7.0432825,5.970052,5.98318,8.864821,20.401232,28.081232,37.80595,50.018467,59.72021,55.522465,51.79077,49.39816,46.562466,38.846363,26.850464,24.425028,23.827694,21.953642,20.355284,23.04,23.18113,22.281847,20.555489,16.905848,20.982155,20.683489,15.619284,9.419488,9.750975,8.723693,7.8014364,6.8233852,5.5171285,3.4789746,3.2000003,3.82359,4.269949,4.4012313,5.034667,7.525744,8.395488,7.637334,6.052103,5.2348723,6.5903597,6.73477,8.041026,9.796924,8.208411,5.402257,8.802463,12.721231,13.426873,9.156924,15.235283,13.833847,11.277129,9.714872,7.125334,8.198565,4.7524104,1.8707694,1.2373334,1.1126155,1.4933335,1.1749744,1.0666667,2.986667,9.688616,6.3212314,6.997334,7.125334,5.182359,2.7175386,3.6069746,4.634257,4.8311796,3.7842054,1.6475899,2.477949,5.330052,10.184206,13.515489,8.316719,3.82359,2.2153847,2.9111798,4.923077,6.8496413,4.240411,3.9811285,5.2315903,5.865026,2.4713848,1.9593848,2.8488207,3.6890259,4.0336413,4.4242053,2.8389745,2.8356924,3.0785644,2.7831798,1.7099489,1.5753847,1.4145643,1.4572309,1.6968206,1.8904617,2.0644104,2.802872,3.5413337,4.309334,5.737026,4.1747694,3.7284105,3.6004105,3.5314875,3.8006158,3.3608208,3.7185643,3.820308,3.4724104,3.3280003,3.117949,2.7569232,2.5862565,2.5140514,2.0151796,2.2088206,1.1881026,0.56451285,0.67282057,0.56451285,0.30851284,0.36430773,0.6432821,1.020718,1.3128207,1.8379488,1.6935385,1.2406155,0.9517949,1.404718,1.6968206,1.4867693,1.3883078,1.8379488,3.0818465,3.0227695,2.7142565,2.4746668,2.4516926,2.609231,2.8291285,3.1048207,3.4625645,3.751385,3.6168208,4.397949,4.135385,3.4527183,2.7766156,2.349949,1.8609232,1.1618463,0.5874872,0.38400003,0.702359,1.5556924,2.5764105,2.556718,1.5195899,0.702359,0.34789747,0.63343596,1.2996924,1.7985642,1.2964103,1.467077,2.1333334,2.9997952,3.3280003,1.9364104,0.79097444,0.7515898,1.1716924,1.3489232,0.51856416,0.190359,0.12471796,0.20348719,0.318359,0.36758977,0.24287182,0.23958977,0.38728207,0.58420515,0.5940513,0.2297436,0.072205134,0.036102567,0.108307704,0.36758977,0.39056414,0.48902568,0.51856416,0.4660513,0.44307697,0.636718,0.5874872,0.45292312,0.3249231,0.2297436,0.20348719,0.17066668,0.23958977,0.380718,0.44307697,0.56451285,0.35774362,0.15097436,0.07548718,0.07548718,0.25928208,0.18707694,0.07548718,0.049230773,0.12143591,0.32820517,0.23630771,0.118153855,0.0951795,0.108307704,0.108307704,0.16082053,0.23958977,0.318359,0.36758977,0.37743592,0.45620516,0.48574364,0.4594872,0.47261542,0.48574364,0.7089231,0.7581539,0.67282057,0.9321026,0.4660513,0.56123084,1.079795,1.4112822,0.45620516,0.3117949,0.24615386,0.3249231,0.446359,0.33476925,0.22646156,0.21661541,0.14441027,0.013128206,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.016410258,0.016410258,0.009846155,0.016410258,0.07548718,0.27241027,0.36758977,0.43323082,0.47589746,0.4266667,0.47589746,0.43323082,0.3249231,0.18051283,0.04594872,0.13128206,0.24287182,0.21333335,0.07548718,0.07548718,0.3446154,0.6235898,1.3686155,1.8379488,0.09189744,0.1148718,0.10502565,0.12143591,0.23302566,0.48902568,0.45292312,0.39712822,0.36102566,0.36102566,0.39712822,0.41025645,0.4135385,0.4660513,0.5874872,0.74830776,0.5284103,0.45620516,0.42338464,0.37743592,0.3052308,0.45292312,0.5513847,0.42338464,0.13784617,0.016410258,0.016410258,0.016410258,0.059076928,0.15097436,0.25928208,0.35774362,0.46276927,0.512,0.48574364,0.4135385,0.508718,0.63343596,0.77456415,0.8533334,0.7318975,0.7089231,0.60061544,0.636718,0.7975385,0.80738467,0.77128214,0.86317956,0.85005134,0.73517954,0.74830776,0.636718,0.6465641,0.7089231,0.7515898,0.702359,0.761436,0.8598975,0.9944616,1.0436924,0.761436,0.77456415,0.8041026,0.88615394,0.9747693,0.9616411,0.79097444,0.8566154,0.9485129,0.9517949,0.8533334,0.96492314,1.083077,1.2176411,1.4145643,1.7558975,1.657436,1.6705642,1.7558975,1.8346668,1.785436,2.028308,2.3926156,2.294154,1.7624617,1.4342566,1.8379488,2.1202054,2.0644104,1.7887181,1.7394873,1.847795,1.8412309,1.9364104,2.0250258,1.6475899,1.3784616,1.7165129,2.2514873,2.5632823,2.1956925,2.868513,3.0654361,3.2787695,3.4822567,3.1277952,3.3247182,3.370667,3.6102567,3.8629746,3.4494362,3.7185643,5.156103,6.0849237,6.2096415,6.636308,6.4065647,5.651693,5.097026,4.8607183,4.4701543,4.201026,4.023795,4.023795,3.9942567,3.4330258,2.993231,2.737231,2.412308,2.0086155,1.7394873,1.3718976,1.3193847,1.5556924,1.9364104,2.166154,1.8970258,1.591795,1.3620514,1.1979488,0.97805136,1.1093334,1.5556924,1.8970258,2.100513,2.5009232,2.4057438,2.297436,2.1202054,2.103795,2.7634873,3.2623591,3.7907696,3.889231,3.43959,2.6715899,2.487795,2.294154,2.5632823,3.2262566,3.6758976,4.0303593,4.092718,4.3060517,4.522667,3.9975388,3.7907696,3.6758976,3.4592824,3.0785644,2.5796926,1.9922053,2.3762052,2.7306669,2.7208207,2.6847181,2.3926156,2.100513,1.847795,1.7427694,1.9364104,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.052512825,0.2100513,0.42338464,0.51856416,1.3620514,2.6223593,3.370667,3.2000003,2.2088206,2.0906668,2.284308,2.9078977,4.2535386,6.7840004,9.53436,12.002462,13.495796,14.181745,15.120412,18.294155,20.969027,20.292925,17.158566,16.193642,13.965129,11.585642,11.510155,13.545027,14.831591,12.028719,11.651283,13.046155,13.915898,10.315488,8.214975,7.64718,7.722667,8.3823595,10.423796,11.067078,10.955488,10.9226675,11.575796,13.29559,15.363283,17.329231,18.110361,17.58195,16.584206,14.946463,13.994668,12.704822,11.585642,12.635899,12.947693,12.553847,12.652308,13.942155,16.630156,20.821335,22.478771,22.62318,21.136412,16.722052,18.563284,21.556515,24.576002,26.112001,24.247797,24.139488,25.668924,26.43036,25.393232,22.882463,18.336823,14.477129,11.83836,10.338462,9.252103,9.068309,10.515693,12.727796,14.41477,13.866668,17.322668,27.418259,35.22954,35.856415,28.409437,25.938053,27.43795,26.65354,24.129642,27.237745,28.504618,26.788105,23.007181,18.81272,16.594053,13.098668,14.854566,17.227488,17.191385,13.308719,11.900719,13.75836,16.955078,19.876104,21.221745,18.819284,17.929848,17.493334,17.778873,20.38154,26.768412,29.80431,30.073439,29.863386,33.158566,32.256004,28.599796,24.195284,19.15077,11.67754,8.234667,6.6494365,5.976616,5.5565133,5.024821,4.6145644,3.9712822,3.4822567,3.4297438,4.007385,4.069744,4.197744,3.8071797,3.1770258,3.436308,3.8728209,3.7874875,3.3509746,2.8422565,2.665026,2.7306669,3.259077,4.0008206,4.9526157,6.3343596,6.669129,6.189949,6.47877,7.830975,9.232411,8.237949,8.43159,9.370257,11.227899,14.815181,18.12349,18.22195,21.924105,30.355694,38.95467,27.913849,16.298668,9.107693,7.3025646,7.8145647,10.9686165,13.650052,14.792206,14.532925,14.221129,14.431181,14.221129,16.508718,21.658258,27.460926,25.1799,19.265642,15.163078,13.945437,12.324103,9.097847,7.3025646,6.4722056,6.311385,6.685539,6.7971287,7.3419495,7.4436927,7.1154876,7.259898,7.7259493,9.475283,12.373334,15.199181,15.66195,13.492514,13.791181,16.984617,21.671387,24.605541,24.628515,28.580105,30.67077,29.062567,25.875694,23.292719,20.949335,17.440823,14.293334,15.9573345,18.451694,18.274464,17.302977,17.306257,19.974566,18.888206,14.907078,9.819899,5.8486156,5.6418467,10.226872,15.42236,24.136208,37.632004,55.54872,65.93642,70.67242,72.2478,71.552,67.84985,53.91754,43.063797,36.03036,32.213337,29.669746,30.030771,24.74995,21.78954,21.766565,17.920002,15.543797,17.483488,17.05354,13.29559,10.95877,9.816616,9.498257,10.41395,11.277129,9.130668,7.834257,9.222565,9.586872,7.896616,5.8157954,7.8080006,9.229129,8.763078,7.571693,9.275078,13.764924,14.040616,11.418258,8.480822,9.101129,10.443488,11.812103,13.049437,12.166565,5.333334,4.850872,4.9394875,4.7983594,4.397949,4.4767184,5.504,3.8859491,2.7109745,2.7437952,2.4549747,2.2777438,1.5360001,1.3522053,2.1464617,3.623385,2.9407182,3.0720003,3.0785644,2.858667,3.1540515,4.886975,5.398975,5.2578464,4.3684106,1.9889232,2.1169233,3.879385,7.00718,9.271795,6.485334,3.8498464,2.989949,3.5478978,4.6966157,5.142975,5.2447186,4.630975,5.2480006,6.2129235,3.8137438,2.5698464,3.5807183,4.2535386,3.9318976,3.9122055,2.9997952,2.878359,2.8947694,2.556718,1.5491283,1.3095386,1.4342566,1.8281027,2.3072822,2.5993848,2.2153847,2.353231,2.6157951,3.1606157,4.6867695,3.876103,3.8038976,4.2896414,4.7360005,4.1058464,2.5895386,2.4385643,2.8488207,3.1803079,2.937436,3.4231799,3.1967182,2.2580514,1.0896411,0.6465641,0.67610264,0.74830776,0.8467693,0.9124103,0.8205129,0.92553854,1.0338463,0.9353847,0.6629744,0.50543594,0.7089231,1.0568206,1.1749744,1.0338463,0.93866676,1.7690258,2.103795,2.03159,1.9823592,2.7273848,2.9013336,2.5796926,2.3860514,2.6617439,3.4625645,4.141949,4.8114877,5.2742567,5.1626673,3.9351797,3.7874875,3.5052311,3.2065644,3.0982566,3.4592824,3.5282054,3.2098465,2.0742567,0.67938465,0.5677949,1.2274873,1.6344616,1.4572309,0.8598975,0.48246157,0.3708718,0.7778462,1.4342566,1.8281027,1.1979488,0.8041026,0.8598975,1.2800001,1.723077,1.5721027,1.0896411,0.98133343,1.2504616,1.4539489,0.702359,0.33476925,0.34133336,0.5316923,0.7778462,1.014154,0.71548724,0.77128214,0.8402052,0.7417436,0.4594872,0.14441027,0.036102567,0.02297436,0.07548718,0.24287182,0.25928208,0.84348726,1.1093334,0.81394875,0.3708718,1.0338463,1.024,0.8730257,0.9682052,1.585231,0.60389745,0.18379489,0.08533334,0.16082053,0.35774362,0.5481026,0.5973334,0.49230772,0.27569234,0.052512825,0.07876924,0.12143591,0.09189744,0.02297436,0.049230773,0.14769232,0.14441027,0.14112821,0.190359,0.28882053,0.28882053,0.24287182,0.2100513,0.21661541,0.256,0.34789747,0.49230772,0.54482055,0.50543594,0.54482055,0.42994875,0.3446154,0.67282057,1.1355898,0.7975385,0.51856416,0.92225647,1.4802053,1.6213335,0.7253334,0.35446155,0.21333335,0.3511795,0.56123084,0.38400003,0.4397949,0.9714873,0.8598975,0.13784617,0.0,0.0,0.13784617,0.16410258,0.049230773,0.0032820515,0.0032820515,0.0032820515,0.0032820515,0.006564103,0.026256412,0.1148718,0.23302566,0.35446155,0.44307697,0.46276927,0.58092314,0.7253334,0.62030774,0.318359,0.19364104,0.13128206,0.118153855,0.2297436,0.34133336,0.13784617,0.23958977,0.5940513,0.7417436,0.5284103,0.09189744,0.08533334,0.0951795,0.13784617,0.27569234,0.6104616,0.574359,0.48246157,0.40697438,0.36430773,0.3249231,0.37415388,0.40369233,0.4135385,0.4135385,0.40697438,0.4594872,0.47589746,0.446359,0.37743592,0.29210258,0.4004103,0.5415385,0.45292312,0.17066668,0.03938462,0.029538464,0.01969231,0.029538464,0.07876924,0.19692309,0.43323082,0.6170257,0.6826667,0.6268718,0.5349744,0.39712822,0.43323082,0.62030774,0.82379496,0.8172308,0.8730257,0.8566154,0.78769237,0.7384616,0.8566154,0.9485129,0.81394875,0.69907695,0.6826667,0.6859488,0.5677949,0.508718,0.49230772,0.50543594,0.5546667,0.7056411,0.7220513,0.78769237,0.9353847,1.0568206,0.8533334,0.73517954,0.67282057,0.65312827,0.67938465,0.71548724,0.827077,0.9616411,1.0043077,0.7811283,0.73517954,0.8730257,1.0502565,1.2898463,1.7788719,1.7887181,1.5064616,1.3259488,1.4276924,1.7493335,1.7788719,1.8904617,1.8904617,1.7296412,1.5064616,1.6869745,1.9659488,1.9003079,1.5360001,1.4112822,1.5688206,1.8871796,1.9790771,1.785436,1.5622566,1.5688206,1.6410258,1.8084104,2.038154,2.2580514,2.6453335,2.7798977,2.8553848,3.0030773,3.2754874,3.5577438,3.3936412,3.2032824,3.0162053,2.484513,3.9056413,4.785231,5.0674877,4.9493337,4.8804107,4.4438977,4.588308,4.8049235,4.706462,4.0434875,3.82359,3.4100516,3.2787695,3.3608208,3.0424619,2.553436,2.1825643,1.8806155,1.6508719,1.5688206,1.3292309,1.3587693,1.5064616,1.6869745,1.8609232,1.6705642,1.4145643,1.1782565,0.9682052,0.7187693,1.0896411,1.4244103,1.6935385,1.8576412,1.8806155,1.723077,1.8084104,1.8543591,1.9298463,2.4320002,2.6387694,2.917744,3.0326157,2.8717952,2.4615386,2.3958976,2.7602053,3.2000003,3.501949,3.5905645,4.1222568,4.020513,3.948308,3.879385,3.117949,3.058872,2.6486156,2.5862565,2.7634873,2.2613335,2.0742567,2.1497438,2.3860514,2.6354873,2.6978464,2.297436,2.0808206,1.9035898,1.7952822,1.9626669,0.0,0.029538464,0.06564103,0.07548718,0.08861539,0.19364104,0.18379489,0.20348719,0.3117949,0.44307697,0.4135385,0.8205129,1.2865642,1.6475899,1.7985642,1.6804104,1.9331284,2.674872,4.023795,5.720616,7.138462,10.220308,13.167591,14.772514,15.963899,19.8039,27.556105,28.724516,26.151386,22.212925,18.819284,16.915693,14.460719,13.482668,13.952001,13.761642,11.523283,11.250873,11.218052,10.259693,7.781744,8.674462,8.057437,7.7259493,8.300308,9.219283,9.984001,10.354873,10.9915905,12.360206,14.713437,15.688207,16.272411,15.996719,14.907078,13.548308,11.634872,10.985026,10.315488,9.8363085,11.260718,11.296822,11.96636,14.27036,17.637745,19.908924,21.993027,22.57395,21.832207,20.01395,17.427694,18.310566,20.614565,22.90872,23.926155,22.577232,25.025642,26.2039,24.986258,21.53354,17.302977,13.794462,10.994873,9.344001,8.687591,8.28718,11.556104,14.946463,15.960617,14.762668,14.188309,20.634258,28.324104,36.069748,41.00267,38.583797,32.354465,31.917952,30.79549,27.700516,26.532104,24.802464,23.06954,21.10031,18.786463,16.118155,14.588719,15.27795,15.9343605,15.507693,14.168616,15.66195,15.415796,15.432206,16.534975,18.379488,16.94195,16.469334,16.354464,17.02072,19.91877,25.711592,27.539694,27.418259,27.680822,30.976002,30.611694,26.919386,20.594873,13.206975,7.194257,6.2129235,5.356308,4.670359,4.20759,4.023795,4.4438977,4.4865646,4.089436,3.56759,3.5938463,3.8038976,3.7284105,3.373949,2.9833848,3.0523078,3.3345644,3.639795,3.629949,3.314872,3.058872,3.629949,3.95159,4.0369234,4.4898467,6.5017443,7.312411,7.276308,8.211693,10.154668,11.372309,10.640411,9.370257,9.26195,11.027693,14.385232,17.135592,18.176,20.995283,25.586874,28.484924,20.95918,13.604104,9.284924,8.4512825,9.124104,11.493745,14.057027,15.169642,14.706873,14.070155,15.80636,17.91672,22.354053,28.228926,31.799797,28.051695,21.99631,17.667284,15.330462,11.493745,8.113232,6.803693,6.51159,6.567385,6.695385,6.9382567,7.430565,7.6701546,7.5913854,7.571693,8.795898,10.233437,12.678565,15.599591,17.125746,14.523078,15.816206,20.09272,24.687592,25.16677,25.271797,32.8599,42.87672,50.45826,50.95057,46.15877,45.18072,43.520004,39.83754,35.971283,32.938667,28.46195,24.342976,21.687796,20.90995,17.792002,12.747488,7.522462,3.6824617,2.6026669,3.9909747,7.5520005,14.985847,26.689644,41.750977,54.114464,58.85375,62.57231,66.816,68.07303,59.838364,55.085953,52.978874,51.37395,46.80862,42.400826,35.561028,29.417028,24.352823,18.028309,14.8480015,15.002257,15.330462,14.102976,11.004719,10.322052,10.84718,11.332924,11.099898,10.039796,10.555078,11.45436,10.55836,8.073847,6.5969234,7.827693,11.405129,15.970463,17.99549,11.805539,15.524104,17.253744,15.327181,10.952206,8.198565,12.130463,15.872002,17.969233,16.764719,10.384411,9.770667,7.9885135,5.5926156,3.5807183,3.4034874,4.6572313,3.6594875,10.04636,18.011898,6.3179493,5.9569235,3.442872,2.0939488,2.3827693,1.9331284,1.6771283,1.657436,1.6410258,1.8182565,2.7995899,4.5554876,4.457026,3.820308,3.0358977,1.5622566,2.0545642,2.8389745,3.8498464,4.644103,4.4077954,3.889231,4.522667,5.0051284,4.850872,4.3684106,5.1987696,5.674667,6.363898,7.3353853,8.15918,5.297231,4.201026,3.757949,3.3476925,2.858667,2.7536411,3.1474874,3.1671798,2.550154,1.657436,1.7690258,1.9856411,2.0841026,2.034872,2.0086155,2.156308,2.2678976,2.2219489,2.4385643,3.8859491,3.4756925,3.1671798,3.190154,3.3280003,2.92759,2.5009232,2.6190772,2.858667,2.9144619,2.609231,2.8947694,2.4385643,1.5556924,0.69251287,0.43323082,0.8172308,1.0896411,1.1224617,0.97805136,0.9321026,1.4178462,1.5097437,1.1749744,0.64000005,0.38728207,0.40697438,0.8402052,1.1552821,1.1388719,0.90584624,1.4309745,1.8510771,2.0020514,2.0020514,2.2646155,2.5271797,2.6289232,2.674872,2.9801028,4.0992823,5.110154,5.356308,5.658257,5.970052,5.3760004,4.2896414,3.6529233,3.511795,3.7743592,4.2338467,4.95918,4.827898,3.4691284,1.6016412,1.0371283,1.083077,1.020718,0.8369231,0.61374366,0.53825647,0.6498462,1.1913847,1.6607181,1.7165129,1.1749744,0.7122052,0.7187693,1.0666667,1.4408206,1.3522053,1.0338463,0.892718,0.97805136,1.0404103,0.5284103,0.34789747,0.3052308,0.35774362,0.446359,0.5152821,0.36430773,0.39384618,0.4135385,0.34133336,0.19692309,0.068923086,0.029538464,0.029538464,0.055794876,0.12143591,0.17066668,0.92225647,1.2176411,0.8336411,0.45292312,0.99774367,1.1093334,1.0010257,0.96492314,1.3653334,0.6498462,0.27569234,0.19692309,0.2986667,0.39056414,0.52512825,0.58420515,0.56451285,0.44307697,0.18379489,0.07548718,0.07876924,0.06564103,0.016410258,0.02297436,0.059076928,0.06564103,0.07548718,0.14112821,0.3446154,0.4266667,0.35446155,0.3052308,0.3117949,0.27569234,0.3052308,0.4594872,0.5874872,0.65641034,0.74830776,0.45620516,0.25271797,0.3511795,0.6071795,0.5513847,0.5021539,0.9321026,1.2077949,1.0633847,0.60061544,0.42338464,0.7778462,1.0732309,1.0436924,0.75487185,0.86646163,0.99774367,0.7778462,0.28225642,0.009846155,0.0032820515,0.068923086,0.08205129,0.02297436,0.0,0.036102567,0.02297436,0.01969231,0.029538464,0.006564103,0.059076928,0.0951795,0.17723078,0.30851284,0.41682056,0.5874872,0.7384616,0.7253334,0.54482055,0.3117949,0.20676924,0.12471796,0.15753847,0.25271797,0.21661541,0.16082053,0.4266667,0.46933338,0.2231795,0.08205129,0.068923086,0.08533334,0.13128206,0.23302566,0.44964105,0.44964105,0.43323082,0.41682056,0.39056414,0.31507695,0.3446154,0.39384618,0.45292312,0.48902568,0.4397949,0.52512825,0.4955898,0.446359,0.41682056,0.39056414,0.37743592,0.48246157,0.45620516,0.27241027,0.108307704,0.04594872,0.026256412,0.02297436,0.04594872,0.14769232,0.38728207,0.54482055,0.5874872,0.51856416,0.4004103,0.29210258,0.32820517,0.5218462,0.7778462,0.90256417,0.8533334,0.8533334,0.81066674,0.75487185,0.85005134,0.85005134,0.7122052,0.6268718,0.65312827,0.7253334,0.5907693,0.508718,0.45620516,0.44964105,0.574359,0.6498462,0.69251287,0.7318975,0.8041026,0.9747693,0.8795898,0.7515898,0.6826667,0.7253334,0.892718,0.8336411,0.8730257,0.9714873,1.0075898,0.80738467,0.8336411,0.8730257,0.94523084,1.1060513,1.4473847,1.3226668,1.1454359,1.0535386,1.1290257,1.3915899,1.6082052,1.8215386,1.8445129,1.7033848,1.6640002,1.6607181,1.8740515,1.8412309,1.5360001,1.3718976,1.4211283,1.5622566,1.595077,1.5163078,1.522872,1.785436,1.9626669,2.1300514,2.359795,2.7503593,2.7667694,2.7306669,2.9440002,3.1967182,2.7536411,3.3575387,3.2754874,2.934154,2.6223593,2.5074873,3.623385,4.164923,4.1189747,3.6660516,3.1770258,3.2886157,3.7448208,4.1124105,4.092718,3.5446157,3.3936412,3.006359,2.7142565,2.5829747,2.4155898,1.972513,1.7066668,1.6344616,1.6771283,1.6640002,1.4834872,1.4802053,1.4703591,1.404718,1.3653334,1.2438976,1.1454359,0.9911796,0.79097444,0.6301539,0.9911796,1.3686155,1.5786668,1.5524104,1.339077,1.2570257,1.4112822,1.4375386,1.3554872,1.5721027,1.8445129,2.2219489,2.4024618,2.3663592,2.3926156,2.1136413,2.537026,3.0654361,3.4231799,3.6332312,3.636513,3.511795,3.5249233,3.5807183,3.245949,2.7109745,2.1858463,2.2153847,2.5731285,2.300718,2.048,1.9364104,2.2482052,2.7963078,2.9013336,2.4681027,2.4713848,2.412308,2.231795,2.3269746,0.0,0.118153855,0.13784617,0.14112821,0.19364104,0.3511795,0.39384618,0.36430773,0.3314872,0.3249231,0.32820517,0.54482055,0.7122052,1.0305642,1.4605129,1.7165129,2.281026,3.18359,4.453744,5.9536414,7.387898,11.293539,14.864411,16.49231,17.28,21.041233,28.90831,31.30749,29.32513,24.776207,20.230566,18.051283,16.15754,15.126975,14.457437,12.583385,11.881026,11.392001,10.292514,8.569437,7.020308,7.860513,7.394462,7.250052,7.716103,7.762052,8.280616,8.858257,9.895386,11.451077,13.223386,13.013334,12.560411,11.956513,11.208206,10.240001,9.278359,9.567181,9.38995,8.907488,10.161232,10.738873,13.092104,17.975796,23.394463,24.635078,23.286156,22.255592,20.427488,18.120207,17.092924,17.618053,18.865232,20.660515,22.501745,23.542156,25.573746,24.923899,21.851898,17.463797,13.702565,11.933539,10.761847,10.624001,11.539693,13.121642,19.419899,21.625437,19.06872,15.035078,16.75159,24.07713,29.59426,41.06831,54.501747,54.15385,38.902157,33.430977,33.08636,33.08308,28.521029,24.004925,21.664822,20.158361,18.743795,17.28,17.795284,17.115898,15.944206,15.048206,15.291079,16.89272,14.818462,13.174155,13.456411,14.536206,14.03077,14.585437,15.547078,16.633438,17.952822,21.54995,22.127592,22.3639,24.136208,28.534157,28.100925,23.666874,16.643284,9.787078,7.1876926,6.2884107,5.024821,4.1813335,4.135385,4.854154,5.2611284,4.8114877,4.0369234,3.383795,3.2164104,3.9778464,3.9548721,3.5413337,3.0916924,2.930872,3.121231,3.7382567,4.276513,4.519385,4.5456414,4.9887185,4.7327185,4.6244106,5.362872,7.4732313,8.146052,8.211693,8.887795,10.164514,10.8307705,10.512411,9.078155,8.644924,9.892103,12.035283,14.424617,16.682669,19.400208,21.638565,20.94277,15.8654375,11.835078,9.632821,9.216001,9.711591,11.34277,13.059283,14.171899,14.677335,15.268104,19.849848,26.417233,33.237335,37.75672,36.62113,29.239798,23.007181,18.353231,14.628103,10.069334,7.325539,6.564103,6.6527185,6.882462,6.9710774,7.1089234,7.328821,7.4404106,7.456821,7.5881033,8.753231,10.725744,14.880821,19.961437,22.068514,16.154257,15.258258,17.545847,20.240412,19.61354,21.497438,31.4519,46.15221,59.19508,61.072414,55.3879,55.076107,54.43939,50.4878,42.93908,36.417645,30.001232,24.165745,19.11795,14.795488,10.712616,6.8299494,3.8071797,1.9068719,0.99774367,1.1848207,3.4756925,9.170052,17.959387,27.946669,36.614567,39.811287,45.17744,52.368416,53.041233,49.7559,51.659492,55.473236,57.389954,53.054363,46.664207,41.124107,33.683697,25.071592,19.505232,16.262566,14.102976,13.919181,14.319591,11.628308,10.932513,12.2617445,13.174155,12.977232,12.708103,14.41477,14.053744,11.923694,9.196308,7.939283,8.116513,13.925745,20.52595,22.948105,16.088617,20.624413,20.394669,17.844515,14.086565,8.891078,11.32636,15.766975,18.034874,17.132309,15.248411,14.057027,10.607591,6.7216415,3.826872,2.9440002,4.315898,3.6430771,15.087591,28.258463,8.198565,8.3823595,4.7556925,2.5042052,2.7109745,2.353231,1.5163078,1.8707694,2.1103592,2.048,2.5862565,3.4527183,2.8225644,2.0086155,1.4966155,0.94523084,1.7952822,2.4746668,2.428718,2.0053334,2.4484105,3.1934361,4.9329233,5.605744,4.7622566,3.56759,4.240411,5.277539,6.419693,7.9425645,10.686359,7.719385,5.037949,3.442872,2.8225644,2.1398976,2.4713848,3.1409233,3.255795,2.6486156,1.8838975,2.0873847,2.1366155,1.9561027,1.6278975,1.3915899,1.6836925,1.7952822,1.8051283,2.0578463,3.190154,2.9801028,2.5009232,2.0873847,1.8674873,1.7723079,2.4484105,2.9472823,2.9768207,2.6387694,2.409026,2.0578463,1.595077,1.1093334,0.74830776,0.71548724,1.4867693,1.4244103,1.083077,0.8369231,0.88287187,1.2931283,1.3259488,1.014154,0.5874872,0.48574364,0.47917953,0.8467693,1.2865642,1.5458462,1.401436,1.5163078,1.7920002,1.972513,1.9889232,1.9823592,2.1267693,2.4484105,2.6518977,2.865231,3.629949,5.1298466,5.464616,5.9930263,6.813539,6.744616,4.893539,4.092718,4.010667,4.315898,4.6966157,5.7764106,5.5762057,4.273231,2.6289232,1.9823592,1.5327181,1.1388719,0.95835906,0.94523084,0.8730257,1.086359,1.7887181,2.3138463,2.3368206,1.8510771,1.1158975,0.8763078,1.1290257,1.5130258,1.3095386,0.86646163,0.67938465,0.65312827,0.6104616,0.30851284,0.24943592,0.17394873,0.12143591,0.0951795,0.052512825,0.036102567,0.036102567,0.032820515,0.026256412,0.026256412,0.036102567,0.08533334,0.128,0.128,0.06564103,0.11158975,0.63343596,0.88287187,0.69579494,0.48246157,0.86646163,1.2471796,1.3161026,1.0765129,0.8467693,0.512,0.30851284,0.28225642,0.36758977,0.39056414,0.48246157,0.46276927,0.4594872,0.4594872,0.3249231,0.15753847,0.0951795,0.06235898,0.029538464,0.016410258,0.02297436,0.036102567,0.03938462,0.08861539,0.31507695,0.43323082,0.380718,0.36102566,0.39384618,0.318359,0.25271797,0.3314872,0.49887183,0.67610264,0.761436,0.47589746,0.26912823,0.15753847,0.16738462,0.3511795,0.38400003,0.63343596,0.6826667,0.48574364,0.380718,0.47589746,0.9944616,1.3029745,1.2635899,1.211077,1.0601027,0.90912825,0.77128214,0.5874872,0.2100513,0.04266667,0.0,0.0,0.0,0.0,0.036102567,0.029538464,0.055794876,0.08861539,0.0,0.029538464,0.013128206,0.052512825,0.17066668,0.32164106,0.48246157,0.5940513,0.6465641,0.60389745,0.4266667,0.32820517,0.26256412,0.23302566,0.2231795,0.20348719,0.118153855,0.34789747,0.446359,0.28882053,0.068923086,0.052512825,0.059076928,0.101743594,0.18051283,0.28225642,0.318359,0.36102566,0.39384618,0.4004103,0.3446154,0.3511795,0.38400003,0.4594872,0.5284103,0.47589746,0.49887183,0.46933338,0.46276927,0.48246157,0.46933338,0.3708718,0.41025645,0.446359,0.38728207,0.18379489,0.07548718,0.032820515,0.02297436,0.036102567,0.098461546,0.30851284,0.5152821,0.60389745,0.5481026,0.39384618,0.2855385,0.27241027,0.42338464,0.6859488,0.86646163,0.81394875,0.8205129,0.80738467,0.79097444,0.85005134,0.77456415,0.6629744,0.58420515,0.58092314,0.6892308,0.6301539,0.52512825,0.42338464,0.39712822,0.5481026,0.61374366,0.6498462,0.6498462,0.65969235,0.79097444,0.8992821,0.8205129,0.74830776,0.7975385,1.0108719,0.93866676,0.9156924,0.95835906,0.9878975,0.8402052,0.8795898,0.8960001,0.88287187,0.9124103,1.1224617,0.9682052,0.9419488,0.98461545,1.0765129,1.2504616,1.4867693,1.6377437,1.6049232,1.5195899,1.7165129,1.6902566,1.723077,1.6672822,1.5064616,1.3489232,1.2865642,1.3062565,1.3489232,1.4112822,1.5425643,1.7952822,1.9429746,2.1300514,2.4155898,2.7733335,2.8455386,2.6157951,2.674872,2.868513,2.300718,2.7733335,2.7700515,2.5829747,2.5173335,2.8750772,3.2722054,3.4756925,3.3050258,2.806154,2.2416413,2.6912823,3.239385,3.5478978,3.501949,3.1967182,3.0818465,2.7766156,2.428718,2.1366155,1.9495386,1.6640002,1.522872,1.5360001,1.6180514,1.6147693,1.529436,1.463795,1.3193847,1.1027694,0.9321026,0.8795898,0.88943595,0.827077,0.69579494,0.6301539,1.0010257,1.2471796,1.3128207,1.204513,0.99774367,0.9944616,1.1191796,1.0896411,0.95835906,1.1191796,1.404718,1.8838975,2.1103592,2.0939488,2.2777438,2.1103592,2.3105643,2.6978464,3.0982566,3.3542566,3.170462,3.006359,2.9505644,3.0326157,3.2295387,2.3991797,2.0808206,2.2547693,2.5993848,2.5009232,2.1366155,1.9823592,2.428718,3.1540515,3.1343591,2.7831798,2.6518977,2.4648206,2.2547693,2.3860514,0.0,0.17723078,0.14769232,0.14441027,0.24287182,0.35446155,0.50543594,0.49887183,0.34789747,0.190359,0.2855385,0.5513847,0.8008206,1.1979488,1.6738462,1.9200002,2.7044106,3.629949,4.640821,6.0619493,8.618668,12.327386,16.351181,18.58954,18.793028,18.550156,21.4679,26.916105,28.255182,24.644924,21.064207,17.575386,16.787693,17.08636,16.971489,15.051488,14.129231,12.6063595,11.162257,9.793642,7.830975,6.262154,6.242462,6.6428723,6.87918,6.928411,7.128616,7.322257,7.857231,8.677744,9.340718,9.048616,8.438154,7.9458466,7.7423596,7.706257,8.027898,9.344001,9.668923,9.02236,9.442462,11.293539,15.826053,23.151592,30.168617,30.58872,26.003695,23.171284,19.941746,16.531694,15.524104,17.243898,18.389336,20.17477,22.659285,24.746668,23.27631,20.804924,17.782156,14.838155,12.76718,11.723488,12.389745,14.267078,17.11918,21.001848,27.204926,25.632822,19.754667,15.176207,19.610258,25.718155,31.7079,49.414566,70.63303,67.09826,42.505848,30.280207,29.390772,32.79426,27.431387,21.622156,18.422155,18.005335,19.252514,19.754667,19.01949,18.304,16.984617,15.435489,15.031796,14.585437,12.514462,11.08677,10.633847,9.590155,9.997129,12.908309,16.210052,18.195694,17.56554,19.849848,19.718565,20.004105,22.226053,26.624002,24.33313,18.87836,12.99036,8.835282,7.9950776,5.973334,4.8016415,4.713026,5.4514875,6.2916927,5.579488,4.092718,3.0818465,2.993231,3.4494362,4.4274874,4.4340515,3.826872,3.1113849,2.934154,3.314872,4.1714873,5.080616,5.7534366,6.0291286,5.467898,4.7556925,5.1856413,6.8332314,8.55959,8.464411,8.136206,7.893334,7.9163084,8.2445135,7.90318,7.5946674,7.6603084,8.198565,9.078155,11.323078,14.208001,16.918976,18.228514,16.515284,12.586668,10.505847,9.498257,9.15036,9.40636,10.765129,11.661129,13.4859495,16.738462,21.014977,29.302156,39.79159,46.966156,47.4519,40.018055,27.831797,21.497438,16.922258,12.435693,8.786052,7.0925136,6.770872,6.9809237,7.2303596,7.394462,7.181129,7.1614366,6.9087186,6.567385,6.8233852,7.256616,9.957745,16.896002,25.110977,26.696207,16.715488,12.104206,10.8996935,11.237744,11.319796,14.70359,23.361643,34.71754,43.83508,43.428104,39.04985,38.85621,38.20308,34.724106,28.327387,23.584822,19.373951,15.156514,10.7848215,6.488616,3.3312824,1.785436,1.5261539,1.7526156,1.1848207,0.764718,1.9561027,5.687795,11.703795,18.556719,23.24677,25.600002,31.72431,39.089233,36.529232,33.00103,35.53477,40.677746,44.50462,42.627285,39.683285,36.83118,31.176207,24.49395,23.210669,19.538054,15.524104,14.368821,15.570052,14.890668,13.272616,14.890668,17.26031,18.65518,18.103796,19.045746,17.27672,14.63795,12.028719,9.426052,8.493949,15.474873,20.010668,19.96472,21.448206,29.18072,24.654772,19.419899,17.030565,13.036308,10.240001,12.343796,13.144616,12.435693,15.973744,14.500104,10.555078,6.688821,4.516103,4.71959,4.650667,3.892513,15.730873,28.816412,7.1647186,8.251078,4.818052,2.3762052,2.605949,3.3411283,1.6508719,2.6026669,3.3444104,3.0785644,3.0523078,2.8389745,1.7788719,1.0633847,0.92225647,0.6071795,1.2012309,2.2646155,2.477949,1.8051283,1.4966155,2.166154,3.8662567,4.6933336,4.0303593,2.540308,2.8127182,3.4297438,4.7294364,6.7610264,9.275078,7.893334,5.4482055,3.5774362,2.733949,2.166154,2.7076926,3.4724104,3.8662567,3.6102567,2.740513,2.4549747,1.9922053,1.6508719,1.4736412,1.2274873,1.0404103,1.0732309,1.3784616,1.9167181,2.5731285,2.4155898,2.034872,1.6443079,1.401436,1.4211283,2.3630772,2.8488207,2.7503593,2.3040001,2.1103592,1.3161026,1.1224617,1.0010257,0.86317956,1.0633847,1.7887181,1.3686155,0.82379496,0.65312827,0.8205129,0.75487185,0.7220513,0.60061544,0.45620516,0.54482055,0.62030774,0.9124103,1.4309745,1.9495386,2.0118976,2.0545642,2.169436,2.162872,2.034872,1.9856411,1.8707694,2.0906668,2.28759,2.3729234,2.546872,4.4800005,5.533539,6.6428723,7.584821,6.9842057,4.6112823,3.8367183,3.767795,3.9220517,4.20759,5.093744,4.7655387,3.948308,3.2754874,3.308308,2.7306669,2.0578463,1.7165129,1.6672822,1.4112822,1.5721027,2.3729234,3.170462,3.4560003,2.8521028,1.654154,0.9419488,0.9747693,1.4080001,1.2832822,0.65312827,0.4266667,0.380718,0.33805132,0.17066668,0.108307704,0.052512825,0.02297436,0.016410258,0.016410258,0.016410258,0.006564103,0.0032820515,0.0,0.0,0.029538464,0.13784617,0.2297436,0.2297436,0.0951795,0.0951795,0.19692309,0.35774362,0.47261542,0.39056414,0.75487185,1.394872,1.6771283,1.3653334,0.6301539,0.36102566,0.2986667,0.27897438,0.25271797,0.28225642,0.37415388,0.3314872,0.30851284,0.34789747,0.36758977,0.2297436,0.13784617,0.08533334,0.055794876,0.02297436,0.016410258,0.03938462,0.04594872,0.068923086,0.22646156,0.32820517,0.30194873,0.2986667,0.33805132,0.31507695,0.2231795,0.18051283,0.3052308,0.5218462,0.56451285,0.46933338,0.33805132,0.23302566,0.20348719,0.26584616,0.2297436,0.25928208,0.26912823,0.24615386,0.26912823,0.508718,0.69907695,0.8795898,1.1618463,1.7296412,1.1257436,0.95835906,1.0075898,1.0010257,0.5940513,0.256,0.1148718,0.049230773,0.006564103,0.0,0.0,0.013128206,0.072205134,0.118153855,0.0,0.0,0.0,0.01969231,0.07876924,0.19692309,0.29538465,0.4004103,0.4594872,0.48246157,0.5152821,0.446359,0.4397949,0.43323082,0.36102566,0.17394873,0.14769232,0.36430773,0.47261542,0.33805132,0.06564103,0.03938462,0.029538464,0.072205134,0.15097436,0.2231795,0.27897438,0.32164106,0.36758977,0.40369233,0.40369233,0.40369233,0.39712822,0.446359,0.508718,0.44964105,0.4201026,0.45292312,0.51856416,0.56451285,0.5316923,0.446359,0.4135385,0.45620516,0.47589746,0.28225642,0.15753847,0.06564103,0.026256412,0.036102567,0.055794876,0.22646156,0.5349744,0.7253334,0.69907695,0.512,0.3446154,0.24943592,0.33476925,0.5546667,0.73517954,0.78769237,0.8041026,0.8205129,0.8730257,0.98133343,0.8598975,0.69907695,0.55794877,0.4955898,0.5677949,0.64000005,0.5284103,0.37743592,0.3052308,0.4135385,0.5481026,0.5415385,0.512,0.54482055,0.67610264,0.9156924,0.9124103,0.827077,0.7844103,0.8533334,0.9156924,0.892718,0.8992821,0.92553854,0.8369231,0.77128214,0.84348726,0.8402052,0.79425645,0.955077,0.9189744,0.9517949,1.0633847,1.2406155,1.4441026,1.4473847,1.3423591,1.2242053,1.2373334,1.5655385,1.6607181,1.5064616,1.4112822,1.4145643,1.2570257,1.1716924,1.2537436,1.3718976,1.4703591,1.5688206,1.7001027,1.6902566,1.8051283,2.0808206,2.3302567,2.7011285,2.3204105,1.9331284,1.8740515,2.0775387,2.1169233,2.1103592,2.166154,2.412308,3.006359,2.937436,2.7733335,2.5961027,2.3991797,2.0808206,2.4320002,2.9801028,3.2032824,3.0490258,2.9243078,2.8356924,2.5895386,2.3401027,2.1136413,1.8051283,1.6836925,1.5589745,1.4375386,1.3522053,1.3718976,1.3456411,1.2340513,1.0502565,0.84348726,0.6892308,0.7122052,0.7253334,0.7089231,0.67282057,0.6859488,1.0929232,1.0535386,0.92553854,0.8566154,0.8041026,0.8205129,0.8730257,0.8533334,0.84348726,1.1323078,1.3161026,1.7755898,2.038154,2.0151796,1.9987694,2.156308,2.231795,2.4385643,2.733949,2.8160002,2.8553848,2.6715899,2.4615386,2.412308,2.7076926,2.041436,2.0578463,2.3630772,2.6518977,2.7076926,2.5435898,2.4648206,2.868513,3.4724104,3.2918978,2.9702566,2.4943593,2.0808206,1.9003079,2.0676925,0.0,0.0,0.0,0.06235898,0.15753847,0.18379489,0.45292312,0.6301539,0.48246157,0.15097436,0.15097436,0.4955898,1.2832822,1.9561027,2.2121027,2.028308,2.4320002,4.1813335,6.7610264,9.764103,12.87877,16.246155,20.404514,23.56513,24.021336,20.12554,18.881643,19.98113,21.763283,22.810259,21.940514,18.658463,19.065437,20.857437,22.66913,24.047592,18.615797,15.041642,12.619488,10.371283,7.0498466,6.183385,6.2227697,5.8256416,5.2545643,6.377026,6.2063594,5.717334,5.356308,5.654975,7.2172313,9.317744,8.907488,7.4141545,6.193231,6.547693,6.547693,7.1220517,8.470975,10.089026,10.771693,12.225642,17.696821,26.69949,35.029335,34.773335,29.72226,25.967592,21.218464,16.196924,14.634667,18.208822,21.576206,22.4919,20.450462,16.679386,11.625027,9.07159,8.484103,8.887795,8.851693,9.5835905,12.868924,16.311796,19.377232,23.40759,22.294975,17.926565,14.276924,13.725539,17.060104,23.62749,32.850056,52.594875,73.15365,67.24596,45.01662,30.926771,25.501541,24.024618,16.54154,14.647796,13.53518,15.82277,20.266668,21.743591,18.264616,16.315079,14.647796,13.177437,12.970668,11.506873,10.883283,10.151385,9.330873,9.429334,11.027693,15.842463,20.41436,22.373745,20.447182,21.461334,21.474463,21.792822,21.910976,19.531488,16.577642,13.210258,10.31877,7.6668725,3.9056413,3.7973337,3.82359,4.44718,5.290667,5.156103,3.9844105,3.5905645,3.6463592,3.9975388,4.670359,4.7294364,4.3618464,3.7185643,3.1803079,3.3280003,3.754667,4.821334,5.4153852,5.1987696,4.637539,3.0391798,3.4166157,4.8344617,6.413129,7.3386674,8.425026,8.129642,7.64718,7.427283,7.171283,6.7216415,6.488616,6.3967185,6.626462,7.6143594,9.895386,12.281437,13.860104,13.745232,11.047385,8.973129,8.123077,8.369231,9.245539,9.980719,10.627283,11.913847,15.642258,23.213951,35.62667,48.738464,56.96985,58.19734,51.52821,37.30708,23.588104,17.785437,14.739694,11.861334,9.140513,7.748924,7.4830775,7.64718,7.834257,7.9195905,7.2960005,7.1122055,6.3507695,5.077334,4.457026,4.713026,6.9743595,12.937847,19.764515,20.079592,11.684103,7.6701546,5.904411,5.32677,5.937231,7.522462,9.734565,12.137027,13.581129,12.179693,10.164514,9.91836,10.630565,10.896411,8.697436,5.733744,3.892513,2.7864618,2.0808206,1.4966155,0.8960001,0.5907693,1.6672822,3.2722054,2.6256413,1.1585642,1.5360001,3.764513,7.6570263,12.832822,17.033848,16.846771,20.709745,28.704823,32.561234,23.079386,21.044514,22.121027,23.256617,22.705233,28.688412,27.986053,26.551796,26.994873,28.593233,26.837336,19.879387,16.308514,18.615797,23.194258,19.93518,20.630976,22.636309,23.6439,21.668104,20.667078,18.090668,15.875283,13.833847,9.659078,8.070564,14.450873,18.320412,18.530462,23.253336,32.679386,28.39631,22.87918,21.17908,20.932924,12.425847,12.504617,12.566976,11.10318,13.702565,20.598156,15.750566,9.452309,7.8473854,12.924719,7.3452315,4.9526157,16.561232,29.151182,5.858462,7.0793853,4.46359,2.103795,1.9987694,4.073026,1.4867693,2.5435898,3.761231,3.9778464,4.332308,4.394667,2.8521028,1.9692309,1.9364104,0.8992821,0.49887183,0.90912825,1.7329233,2.556718,2.9604106,2.3630772,2.477949,2.6354873,2.4549747,1.8313848,1.6836925,1.9331284,2.0841026,2.5238976,4.5029745,4.332308,3.820308,3.4592824,3.2886157,2.8980515,4.194462,5.861744,7.0531287,7.072821,5.402257,4.1189747,2.681436,1.8412309,1.591795,1.1913847,0.94523084,1.1323078,1.5031796,1.8773335,2.1202054,1.8149745,1.5458462,1.401436,1.4834872,1.9232821,2.7175386,2.484513,2.1169233,1.8412309,1.204513,0.9616411,0.8369231,0.761436,0.83035904,1.2832822,1.0633847,0.9616411,0.85005134,0.7975385,1.0535386,0.7220513,0.6301539,0.58420515,0.51856416,0.51856416,0.65312827,0.92553854,1.1979488,1.4605129,1.8149745,2.281026,2.3958976,2.3335385,2.231795,2.1825643,1.8412309,2.0939488,2.1924105,2.1464617,2.7306669,4.3290257,5.6451287,6.9382567,7.4141545,5.2020516,2.4681027,1.3817437,1.2603078,1.4736412,1.4506668,1.5360001,1.4834872,1.9035898,3.0752823,4.9427695,4.588308,3.511795,2.6322052,2.2383592,1.9823592,1.972513,2.6453335,3.4592824,3.757949,2.793026,1.6804104,0.98133343,0.8598975,1.0666667,0.9321026,0.30851284,0.108307704,0.068923086,0.06235898,0.06235898,0.036102567,0.02297436,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.009846155,0.0,0.0,0.0,0.036102567,0.10502565,0.16738462,0.16738462,0.16738462,0.13128206,0.101743594,0.12143591,0.24287182,0.5481026,1.0272821,1.3161026,1.2012309,0.64000005,0.38400003,0.4135385,0.35774362,0.16082053,0.07548718,0.13784617,0.22646156,0.26256412,0.24287182,0.24287182,0.19692309,0.108307704,0.06564103,0.072205134,0.06235898,0.02297436,0.032820515,0.03938462,0.04266667,0.09189744,0.21333335,0.19692309,0.13128206,0.108307704,0.2297436,0.25271797,0.16738462,0.18051283,0.32164106,0.44307697,0.45620516,0.5021539,0.49887183,0.4135385,0.28882053,0.20348719,0.23958977,0.28225642,0.3052308,0.36758977,0.53825647,0.54482055,0.6892308,1.2537436,2.487795,1.7165129,1.0305642,0.96492314,1.2800001,0.9616411,0.8763078,0.571077,0.24615386,0.036102567,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016410258,0.07548718,0.12471796,0.23958977,0.3249231,0.380718,0.5021539,0.49230772,0.44307697,0.45620516,0.49230772,0.380718,0.29538465,0.26584616,0.25928208,0.22646156,0.09189744,0.04266667,0.029538464,0.06235898,0.12471796,0.19692309,0.28225642,0.34133336,0.39712822,0.45292312,0.48902568,0.49887183,0.5021539,0.571077,0.65641034,0.5940513,0.5940513,0.5874872,0.6170257,0.67610264,0.702359,0.761436,0.6235898,0.5316923,0.53825647,0.48902568,0.35446155,0.16410258,0.049230773,0.029538464,0.029538464,0.10502565,0.36102566,0.5546667,0.56123084,0.36758977,0.3052308,0.28882053,0.31507695,0.41682056,0.6859488,0.6629744,0.6662565,0.82379496,1.1290257,1.4342566,1.0666667,0.7581539,0.5677949,0.50543594,0.51856416,0.58092314,0.5874872,0.46276927,0.28225642,0.24287182,0.32820517,0.40697438,0.45620516,0.51856416,0.702359,0.8730257,0.99774367,1.017436,0.90256417,0.67282057,0.7318975,0.77456415,0.761436,0.7384616,0.82379496,0.702359,0.69907695,0.764718,0.8467693,0.86974365,0.8336411,0.92553854,1.1454359,1.4309745,1.6640002,1.5786668,1.5097437,1.339077,1.1388719,1.1749744,1.4080001,1.3357949,1.3620514,1.463795,1.2209232,1.1848207,1.2570257,1.3850257,1.4966155,1.4966155,1.9593848,2.156308,2.2121027,2.2350771,2.3204105,2.3696413,1.913436,1.3587693,1.1257436,1.6640002,1.9561027,2.0217438,1.9298463,1.9200002,2.3958976,2.3958976,1.9823592,1.8543591,2.0578463,1.9823592,2.3269746,2.6584618,2.7011285,2.484513,2.349949,2.3991797,2.2449234,2.1956925,2.2088206,1.8904617,1.7099489,1.4605129,1.2176411,1.0929232,1.2504616,1.020718,0.86974365,0.7844103,0.7253334,0.64000005,0.7515898,0.71548724,0.6465641,0.6498462,0.80738467,1.0272821,0.9353847,0.72861546,0.55794877,0.5349744,0.5218462,0.54482055,0.5874872,0.65641034,0.7778462,1.0601027,1.4769232,1.8116925,1.8773335,1.5097437,1.3161026,1.8970258,2.4484105,2.6322052,2.609231,2.3663592,2.3958976,2.609231,2.6945643,2.1202054,1.8281027,1.782154,1.9364104,2.2678976,2.793026,3.43959,3.4822567,3.3608208,3.3050258,3.3411283,2.609231,2.353231,2.2186668,2.044718,1.8609232,0.0,0.0,0.0,0.013128206,0.052512825,0.14769232,0.30851284,0.33476925,0.26912823,0.20020515,0.24943592,0.36758977,0.83035904,1.1782565,1.3128207,1.4933335,2.6190772,5.293949,8.641642,11.562668,12.731078,11.579078,11.992617,12.786873,12.931283,11.559385,13.252924,15.474873,18.924309,23.000618,25.77395,23.936003,27.464207,34.258053,40.49067,40.598976,27.864618,19.554462,14.395078,11.10318,8.4283085,7.824411,7.857231,7.8506675,7.4075904,6.4032826,6.2129235,6.997334,6.514872,4.886975,4.604718,4.2830772,3.9647183,3.5840003,3.4100516,4.056616,5.356308,6.62318,8.385642,10.456616,11.920411,14.339283,17.673847,22.721643,27.152412,25.498259,24.086977,22.268719,19.400208,16.23631,14.9398985,17.939693,19.321438,17.772308,13.853539,10.013539,8.044309,7.207385,6.6560006,6.373744,7.177847,9.219283,11.388719,13.51877,15.412514,16.853334,15.186052,13.525334,13.410462,15.409232,19.121233,23.893335,29.758362,37.796104,48.850056,63.533955,52.02708,38.12103,31.287798,30.32944,23.364925,21.129848,19.426462,18.582975,18.30072,17.618053,16.708925,14.989129,12.849232,11.067078,10.820924,11.798975,11.332924,10.774975,11.201642,13.410462,15.963899,19.977848,23.492926,24.740105,22.107899,24.136208,24.398771,24.260925,23.266464,19.127796,18.008617,13.190565,8.306872,5.097026,3.4067695,3.4133337,4.1878977,4.450462,3.9056413,3.2525132,3.498667,3.620103,3.8531284,4.2207184,4.5095387,3.7218463,3.639795,3.5872824,3.4198978,3.498667,3.8367183,4.0467696,4.0008206,3.6562054,3.0752823,3.5380516,4.2994876,5.2020516,5.9995904,6.3507695,6.422975,6.633026,6.701949,6.619898,6.6461544,6.488616,6.695385,7.1154876,7.515898,7.578257,8.825437,10.003693,10.410667,9.77395,8.277334,7.568411,7.2237954,7.604513,8.973129,11.493745,14.706873,20.233849,30.01108,43.20821,56.208416,62.6117,62.98257,57.373543,45.73867,27.93354,17.522873,13.50236,11.408411,9.43918,8.457847,8.139488,8.214975,7.824411,6.889026,6.124308,6.226052,6.5969234,6.3212314,5.2348723,3.9187696,3.754667,4.2929235,5.7796926,7.318975,6.885744,4.7655387,3.7218463,3.2853336,3.255795,3.6890259,4.3585644,4.890257,5.218462,5.225026,4.7294364,3.6824617,3.31159,3.2918978,3.2229745,2.6190772,1.7526156,1.1684103,0.8402052,0.69251287,0.60389745,0.43651286,0.35446155,0.77128214,1.5721027,2.1366155,1.5195899,1.529436,2.4976413,5.1659493,10.683078,21.697643,18.668308,20.151796,27.90072,26.886566,25.488413,21.786259,20.667078,22.777437,24.51036,23.45354,25.252104,24.654772,21.156105,19.026052,25.363695,26.74872,26.28267,29.568003,44.711388,45.377644,44.11077,41.734566,37.920822,31.189335,28.918156,23.138464,19.521643,17.732924,11.441232,9.970873,11.339488,13.925745,18.776617,29.61395,30.785643,31.59631,27.329643,20.906668,22.898874,16.305231,14.306462,14.857847,17.47036,23.223797,31.16308,23.712822,13.899488,9.419488,12.642463,7.6307697,4.896821,6.6527185,9.442462,4.138667,6.550975,3.7054362,1.2800001,1.273436,2.0118976,1.913436,3.1606157,3.5347695,3.6135387,6.75118,6.439385,3.1967182,1.3883078,1.9167181,2.2186668,0.8992821,0.6498462,0.9682052,1.4998976,2.0217438,1.9200002,1.7362052,1.404718,1.086359,1.148718,1.332513,1.4572309,1.3850257,1.522872,2.8160002,4.1878977,4.0434875,4.4734364,5.602462,5.5729237,8.12636,11.523283,14.555899,15.753847,13.397334,12.2617445,8.950154,5.3825645,2.6880002,1.1913847,0.9747693,1.0732309,1.1979488,1.2603078,1.3883078,1.3751796,1.6508719,2.1136413,2.4549747,2.1431797,1.5195899,1.3062565,1.276718,1.2898463,1.2800001,1.0338463,0.9321026,0.86317956,0.90256417,1.3062565,1.1158975,0.764718,0.72861546,1.0601027,1.394872,0.93866676,1.0338463,1.0338463,0.8041026,0.7253334,0.761436,1.1848207,1.6114873,1.8642052,1.975795,2.1858463,2.0250258,2.0939488,2.3762052,2.2186668,1.7985642,1.6869745,1.5556924,1.5819489,2.4516926,2.740513,2.9965131,3.3542566,3.436308,2.359795,1.0108719,0.50543594,0.56123084,0.7450257,0.48574364,0.58092314,0.79425645,1.0436924,1.463795,2.3926156,2.4681027,2.166154,1.5983591,1.1355898,1.3981539,2.5074873,3.6036925,3.8432825,3.1737437,2.3171284,1.6344616,1.1158975,0.73517954,0.508718,0.49230772,0.38728207,0.17394873,0.06564103,0.17723078,0.5481026,0.20348719,0.08533334,0.049230773,0.026256412,0.016410258,0.006564103,0.009846155,0.009846155,0.0,0.0,0.0,0.02297436,0.03938462,0.049230773,0.059076928,0.098461546,0.08533334,0.055794876,0.052512825,0.14769232,0.3249231,0.5152821,0.5677949,0.48246157,0.41025645,0.5152821,0.65312827,0.5546667,0.24615386,0.052512825,0.04594872,0.06564103,0.101743594,0.14441027,0.18379489,0.17394873,0.128,0.07548718,0.03938462,0.036102567,0.03938462,0.04266667,0.04594872,0.03938462,0.01969231,0.37415388,0.4266667,0.3249231,0.2100513,0.20348719,0.5907693,0.37415388,0.23630771,0.38400003,0.56451285,0.508718,0.7089231,0.7450257,0.53825647,0.33805132,0.15425642,0.15097436,0.17723078,0.18051283,0.18379489,0.3446154,0.53825647,0.7515898,1.079795,1.7066668,1.8051283,1.1684103,0.6432821,0.512,0.49887183,0.77456415,1.1881026,0.9682052,0.23302566,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.026256412,0.098461546,0.18051283,0.256,0.35774362,0.48246157,0.5021539,0.43651286,0.3511795,0.3708718,0.4594872,0.42994875,0.4660513,0.5513847,0.446359,0.14441027,0.04594872,0.04266667,0.09189744,0.2231795,0.27897438,0.3511795,0.4004103,0.43323082,0.48902568,0.49230772,0.65312827,0.8205129,0.88287187,0.75487185,0.6170257,0.54482055,0.52512825,0.5481026,0.5907693,0.56451285,0.5940513,0.6432821,0.6432821,0.47589746,0.4397949,0.23958977,0.072205134,0.01969231,0.029538464,0.07548718,0.30851284,0.46933338,0.5021539,0.56123084,0.6268718,0.41682056,0.256,0.3052308,0.56451285,0.512,0.6104616,0.9156924,1.2996924,1.4572309,0.92553854,0.64000005,0.48574364,0.4266667,0.50543594,0.6268718,0.6170257,0.508718,0.35774362,0.24287182,0.30851284,0.36102566,0.44307697,0.56451285,0.6892308,0.77128214,0.8467693,0.92225647,0.9485129,0.79425645,0.8041026,0.8795898,0.8205129,0.65969235,0.67610264,0.8566154,0.9156924,0.86646163,0.76800007,0.7220513,0.71548724,0.77128214,0.955077,1.3029745,1.8084104,1.6935385,1.5556924,1.4375386,1.3423591,1.211077,1.2373334,1.3161026,1.3292309,1.2438976,1.0994873,1.1093334,1.394872,1.5425643,1.4966155,1.5425643,1.7165129,2.0086155,2.556718,3.0194874,2.5862565,1.9429746,1.8215386,1.8018463,1.6935385,1.5163078,1.7690258,1.6869745,1.7099489,1.8674873,1.7362052,1.8838975,2.041436,2.1300514,2.2580514,2.740513,2.9440002,2.5337439,2.1136413,1.8871796,1.654154,1.5458462,1.654154,1.8018463,1.8412309,1.6607181,1.3883078,1.1355898,1.0404103,1.0994873,1.142154,0.86974365,0.7253334,0.69907695,0.7318975,0.71548724,0.6859488,0.7056411,0.7089231,0.7253334,0.8467693,0.8402052,0.6629744,0.446359,0.3117949,0.37415388,0.42338464,0.46933338,0.52512825,0.6104616,0.7417436,1.0502565,1.4473847,1.5491283,1.3423591,1.1815386,1.1224617,1.585231,1.9987694,2.1267693,2.0841026,1.8215386,1.7723079,1.8904617,2.038154,2.0118976,2.3433847,2.2777438,2.4746668,2.8947694,2.806154,3.3050258,3.3476925,3.308308,3.3378465,3.3542566,2.3762052,2.2416413,2.356513,2.359795,2.1169233,0.0,0.0,0.0,0.0,0.016410258,0.08205129,0.14441027,0.118153855,0.17066668,0.34133336,0.5415385,0.57764107,0.7417436,0.92553854,1.0699488,1.148718,1.6410258,3.3411283,5.4613338,7.200821,7.762052,6.9710774,6.885744,7.2205133,7.8441033,8.78277,12.114052,15.382976,19.652925,24.802464,29.535181,28.928001,34.87836,44.097645,50.93744,47.382977,31.409233,22.114464,17.14872,14.401642,11.995898,13.033027,13.755078,13.607386,12.045129,8.513641,7.6668725,7.2631803,6.0192823,4.1878977,3.5774362,2.868513,2.7044106,2.7798977,3.0162053,3.5610259,4.768821,6.170257,8.008205,9.954462,11.109744,14.838155,19.24595,22.856207,24.116514,21.376001,20.391386,19.666052,17.7559,14.979283,13.4400015,16.324924,16.193642,13.702565,10.203898,7.762052,6.770872,6.626462,6.5083084,6.491898,7.565129,9.977437,12.045129,13.3251295,13.66318,13.190565,12.642463,12.1238985,13.170873,16.114874,20.07631,23.03672,25.465437,28.92472,38.403286,62.303185,66.50093,59.43139,49.782158,40.933746,30.95631,25.524515,21.382566,18.084105,15.579899,14.244103,13.387488,11.388719,9.82318,10.180923,13.863386,15.625848,14.821745,15.510976,18.215385,19.889233,19.649643,20.299488,21.225027,22.144001,23.108925,27.369028,27.80554,26.427078,24.293745,21.51713,16.361027,10.47959,6.0291286,3.7316926,2.868513,2.8849232,3.7120004,4.2240005,4.161641,4.1517954,3.9220517,3.8695388,3.8662567,3.8695388,3.948308,3.6660516,3.6135387,3.446154,3.2229745,3.4034874,3.3542566,3.308308,3.3017437,3.2722054,3.062154,3.82359,4.309334,4.7425647,5.10359,5.152821,5.182359,5.5630774,5.8125134,5.83877,5.930667,5.835488,5.651693,5.661539,5.910975,6.2227697,6.99077,7.9917955,8.300308,7.7292314,6.8332314,7.315693,8.474257,10.6469755,13.99795,18.517334,24.822155,33.506466,43.779285,53.943798,61.40062,61.89949,57.58031,48.49231,35.44944,20.01395,13.200411,10.463181,8.966565,7.8539495,8.247795,8.008205,7.4699492,6.76759,6.1078978,5.7764106,6.1308722,7.522462,7.712821,6.409847,5.2480006,8.487385,8.034462,5.8912826,3.6824617,2.6322052,2.5173335,2.609231,2.537026,2.878359,5.152821,12.07795,15.655386,21.008411,26.446772,23.476515,19.922052,15.619284,10.755282,6.8397956,6.7282057,2.8192823,1.0108719,0.6170257,1.0601027,1.8740515,2.28759,2.0151796,1.3784616,0.9747693,1.657436,1.5556924,2.789744,3.4330258,3.5840003,5.3398976,11.323078,9.846154,12.045129,21.454771,33.99877,27.421541,21.871592,20.59159,22.229336,20.808207,18.668308,19.34113,18.169437,17.332514,25.869131,36.67036,49.06667,65.19795,85.68452,109.64349,104.635086,94.24411,78.56575,60.353645,45.0199,36.818054,28.498053,25.80677,25.678772,16.226463,13.371078,11.510155,11.648001,15.176207,23.834259,21.93395,28.310976,26.745438,18.28431,21.257847,18.34995,15.261539,15.00554,18.871796,26.41067,27.743181,22.757746,15.556924,9.603283,7.702975,5.8190775,6.560821,9.232411,10.496001,4.3585644,4.460308,3.9712822,4.31918,4.647385,1.8051283,3.0194874,5.973334,6.47877,5.159385,7.4469748,4.1058464,1.8051283,1.0371283,1.3850257,1.522872,1.086359,2.0578463,2.3696413,1.8904617,2.4155898,2.1792822,1.8248206,1.2209232,0.6859488,1.014154,0.94523084,0.86646163,0.8205129,1.0699488,2.1103592,2.9833848,3.255795,4.2535386,5.579488,5.106872,7.0137444,10.676514,14.486976,17.51959,19.524925,18.901335,14.290052,8.736821,4.201026,1.5392822,1.2931283,1.3062565,1.3062565,1.2242053,1.1946667,1.273436,1.4933335,1.782154,1.9265642,1.5655385,0.9616411,0.88287187,0.98133343,1.0699488,1.1126155,1.0666667,0.9485129,0.7975385,0.761436,1.1027694,1.2931283,1.0994873,1.1815386,1.7394873,2.5337439,1.8182565,1.5130258,1.719795,1.9068719,0.9156924,0.86317956,1.1782565,1.5622566,1.8707694,2.1234872,2.176,1.8609232,1.8182565,2.1103592,2.228513,1.8379488,1.6738462,1.4933335,1.3653334,1.6377437,1.6836925,1.5031796,1.4178462,1.4211283,1.1520001,0.4955898,0.4660513,1.0075898,1.5064616,0.7581539,0.4004103,0.69251287,0.9419488,0.94523084,1.0043077,1.2012309,1.2832822,1.0436924,0.69907695,0.88615394,2.041436,2.9636924,3.3772311,3.1507695,2.3072822,1.7394873,1.3423591,0.84348726,0.33476925,0.25271797,0.32164106,0.20020515,0.08861539,0.128,0.42338464,0.37743592,0.2100513,0.072205134,0.01969231,0.016410258,0.0032820515,0.0032820515,0.0032820515,0.0,0.0,0.0,0.006564103,0.009846155,0.006564103,0.013128206,0.032820515,0.029538464,0.016410258,0.016410258,0.059076928,0.14441027,0.23958977,0.36430773,0.52512825,0.69907695,0.5349744,0.4594872,0.35774362,0.21661541,0.128,0.04594872,0.02297436,0.032820515,0.059076928,0.0951795,0.07876924,0.055794876,0.029538464,0.02297436,0.059076928,0.055794876,0.059076928,0.055794876,0.03938462,0.009846155,0.33476925,0.48574364,0.50543594,0.43323082,0.318359,0.73517954,0.636718,0.4201026,0.2986667,0.3117949,0.2297436,0.3511795,0.4201026,0.3511795,0.24943592,0.13784617,0.098461546,0.101743594,0.118153855,0.09189744,0.190359,0.37415388,0.49887183,0.56123084,0.6859488,0.77128214,0.508718,0.24615386,0.14769232,0.20676924,0.37743592,0.7778462,1.0075898,0.8598975,0.33805132,0.068923086,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.026256412,0.07876924,0.14769232,0.20020515,0.31507695,0.38400003,0.34789747,0.256,0.23958977,0.36430773,0.40369233,0.47917953,0.6071795,0.7089231,0.37743592,0.15425642,0.049230773,0.068923086,0.20020515,0.27897438,0.34133336,0.39712822,0.45292312,0.50543594,0.5349744,0.6235898,0.7384616,0.81394875,0.7581539,0.65969235,0.6498462,0.702359,0.7318975,0.58420515,0.47589746,0.508718,0.5940513,0.6235898,0.46276927,0.47261542,0.29210258,0.12143591,0.049230773,0.03938462,0.06235898,0.23302566,0.42338464,0.57764107,0.69251287,0.5481026,0.36102566,0.24615386,0.26256412,0.42338464,0.5546667,0.81066674,0.98133343,1.024,1.079795,0.85005134,0.7220513,0.61374366,0.508718,0.4660513,0.55794877,0.5349744,0.48246157,0.42994875,0.35446155,0.28225642,0.28882053,0.35446155,0.4594872,0.57764107,0.75487185,0.99774367,1.2603078,1.4244103,1.3193847,0.8730257,0.81066674,0.8402052,0.8172308,0.761436,0.71548724,0.7811283,0.81066674,0.78769237,0.8041026,0.75487185,0.86317956,1.024,1.1815386,1.3522053,1.3259488,1.3653334,1.4211283,1.4145643,1.2668719,1.1749744,1.3062565,1.3686155,1.2832822,1.1585642,1.2209232,1.3883078,1.4703591,1.4539489,1.5392822,1.6344616,1.8642052,2.5009232,3.0424619,2.2153847,2.1825643,2.1956925,2.097231,1.847795,1.5163078,1.5786668,1.463795,1.5589745,1.8084104,1.7165129,1.6902566,1.9003079,1.9889232,2.0053334,2.409026,2.4746668,1.9856411,1.5885129,1.4867693,1.3981539,1.2209232,1.2898463,1.4736412,1.6246156,1.5753847,1.2832822,1.1257436,1.1257436,1.1749744,1.0404103,0.86974365,0.8730257,0.90256417,0.8795898,0.8041026,0.9288206,1.0371283,0.9878975,0.8172308,0.73517954,0.6170257,0.4397949,0.2986667,0.23958977,0.28882053,0.36430773,0.44307697,0.512,0.57764107,0.65969235,0.8533334,1.1224617,1.2832822,1.3522053,1.5556924,1.401436,1.4539489,1.6508719,1.8576412,1.8904617,1.7296412,1.7624617,2.028308,2.4057438,2.5862565,2.9505644,2.8488207,2.8455386,3.0030773,2.8914874,3.3017437,3.3969233,3.3214362,3.1409233,2.8521028,2.4910772,2.5107694,2.4976413,2.425436,2.6683078,0.0,0.0,0.0,0.0,0.006564103,0.026256412,0.036102567,0.068923086,0.16082053,0.318359,0.5284103,0.5316923,0.7220513,0.9878975,1.1323078,0.8730257,0.9321026,1.7690258,2.8816411,3.8564105,4.3618464,4.378257,4.453744,4.8738465,5.976616,8.172308,11.923694,15.356719,18.960411,22.938257,27.221336,28.038567,34.067696,41.934772,46.900517,42.85703,31.209028,24.103386,19.99754,17.673847,16.226463,18.162872,19.177027,18.674873,16.210052,11.500309,9.957745,8.835282,7.7259493,6.5050263,5.3169236,4.6572313,4.4800005,4.594872,4.903385,5.398975,6.491898,7.962257,9.780514,11.546257,12.481642,15.816206,20.437334,23.712822,24.054155,20.93949,19.938463,19.058874,17.45395,15.323898,13.909334,16.278976,16.032822,13.889642,11.178667,9.82318,8.759795,8.379078,8.582564,9.344001,10.70277,12.084514,14.36554,15.402668,14.280207,11.316514,11.277129,11.831796,14.132514,18.021746,22.042257,24.214975,25.366976,28.708105,38.79713,61.541748,78.19488,77.84698,64.925545,46.326157,31.428925,24.159182,19.977848,16.777847,13.843694,11.83836,10.28595,9.03877,9.3768215,12.068104,17.378464,18.668308,18.747078,20.368412,22.856207,22.117744,19.88595,18.497643,18.537027,20.404514,24.323284,29.213541,29.29231,26.932514,23.67672,20.243694,13.00677,7.8145647,4.8049235,3.5478978,3.045744,3.5872824,4.096,4.44718,4.670359,4.926359,4.57518,4.4242053,4.141949,3.7776413,3.7776413,3.8596926,3.69559,3.3345644,3.0523078,3.3411283,3.2131286,3.117949,3.2853336,3.6004105,3.5741541,3.889231,3.9614363,4.1058464,4.312616,4.266667,4.3684106,4.604718,4.7622566,4.821334,4.9460516,4.8147697,4.5029745,4.3684106,4.713026,5.7764106,6.5739493,7.5979495,8.257642,8.605539,9.340718,11.270565,13.344822,15.881847,19.18031,23.529028,30.20472,39.476517,48.590775,55.397747,58.354877,55.318977,47.661953,36.48985,23.955694,13.2562065,9.924924,8.490667,7.686565,7.27959,8.067283,7.781744,6.9645133,6.380308,6.232616,6.1440005,6.232616,7.8769236,8.372514,7.210667,6.0849237,8.979693,8.257642,5.730462,3.1967182,2.4320002,3.0523078,4.2502565,4.7556925,5.2512827,8.372514,15.8654375,19.731693,25.642668,31.30749,26.512413,23.43713,18.707693,12.950975,8.553026,9.672206,6.0849237,3.8990772,2.7831798,3.0326157,5.5597954,5.2053337,4.3552823,2.8258464,1.3522053,1.5885129,1.2373334,2.4648206,3.3411283,3.2722054,3.0030773,5.8880005,4.97559,5.792821,12.547283,28.1239,19.91549,17.532719,20.020514,23.056412,18.944002,18.628925,20.453745,18.901335,20.276514,42.68308,53.89457,67.34113,90.19406,121.49827,152.19858,137.92493,119.90319,97.30955,72.917336,53.090466,41.20944,31.730875,28.35036,27.894156,20.322464,16.09518,12.521027,10.817642,11.867898,16.187078,16.36431,26.535387,26.463182,16.66954,18.41559,18.294155,15.317334,14.670771,19.183592,29.315285,26.57149,21.572926,15.770258,10.197334,5.4875903,4.46359,6.229334,10.9226675,13.59754,4.2174363,2.8488207,3.1343591,4.450462,5.182359,2.7109745,6.961231,8.582564,8.79918,8.549745,8.484103,2.3762052,0.8205129,0.86974365,1.0765129,1.5163078,1.0404103,2.7044106,3.3805132,2.6322052,2.6847181,2.3696413,2.3433847,2.1924105,1.7624617,1.1782565,0.99774367,0.65641034,0.49887183,0.86317956,2.0873847,2.1956925,2.7798977,3.754667,4.5522056,4.1222568,5.4416413,7.4765134,9.938052,13.190565,18.251488,20.785233,17.637745,11.82195,5.9503593,2.228513,1.5786668,1.4966155,1.4473847,1.276718,1.1946667,1.2274873,1.2898463,1.4244103,1.4998976,1.204513,0.9156924,0.9911796,1.142154,1.2504616,1.3883078,1.2635899,1.1552821,1.0108719,0.92225647,1.1191796,1.404718,1.4539489,1.8182565,2.6026669,3.4789746,2.412308,1.719795,1.9626669,2.4320002,1.148718,0.9682052,1.1618463,1.4998976,1.847795,2.1924105,2.2186668,1.9003079,1.7066668,1.8543591,2.284308,1.9626669,1.6705642,1.4605129,1.3620514,1.3817437,1.4703591,1.1782565,1.0338463,1.1290257,1.1355898,0.9714873,0.86974365,1.5360001,2.3269746,1.214359,0.62030774,0.85005134,1.2209232,1.2898463,0.8402052,0.85005134,0.98461545,0.9321026,0.79097444,1.079795,1.467077,1.785436,2.231795,2.5304618,1.910154,1.4572309,1.2274873,0.827077,0.30194873,0.15097436,0.22646156,0.2231795,0.13784617,0.06235898,0.19364104,0.3249231,0.19692309,0.059076928,0.02297436,0.026256412,0.009846155,0.006564103,0.006564103,0.0032820515,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.009846155,0.02297436,0.016410258,0.03938462,0.09189744,0.24943592,0.5415385,0.955077,0.6662565,0.33805132,0.15097436,0.13456412,0.15753847,0.08205129,0.036102567,0.016410258,0.013128206,0.026256412,0.013128206,0.0032820515,0.0032820515,0.016410258,0.059076928,0.06564103,0.07548718,0.07548718,0.055794876,0.016410258,0.17723078,0.37743592,0.56123084,0.61374366,0.32820517,0.5874872,0.5940513,0.44964105,0.2986667,0.33476925,0.17066668,0.13456412,0.14769232,0.16738462,0.15753847,0.18707694,0.118153855,0.07548718,0.08533334,0.06564103,0.08861539,0.18379489,0.21989745,0.17066668,0.101743594,0.06564103,0.068923086,0.06564103,0.055794876,0.07876924,0.101743594,0.256,0.5513847,0.74830776,0.33805132,0.068923086,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02297436,0.059076928,0.072205134,0.12471796,0.190359,0.2100513,0.17394873,0.12143591,0.20020515,0.26256412,0.36102566,0.5284103,0.79425645,0.6498462,0.33805132,0.108307704,0.06564103,0.190359,0.2855385,0.34133336,0.40369233,0.48246157,0.5481026,0.574359,0.58420515,0.65312827,0.76800007,0.84348726,0.8533334,0.88615394,0.90584624,0.84348726,0.6268718,0.5284103,0.508718,0.5284103,0.5284103,0.43323082,0.44964105,0.2986667,0.14769232,0.06564103,0.03938462,0.052512825,0.16738462,0.36430773,0.571077,0.6859488,0.4594872,0.3052308,0.23958977,0.256,0.30851284,0.58420515,0.8467693,0.88943595,0.78769237,0.892718,0.86646163,0.7811283,0.67938465,0.58092314,0.48574364,0.5218462,0.55794877,0.5546667,0.508718,0.45292312,0.28882053,0.256,0.30194873,0.38728207,0.47917953,0.6662565,0.9682052,1.2570257,1.4441026,1.4966155,1.1815386,1.0371283,1.0043077,1.0075898,0.9419488,0.636718,0.6071795,0.6892308,0.7778462,0.8369231,0.761436,0.9156924,1.0502565,1.0699488,1.0404103,1.0765129,1.2242053,1.3489232,1.3587693,1.2307693,1.0896411,1.211077,1.3128207,1.3062565,1.276718,1.2635899,1.2504616,1.2898463,1.3653334,1.3850257,1.4834872,1.7099489,2.2055387,2.5731285,1.8609232,2.162872,2.2514873,2.169436,1.9692309,1.7066668,1.595077,1.5655385,1.6640002,1.782154,1.657436,1.4703591,1.5983591,1.6738462,1.6804104,1.9561027,1.8871796,1.5195899,1.2865642,1.3095386,1.3981539,1.3620514,1.2471796,1.2832822,1.4408206,1.4342566,1.1913847,1.1881026,1.2438976,1.1946667,0.8992821,0.955077,1.0108719,1.014154,0.9682052,0.96492314,1.0765129,1.1520001,1.083077,0.8763078,0.62030774,0.4660513,0.33805132,0.26912823,0.25928208,0.28225642,0.37415388,0.47261542,0.571077,0.63343596,0.60389745,0.6859488,0.9353847,1.1355898,1.2865642,1.5983591,1.4473847,1.3489232,1.4145643,1.6377437,1.8904617,1.7887181,1.8642052,2.1333334,2.5074873,2.7831798,3.0162053,2.9604106,2.9440002,3.0391798,3.0720003,3.3772311,3.4625645,3.3280003,3.0194874,2.6322052,2.7766156,2.809436,2.612513,2.3926156,2.678154,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.12471796,0.17066668,0.13456412,0.23958977,0.23630771,0.67938465,1.086359,1.1257436,0.62030774,0.82379496,1.5491283,2.540308,3.4756925,3.9614363,3.7087183,3.5938463,3.9876926,5.182359,7.381334,10.640411,13.400617,15.412514,17.03713,19.209848,21.32677,25.554052,29.600822,31.809643,31.153233,28.018873,24.178873,20.785233,18.822565,19.131079,20.647387,21.136412,20.132105,17.545847,13.656616,11.956513,11.674257,11.628308,11.07036,9.691898,9.38995,9.281642,9.55077,10.056206,10.322052,11.628308,13.321847,14.8939495,16.059078,16.761436,17.509745,20.575182,23.88677,25.173336,21.976618,21.986464,20.824617,19.590565,18.678156,17.785437,19.285336,20.079592,19.259079,17.319386,16.134565,13.879796,12.35036,12.048411,12.980514,14.660924,14.818462,17.227488,17.979078,15.488001,10.509129,10.791386,12.885334,16.902565,21.979898,26.262976,27.75631,29.522053,34.21867,43.267284,56.82216,76.39632,78.299904,64.08862,41.49826,24.451284,18.678156,16.856617,15.616001,13.456411,10.765129,8.812308,9.357129,11.861334,15.350155,18.392616,19.27877,20.929642,22.272001,22.09477,19.049026,17.457232,17.106052,18.454975,21.471182,25.622976,28.468515,27.224617,24.274054,20.292925,14.227694,9.32759,6.173539,4.670359,4.2863593,4.0369234,5.3398976,5.3037953,5.0149746,4.955898,5.0182567,5.024821,4.900103,4.5456414,4.096,3.9089234,3.7842054,3.6069746,3.3509746,3.1803079,3.442872,3.5741541,3.564308,3.876103,4.3684106,4.2830772,4.135385,3.9745643,4.0434875,4.2272825,4.0434875,3.7809234,3.6758976,3.6496413,3.6857438,3.8498464,3.895795,4.279795,4.788513,5.7009234,7.785026,9.409642,10.735591,11.795693,13.121642,15.744001,18.6519,20.486567,21.602463,22.869335,25.672207,30.818464,38.63959,46.286774,51.33785,51.797337,46.306465,36.31262,24.6679,14.332719,8.379078,7.7292314,7.4371285,7.253334,7.197539,7.5520005,7.276308,6.8397956,6.7183595,6.882462,6.803693,6.8594875,7.972103,8.385642,7.53559,6.0291286,4.647385,3.9548721,3.4231799,3.0654361,3.442872,4.4767184,6.6395903,7.7259493,7.958975,10.006975,11.940104,13.019898,14.129231,14.329437,10.850462,12.347078,11.506873,9.990565,9.298052,10.765129,10.880001,9.127385,6.8594875,6.0685134,9.38995,7.3485136,5.651693,3.7874875,2.100513,1.8018463,0.90912825,0.892718,2.044718,3.6562054,4.013949,8.208411,6.7872825,4.84759,5.677949,10.765129,8.438154,12.150155,19.275488,24.65149,20.555489,23.095797,27.369028,26.056208,27.339489,54.90544,67.81703,74.02667,88.270775,113.86749,142.74626,126.87755,110.73642,93.56473,75.8318,59.2279,47.40267,36.870567,29.449848,25.24554,22.639591,17.51631,13.538463,11.234463,10.788103,12.045129,16.085335,26.482874,26.811079,17.683693,16.7319,16.932104,14.788924,14.503386,19.643078,33.14544,32.59077,25.616413,18.993233,14.605129,9.43918,5.730462,4.46359,7.5881033,10.748719,3.308308,2.300718,1.3259488,1.2307693,2.100513,3.2722054,9.813334,8.418462,8.5202055,11.168821,9.035488,2.349949,0.90912825,1.020718,1.2274873,2.3105643,0.80738467,2.225231,3.9712822,4.3585644,2.5862565,3.2328207,3.4724104,3.698872,3.5610259,1.9692309,1.6082052,0.955077,0.5481026,0.8467693,2.2219489,2.1398976,2.865231,3.43959,3.6168208,3.8695388,5.221744,4.9526157,5.1265645,6.957949,10.843898,16.09518,16.272411,12.553847,7.066257,2.8816411,1.6246156,1.4375386,1.404718,1.2242053,1.214359,1.1520001,1.204513,1.4703591,1.7066668,1.3095386,1.1684103,1.394872,1.6049232,1.7493335,2.097231,1.6607181,1.5425643,1.5097437,1.467077,1.467077,1.463795,1.5753847,2.162872,3.0358977,3.4592824,2.3105643,1.5688206,1.6344616,2.03159,1.401436,1.0601027,1.1454359,1.4441026,1.7887181,2.028308,2.2350771,2.1202054,1.9167181,1.8773335,2.2678976,2.028308,1.5983591,1.3686155,1.4998976,1.9396925,2.0151796,1.6869745,1.5753847,1.7657437,1.8051283,1.9462565,1.4112822,1.6738462,2.3926156,1.4112822,0.9353847,0.9911796,1.4375386,1.8281027,1.3883078,1.1224617,1.1749744,1.1684103,1.1782565,1.7394873,1.3095386,0.9353847,1.014154,1.3357949,1.0699488,0.7975385,0.8041026,0.636718,0.27897438,0.12143591,0.15425642,0.2100513,0.15425642,0.036102567,0.072205134,0.09189744,0.055794876,0.03938462,0.055794876,0.06564103,0.026256412,0.01969231,0.026256412,0.026256412,0.016410258,0.016410258,0.006564103,0.0,0.0,0.0,0.0,0.0,0.01969231,0.04266667,0.013128206,0.0032820515,0.01969231,0.07876924,0.29210258,0.86646163,0.82379496,0.40369233,0.0951795,0.055794876,0.11158975,0.101743594,0.059076928,0.02297436,0.0032820515,0.0,0.0032820515,0.006564103,0.013128206,0.01969231,0.029538464,0.06564103,0.07876924,0.08533334,0.07548718,0.029538464,0.01969231,0.17066668,0.43323082,0.58420515,0.21661541,0.256,0.26584616,0.27569234,0.3511795,0.60389745,0.37415388,0.25271797,0.16738462,0.10502565,0.101743594,0.26912823,0.18051283,0.08533334,0.07548718,0.08861539,0.04594872,0.052512825,0.068923086,0.07876924,0.08205129,0.0951795,0.1148718,0.128,0.118153855,0.055794876,0.108307704,0.072205134,0.02297436,0.0,0.0,0.006564103,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0,0.029538464,0.068923086,0.09189744,0.06235898,0.072205134,0.0951795,0.19364104,0.39712822,0.69579494,0.8730257,0.5513847,0.2100513,0.08205129,0.18379489,0.29538465,0.36102566,0.4135385,0.48574364,0.58420515,0.57764107,0.60061544,0.69251287,0.85005134,1.024,1.0666667,1.0732309,0.9714873,0.79097444,0.6859488,0.6629744,0.574359,0.47917953,0.41025645,0.37743592,0.39384618,0.2986667,0.17066668,0.068923086,0.036102567,0.04266667,0.13128206,0.27241027,0.43651286,0.56451285,0.48574364,0.32164106,0.24943592,0.28882053,0.30194873,0.61374366,0.7220513,0.7384616,0.79097444,1.0305642,0.9321026,0.7778462,0.65641034,0.5973334,0.5513847,0.5349744,0.65969235,0.67282057,0.5513847,0.48574364,0.3446154,0.28225642,0.30194873,0.37415388,0.42338464,0.512,0.7122052,0.86974365,0.9878975,1.2274873,1.4966155,1.4276924,1.2406155,1.086359,1.024,0.67282057,0.5218462,0.5513847,0.67938465,0.7417436,0.702359,0.8598975,0.98133343,1.014154,1.0896411,1.148718,1.2373334,1.273436,1.2209232,1.0929232,0.9616411,1.0469744,1.1520001,1.211077,1.2996924,1.1913847,1.1158975,1.1716924,1.273436,1.1881026,1.2668719,1.5360001,1.8051283,1.9035898,1.6508719,1.7329233,1.8806155,2.044718,2.1234872,1.9429746,1.7526156,1.7887181,1.8149745,1.7033848,1.4342566,1.273436,1.3522053,1.4408206,1.5163078,1.7690258,1.5983591,1.3456411,1.214359,1.2865642,1.4998976,1.6705642,1.404718,1.2570257,1.3226668,1.2668719,1.0929232,1.1848207,1.2537436,1.1355898,0.78769237,1.0469744,1.0535386,1.0043077,1.020718,1.1323078,1.0404103,0.9682052,0.9321026,0.8533334,0.54482055,0.41025645,0.34133336,0.31507695,0.32820517,0.38728207,0.52512825,0.6301539,0.7318975,0.77456415,0.6268718,0.6268718,0.892718,1.0338463,1.020718,1.1782565,1.1651284,1.211077,1.2603078,1.404718,1.8806155,1.7591796,1.8642052,1.9692309,2.0644104,2.3663592,2.5074873,2.6157951,2.8225644,3.117949,3.3509746,3.5216413,3.5216413,3.3805132,3.1409233,2.8553848,2.9801028,2.878359,2.609231,2.284308,2.0873847,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08205129,0.08205129,0.04266667,0.21333335,0.2986667,0.71548724,0.86646163,0.6432821,0.4135385,0.55794877,1.1716924,2.0250258,2.789744,3.0227695,2.8389745,2.7470772,3.058872,3.9286156,5.356308,7.7357955,9.878975,11.136001,11.631591,12.251899,14.536206,17.624617,19.206566,19.666052,22.09477,21.362873,18.251488,16.065641,16.226463,18.264616,19.009642,18.379488,16.561232,14.280207,12.803283,12.022155,13.380924,13.833847,13.413745,15.258258,16.968206,17.742771,19.114668,20.565334,19.515078,20.663797,22.708515,23.292719,22.180105,21.241438,18.297438,20.273232,23.985233,25.770668,21.50072,23.758772,24.835283,25.176617,24.976412,24.169027,25.426054,26.985027,28.04185,28.035284,26.656822,20.89354,17.266872,14.710155,13.426873,14.8939495,16.515284,18.84554,17.831387,13.59754,10.436924,13.988104,17.631182,22.130873,27.520002,33.112617,31.159798,32.63672,36.89354,41.30462,41.3079,49.91344,47.6718,38.094772,25.954464,17.273438,16.039387,14.762668,14.024206,13.4170265,11.536411,9.826463,11.661129,14.17518,15.681643,15.671796,18.491077,19.59713,19.085129,17.401438,15.350155,16.131283,19.495386,22.088207,23.424002,25.878977,24.684309,20.74913,16.817232,13.203693,7.781744,6.7216415,4.7524104,4.3716927,5.464616,5.293949,6.380308,5.5893335,5.0477953,5.481026,6.226052,5.0904617,4.466872,4.3651285,4.312616,3.370667,3.0916924,3.387077,3.6693337,3.7120004,3.6627696,3.8334363,4.315898,4.955898,5.4908724,5.540103,5.3924108,5.284103,5.412103,5.47118,4.6539493,3.3476925,2.930872,2.8882053,2.934154,3.006359,3.9811285,5.901129,7.6603084,9.517949,13.108514,16.97477,19.876104,21.225027,21.714052,23.299284,24.848412,25.721437,26.010258,26.916105,30.762669,37.366158,44.24534,48.90585,49.34236,44.022156,33.010876,22.787283,14.6871805,9.429334,7.1122055,7.3682055,7.194257,6.764308,6.380308,6.4557953,5.7107697,5.661539,5.979898,6.5837955,7.643898,9.43918,10.436924,10.095591,8.556309,6.6527185,4.273231,3.045744,2.7602053,3.3444104,4.8836927,4.8836927,5.835488,5.907693,5.113436,5.293949,7.5913854,9.645949,10.384411,10.499283,12.452104,18.369642,20.04349,22.180105,24.1559,20.017233,18.724104,14.811898,11.211488,9.232411,8.55959,6.314667,3.6660516,2.2744617,2.1431797,1.6180514,1.2635899,1.585231,2.4418464,3.2196925,2.8521028,3.9154875,6.1407185,6.7150774,6.636308,10.725744,12.924719,16.256,20.883694,24.339695,21.546669,27.30667,27.457644,26.217028,28.488207,39.840824,66.85539,73.54421,76.31754,82.00206,87.8638,94.55262,97.18483,94.36883,87.58482,81.17498,69.162674,54.432823,40.113235,29.233232,24.704002,18.563284,15.333745,13.161027,11.654565,11.88759,14.854566,20.594873,23.095797,21.188925,18.54031,16.121437,14.355694,14.148924,18.852104,34.254772,39.443695,37.097027,32.797543,27.808823,19.058874,11.405129,6.11118,4.33559,4.663795,3.1113849,1.9396925,0.9517949,0.5677949,0.8172308,1.3423591,1.5753847,2.7503593,5.477744,7.8408213,5.3858466,1.2471796,1.2668719,1.8215386,1.5655385,1.4178462,0.49230772,2.3466668,6.6428723,9.419488,3.0982566,7.017026,5.973334,4.3716927,4.056616,4.2863593,2.5435898,1.5195899,1.0994873,1.1946667,1.7690258,1.9528207,2.674872,3.2754874,3.636513,4.210872,5.408821,5.0215387,5.3858466,6.373744,5.3858466,4.44718,5.8223596,6.8660517,6.0061545,2.7470772,1.3423591,1.0469744,1.1027694,1.1520001,1.2504616,1.1290257,1.3259488,1.7657437,2.028308,1.3587693,1.4309745,1.8051283,2.1366155,2.3269746,2.546872,2.1202054,1.8215386,1.8510771,2.0545642,1.9068719,1.6869745,1.467077,1.6443079,2.044718,1.9232821,1.6410258,1.2340513,1.148718,1.401436,1.5721027,1.0962052,0.90256417,1.014154,1.2832822,1.4178462,2.103795,2.5107694,2.5731285,2.3171284,1.8773335,1.7558975,1.6705642,1.5885129,1.7690258,2.7470772,2.8324106,2.3236926,1.913436,1.9856411,2.609231,2.4024618,1.8642052,1.5425643,1.5327181,1.4966155,1.1290257,0.90912825,1.0732309,1.4736412,1.5721027,1.3653334,1.5425643,1.6016412,1.5195899,1.7394873,1.7394873,1.0994873,0.7384616,0.7778462,0.5349744,0.33805132,0.54482055,0.5513847,0.26912823,0.12143591,0.08533334,0.059076928,0.032820515,0.013128206,0.0,0.0,0.009846155,0.068923086,0.15097436,0.15097436,0.04266667,0.04266667,0.072205134,0.08861539,0.07548718,0.026256412,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.026256412,0.032820515,0.08533334,0.36758977,0.6465641,0.38728207,0.11158975,0.03938462,0.07548718,0.07548718,0.059076928,0.032820515,0.013128206,0.0,0.02297436,0.03938462,0.03938462,0.029538464,0.029538464,0.055794876,0.052512825,0.059076928,0.07876924,0.09189744,0.029538464,0.016410258,0.0951795,0.20348719,0.16738462,0.068923086,0.055794876,0.072205134,0.15097436,0.39712822,0.3708718,0.40369233,0.2986667,0.08861539,0.016410258,0.27241027,0.19692309,0.108307704,0.11158975,0.13784617,0.07548718,0.032820515,0.06564103,0.15425642,0.2297436,0.19364104,0.15425642,0.18051283,0.20020515,0.029538464,0.2986667,0.21989745,0.072205134,0.0,0.0,0.036102567,0.01969231,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.07876924,0.256,0.48902568,0.97805136,0.71548724,0.318359,0.108307704,0.12143591,0.29210258,0.3708718,0.40369233,0.43651286,0.5349744,0.55794877,0.6465641,0.78769237,0.9517949,1.0994873,0.9156924,0.85005134,0.8205129,0.7844103,0.74830776,0.7220513,0.5349744,0.37415388,0.318359,0.3052308,0.37743592,0.37743592,0.27569234,0.12143591,0.06235898,0.049230773,0.101743594,0.18051283,0.28225642,0.44307697,0.49230772,0.36758977,0.318359,0.4135385,0.5349744,0.86317956,0.892718,0.8795898,0.9714873,1.1913847,0.9353847,0.84348726,0.761436,0.6498462,0.56451285,0.47917953,0.5481026,0.5481026,0.4594872,0.47261542,0.4594872,0.34789747,0.27569234,0.28882053,0.3511795,0.44964105,0.6301539,0.7811283,0.8960001,1.0666667,1.1060513,1.2242053,1.1979488,0.9878975,0.7318975,0.5874872,0.44964105,0.40697438,0.48574364,0.65641034,0.7056411,0.86317956,1.0043077,1.0896411,1.1749744,1.3226668,1.3292309,1.2438976,1.1060513,0.94523084,0.8730257,0.9353847,1.017436,1.0568206,1.0666667,1.1520001,1.276718,1.3259488,1.2832822,1.2373334,1.2471796,1.3522053,1.3883078,1.3095386,1.1749744,1.4933335,1.654154,1.8674873,2.0676925,1.9068719,1.6738462,1.5261539,1.4145643,1.3718976,1.4966155,1.5195899,1.5425643,1.5688206,1.5983591,1.6475899,1.4769232,1.3620514,1.2504616,1.2406155,1.5721027,1.595077,1.4276924,1.3850257,1.4605129,1.3259488,1.1454359,1.0699488,1.0765129,1.0666667,0.88615394,1.0666667,1.142154,1.2209232,1.2800001,1.1454359,1.020718,0.892718,0.79425645,0.69251287,0.47261542,0.37415388,0.36102566,0.38400003,0.4594872,0.65641034,0.9485129,1.0601027,1.0272821,0.90584624,0.74830776,0.60061544,0.574359,0.69579494,0.90912825,1.0666667,1.0568206,1.0699488,1.0962052,1.2077949,1.5885129,1.463795,1.8281027,1.9626669,1.8051283,1.9364104,2.0118976,2.359795,2.681436,3.0096412,3.692308,3.764513,3.7185643,3.6758976,3.5511796,3.0523078,2.733949,2.553436,2.3269746,1.9889232,1.5885129,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016410258,0.03938462,0.08533334,0.190359,0.20676924,0.35446155,0.42338464,0.38400003,0.38728207,0.58420515,1.1126155,1.6508719,2.0118976,2.1530259,2.353231,2.3204105,2.546872,3.2295387,4.2568207,4.969026,6.377026,7.578257,8.103385,7.9425645,9.924924,13.098668,15.448617,15.780104,13.696001,11.352616,9.846154,9.69518,10.610872,11.477334,12.809847,12.891898,12.576821,12.097642,11.080206,10.417232,11.244308,13.571283,17.204514,21.753437,23.850668,24.943592,25.98072,27.050669,27.375591,29.472822,31.72431,32.50544,30.739695,25.91508,22.564104,23.922874,25.317745,23.72595,17.765745,19.055592,22.28513,24.694157,25.350567,25.170053,26.673233,29.889643,36.50626,44.786877,49.57867,40.352825,33.079796,25.078156,17.631182,15.990155,16.423386,16.512001,14.372104,12.370052,17.138874,23.45354,21.950361,20.722874,23.112207,27.716925,31.681643,39.223797,44.097645,43.716927,39.158157,37.9799,32.705643,25.242258,18.871796,18.248207,17.289848,15.209026,13.984821,13.689437,12.461949,11.398565,12.931283,14.700309,15.225437,13.912617,16.20677,18.46154,18.46154,16.09518,13.361232,15.547078,18.025026,20.033642,21.431797,22.692104,19.27877,15.130258,11.237744,7.906462,4.7425647,5.5269747,5.1922054,5.080616,5.4580517,5.5007186,5.622154,5.35959,5.0543594,4.8836927,4.857436,5.3431797,5.7140517,5.398975,4.5522056,4.0434875,4.2601027,4.7261543,4.7556925,4.4373336,4.6145644,4.9427695,5.4482055,5.986462,6.2162056,5.5991797,4.8377438,3.9089234,3.3378465,3.186872,3.0424619,2.7241027,2.6978464,2.8389745,3.245949,4.2272825,6.052103,7.7456417,9.370257,11.083488,13.11836,15.593027,17.585232,18.06113,17.772308,19.259079,23.240208,27.936823,32.02626,35.86954,41.50154,45.57785,46.273643,41.849438,33.335796,24.516926,18.691284,13.90277,10.709334,9.002667,8.001641,7.525744,7.8047185,7.9261546,7.276308,5.5630774,5.717334,6.47877,7.9130263,9.7673855,11.45436,11.9860525,11.667693,10.006975,7.499488,5.61559,4.7491283,4.3618464,4.2929235,4.7524104,6.298257,5.353026,5.3136415,6.009436,7.9130263,12.117334,10.906258,11.32636,10.857026,9.383386,9.179898,10.092308,12.488206,14.565744,14.884104,12.36677,15.123693,14.736411,11.608616,8.674462,11.392001,12.612924,7.4404106,3.748103,3.4133337,2.300718,1.847795,2.28759,2.7569232,2.8488207,2.609231,1.9331284,3.3641028,4.71959,5.287385,5.832206,9.202872,10.029949,12.278154,16.324924,18.95713,29.669746,37.700928,43.080208,46.69375,50.264618,69.4679,72.18216,65.35549,56.28062,52.608006,60.314262,69.53683,77.653336,81.95283,79.625854,82.42873,81.13232,65.65744,41.793644,31.209028,23.82113,19.96472,17.365335,15.763694,16.902565,19.078566,20.26995,22.186668,24.037745,22.531284,20.250257,18.83241,17.555695,18.976822,28.934566,36.066463,37.120003,38.71508,40.320004,34.241642,18.835693,9.6,5.2348723,4.2469745,4.9329233,3.05559,1.4605129,0.69907695,0.76800007,1.086359,1.2800001,2.7306669,3.367385,2.7011285,1.8084104,0.6892308,0.7581539,1.1323078,1.5983591,2.6157951,1.1323078,1.4572309,4.7950773,7.9327188,3.2196925,6.7282057,9.015796,7.9097443,5.169231,6.485334,2.9997952,1.4572309,1.1323078,1.3489232,1.4539489,1.148718,1.6475899,2.6289232,3.8531284,5.139693,5.58277,6.9120007,12.488206,23.013746,36.535797,20.929642,8.92718,3.623385,3.31159,1.4900514,0.76800007,0.98133343,1.1782565,1.1126155,1.2406155,1.4966155,1.6508719,1.6869745,1.5688206,1.2471796,1.4276924,1.3489232,1.6640002,2.1956925,1.9265642,1.7033848,1.8215386,2.0676925,2.231795,2.1136413,2.2646155,1.9856411,1.6836925,1.522872,1.4112822,1.4605129,1.1651284,1.014154,1.1979488,1.585231,1.1749744,0.95835906,1.0075898,1.2209232,1.2964103,1.4834872,2.1464617,2.678154,2.6026669,1.595077,1.5524104,2.1891284,2.2383592,1.8018463,2.3696413,3.255795,2.7700515,2.3204105,2.228513,1.719795,1.7066668,1.913436,1.9035898,1.6311796,1.4473847,1.2964103,0.88615394,0.79425645,0.9714873,0.764718,0.6465641,0.7581539,0.84348726,0.94523084,1.4112822,1.7033848,1.0338463,0.5546667,0.56451285,0.48574364,0.2231795,0.19364104,0.23302566,0.21333335,0.049230773,0.052512825,0.03938462,0.02297436,0.0032820515,0.0,0.0,0.0032820515,0.013128206,0.032820515,0.04266667,0.01969231,0.013128206,0.013128206,0.016410258,0.016410258,0.006564103,0.0,0.0032820515,0.009846155,0.0,0.0,0.0,0.009846155,0.01969231,0.0,0.0,0.13784617,0.33805132,0.5677949,0.8172308,0.56123084,0.256,0.098461546,0.101743594,0.08861539,0.08861539,0.09189744,0.06235898,0.013128206,0.0,0.09189744,0.08205129,0.055794876,0.07548718,0.15097436,0.08861539,0.06564103,0.04594872,0.03938462,0.07876924,0.10502565,0.055794876,0.026256412,0.049230773,0.08205129,0.16082053,0.15097436,0.128,0.118153855,0.128,0.13456412,0.21333335,0.23302566,0.15097436,0.03938462,0.101743594,0.0951795,0.11158975,0.15097436,0.13784617,0.0951795,0.049230773,0.032820515,0.07548718,0.21661541,0.16082053,0.07548718,0.036102567,0.04266667,0.01969231,0.072205134,0.049230773,0.01969231,0.009846155,0.0,0.006564103,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016410258,0.07548718,0.21989745,0.512,0.6268718,0.512,0.29210258,0.256,0.32820517,0.39056414,0.42338464,0.4397949,0.49887183,0.5415385,0.6432821,0.761436,0.90912825,1.1224617,0.97805136,0.92553854,0.9878975,1.0962052,1.0896411,0.97805136,0.67938465,0.43651286,0.35446155,0.39056414,0.34789747,0.3249231,0.24943592,0.13456412,0.072205134,0.052512825,0.06564103,0.14441027,0.32164106,0.636718,0.6268718,0.43651286,0.32820517,0.4135385,0.6432821,0.574359,0.6629744,0.7515898,0.761436,0.6892308,0.77456415,0.9156924,0.86646163,0.6695385,0.6629744,0.5973334,0.5316923,0.49230772,0.49887183,0.55794877,0.508718,0.4201026,0.32820517,0.2855385,0.37415388,0.512,0.52512825,0.6432821,0.90256417,1.142154,1.3161026,1.394872,1.3620514,1.204513,0.93866676,0.65641034,0.49887183,0.47589746,0.5546667,0.65641034,0.73517954,0.86974365,1.0601027,1.2898463,1.5425643,1.3850257,1.2964103,1.332513,1.3850257,1.1782565,1.086359,0.9682052,0.94523084,1.0404103,1.1782565,1.1946667,1.2996924,1.3620514,1.3653334,1.394872,1.6114873,1.657436,1.5097437,1.339077,1.5163078,1.5524104,1.5261539,1.4834872,1.4506668,1.4178462,1.3226668,1.332513,1.273436,1.1651284,1.2406155,1.4408206,1.5163078,1.5392822,1.5819489,1.7099489,1.5392822,1.3357949,1.2832822,1.4112822,1.585231,1.6771283,1.4244103,1.4342566,1.7132308,1.657436,1.2898463,1.0305642,1.0108719,1.1290257,1.0436924,1.1290257,1.0108719,0.9878975,1.0765129,1.0108719,1.0338463,1.0043077,0.88943595,0.702359,0.5218462,0.571077,0.7975385,0.8402052,0.7089231,0.7778462,0.9747693,0.8598975,0.69907695,0.6268718,0.6629744,0.58420515,0.55794877,0.6432821,0.7811283,0.82379496,0.85005134,1.014154,1.1815386,1.2832822,1.3292309,1.3751796,1.5163078,1.6508719,1.6640002,1.4375386,1.9003079,2.1202054,2.2514873,2.6387694,3.8038976,3.3378465,2.8521028,2.7798977,3.0818465,3.2361028,2.556718,2.1989746,1.9331284,1.6443079,1.3193847,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.04594872,0.108307704,0.190359,0.23302566,0.26584616,0.33805132,0.508718,0.761436,0.9353847,1.2274873,1.6114873,1.8281027,1.9528207,1.9954873,2.2186668,2.6256413,2.9669745,2.7831798,3.5544617,4.4964104,5.1659493,5.4941545,6.672411,8.402052,9.603283,9.472001,7.4765134,6.0619493,5.865026,6.3245134,6.961231,7.3747697,9.596719,11.257437,12.186257,12.534155,12.763899,13.059283,14.221129,17.250463,21.720617,25.767387,26.98831,28.212515,29.728823,31.56349,33.47036,38.065235,47.005543,53.687798,52.07303,36.68677,28.845951,26.932514,25.577028,22.272001,17.38831,18.343386,20.440617,22.4919,24.113234,25.72472,28.803284,32.65313,43.346054,60.28472,76.21252,67.87611,58.624004,46.483696,33.280003,24.625233,21.822361,17.83795,14.998976,16.216616,25.012514,28.655592,26.60431,25.232412,26.791388,29.397335,33.12903,38.744617,39.67672,35.186874,30.38195,27.766155,23.45354,20.420925,19.334566,18.520617,17.375181,16.521847,14.690463,12.015591,10.029949,10.512411,12.317539,13.410462,13.423591,13.6467705,16.239592,16.850052,15.711181,13.843694,13.056001,16.41354,18.261335,19.213129,19.561028,19.249231,16.915693,12.596514,9.531077,8.388924,7.269744,7.75877,7.066257,6.1374364,5.435077,4.9329233,4.5817437,4.5587697,4.4898467,4.2371287,3.8859491,4.59159,5.024821,4.8804107,4.4996924,4.8804107,5.221744,5.169231,4.7261543,4.2207184,4.276513,4.027077,3.9023592,3.9122055,3.9089234,3.5840003,3.2689233,2.8160002,2.5107694,2.4516926,2.546872,2.5862565,2.8455386,2.917744,2.993231,3.8728209,5.546667,6.9645133,8.664616,10.587898,12.06154,13.036308,14.01436,14.5263605,15.300924,18.267899,23.794874,30.198156,34.648617,36.28636,36.197746,33.64103,31.044926,26.095592,19.360823,14.283488,12.176412,10.59118,9.252103,8.165744,7.6110773,6.987488,6.744616,6.5706673,6.232616,5.549949,5.7468724,7.3583593,9.107693,10.482873,11.720206,12.832822,12.0549755,9.780514,7.0925136,5.7403083,6.439385,6.183385,5.6352825,5.5630774,6.872616,5.2644105,4.9920006,5.5138464,6.9152827,9.924924,11.556104,14.336001,15.570052,14.834873,13.965129,11.536411,13.042872,15.176207,15.186052,10.893129,14.569027,15.258258,13.062565,10.167795,10.8537445,11.155693,8.2215395,5.4383593,4.135385,3.5872824,2.556718,2.3663592,2.2219489,2.0053334,2.2744617,1.6672822,8.300308,9.672206,4.7655387,4.059898,6.6428723,8.15918,11.474052,15.704617,16.196924,24.001642,44.872208,64.72205,74.909546,72.270775,68.30934,59.72021,48.771286,38.85949,34.47467,35.981133,42.870155,53.192207,62.6117,64.416824,70.6757,65.86421,53.38585,38.97436,30.687181,25.685335,26.512413,28.074669,28.038567,26.82749,27.648003,25.53436,25.80677,28.196104,26.843899,23.578259,22.032412,20.690052,21.733746,31.044926,37.103592,34.22195,32.01313,32.416824,29.718977,15.655386,7.460103,4.453744,4.7392826,5.1954875,3.2164104,1.7099489,1.024,1.083077,1.3784616,1.782154,2.1530259,1.8740515,1.3161026,1.847795,2.428718,1.7624617,1.6738462,2.487795,3.0326157,1.5786668,2.2547693,5.533539,8.208411,3.387077,5.920821,9.501539,8.631796,4.673641,5.8453336,4.4242053,3.1081028,2.0808206,1.595077,1.9856411,1.5458462,1.142154,1.4244103,3.045744,6.672411,8.664616,9.3768215,12.576821,20.54236,34.07426,17.545847,7.0367184,4.332308,5.7403083,2.100513,0.7515898,1.0010257,1.2931283,1.142154,1.1454359,1.3095386,1.3883078,1.4178462,1.4276924,1.4211283,1.2635899,1.1520001,1.5360001,2.1858463,2.1825643,1.8510771,2.0611284,2.1202054,1.8707694,1.6738462,2.0644104,1.6836925,1.2438976,1.086359,1.1913847,1.3522053,1.086359,0.8598975,0.9485129,1.4408206,1.211077,1.0535386,1.1224617,1.3587693,1.4867693,1.4966155,2.041436,2.5206156,2.4746668,1.5885129,1.4703591,1.8838975,2.044718,2.038154,2.8225644,4.164923,3.9811285,3.259077,2.4451284,1.4309745,1.4309745,1.9035898,1.8937438,1.2996924,0.86646163,1.0338463,0.8533334,0.90912825,1.1323078,0.7844103,0.446359,0.37415388,0.39712822,0.46276927,0.6498462,0.78769237,0.48246157,0.25271797,0.25271797,0.28225642,0.13128206,0.072205134,0.07548718,0.08861539,0.013128206,0.02297436,0.01969231,0.009846155,0.006564103,0.0,0.0,0.006564103,0.006564103,0.0,0.006564103,0.006564103,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0032820515,0.009846155,0.0,0.0,0.07548718,0.30851284,0.6071795,0.7122052,0.56123084,0.3314872,0.16738462,0.12143591,0.15425642,0.08205129,0.08533334,0.07876924,0.04594872,0.01969231,0.1148718,0.098461546,0.06235898,0.08205129,0.20020515,0.1148718,0.118153855,0.0951795,0.036102567,0.049230773,0.10502565,0.08861539,0.04594872,0.013128206,0.032820515,0.08205129,0.09189744,0.13128206,0.18379489,0.14441027,0.08861539,0.17723078,0.21989745,0.15753847,0.06564103,0.04594872,0.03938462,0.06235898,0.118153855,0.21989745,0.24287182,0.15425642,0.07548718,0.055794876,0.10502565,0.108307704,0.049230773,0.006564103,0.0,0.006564103,0.006564103,0.0032820515,0.029538464,0.06235898,0.026256412,0.026256412,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01969231,0.098461546,0.16738462,0.32820517,0.38728207,0.318359,0.28882053,0.3314872,0.39384618,0.43323082,0.44964105,0.4594872,0.5316923,0.6695385,0.8467693,1.0305642,1.1749744,0.93866676,0.88943595,1.020718,1.1946667,1.1290257,1.148718,0.86646163,0.5546667,0.38728207,0.4201026,0.37743592,0.34133336,0.25928208,0.14769232,0.08533334,0.06235898,0.068923086,0.20348719,0.446359,0.6695385,0.6498462,0.58420515,0.47261542,0.4201026,0.6268718,0.46276927,0.5513847,0.8533334,1.079795,0.69251287,0.6301539,0.764718,0.7778462,0.65312827,0.65969235,0.71548724,0.67938465,0.60061544,0.5152821,0.43323082,0.51856416,0.9911796,0.9419488,0.40697438,0.3708718,0.4397949,0.46276927,0.5973334,0.8467693,1.0601027,1.3095386,1.3686155,1.2603078,1.0502565,0.86317956,0.8041026,0.5940513,0.46276927,0.51856416,0.7581539,0.65969235,0.7384616,0.9616411,1.2668719,1.5688206,1.4966155,1.3489232,1.3128207,1.3784616,1.3259488,1.273436,1.1454359,1.086359,1.148718,1.3062565,1.0994873,1.1716924,1.2931283,1.3653334,1.4080001,1.5655385,1.7558975,1.8051283,1.6607181,1.3817437,1.5130258,1.5163078,1.3915899,1.2307693,1.2242053,1.148718,1.083077,1.0601027,1.079795,1.1093334,1.2438976,1.1848207,1.1913847,1.3587693,1.6147693,1.5458462,1.2635899,1.1913847,1.3817437,1.522872,1.4506668,1.2898463,1.2438976,1.3456411,1.4473847,1.0962052,0.8730257,0.90584624,1.1191796,1.2570257,1.2307693,1.1224617,1.0633847,1.0535386,0.9682052,0.99774367,0.92225647,0.81394875,0.71548724,0.6170257,0.60061544,0.75487185,0.80738467,0.7220513,0.7089231,0.90912825,0.8960001,0.7811283,0.65969235,0.61374366,0.5973334,0.60389745,0.6629744,0.7220513,0.6629744,0.8008206,1.0272821,1.204513,1.2964103,1.3751796,1.5786668,1.5556924,1.5589745,1.6246156,1.5885129,1.591795,1.719795,1.8510771,2.2186668,3.4264617,2.8291285,2.4549747,2.553436,2.9210258,2.9243078,2.1398976,1.657436,1.3751796,1.2242053,1.1585642,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.036102567,0.18707694,0.20348719,0.23958977,0.37415388,0.6071795,0.7515898,0.81066674,1.079795,1.5327181,1.8281027,1.7624617,1.7099489,1.7624617,1.8576412,1.7887181,1.4966155,1.8970258,2.4516926,2.9505644,3.501949,3.9220517,4.46359,4.6966157,4.568616,4.4012313,3.876103,4.2436924,4.7294364,5.07077,5.5171285,7.9852314,10.469745,12.347078,13.761642,15.616001,18.5239,21.464617,23.108925,23.80472,25.590157,26.735592,28.842669,31.10072,33.736206,38.048824,45.505646,64.52513,80.600624,81.14873,55.52903,39.25662,31.944208,28.17313,25.133951,22.642874,22.249027,21.274258,21.369438,22.882463,24.868105,28.327387,31.537233,40.067284,54.176826,68.81149,63.10729,57.248825,48.92226,38.73149,30.198156,25.816618,20.260103,18.884924,23.223797,30.962873,31.478157,30.848001,30.431181,30.611694,30.782362,33.736206,35.807182,33.614773,28.038567,24.234669,22.921848,21.523693,21.845335,22.787283,20.329027,18.921026,17.641027,14.723283,10.8767185,9.291488,10.725744,13.590976,14.946463,14.598565,15.110565,16.83036,15.878566,14.339283,13.745232,15.067899,19.272207,20.214155,19.495386,17.864206,15.209026,13.90277,10.952206,9.248821,9.258667,9.02236,8.950154,7.968821,6.521436,5.0904617,4.1813335,3.6693337,3.6069746,3.5971284,3.4789746,3.3247182,3.8564105,4.309334,4.417641,4.417641,5.0642056,4.965744,4.667077,4.1878977,3.761231,3.817026,3.3936412,2.9538465,2.5796926,2.349949,2.3269746,2.3335385,2.359795,2.356513,2.3630772,2.5173335,2.7044106,2.9768207,3.1409233,3.4100516,4.414359,5.910975,7.381334,9.097847,10.8996935,12.20595,12.242052,12.800001,13.781334,15.570052,19.029335,23.200823,27.3559,29.154465,28.009027,25.088001,20.598156,17.956104,15.520822,12.928001,11.109744,10.354873,9.826463,9.088,8.178872,7.6242056,7.128616,6.5017443,6.232616,6.436103,6.8397956,7.8014364,10.220308,11.933539,12.481642,13.115078,13.640206,12.977232,10.962052,8.5891285,8.004924,8.79918,8.083693,7.1154876,7.0334363,8.848411,8.900924,10.912822,14.54277,20.936207,32.705643,46.185028,45.026466,34.208824,21.047796,15.199181,11.815386,12.268309,14.624822,15.924514,12.1928215,13.587693,13.387488,11.910565,10.006975,9.048616,7.90318,7.0137444,6.2851286,5.654975,5.110154,4.57518,3.7874875,2.5173335,1.3784616,1.8215386,3.6660516,10.292514,10.180923,4.023795,4.7294364,5.904411,7.381334,11.736616,16.544823,14.358975,16.577642,39.168003,67.1278,86.52473,84.496414,61.00021,44.307697,33.828106,28.258463,25.593437,22.544413,25.728003,33.539284,42.663387,48.08534,53.566364,49.618053,43.62831,38.948105,34.89477,33.05026,37.72062,45.16103,51.744823,53.95693,50.113644,40.12308,33.48021,32.48903,32.262566,27.608618,25.429335,23.768618,24.175592,31.734156,36.47344,30.802053,24.6679,21.943796,20.447182,10.811078,4.896821,3.2328207,4.1813335,3.9056413,2.6223593,1.7558975,1.394872,1.4769232,1.8018463,1.8773335,1.7296412,1.5130258,1.7591796,3.4067695,5.989744,8.001641,6.889026,4.378257,6.4754877,2.609231,4.1091285,7.6110773,9.248821,4.663795,3.8662567,5.7665644,5.3398976,3.1606157,5.3792825,6.166975,4.601436,2.6945643,1.8215386,2.7241027,2.3269746,1.5097437,1.1224617,2.0644104,5.2742567,7.529026,7.5487185,8.103385,11.040821,17.283283,8.073847,5.83877,8.01477,9.43918,2.3860514,1.0436924,1.0962052,1.1913847,0.9714873,1.0699488,0.955077,0.97805136,1.0929232,1.2438976,1.3620514,1.0666667,1.0994873,1.4473847,1.9167181,2.1333334,1.8149745,1.975795,1.910154,1.591795,1.6410258,2.1924105,1.6836925,1.1651284,1.0305642,1.0305642,1.1618463,0.98133343,0.764718,0.7581539,1.1585642,1.1552821,1.020718,1.024,1.2176411,1.4375386,1.3981539,1.6902566,1.9528207,1.9593848,1.6082052,1.3554872,1.394872,1.4900514,1.7066668,2.4155898,3.820308,4.013949,3.383795,2.3236926,1.2406155,1.4080001,1.910154,1.8674873,1.211077,0.69579494,0.8730257,0.8467693,0.93866676,1.0732309,0.79097444,0.5349744,0.34133336,0.2297436,0.17723078,0.13128206,0.12471796,0.08861539,0.055794876,0.052512825,0.098461546,0.06235898,0.032820515,0.013128206,0.006564103,0.0,0.013128206,0.006564103,0.006564103,0.013128206,0.0,0.0,0.006564103,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.009846155,0.14441027,0.34133336,0.3708718,0.7581539,0.48574364,0.2100513,0.17066668,0.20348719,0.072205134,0.06235898,0.07876924,0.06564103,0.01969231,0.098461546,0.09189744,0.068923086,0.0951795,0.24943592,0.15425642,0.19692309,0.18707694,0.101743594,0.07876924,0.10502565,0.15753847,0.128,0.03938462,0.032820515,0.01969231,0.036102567,0.10502565,0.18379489,0.18051283,0.13456412,0.21333335,0.24287182,0.17723078,0.0951795,0.04266667,0.016410258,0.016410258,0.055794876,0.17066668,0.23630771,0.2100513,0.13128206,0.052512825,0.01969231,0.049230773,0.026256412,0.006564103,0.006564103,0.029538464,0.0951795,0.055794876,0.04266667,0.072205134,0.026256412,0.06564103,0.029538464,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.036102567,0.006564103,0.101743594,0.20020515,0.24943592,0.26584616,0.30194873,0.37743592,0.4397949,0.46933338,0.4594872,0.5316923,0.65969235,0.8533334,1.0699488,1.2176411,0.9353847,0.9682052,1.0896411,1.1454359,1.0305642,1.0896411,0.9124103,0.67938465,0.512,0.48902568,0.43323082,0.36102566,0.25928208,0.14769232,0.09189744,0.06235898,0.06564103,0.18707694,0.38728207,0.5284103,0.571077,0.58420515,0.4955898,0.41025645,0.62030774,0.4660513,0.47589746,0.7778462,1.0929232,0.75487185,0.5546667,0.6662565,0.7450257,0.6859488,0.60389745,0.7450257,0.77128214,0.67938465,0.50543594,0.33476925,0.49887183,1.3062565,1.3128207,0.5415385,0.48902568,0.446359,0.47589746,0.57764107,0.7384616,0.9353847,1.1782565,1.2996924,1.214359,0.96492314,0.75487185,0.7811283,0.5973334,0.446359,0.47589746,0.77456415,0.6826667,0.69907695,0.8172308,1.0305642,1.2996924,1.3751796,1.273436,1.2012309,1.2373334,1.3259488,1.3423591,1.2307693,1.2077949,1.3062565,1.3850257,1.1224617,1.1257436,1.2668719,1.3751796,1.2668719,1.4309745,1.7460514,1.8740515,1.7066668,1.3686155,1.6344616,1.5491283,1.2964103,1.0699488,1.0601027,1.0371283,0.9747693,0.9747693,1.0371283,1.0732309,1.0994873,1.020718,1.0305642,1.1913847,1.4441026,1.522872,1.3489232,1.2570257,1.3193847,1.339077,1.1946667,1.1684103,1.2406155,1.3095386,1.1848207,0.9321026,0.8205129,0.8795898,1.079795,1.3489232,1.2832822,1.2176411,1.1618463,1.1323078,1.1388719,1.0732309,0.9353847,0.8336411,0.77456415,0.67610264,0.5973334,0.6498462,0.6826667,0.65312827,0.6235898,0.74830776,0.8205129,0.8205129,0.7581539,0.6859488,0.69251287,0.6498462,0.6498462,0.67938465,0.62030774,0.78769237,0.99774367,1.1651284,1.2964103,1.4802053,1.5753847,1.5261539,1.4933335,1.4998976,1.4539489,1.3883078,1.5195899,1.5622566,1.7132308,2.6289232,2.3991797,2.2219489,2.3433847,2.612513,2.484513,1.6869745,1.2209232,1.0108719,0.9714873,1.0305642,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.016410258,0.01969231,0.0,0.15425642,0.18379489,0.24615386,0.39712822,0.5874872,0.5546667,0.77456415,1.148718,1.5392822,1.782154,1.5721027,1.3029745,1.0962052,0.9944616,0.9616411,0.9878975,1.2209232,1.4080001,1.4998976,1.6508719,1.591795,1.7723079,1.9856411,2.4681027,3.8728209,3.446154,3.620103,3.9253337,4.2601027,4.9132314,6.7282057,9.284924,12.117334,15.094155,18.46154,24.67118,29.472822,28.537437,23.670156,22.826668,25.055182,28.399591,31.159798,34.162876,40.759796,49.591797,74.545235,96.98462,100.91652,73.00267,49.772312,37.66482,32.774567,32.022976,33.174976,30.71672,25.531078,22.465643,22.537848,22.95795,25.294771,27.040823,29.095387,31.583181,33.86421,31.136824,31.622566,31.783386,30.496822,29.075695,26.706053,23.299284,24.556309,29.912617,32.544823,31.583181,32.210052,31.9639,30.395079,29.056002,32.94195,33.83467,31.632412,27.546259,24.09354,23.85395,24.943592,25.944618,25.544207,22.52472,20.716309,17.398155,13.774771,11.241027,11.378873,12.35036,15.809642,18.139898,18.244925,17.54913,17.043694,15.501129,14.644514,15.37313,17.765745,21.782976,21.664822,19.472412,16.114874,11.34277,10.187488,9.616411,9.314463,9.035488,8.576,8.2904625,7.5618467,6.183385,4.5390773,3.6102567,3.2722054,3.1573336,3.045744,3.006359,3.383795,3.692308,4.1878977,4.4373336,4.4242053,4.525949,3.9187696,3.9614363,3.9876926,3.8728209,4.0467696,3.9614363,3.757949,3.4100516,3.0916924,3.1671798,2.9538465,2.8849232,2.8849232,3.0030773,3.4133337,3.6627696,3.8334363,4.3290257,5.3103595,6.7117953,8.067283,9.55077,10.994873,12.324103,13.545027,13.61395,14.477129,15.8654375,17.700104,20.086155,21.047796,21.014977,19.771078,17.900309,16.774565,15.163078,14.204719,13.984821,13.945437,12.911591,12.274873,11.785847,11.270565,10.57477,9.563898,9.042052,8.54318,8.595693,9.147078,9.573745,11.569232,14.106257,15.507693,15.648822,15.947489,15.113848,14.55918,13.049437,11.155693,11.23118,11.575796,10.916103,10.400822,11.076924,13.88636,17.122463,23.11877,32.43323,47.570053,72.99611,96.3315,84.30606,53.48103,22.166977,10.407386,8.36595,7.9852314,10.020103,12.934566,12.908309,11.490462,10.154668,9.193027,8.641642,8.303591,6.987488,6.042257,6.3310776,7.138462,6.1768208,6.567385,5.4843082,3.3772311,1.4441026,1.6344616,5.9569235,6.889026,5.3924108,3.9975388,6.7807183,6.685539,6.9809237,10.834052,16.118155,15.415796,13.774771,24.769644,47.829338,72.58257,78.89067,49.572105,31.583181,23.59467,21.753437,19.702156,16.676104,18.530462,23.174566,28.842669,34.090668,37.858463,43.559387,46.23754,45.47939,45.397335,47.30749,52.4439,64.1477,79.163086,87.617645,78.05047,58.581337,42.646976,36.135387,37.376003,32.295387,29.479387,27.188515,26.049643,29.059284,32.4759,27.890875,21.651693,17.191385,15.018668,9.32759,4.519385,2.428718,2.556718,2.0742567,1.7394873,1.5622566,1.5458462,1.6771283,1.9593848,1.3357949,1.5425643,1.7887181,2.2514873,4.059898,8.218257,15.632411,13.74195,6.294975,13.351386,4.8311796,5.293949,8.185436,9.540924,7.962257,2.4549747,1.3554872,1.467077,2.0873847,4.9788723,6.6560006,4.7360005,2.553436,1.975795,3.4231799,3.0030773,2.4155898,1.9495386,1.8412309,2.2908719,2.930872,3.3214362,3.7152824,3.9614363,3.508513,1.5524104,5.7632823,10.299078,10.31877,2.0118976,1.4834872,1.3095386,1.0371283,0.8008206,1.3161026,0.8763078,0.8533334,0.9714873,1.0469744,1.0043077,0.88287187,1.0010257,1.1749744,1.3357949,1.5097437,1.4145643,1.5195899,1.6016412,1.7558975,2.422154,3.1245131,2.5042052,1.7755898,1.3587693,0.8730257,0.88615394,0.8533334,0.7417436,0.6695385,0.9124103,1.083077,0.892718,0.7450257,0.8172308,1.0666667,1.0601027,1.1355898,1.2242053,1.3357949,1.5425643,1.2209232,1.1454359,1.1060513,1.0601027,1.1093334,2.0808206,2.5042052,2.3958976,1.8412309,1.0010257,1.3587693,1.7624617,1.7657437,1.3751796,1.0732309,0.90256417,0.8402052,0.78769237,0.7122052,0.636718,0.65312827,0.44964105,0.23302566,0.0951795,0.026256412,0.026256412,0.036102567,0.029538464,0.013128206,0.013128206,0.013128206,0.006564103,0.0032820515,0.0,0.0,0.08861539,0.052512825,0.013128206,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.02297436,0.06564103,0.9616411,0.6826667,0.3117949,0.24287182,0.20676924,0.06235898,0.03938462,0.055794876,0.052512825,0.0,0.06235898,0.07876924,0.08205129,0.12471796,0.26584616,0.17723078,0.24615386,0.26584616,0.19364104,0.14441027,0.11158975,0.2100513,0.20348719,0.08533334,0.06235898,0.02297436,0.03938462,0.068923086,0.098461546,0.13784617,0.16410258,0.21989745,0.23630771,0.19692309,0.13456412,0.068923086,0.02297436,0.0032820515,0.006564103,0.016410258,0.072205134,0.15753847,0.15425642,0.06235898,0.0032820515,0.0,0.0,0.0,0.016410258,0.07548718,0.19364104,0.11158975,0.03938462,0.032820515,0.013128206,0.08533334,0.04266667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.032820515,0.07876924,0.13784617,0.20020515,0.24943592,0.34133336,0.42338464,0.46933338,0.47917953,0.53825647,0.62030774,0.764718,0.95835906,1.1651284,0.9616411,1.0896411,1.142154,1.024,0.9419488,0.9419488,0.8533334,0.7581539,0.67610264,0.57764107,0.46276927,0.3511795,0.24287182,0.14769232,0.0951795,0.059076928,0.04594872,0.08861539,0.18379489,0.32164106,0.446359,0.46933338,0.41682056,0.40369233,0.64000005,0.50543594,0.40697438,0.512,0.7384616,0.761436,0.55794877,0.6629744,0.7778462,0.7515898,0.5677949,0.71548724,0.76800007,0.6826667,0.4955898,0.35774362,0.46933338,1.1388719,1.2471796,0.7811283,0.8336411,0.64000005,0.574359,0.56123084,0.6170257,0.83035904,1.0272821,1.2307693,1.2340513,1.020718,0.7318975,0.63343596,0.5349744,0.4660513,0.48574364,0.67610264,0.7450257,0.761436,0.72861546,0.7318975,0.92553854,1.086359,1.0929232,1.0469744,1.0436924,1.1585642,1.2340513,1.148718,1.2012309,1.3686155,1.332513,1.2274873,1.1848207,1.2996924,1.4244103,1.1585642,1.3686155,1.6213335,1.6311796,1.4802053,1.6016412,1.7985642,1.4933335,1.1323078,0.9419488,0.955077,0.97805136,0.99774367,0.9944616,0.9878975,1.0535386,1.0568206,1.0929232,1.1191796,1.1585642,1.2865642,1.4769232,1.4998976,1.404718,1.2570257,1.1290257,1.142154,1.1749744,1.3981539,1.5885129,1.0994873,0.9517949,0.9517949,0.99774367,1.0732309,1.2340513,1.2438976,1.2406155,1.1979488,1.1881026,1.3686155,1.2274873,1.0633847,0.9485129,0.86646163,0.702359,0.6268718,0.65641034,0.6629744,0.6268718,0.6498462,0.6268718,0.65641034,0.72861546,0.7975385,0.7844103,0.7975385,0.6662565,0.5940513,0.6170257,0.63343596,0.7384616,0.88943595,1.079795,1.2931283,1.4834872,1.3193847,1.3259488,1.3686155,1.2996924,0.9616411,1.3489232,1.5622566,1.4867693,1.3686155,1.8215386,2.03159,1.9003079,1.9035898,2.0808206,2.0545642,1.3423591,1.0338463,0.93866676,0.92553854,0.8992821,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.036102567,0.08533334,0.098461546,0.0,0.08533334,0.14441027,0.23630771,0.35774362,0.44307697,0.5152821,0.7253334,1.0010257,1.2077949,1.1585642,0.84348726,0.52512825,0.36758977,0.42338464,0.65641034,0.69251287,0.702359,0.7318975,0.761436,0.6859488,0.39384618,0.37415388,0.9353847,2.1267693,3.7382567,3.7021542,3.3444104,3.1540515,3.373949,3.9975388,4.71959,8.247795,12.655591,16.971489,21.195488,28.665438,32.098465,30.102976,24.914053,22.400002,25.537643,28.711388,31.304207,34.37621,40.64821,46.87426,61.587696,76.537445,82.29088,68.25354,50.248207,38.862774,35.27877,38.63303,46.004517,42.98831,32.71549,25.261951,23.213951,21.651693,23.27631,23.893335,23.758772,23.095797,22.09477,22.534565,23.752207,23.863796,23.253336,24.582565,27.976208,28.55713,29.856823,31.248413,27.953234,26.427078,26.496002,26.338463,25.711592,25.954464,31.376413,35.045746,35.167183,31.917952,27.451078,27.720207,28.153439,27.37231,24.782772,20.585028,17.690258,14.506668,12.649027,12.563693,13.50236,12.455385,13.289026,16.000002,19.016207,19.209848,16.78113,14.506668,13.709129,14.785643,17.227488,18.71754,18.162872,16.485744,13.820719,9.537642,9.3768215,9.639385,10.043077,10.161232,9.429334,8.635077,7.6143594,6.0685134,4.3290257,3.3411283,3.757949,4.1091285,3.9417439,3.6529233,4.4701543,4.201026,3.9876926,4.1714873,4.46359,3.95159,3.95159,4.59159,5.2020516,5.4613338,5.402257,5.2676926,5.3431797,5.3924108,5.474462,5.9503593,5.32677,4.716308,4.6900516,5.4547696,6.820103,6.8332314,7.282872,8.103385,9.104411,9.993847,10.384411,10.738873,11.47077,12.603078,13.764924,14.995693,16.485744,17.719797,18.67159,19.80718,19.830154,19.524925,19.682463,19.826874,18.202257,15.701335,14.76595,15.320617,16.718771,17.746052,19.15077,19.840002,19.144207,17.168411,14.8020525,13.5548725,13.308719,13.499078,13.699283,13.627078,14.418053,15.14995,15.691488,16.009848,16.144411,16.997746,15.665232,13.499078,11.851488,12.084514,14.795488,16.817232,18.464823,20.28308,23.056412,27.365746,35.67262,47.717747,63.20575,81.8478,88.40534,67.62339,37.116722,12.274873,6.2555904,6.9382567,5.2709746,4.965744,7.026872,9.734565,10.358154,10.633847,10.650257,10.683078,11.185231,10.709334,8.759795,6.7314878,5.579488,5.799385,4.6769233,3.3608208,2.5862565,2.4648206,2.5009232,4.0402055,3.820308,4.9920006,7.634052,8.759795,7.7456417,8.802463,11.047385,14.930053,22.216208,22.058668,19.866259,25.875694,41.767387,60.70154,40.484104,24.654772,16.951796,15.369847,12.1468725,10.742155,13.587693,18.49436,21.494156,16.83036,17.394873,28.95754,40.556313,47.924515,53.526978,62.352413,65.6476,76.202675,91.58565,94.162056,85.04452,66.25806,48.672825,38.754463,38.55754,36.069748,33.604927,31.524105,29.791182,27.986053,27.789131,25.140514,20.923079,16.886156,15.638975,12.294565,6.3507695,2.5042052,1.8182565,1.7099489,1.3062565,1.0305642,1.1060513,1.4112822,1.4966155,0.90912825,1.0469744,1.211077,1.1552821,1.0699488,3.2656412,13.236514,12.71795,6.1505647,20.673643,8.687591,2.9833848,2.8225644,7.0465646,14.053744,6.2030773,5.028103,5.0838976,3.7809234,1.3883078,3.3903592,2.993231,2.0545642,2.0808206,4.240411,3.4002054,2.868513,2.9046156,3.4133337,3.95159,3.4888208,5.3694363,6.2588725,6.1078978,8.149334,2.2646155,1.9659488,3.4198978,4.0369234,2.487795,1.9987694,1.7296412,1.394872,1.3029745,2.3663592,1.5360001,1.4375386,1.4605129,1.2603078,0.74830776,0.67282057,0.5907693,0.5907693,0.7187693,0.9616411,1.0108719,1.1684103,1.6213335,2.4713848,3.754667,4.670359,4.0369234,2.8914874,1.7887181,0.82379496,0.702359,0.7450257,0.71548724,0.67938465,1.020718,1.1946667,0.9156924,0.6826667,0.67282057,0.74830776,0.9682052,0.95835906,0.9714873,1.1257436,1.4178462,1.2373334,1.3554872,1.5064616,1.3653334,0.5349744,0.42338464,0.67282057,1.0502565,1.2570257,0.9156924,0.892718,1.0404103,1.1191796,1.1355898,1.3423591,0.7811283,0.71548724,0.7515898,0.761436,0.86974365,0.5021539,0.32820517,0.21989745,0.11158975,0.016410258,0.016410258,0.052512825,0.04594872,0.0,0.0,0.0,0.009846155,0.009846155,0.0,0.0,0.39056414,0.23302566,0.04266667,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.6859488,0.9911796,0.761436,0.256,0.18379489,0.049230773,0.006564103,0.006564103,0.013128206,0.0,0.02297436,0.059076928,0.108307704,0.14441027,0.108307704,0.108307704,0.190359,0.23958977,0.20348719,0.108307704,0.04594872,0.12143591,0.17066668,0.13456412,0.06235898,0.02297436,0.032820515,0.059076928,0.07548718,0.07548718,0.06564103,0.08861539,0.0951795,0.098461546,0.18379489,0.14769232,0.06564103,0.016410258,0.016410258,0.016410258,0.0032820515,0.026256412,0.08205129,0.11158975,0.016410258,0.0032820515,0.0,0.0,0.016410258,0.07548718,0.026256412,0.006564103,0.006564103,0.02297436,0.06235898,0.036102567,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.036102567,0.01969231,0.0,0.01969231,0.09189744,0.17723078,0.28225642,0.35446155,0.39384618,0.44307697,0.5415385,0.62030774,0.7187693,0.82379496,0.88615394,0.8467693,0.8763078,0.892718,0.90584624,0.9911796,1.1257436,0.93866676,0.7581539,0.67282057,0.56451285,0.380718,0.28882053,0.23630771,0.18051283,0.108307704,0.068923086,0.052512825,0.08205129,0.16082053,0.25928208,0.39384618,0.49887183,0.50543594,0.46933338,0.58092314,0.48246157,0.35774362,0.44307697,0.7220513,0.9321026,0.60061544,0.56451285,0.65641034,0.7253334,0.64000005,0.78769237,0.8041026,0.7089231,0.5513847,0.44307697,0.4660513,0.79425645,1.1651284,1.4178462,1.4802053,1.0043077,0.7187693,0.5677949,0.5481026,0.7318975,0.9878975,1.079795,1.0371283,0.9156924,0.79425645,0.6826667,0.5907693,0.54482055,0.54482055,0.58092314,0.51856416,0.7220513,0.79097444,0.69251287,0.7778462,1.0469744,1.0502565,0.9288206,0.8172308,0.8533334,0.93866676,0.9878975,1.0666667,1.1388719,1.0535386,1.1126155,1.148718,1.2865642,1.4769232,1.463795,1.3784616,1.2668719,1.3259488,1.5524104,1.723077,1.529436,1.1881026,1.0338463,1.1257436,1.2373334,1.0666667,0.93866676,0.892718,0.90584624,0.9321026,1.0535386,1.0732309,1.086359,1.142154,1.2504616,1.4112822,1.3292309,1.1782565,1.079795,1.1290257,1.4966155,1.394872,1.2242053,1.1585642,1.1585642,1.1093334,1.1979488,1.2603078,1.1848207,0.9156924,1.1224617,1.3587693,1.2898463,1.0502565,1.2209232,1.2570257,1.0568206,0.92225647,0.8960001,0.761436,0.67610264,0.7187693,0.7450257,0.74830776,0.86974365,0.80738467,0.7844103,0.8041026,0.7975385,0.6268718,0.6859488,0.6662565,0.5874872,0.512,0.5481026,0.63343596,0.7581539,0.98133343,1.2406155,1.3128207,1.2274873,1.1881026,1.2242053,1.2176411,0.8992821,1.2800001,1.585231,1.7165129,1.723077,1.785436,1.5163078,1.3029745,1.3817437,1.6278975,1.5425643,1.211077,1.0929232,1.014154,0.8992821,0.7778462,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.098461546,0.2231795,0.19692309,0.13456412,0.14769232,0.18707694,0.256,0.41682056,0.5316923,0.6268718,0.6235898,0.58420515,0.7187693,0.6662565,0.5481026,0.4660513,0.44964105,0.43651286,0.46276927,0.380718,0.40697438,0.5218462,0.47917953,0.3708718,0.39384618,1.1848207,2.605949,3.7382567,3.6036925,3.5511796,3.3641028,3.0162053,2.6912823,3.8498464,8.129642,13.499078,18.65518,23.026873,30.79877,33.713234,32.768,29.449848,25.744411,25.668924,27.526566,30.608412,34.12021,37.169235,45.272617,62.260517,79.277954,86.57395,73.51467,49.631184,37.63857,33.775593,35.94831,43.72349,36.978874,28.678566,23.850668,23.292719,23.555285,23.880207,22.130873,21.12,21.697643,22.71836,19.787489,18.691284,19.538054,22.025848,25.4359,27.093336,26.098873,24.425028,23.158155,22.498463,24.585848,25.61313,26.69949,28.02872,28.85908,30.63795,30.995695,30.083284,27.654566,23.079386,24.326567,26.548515,26.617437,24.395489,22.744617,19.508514,15.8884115,14.319591,15.061335,16.177233,16.288822,17.371899,17.913437,17.227488,15.451899,14.624822,12.888617,12.57354,13.853539,14.762668,16.239592,16.190361,13.653335,9.724719,7.5585647,7.604513,7.4863596,7.9524107,8.5202055,7.463385,5.664821,4.7491283,4.1189747,4.007385,5.477744,5.865026,5.664821,5.6418467,5.832206,5.5565133,6.314667,7.4765134,8.054154,7.9491286,7.9425645,7.7292314,7.2303596,6.7085133,6.4295387,6.672411,6.75118,7.138462,7.7390776,8.228104,8.050873,7.3780518,8.421744,10.400822,12.268309,12.727796,12.087796,10.154668,8.907488,8.815591,8.848411,8.057437,8.523488,9.803488,11.513436,13.348104,15.576616,17.929848,19.705437,20.683489,21.123283,21.412104,20.903387,20.158361,19.177027,17.385027,16.768002,14.441027,12.891898,13.197129,15.025232,20.722874,21.19877,19.974566,19.652925,21.904411,22.583797,20.926361,18.33354,15.849027,14.162052,14.5952835,15.665232,16.65313,17.184822,17.243898,17.168411,17.667284,18.034874,18.097233,18.212105,23.049849,27.319798,28.074669,25.974155,25.27836,28.071386,33.762463,40.004925,44.419285,44.58339,38.16041,28.832823,19.062155,11.749744,10.223591,8.864821,7.197539,5.4383593,4.1485133,4.2305646,4.637539,5.428513,6.678975,8.2904625,10.000411,12.160001,11.910565,11.030975,10.134975,8.65477,7.4830775,5.2020516,3.564308,3.2164104,3.7120004,4.4767184,6.8693337,9.321027,11.237744,12.993642,13.456411,13.495796,12.251899,10.397539,10.157949,16.032822,17.168411,17.398155,21.284103,34.103798,26.417233,17.972515,13.128206,12.389745,12.438975,13.272616,14.358975,19.459284,26.36472,26.925951,22.370462,27.690668,38.32123,49.03385,53.943798,66.49764,71.06298,80.23959,94.1358,100.374985,97.01744,80.97478,62.427902,48.695797,44.23549,40.953438,36.8279,33.847797,32.617027,32.354465,32.617027,28.442259,23.77518,20.522669,18.546873,15.113848,8.310155,3.9286156,3.1606157,2.5993848,1.913436,1.4211283,1.4080001,1.6410258,1.3850257,3.767795,2.281026,1.2996924,1.972513,2.228513,2.4320002,10.482873,10.850462,5.3005133,12.911591,10.230155,4.8016415,2.7634873,4.7392826,5.83877,5.986462,6.4295387,7.1089234,7.315693,5.684513,5.5204105,4.903385,3.3411283,2.2711797,5.0477953,4.2436924,3.3345644,3.5577438,4.5587697,4.4045134,2.4451284,2.9768207,4.273231,5.98318,9.124104,4.6080003,4.768821,4.565334,2.556718,0.8992821,1.8871796,1.7657437,1.4736412,1.4900514,1.8281027,1.339077,1.4309745,1.4539489,1.2176411,0.9682052,0.8566154,0.9517949,1.0010257,0.88943595,0.6432821,0.8008206,0.9485129,1.2800001,1.7526156,2.1169233,2.3105643,2.0841026,1.6114873,1.0338463,0.46933338,0.4660513,0.508718,0.56123084,0.67610264,0.99774367,1.2176411,1.0535386,0.764718,0.5546667,0.5874872,0.5940513,0.5973334,0.81066674,1.1027694,1.017436,0.92225647,1.0043077,1.2242053,1.2865642,0.6301539,0.2986667,0.4004103,0.6432821,0.74830776,0.46276927,0.4594872,0.636718,0.80738467,0.93866676,1.1355898,0.8960001,0.6826667,0.571077,0.5513847,0.5152821,0.26584616,0.15097436,0.0951795,0.055794876,0.016410258,0.016410258,0.13128206,0.16082053,0.068923086,0.0,0.01969231,0.068923086,0.06564103,0.009846155,0.0,0.44964105,0.34133336,0.118153855,0.0032820515,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.19692309,0.67282057,0.76800007,0.41025645,0.12143591,0.06564103,0.01969231,0.0,0.0032820515,0.0,0.0032820515,0.013128206,0.02297436,0.029538464,0.02297436,0.02297436,0.04594872,0.07548718,0.08205129,0.032820515,0.02297436,0.101743594,0.17066668,0.15753847,0.036102567,0.01969231,0.026256412,0.04594872,0.08205129,0.16082053,0.08205129,0.052512825,0.052512825,0.06235898,0.049230773,0.052512825,0.029538464,0.016410258,0.013128206,0.0032820515,0.0,0.006564103,0.016410258,0.02297436,0.0032820515,0.01969231,0.016410258,0.013128206,0.016410258,0.026256412,0.006564103,0.009846155,0.013128206,0.032820515,0.098461546,0.032820515,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.0032820515,0.0,0.0032820515,0.01969231,0.036102567,0.15753847,0.2855385,0.380718,0.47917953,0.53825647,0.5415385,0.56451285,0.6498462,0.8008206,0.85005134,0.9288206,1.017436,1.142154,1.3817437,1.5360001,1.3259488,1.0535386,0.8467693,0.6498462,0.45620516,0.3052308,0.19692309,0.13128206,0.108307704,0.059076928,0.055794876,0.07548718,0.12471796,0.2231795,0.41682056,0.84348726,0.88615394,0.5513847,0.50543594,0.32164106,0.20348719,0.3117949,0.6268718,0.9321026,0.65969235,0.5284103,0.512,0.54482055,0.51856416,0.69579494,0.6629744,0.6071795,0.571077,0.44307697,0.4955898,0.508718,0.77128214,1.211077,1.3686155,1.2570257,1.5753847,1.3915899,0.7384616,0.6104616,0.78769237,0.8533334,0.8730257,0.86317956,0.7811283,0.72861546,0.7122052,0.65312827,0.574359,0.5907693,0.7056411,0.73517954,0.7778462,0.83035904,0.7778462,0.99774367,1.0404103,0.9682052,0.88943595,0.96492314,1.0601027,1.0371283,1.0108719,1.0010257,0.955077,1.0371283,1.1257436,1.2668719,1.4211283,1.4769232,1.3915899,1.4605129,1.463795,1.4276924,1.6278975,1.401436,1.1618463,1.0043077,0.9616411,0.9911796,0.95835906,0.93866676,0.90584624,0.9124103,1.1027694,1.0666667,1.0436924,1.0502565,1.1060513,1.214359,1.1979488,1.0896411,1.0666667,1.1355898,1.1060513,1.1093334,1.086359,1.1126155,1.1585642,1.0994873,0.9616411,0.9616411,0.9878975,0.9682052,0.8533334,0.96492314,1.1979488,1.1684103,0.93866676,1.014154,1.1093334,1.024,1.0010257,1.0404103,0.8960001,0.71548724,0.75487185,0.81394875,0.827077,0.88287187,0.69251287,0.6465641,0.6826667,0.7089231,0.57764107,0.49230772,0.46933338,0.48902568,0.5284103,0.574359,0.6892308,0.8402052,0.98133343,1.1060513,1.2274873,1.014154,0.9353847,1.0929232,1.4506668,1.8149745,1.6082052,1.6935385,1.6180514,1.4506668,1.785436,1.5261539,1.3817437,1.2668719,1.2274873,1.4441026,1.142154,0.96492314,0.8566154,0.7811283,0.7187693,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.059076928,0.16410258,0.21661541,0.13456412,0.08533334,0.08861539,0.15753847,0.3117949,0.45620516,0.5284103,0.48246157,0.39384618,0.43651286,0.508718,0.58420515,0.48246157,0.27897438,0.30851284,0.508718,0.61374366,0.72861546,0.84348726,0.83035904,0.8205129,0.77456415,1.2406155,2.0873847,2.5304618,1.8149745,1.7165129,1.8281027,1.9823592,2.2547693,3.5478978,7.571693,13.407181,18.980104,21.057642,25.091284,28.740925,30.5559,30.2999,28.970669,29.088823,30.608412,32.41354,34.225235,36.60144,48.518566,67.46913,84.1518,87.96883,67.039185,45.824005,34.773335,29.1479,27.730053,32.84349,27.88431,23.473232,21.979898,22.78072,22.291695,23.23036,22.554258,21.59918,21.136412,21.379284,18.976822,19.305027,21.431797,23.834259,24.405334,23.64718,25.721437,24.598976,20.598156,20.36513,22.065233,23.2599,24.30359,25.419489,26.702772,25.337439,24.786053,23.988514,23.14831,23.745644,27.542976,29.010054,27.296824,23.945848,22.882463,21.369438,19.15077,17.634462,17.362053,18.018463,18.346668,19.265642,18.287592,15.688207,14.49354,15.048206,13.781334,13.10195,13.5089245,13.587693,14.162052,12.524308,9.974154,7.752206,7.0465646,6.038975,5.9602056,6.813539,7.6734366,6.698667,5.3431797,5.1626673,5.353026,5.674667,6.442667,6.3901544,6.692103,7.213949,7.830975,8.448001,10.194052,11.398565,11.690667,11.142565,10.295795,9.120821,7.9458466,7.2237954,7.1647186,7.7390776,7.5585647,8.52677,9.6065645,10.381129,11.067078,12.901745,15.346873,16.456207,15.314053,12.045129,9.9282055,7.6996927,6.5805135,6.774154,7.4699492,7.6143594,8.904206,10.902975,13.174155,15.284514,17.529438,18.865232,19.498669,19.62995,19.459284,18.65518,16.580925,14.788924,13.804309,13.108514,15.238565,15.432206,12.987078,10.010257,11.414975,15.323898,18.418873,21.11672,23.752207,26.555079,24.969849,22.869335,20.401232,17.792002,15.330462,15.770258,17.371899,19.459284,21.4679,22.944822,26.325335,35.59713,43.805542,44.56698,32.09518,29.19713,28.389746,26.016823,22.695387,23.305847,26.177643,27.552822,28.304413,27.657848,23.187695,17.8839,15.540514,13.239796,10.322052,8.369231,7.4010262,6.7282057,5.5696416,4.2305646,4.1156926,4.279795,5.044513,6.692103,8.549745,8.982975,8.717129,10.555078,12.950975,13.755078,10.200616,8.3823595,6.567385,5.431795,5.1200004,5.277539,6.1341543,8.598975,11.529847,13.8075905,14.319591,15.412514,14.546052,12.822975,11.286975,10.912822,11.21477,14.854566,15.652103,14.611693,19.925335,19.958155,17.946259,16.049232,15.885129,18.54359,22.14072,20.847591,23.568413,30.614977,33.70667,31.629131,35.367386,40.90421,45.843697,49.424416,66.63221,74.223595,88.66462,110.506676,124.41273,117.58934,99.28206,78.336006,61.43672,53.087185,44.65231,40.546463,37.64185,35.679184,37.264412,35.41662,29.827284,25.366976,22.85949,19.078566,14.36554,8.310155,4.532513,3.6036925,3.0326157,2.100513,1.6082052,1.5425643,1.6738462,1.5589745,2.7798977,1.7952822,3.0096412,5.412103,2.5895386,2.2547693,9.435898,10.499283,6.2785645,12.06154,13.243078,6.547693,4.578462,8.828718,9.688616,11.874462,8.621949,7.4765134,9.770667,10.624001,6.5312824,6.6560006,5.612308,3.2032824,4.4242053,5.405539,4.640821,4.640821,5.5302567,5.0477953,3.045744,2.5600002,3.308308,4.9394875,7.026872,3.1343591,6.045539,7.4863596,5.0018463,1.9692309,1.7558975,1.5392822,1.3357949,1.2012309,1.2373334,1.332513,1.3062565,1.1684103,1.024,1.1060513,1.4802053,1.4802053,1.3095386,1.0272821,0.5284103,0.5513847,0.64000005,0.702359,0.7187693,0.764718,0.83035904,0.8041026,0.69251287,0.5415385,0.43651286,0.33476925,0.3052308,0.30851284,0.37415388,0.5874872,1.0272821,1.020718,0.764718,0.48902568,0.4397949,0.5513847,0.50543594,0.6071795,0.92225647,1.273436,1.0666667,0.86646163,0.93866676,1.1093334,0.7581539,0.31507695,0.40369233,0.58420515,0.6498462,0.6170257,0.571077,0.58420515,0.5874872,0.6498462,0.98133343,0.9419488,0.65969235,0.5218462,0.5940513,0.636718,0.3314872,0.15753847,0.098461546,0.08861539,0.04266667,0.013128206,0.072205134,0.11158975,0.08861539,0.009846155,0.013128206,0.14441027,0.20020515,0.12143591,0.0,0.19364104,0.24615386,0.19692309,0.0951795,0.0,0.0,0.0,0.0,0.0,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.029538464,0.29210258,0.47589746,0.42338464,0.13456412,0.17066668,0.072205134,0.0,0.0032820515,0.009846155,0.009846155,0.029538464,0.055794876,0.06235898,0.01969231,0.0032820515,0.009846155,0.02297436,0.029538464,0.006564103,0.013128206,0.049230773,0.07548718,0.06564103,0.013128206,0.02297436,0.016410258,0.03938462,0.0951795,0.16410258,0.059076928,0.026256412,0.04594872,0.06564103,0.006564103,0.009846155,0.009846155,0.006564103,0.0032820515,0.0,0.0,0.009846155,0.032820515,0.04594872,0.009846155,0.049230773,0.055794876,0.032820515,0.009846155,0.02297436,0.072205134,0.098461546,0.098461546,0.22646156,0.7844103,0.21333335,0.032820515,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02297436,0.02297436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.026256412,0.02297436,0.0,0.0,0.036102567,0.08533334,0.18707694,0.31507695,0.39712822,0.4397949,0.46933338,0.5218462,0.5940513,0.6695385,0.7417436,0.8336411,0.9353847,1.0535386,1.1881026,1.4473847,1.6082052,1.4769232,1.1060513,0.8008206,0.5152821,0.31507695,0.18707694,0.118153855,0.098461546,0.055794876,0.049230773,0.055794876,0.08861539,0.18707694,0.35774362,0.67610264,0.827077,0.7515898,0.6432821,0.28882053,0.14769232,0.2231795,0.47589746,0.81066674,0.7450257,0.6695385,0.65312827,0.69251287,0.7089231,0.7581539,0.69251287,0.62030774,0.5907693,0.58092314,0.6268718,0.5546667,0.60389745,0.7975385,0.9682052,1.339077,1.2373334,0.9353847,0.65969235,0.5973334,0.7187693,0.8795898,0.8992821,0.79425645,0.7417436,0.74830776,0.79425645,0.75487185,0.6629744,0.69579494,1.014154,1.0075898,0.9485129,0.90912825,0.7515898,0.9878975,1.1224617,1.0765129,0.9288206,0.9189744,1.0010257,0.9747693,0.9156924,0.88287187,0.90256417,0.9682052,1.0436924,1.1454359,1.2668719,1.3686155,1.2635899,1.5064616,1.6278975,1.5491283,1.5753847,1.3883078,1.1520001,0.9517949,0.83035904,0.7844103,0.9156924,0.9682052,0.9714873,0.98461545,1.0994873,0.8992821,0.84348726,0.8763078,0.9485129,1.014154,1.0633847,1.0404103,1.0568206,1.1290257,1.1913847,0.95835906,0.8467693,0.81394875,0.81394875,0.79097444,0.8598975,0.85005134,0.88287187,0.9944616,1.142154,1.1027694,1.1224617,0.9878975,0.7811283,0.88943595,1.0404103,1.0305642,1.0075898,1.0010257,0.9124103,0.7187693,0.69251287,0.7318975,0.83035904,1.0601027,0.8041026,0.6465641,0.5973334,0.5940513,0.508718,0.39384618,0.39056414,0.4397949,0.49887183,0.571077,0.6859488,0.8041026,0.90256417,0.9616411,0.95835906,0.8467693,0.8172308,0.9616411,1.2996924,1.7690258,1.585231,1.5425643,1.5261539,1.6082052,2.041436,1.5786668,1.3292309,1.2307693,1.276718,1.5195899,1.1257436,0.93866676,0.8369231,0.764718,0.7384616,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01969231,0.072205134,0.18051283,0.12143591,0.04266667,0.029538464,0.101743594,0.23302566,0.45292312,0.5349744,0.446359,0.26912823,0.21661541,0.27897438,0.4135385,0.38728207,0.25928208,0.38728207,0.57764107,0.8566154,1.014154,1.020718,1.020718,1.0633847,0.9189744,0.92225647,1.0896411,1.1191796,0.44307697,0.37415388,0.69579494,1.3357949,2.353231,3.9712822,7.4404106,12.251899,16.922258,18.999796,21.494156,25.34072,28.57026,30.50995,31.766977,34.566566,37.714054,38.268723,36.417645,35.485542,47.222157,64.607185,76.832825,74.91939,51.731697,37.825645,29.489233,24.018053,21.956924,27.11631,25.954464,24.113234,23.302567,23.194258,21.408823,22.12431,22.787283,22.711796,22.212925,22.593643,22.86277,25.439182,27.464207,27.090054,23.463387,21.769848,24.70072,24.454565,20.611284,20.138668,20.361847,21.828924,23.5159,24.868105,25.83631,24.201847,23.3879,22.150566,21.22831,23.361643,27.001438,27.913849,26.020105,22.836515,21.461334,22.029129,21.897848,20.814772,19.360823,18.944002,18.694565,18.12349,16.466053,14.565744,14.8709755,15.734155,14.5263605,13.443283,13.22995,13.177437,12.557129,10.072617,8.090257,7.2631803,6.5083084,5.1922054,5.35959,6.235898,7.0498466,7.059693,6.9087186,6.744616,6.806975,7.072821,7.2369237,7.282872,7.9524107,8.664616,9.344001,10.443488,12.619488,13.922462,14.592001,14.503386,13.157744,10.453334,8.766359,8.162462,8.395488,8.904206,9.40636,11.034257,12.678565,14.024206,15.53395,17.237335,17.51631,15.635694,11.930258,7.7981544,5.6451287,4.4767184,4.3552823,5.149539,6.49518,7.5946674,9.160206,11.067078,13.167591,15.281232,16.899282,17.536001,17.45395,17.060104,16.918976,16.672821,13.243078,10.525539,9.613129,8.786052,12.235488,14.608412,15.143386,13.833847,11.414975,14.293334,19.889233,25.311182,28.327387,27.342772,23.177849,21.523693,20.09272,18.868515,20.09272,22.291695,25.544207,29.522053,33.394875,35.83016,36.8279,49.204517,64.8238,70.610054,48.580925,40.776207,37.49744,31.291079,22.65272,20.033642,26.4599,26.853746,23.371489,18.133335,13.206975,11.812103,12.740924,12.655591,11.23118,11.175385,11.139283,9.593436,7.7423596,6.298257,5.4547696,6.3212314,7.3321033,9.104411,11.030975,11.277129,9.3768215,11.621744,16.36431,19.99754,16.932104,12.593232,10.256411,9.291488,8.989539,8.579283,8.648206,9.747693,12.288001,15.113848,15.520822,16.400412,15.606155,14.27036,13.37436,13.751796,9.947898,11.720206,12.609642,11.510155,12.681848,14.641232,16.86318,19.652925,23.14831,27.303387,28.416002,24.766361,23.341951,25.892105,28.914873,30.82831,35.029335,38.20308,41.330875,49.680412,69.989746,80.04924,96.794266,121.3998,139.27715,125.44985,105.101135,85.4318,71.3157,65.276726,49.19467,43.565952,40.946877,39.30913,42.02667,38.44267,31.291079,26.725746,24.832003,19.639797,13.978257,8.349539,5.0149746,4.132103,3.7349746,2.5632823,1.9331284,1.7887181,1.9068719,1.8642052,2.3630772,2.048,6.2490263,10.804514,2.0611284,2.612513,8.169026,8.920616,5.723898,10.118565,12.25518,6.229334,4.5029745,9.288206,12.540719,14.14236,9.26195,7.522462,10.729027,12.855796,7.5585647,8.277334,8.080411,5.346462,3.754667,5.284103,5.3202057,5.658257,6.422975,6.0980515,3.6562054,2.169436,2.4746668,3.9286156,4.4242053,1.782154,4.571898,6.2851286,4.8771286,2.7667694,1.6410258,1.2931283,1.1323078,0.95835906,0.9485129,1.1520001,0.9714873,0.761436,0.79425645,1.276718,1.7493335,1.7263591,1.4112822,0.955077,0.44964105,0.4594872,0.4594872,0.35446155,0.19364104,0.16738462,0.2231795,0.25271797,0.26256412,0.27569234,0.35774362,0.25271797,0.18707694,0.16082053,0.18707694,0.28882053,0.7450257,0.81394875,0.6301539,0.38400003,0.32820517,0.48246157,0.45620516,0.46276927,0.7318975,1.5031796,1.211077,0.80738467,0.7187693,0.88615394,0.78769237,0.38400003,0.4201026,0.55794877,0.73517954,1.1651284,0.77456415,0.5481026,0.4266667,0.46933338,0.8467693,0.8992821,0.6071795,0.446359,0.57764107,0.8763078,0.61374366,0.318359,0.14441027,0.1148718,0.128,0.059076928,0.032820515,0.03938462,0.052512825,0.009846155,0.03938462,0.13784617,0.19692309,0.16410258,0.036102567,0.029538464,0.11158975,0.16738462,0.14441027,0.04266667,0.009846155,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.01969231,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.08205129,0.25271797,0.39712822,0.256,0.20348719,0.08205129,0.0032820515,0.0032820515,0.016410258,0.009846155,0.03938462,0.08205129,0.11158975,0.06564103,0.013128206,0.07548718,0.190359,0.24943592,0.09189744,0.026256412,0.009846155,0.006564103,0.0,0.0,0.06235898,0.036102567,0.03938462,0.10502565,0.15753847,0.068923086,0.036102567,0.049230773,0.06564103,0.01969231,0.009846155,0.006564103,0.0032820515,0.0,0.0,0.0,0.013128206,0.04266667,0.059076928,0.009846155,0.098461546,0.1148718,0.08205129,0.04594872,0.08533334,0.11158975,0.118153855,0.108307704,0.22646156,0.74830776,0.21989745,0.059076928,0.03938462,0.036102567,0.006564103,0.006564103,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02297436,0.02297436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.026256412,0.02297436,0.0,0.0,0.036102567,0.03938462,0.098461546,0.21989745,0.2986667,0.3511795,0.380718,0.44964105,0.53825647,0.571077,0.7089231,0.80738467,0.90256417,0.9878975,1.0338463,1.2209232,1.6475899,1.7657437,1.4703591,1.0732309,0.5907693,0.318359,0.18707694,0.13128206,0.098461546,0.07548718,0.052512825,0.04266667,0.06564103,0.15097436,0.26256412,0.45292312,0.7089231,0.88943595,0.7187693,0.2986667,0.14112821,0.16738462,0.318359,0.5677949,0.6629744,0.81394875,0.90912825,0.90584624,0.8598975,0.7844103,0.69907695,0.6301539,0.61374366,0.702359,0.69907695,0.6268718,0.55794877,0.54482055,0.62030774,0.98133343,0.69907695,0.4397949,0.446359,0.512,0.62030774,0.7811283,0.82379496,0.7581539,0.7844103,0.77128214,0.8402052,0.8336411,0.7581539,0.79425645,1.142154,1.2012309,1.1158975,0.95835906,0.7318975,0.90912825,1.014154,0.9714873,0.8402052,0.81394875,0.8598975,0.86974365,0.8533334,0.8172308,0.7811283,0.86317956,0.94523084,1.0436924,1.1684103,1.3161026,1.2898463,1.5885129,1.7788719,1.723077,1.5622566,1.3489232,1.0994873,0.92225647,0.8730257,0.9747693,1.0896411,0.9714873,0.88943595,0.9189744,0.9517949,0.69907695,0.6629744,0.7187693,0.78769237,0.8467693,1.024,1.0896411,1.1060513,1.1224617,1.1520001,0.8205129,0.65312827,0.5874872,0.574359,0.57764107,0.76800007,0.7515898,0.76800007,0.90912825,1.1224617,1.1585642,1.1060513,0.94523084,0.79425645,0.9353847,1.014154,0.97805136,0.8992821,0.82379496,0.7844103,0.69251287,0.6695385,0.6695385,0.7220513,0.9189744,0.78769237,0.6465641,0.5513847,0.4955898,0.4004103,0.33805132,0.34133336,0.38400003,0.446359,0.5284103,0.63343596,0.7417436,0.86317956,0.9288206,0.78769237,0.7515898,0.76800007,0.88943595,1.142154,1.4966155,1.5163078,1.4473847,1.4572309,1.595077,1.8051283,1.5819489,1.2373334,1.1027694,1.2340513,1.404718,1.1158975,1.0962052,1.0601027,0.9419488,0.88615394,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.04266667,0.16738462,0.101743594,0.032820515,0.02297436,0.08861539,0.2297436,0.53825647,0.60389745,0.40697438,0.11158975,0.06564103,0.055794876,0.118153855,0.2297436,0.37415388,0.54482055,0.60389745,0.9288206,1.1257436,1.1257436,1.1782565,1.0371283,0.7515898,0.46933338,0.27569234,0.18707694,0.19692309,0.34133336,0.6892308,1.522872,3.3312824,5.293949,8.139488,11.234463,14.614976,18.98995,23.391182,26.564924,29.128208,31.570053,34.274464,40.598976,46.959595,46.788925,39.857235,32.262566,39.37477,51.28862,56.349545,49.664005,33.106052,27.638157,23.364925,20.594873,21.346462,29.331694,31.27467,30.083284,27.736618,24.996105,21.385847,21.241438,22.275284,23.256617,24.201847,26.368002,28.806566,32.07221,32.495594,29.029745,23.23036,23.09908,23.896618,23.509335,22.09477,22.075079,22.081642,24.631796,27.477335,28.983797,28.110771,27.559387,26.246567,24.277336,22.324514,21.622156,23.02031,24.159182,23.808002,22.186668,20.982155,22.567387,23.473232,22.836515,20.98872,19.462566,18.500925,15.894976,14.076719,14.070155,15.504412,15.419078,14.020925,12.868924,12.475078,12.320822,11.053949,9.186462,7.899898,7.0990777,5.421949,4.9985647,5.579488,6.3442054,7.1154876,8.369231,8.966565,8.119796,7.532308,7.7718983,8.283898,8.864821,9.409642,10.06277,10.935796,12.087796,14.503386,16.272411,17.46708,17.631182,15.75713,11.730052,9.908514,9.701744,10.387693,11.132719,13.075693,15.0088215,16.66954,17.929848,18.7799,17.122463,13.282462,8.723693,4.903385,3.2361028,2.5271797,2.6880002,3.4231799,4.5554876,6.0225644,7.4240007,8.756514,9.796924,10.748719,12.2847185,13.590976,14.775796,14.76595,13.922462,14.034052,15.24513,12.025436,9.278359,8.356103,7.059693,10.496001,14.641232,20.86072,24.969849,17.24718,19.62995,24.914053,30.076721,32.577644,30.385233,26.456617,24.802464,22.912003,22.403284,29.003489,31.875284,36.158363,41.199593,45.46298,46.53621,42.207184,50.356518,66.560005,76.26831,54.81354,50.3598,52.66708,47.245132,32.403694,19.249231,28.898464,32.41354,28.317541,19.603693,13.728822,13.948719,14.381949,14.099693,14.25395,18.054565,17.962667,14.260514,11.057232,9.517949,7.8473854,10.31877,10.788103,11.352616,12.914873,15.179488,15.494565,17.046976,21.779694,27.506874,27.910566,22.66913,17.946259,14.549335,12.662155,11.861334,11.572514,11.684103,13.587693,16.551386,17.736206,17.552412,17.985641,17.414566,15.855591,14.972719,12.383181,9.82318,8.533334,8.539898,8.651488,8.904206,12.534155,19.186872,26.994873,32.58421,28.196104,23.14831,18.546873,16.196924,18.609232,22.426258,26.607592,30.880823,38.288414,55.19098,76.73765,88.19529,101.179085,117.63857,129.85437,112.10175,93.74852,80.03939,73.85272,75.67754,53.730465,45.092106,42.164516,41.71816,44.918156,41.439182,32.99118,27.37231,25.288208,20.325745,15.350155,9.764103,6.373744,5.602462,5.504,5.1364107,5.3366156,4.4242053,2.6683078,2.297436,3.1343591,3.0391798,9.636104,16.118155,1.270154,2.7569232,5.7764106,6.012718,4.2174363,6.2227697,7.6570263,4.2962055,2.5140514,4.7655387,9.577026,10.55836,8.749949,8.720411,10.935796,11.739899,8.139488,9.051898,9.573745,7.650462,4.06318,4.1878977,4.9920006,6.5411286,7.9885135,7.565129,3.7743592,1.7132308,1.8084104,3.045744,2.993231,2.2514873,1.9298463,1.7099489,1.657436,2.231795,1.4605129,1.1388719,1.0305642,0.9878975,0.9714873,0.8467693,0.6235898,0.47917953,0.62030774,1.2800001,1.3817437,1.4703591,1.2209232,0.69251287,0.3314872,0.48246157,0.42338464,0.34133336,0.29210258,0.2100513,0.2100513,0.23958977,0.22646156,0.18379489,0.19692309,0.20676924,0.16082053,0.15425642,0.20020515,0.21661541,0.44964105,0.52512825,0.42994875,0.26912823,0.23958977,0.2855385,0.3314872,0.36102566,0.56451285,1.339077,1.0994873,0.7417436,0.58420515,0.6629744,0.7089231,0.4266667,0.3708718,0.446359,0.7581539,1.5885129,0.82379496,0.49887183,0.40697438,0.47261542,0.7318975,0.81394875,0.5874872,0.380718,0.4266667,0.8730257,0.8566154,0.51856416,0.2100513,0.10502565,0.20020515,0.13784617,0.06235898,0.013128206,0.0,0.0,0.101743594,0.09189744,0.08533334,0.108307704,0.108307704,0.059076928,0.032820515,0.059076928,0.11158975,0.101743594,0.02297436,0.009846155,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.036102567,0.029538464,0.013128206,0.0032820515,0.0,0.0,0.0,0.052512825,0.17394873,0.31507695,0.3708718,0.190359,0.072205134,0.013128206,0.0032820515,0.013128206,0.0032820515,0.013128206,0.052512825,0.098461546,0.108307704,0.02297436,0.14112821,0.39056414,0.56123084,0.3117949,0.10502565,0.026256412,0.006564103,0.0,0.0,0.108307704,0.07876924,0.07548718,0.14769232,0.2297436,0.17394873,0.098461546,0.052512825,0.052512825,0.06564103,0.036102567,0.01969231,0.009846155,0.0032820515,0.0,0.0,0.006564103,0.02297436,0.032820515,0.0,0.118153855,0.15753847,0.13784617,0.11158975,0.17394873,0.0951795,0.055794876,0.049230773,0.052512825,0.029538464,0.049230773,0.072205134,0.08861539,0.08861539,0.059076928,0.06564103,0.026256412,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.04266667,0.118153855,0.23302566,0.2986667,0.28225642,0.3249231,0.44307697,0.51856416,0.71548724,0.8205129,0.90256417,0.9911796,1.0633847,1.0765129,1.4769232,1.8051283,1.8084104,1.4112822,0.7417436,0.3708718,0.20348719,0.15425642,0.118153855,0.1148718,0.068923086,0.04594872,0.06564103,0.1148718,0.18051283,0.35446155,0.636718,0.86646163,0.71548724,0.39056414,0.190359,0.13128206,0.18379489,0.28882053,0.4660513,0.8566154,1.0699488,0.9944616,0.8172308,0.7187693,0.65312827,0.6104616,0.6071795,0.6859488,0.6629744,0.62030774,0.5973334,0.57764107,0.49887183,0.4397949,0.43323082,0.35774362,0.256,0.35774362,0.4660513,0.52512825,0.6071795,0.73517954,0.8730257,0.79425645,0.85005134,0.86646163,0.81394875,0.81394875,1.014154,1.1618463,1.1388719,0.9517949,0.7122052,0.74830776,0.71548724,0.6662565,0.65312827,0.7220513,0.7417436,0.79425645,0.83035904,0.78769237,0.62030774,0.73517954,0.8533334,0.97805136,1.1191796,1.2832822,1.4802053,1.782154,1.9462565,1.8674873,1.5556924,1.3259488,1.1158975,0.9911796,1.0305642,1.3128207,1.2898463,0.92225647,0.7056411,0.75487185,0.7975385,0.5973334,0.6071795,0.65969235,0.69251287,0.761436,0.98461545,1.0633847,1.079795,1.0601027,0.9616411,0.6629744,0.55794877,0.56123084,0.5874872,0.5415385,0.6498462,0.62030774,0.6104616,0.67610264,0.77128214,1.0010257,1.0568206,0.98461545,0.90912825,1.020718,0.9353847,0.8205129,0.7089231,0.6268718,0.60061544,0.65641034,0.69579494,0.65312827,0.5513847,0.51856416,0.60061544,0.58092314,0.51856416,0.43651286,0.3117949,0.3249231,0.32164106,0.3446154,0.40369233,0.46276927,0.5415385,0.65641034,0.80738467,0.90256417,0.7581539,0.7220513,0.7844103,0.9485129,1.1815386,1.3981539,1.5163078,1.4605129,1.3423591,1.2176411,1.079795,1.3817437,1.1126155,0.9517949,1.0666667,1.1126155,1.0896411,1.2931283,1.3456411,1.1881026,1.0666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02297436,0.0951795,0.2297436,0.04594872,0.0,0.013128206,0.08205129,0.28882053,0.571077,0.5415385,0.30851284,0.06564103,0.09189744,0.09189744,0.072205134,0.1148718,0.23958977,0.4135385,0.7056411,1.0075898,1.4834872,2.03159,2.28759,1.2865642,0.73517954,0.5513847,0.47917953,0.07548718,0.3708718,0.71548724,1.0962052,2.356513,6.226052,7.6898465,9.613129,12.895181,17.329231,21.592617,27.585644,30.365541,31.744003,33.444103,37.093746,45.380928,54.79713,53.65498,41.137234,27.283695,30.372105,35.347694,35.085133,28.248617,19.288616,20.263386,20.33559,20.680206,23.361643,31.294361,33.736206,33.358772,31.448618,27.588924,19.652925,21.11672,22.298258,23.305847,24.841848,28.199387,28.770464,29.298874,28.297848,25.721437,22.948105,26.78154,27.759592,26.758566,25.810053,28.107489,30.976002,35.892517,38.114464,35.971283,30.867695,27.329643,25.261951,24.507078,24.441439,24.001642,26.601028,27.168823,26.089027,24.841848,26.000412,26.404104,24.986258,23.427284,22.22277,20.660515,20.036924,17.329231,15.02195,14.431181,15.701335,13.906053,12.724514,11.762873,10.660104,9.110975,8.828718,7.680001,6.5378466,5.5696416,4.2272825,4.788513,6.1013336,7.7718983,9.357129,10.345026,9.478565,8.648206,8.5891285,9.173334,9.429334,9.80677,10.203898,11.546257,14.040616,17.165129,20.900105,22.741335,22.20308,19.272207,14.388514,10.617436,9.77395,10.781539,12.964104,16.052513,18.395899,19.623386,19.311592,17.54913,14.923489,10.686359,7.322257,4.5128207,2.4549747,1.8313848,1.8543591,2.1989746,2.9210258,4.056616,5.6320004,7.4141545,9.340718,9.7673855,8.841846,8.500513,11.378873,14.004514,13.466257,10.555078,9.750975,8.822155,8.507077,7.9097443,7.634052,9.780514,14.368821,24.004925,33.588516,37.353027,28.868925,23.975386,23.722668,27.700516,36.02708,49.329235,50.832413,46.116108,39.48308,35.741543,40.221542,35.584003,35.889233,37.79939,38.114464,33.769028,37.16267,43.01785,45.929028,42.27939,30.230976,35.55118,52.480003,61.581135,52.831184,25.632822,28.662155,35.92862,38.6199,34.3959,27.38872,28.097643,23.348515,18.159592,15.711181,17.332514,15.028514,11.933539,11.296822,13.184001,14.464001,18.369642,14.54277,9.892103,9.002667,14.129231,20.78195,23.7719,26.325335,30.01108,34.76021,38.482056,30.194874,18.914463,11.021129,10.240001,14.401642,16.403694,18.763489,21.16595,20.447182,18.346668,20.634258,22.390156,21.35631,17.913437,16.498873,14.486976,11.96636,9.055181,5.904411,6.088206,8.303591,11.191795,15.737437,25.284925,22.636309,18.36636,16.20349,17.890463,23.161438,25.701746,26.942362,30.358976,39.345234,57.206158,79.9836,93.06586,99.58401,100.16493,92.92801,81.85765,71.939285,65.77888,65.729645,73.88226,54.52144,44.737644,40.0279,38.961235,43.19836,41.62298,33.21108,25.317745,20.985437,18.921026,17.332514,13.210258,9.878975,8.726975,9.216001,12.793437,17.385027,13.722258,4.2272825,3.006359,1.9068719,2.3204105,10.492719,17.969233,1.5885129,1.3062565,2.353231,4.33559,6.2818465,6.636308,5.7107697,3.6463592,2.3269746,2.5928206,4.2436924,6.36718,10.246565,12.701539,12.288001,9.324308,6.2096415,7.5388722,8.5202055,7.515898,6.0258465,4.31918,4.338872,7.6734366,11.628308,9.26195,4.023795,2.9440002,2.284308,1.5524104,3.495385,4.0303593,2.537026,1.1388719,0.764718,1.1454359,0.99774367,1.0633847,1.1946667,1.2274873,0.94523084,0.8598975,0.7581539,0.6465641,0.571077,0.5940513,0.62030774,0.7187693,0.6695385,0.44307697,0.19692309,0.30851284,0.3249231,0.380718,0.41682056,0.19692309,0.24615386,0.3249231,0.2855385,0.18707694,0.25928208,0.25928208,0.18707694,0.15425642,0.16738462,0.108307704,0.15425642,0.31507695,0.38728207,0.2986667,0.09189744,0.128,0.13784617,0.16082053,0.30194873,0.7187693,0.69251287,0.61374366,0.5218462,0.48902568,0.6104616,0.37743592,0.34789747,0.34133336,0.45620516,1.0535386,0.6859488,0.7318975,0.7187693,0.5874872,0.67282057,0.7811283,0.75487185,0.54482055,0.2855385,0.27569234,0.6301539,0.5513847,0.30194873,0.09189744,0.09189744,0.16410258,0.108307704,0.036102567,0.0,0.0,0.12143591,0.19692309,0.15425642,0.072205134,0.18379489,0.072205134,0.01969231,0.029538464,0.07548718,0.07548718,0.026256412,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.016410258,0.009846155,0.0,0.0,0.0,0.009846155,0.026256412,0.07548718,0.19692309,0.3314872,0.17394873,0.026256412,0.0,0.0,0.0,0.0,0.0,0.009846155,0.04594872,0.02297436,0.016410258,0.13784617,0.38400003,0.64000005,0.33476925,0.13128206,0.026256412,0.0,0.0,0.049230773,0.108307704,0.19364104,0.31507695,0.47261542,0.44964105,0.23302566,0.055794876,0.026256412,0.13784617,0.08861539,0.03938462,0.016410258,0.013128206,0.0,0.0,0.0,0.013128206,0.02297436,0.0,0.013128206,0.098461546,0.13456412,0.12471796,0.19692309,0.052512825,0.02297436,0.08533334,0.15097436,0.09189744,0.04266667,0.07548718,0.08861539,0.0951795,0.2297436,0.26584616,0.108307704,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.06235898,0.18379489,0.21989745,0.2100513,0.23630771,0.3249231,0.45620516,0.51856416,0.5874872,0.6859488,0.8041026,0.9156924,1.086359,1.3128207,1.6246156,1.847795,1.6180514,1.0666667,0.5907693,0.27569234,0.14441027,0.16738462,0.14441027,0.101743594,0.07548718,0.07876924,0.09189744,0.16410258,0.28225642,0.45620516,0.6662565,0.88615394,0.7253334,0.35774362,0.108307704,0.08205129,0.16738462,0.4594872,0.77128214,0.90584624,0.8172308,0.6104616,0.65969235,0.67938465,0.6071795,0.47917953,0.44307697,0.56451285,0.64000005,0.7450257,0.8041026,0.5940513,0.49887183,0.41025645,0.318359,0.25928208,0.32164106,0.380718,0.39712822,0.46933338,0.6301539,0.82379496,0.77456415,0.80738467,0.81394875,0.764718,0.7187693,0.7778462,0.92225647,0.93866676,0.7975385,0.6268718,0.56451285,0.5218462,0.49887183,0.5284103,0.6859488,0.77128214,0.83035904,0.8041026,0.7056411,0.5940513,0.6432821,0.7581539,0.8730257,0.96492314,1.0371283,1.5392822,2.048,2.2416413,2.0217438,1.4966155,1.5064616,1.4473847,1.270154,1.0436924,0.94523084,0.98133343,0.827077,0.7220513,0.761436,0.86974365,0.69907695,0.7122052,0.72861546,0.6859488,0.6268718,0.7220513,0.7122052,0.7220513,0.7778462,0.7778462,0.65641034,0.6892308,0.7318975,0.6859488,0.5021539,0.4660513,0.4660513,0.5152821,0.60061544,0.6859488,0.761436,0.8041026,0.78769237,0.7417436,0.7778462,0.67938465,0.5546667,0.53825647,0.60061544,0.56451285,0.6498462,0.65312827,0.574359,0.46933338,0.45620516,0.46933338,0.46276927,0.45292312,0.43323082,0.39712822,0.4201026,0.41682056,0.41682056,0.4266667,0.4266667,0.4266667,0.46276927,0.512,0.574359,0.67282057,0.69579494,0.93866676,1.2274873,1.4473847,1.5556924,1.5064616,1.3686155,1.0502565,0.6892308,0.64000005,0.77456415,0.88287187,1.0765129,1.2471796,1.0535386,1.0272821,1.1520001,1.2242053,1.1782565,1.0666667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02297436,0.026256412,0.01969231,0.04594872,0.009846155,0.0,0.006564103,0.059076928,0.21661541,0.3511795,0.29210258,0.15753847,0.049230773,0.04266667,0.032820515,0.032820515,0.04266667,0.08861539,0.2297436,0.65969235,1.1257436,1.5524104,1.8740515,2.03159,1.0994873,0.7975385,0.8369231,0.9124103,0.73517954,0.6465641,0.7318975,1.3161026,3.006359,6.688821,9.373539,11.792411,16.630156,23.433847,28.622772,32.055798,34.103798,35.87282,38.012722,40.694157,47.264824,50.57313,45.952003,35.252514,26.857027,29.971695,30.79549,28.389746,23.588104,18.983387,19.206566,20.4439,22.997335,26.345028,29.121643,30.519796,32.26913,32.298668,29.266054,22.534565,22.806976,23.42072,24.97313,27.359182,29.748514,31.396105,34.888206,36.562054,36.752415,39.781746,47.55036,54.97436,54.6199,45.98154,35.456,38.166977,47.140106,59.05067,66.62565,58.660107,42.436928,31.172926,24.615387,21.507284,19.584002,21.54995,24.198566,25.744411,25.53436,24.047592,22.291695,21.264412,21.382566,21.481028,18.806156,18.09395,16.689232,15.051488,13.584412,12.63918,11.936821,12.324103,11.798975,10.236719,9.38995,9.225847,7.6143594,5.858462,4.6539493,4.092718,4.9362054,6.518154,7.7259493,8.080411,7.722667,8.464411,8.930462,9.314463,9.573745,9.429334,11.155693,13.046155,15.130258,17.168411,18.642054,18.91118,18.048002,16.489027,14.506668,12.1928215,12.130463,13.213539,15.497848,18.372925,20.545643,20.368412,18.891489,16.925539,14.8939495,12.836103,8.677744,6.245744,4.824616,3.7218463,2.2580514,2.2055387,2.7798977,3.9056413,5.612308,8.04759,12.524308,14.027489,12.471796,9.347282,7.706257,7.5881033,7.4797955,7.312411,7.3714876,8.274052,8.789334,13.400617,19.275488,26.016823,35.646362,41.649235,45.16431,46.244106,43.05067,31.872002,28.8919,29.476105,38.590363,58.41067,88.31673,105.51139,97.49006,74.046364,48.705647,38.744617,27.897438,25.573746,27.27713,29.072412,27.579079,27.270567,27.641438,26.157951,22.176823,16.922258,21.582771,32.239594,39.040005,34.94072,15.711181,13.8075905,21.943796,28.17313,29.092104,29.817438,33.650875,29.187284,21.13313,16.06236,22.41313,23.092514,19.413334,13.801026,8.812308,7.1056414,10.210463,11.116308,11.523283,14.54277,24.687592,40.930466,41.22913,37.710773,36.36185,37.01826,43.825233,40.85826,30.276926,17.621334,11.802258,15.826053,17.588514,17.657436,17.391592,18.944002,17.752617,19.35754,22.186668,22.816822,15.986873,19.948309,19.18031,15.714462,11.306667,7.4436927,6.3967185,8.2904625,10.492719,11.848206,12.675283,22.006155,24.82872,23.364925,23.066257,32.597336,34.169437,38.866055,46.03734,53.51713,57.606567,65.34893,75.38216,81.7198,80.764725,71.309135,61.09539,55.53231,54.20308,55.220516,55.233646,44.36677,40.237953,37.113438,34.162876,35.459286,34.31385,28.616207,23.003899,19.029335,15.163078,16.971489,14.621539,12.875488,12.412719,9.826463,10.269539,16.866463,14.470565,3.9876926,2.3958976,1.4834872,1.9200002,4.844308,7.2631803,2.0512822,3.1573336,4.709744,7.3091288,8.854975,4.562052,5.5696416,4.3027697,2.6617439,2.1891284,4.069744,5.6287184,6.8496413,8.283898,10.023385,11.716924,8.651488,6.7905645,6.3376417,7.072821,8.346257,6.2162056,3.95159,4.325744,6.3507695,5.2709746,6.058667,5.648411,3.7448208,1.8871796,3.4592824,3.058872,2.4484105,1.5589745,0.8369231,1.2537436,0.9419488,0.9353847,1.1323078,1.3686155,1.4112822,1.0404103,0.88287187,0.77128214,0.6301539,0.44964105,0.48246157,0.69251287,0.6892308,0.4594872,0.380718,0.3249231,0.24943592,0.33476925,0.47261542,0.28225642,0.21661541,0.3511795,0.54482055,0.6432821,0.49230772,0.2855385,0.17066668,0.118153855,0.098461546,0.04594872,0.055794876,0.118153855,0.16410258,0.16082053,0.09189744,0.108307704,0.15097436,0.14112821,0.13456412,0.31507695,0.8172308,0.65641034,0.5415385,0.7318975,1.0502565,0.7778462,0.827077,0.7384616,0.512,0.60061544,0.42994875,0.42994875,0.43323082,0.41025645,0.47589746,0.53825647,0.6432821,0.7450257,0.74830776,0.5316923,0.39712822,0.32164106,0.26256412,0.18379489,0.06564103,0.052512825,0.06235898,0.049230773,0.009846155,0.0,0.190359,0.20348719,0.14441027,0.10502565,0.14769232,0.07548718,0.03938462,0.049230773,0.08533334,0.07548718,0.036102567,0.01969231,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0032820515,0.006564103,0.016410258,0.03938462,0.15425642,0.12143591,0.049230773,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.0032820515,0.0032820515,0.036102567,0.12143591,0.24943592,0.23958977,0.12143591,0.026256412,0.0,0.0,0.009846155,0.101743594,0.16738462,0.26256412,0.6071795,0.827077,0.508718,0.2100513,0.15097436,0.2100513,0.101743594,0.04594872,0.016410258,0.0032820515,0.0,0.0,0.0,0.006564103,0.013128206,0.0,0.0032820515,0.01969231,0.032820515,0.036102567,0.03938462,0.009846155,0.026256412,0.068923086,0.12471796,0.20020515,0.07548718,0.036102567,0.059076928,0.13456412,0.27897438,0.19692309,0.2231795,0.15425642,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.02297436,0.098461546,0.13456412,0.15425642,0.17723078,0.21989745,0.27569234,0.3446154,0.39712822,0.46933338,0.5973334,0.8041026,1.0436924,1.1552821,1.3456411,1.5556924,1.4703591,1.1552821,0.7975385,0.48574364,0.27569234,0.19364104,0.128,0.07548718,0.06564103,0.0951795,0.128,0.190359,0.30194873,0.512,0.827077,1.2012309,1.1913847,0.6071795,0.16410258,0.08861539,0.15425642,0.3314872,0.4660513,0.53825647,0.5874872,0.7318975,0.8598975,0.7975385,0.65641034,0.5021539,0.3708718,0.5415385,0.69579494,0.7844103,0.79425645,0.75487185,0.636718,0.5152821,0.38400003,0.30194873,0.39384618,0.5415385,0.46933338,0.380718,0.39056414,0.50543594,0.54482055,0.77128214,0.8598975,0.75487185,0.65641034,0.73517954,0.8336411,0.8369231,0.73517954,0.61374366,0.56123084,0.49887183,0.4594872,0.46933338,0.5415385,0.5481026,0.56451285,0.574359,0.5677949,0.54482055,0.6235898,0.72861546,0.8369231,0.9714873,1.2209232,1.5655385,2.1956925,2.5435898,2.3794873,1.8248206,1.4473847,1.3095386,1.1782565,1.0272821,1.0568206,1.1815386,1.0699488,0.8763078,0.7417436,0.77128214,0.6498462,0.69579494,0.8402052,0.9517949,0.8205129,0.702359,0.702359,0.77456415,0.82379496,0.7187693,0.5940513,0.5546667,0.53825647,0.512,0.45620516,0.48574364,0.47261542,0.47917953,0.5218462,0.5874872,0.6235898,0.67282057,0.7089231,0.71548724,0.69251287,0.6826667,0.5284103,0.47261542,0.52512825,0.47917953,0.47589746,0.54482055,0.51856416,0.4201026,0.45620516,0.4201026,0.43323082,0.41025645,0.33805132,0.26256412,0.33476925,0.380718,0.36102566,0.3052308,0.3052308,0.3249231,0.3446154,0.38400003,0.4660513,0.6235898,0.81394875,0.92225647,1.083077,1.270154,1.3128207,1.1257436,1.0699488,0.95835906,0.74830776,0.54482055,0.7450257,0.892718,1.0633847,1.2209232,1.211077,1.2077949,1.3128207,1.3128207,1.2307693,1.3357949,0.009846155,0.016410258,0.01969231,0.029538464,0.04594872,0.04594872,0.059076928,0.04266667,0.016410258,0.0032820515,0.009846155,0.0032820515,0.0,0.006564103,0.049230773,0.190359,0.2297436,0.15097436,0.072205134,0.032820515,0.013128206,0.013128206,0.01969231,0.032820515,0.098461546,0.28225642,0.702359,1.1651284,1.6771283,2.1300514,2.2711797,1.3850257,0.9616411,0.9747693,1.1881026,1.148718,0.86974365,0.81394875,1.3686155,2.930872,5.917539,9.596719,16.150976,22.787283,27.828514,30.70031,30.677336,31.816208,34.38277,38.41313,43.71036,45.469543,41.87898,35.669334,30.214567,29.541746,30.792208,28.45867,24.65149,21.14954,19.400208,18.62236,19.685745,22.583797,25.590157,25.255386,25.652515,27.966362,28.586668,26.482874,23.200823,23.115488,23.30913,24.795898,27.250874,28.973951,34.084106,44.11077,53.83877,59.730057,59.956516,72.29703,85.88144,83.79078,64.6958,42.886566,41.186466,44.36349,52.818054,61.124928,58.033234,42.033234,30.592003,23.995079,20.949335,18.596104,21.904411,25.787079,27.867899,27.631592,26.407387,22.324514,20.903387,21.234873,21.349745,18.212105,17.378464,15.986873,14.8020525,14.145642,13.912617,13.689437,14.227694,13.673027,11.930258,10.650257,10.039796,8.001641,6.052103,4.7655387,3.7842054,4.588308,5.579488,6.091488,6.117744,6.2785645,7.030154,8.109949,8.825437,9.176616,9.878975,11.552821,13.105232,14.434463,15.43877,16.019693,15.369847,14.480412,13.66318,13.206975,13.371078,14.979283,16.022976,17.391592,18.825848,18.921026,17.851078,16.315079,14.880821,13.37436,10.896411,8.293744,6.3507695,4.7458467,3.5380516,3.1606157,5.4383593,7.785026,10.092308,14.139078,23.591387,16.147694,13.4629755,11.648001,9.18318,6.9021544,10.282667,12.58995,13.364513,12.849232,11.995898,14.815181,30.263798,36.10585,31.113848,35.091694,38.104618,37.825645,38.47549,37.120003,23.670156,27.618464,34.63549,44.852516,57.57375,71.26318,90.397545,76.189545,51.92534,32.6039,24.917336,19.370668,18.162872,18.517334,18.553438,17.289848,19.124514,19.344412,16.482462,12.228924,11.418258,13.338258,20.673643,25.311182,23.302567,14.867694,8.4053335,13.627078,18.720821,19.830154,21.034668,30.240824,29.705849,21.910976,13.66318,16.121437,22.514874,21.504002,15.284514,7.857231,5.0543594,6.5312824,7.955693,11.700514,19.59713,32.932106,59.890877,57.98072,47.507694,39.939285,37.910976,38.36062,37.622158,29.761642,17.046976,9.957745,13.15118,16.039387,17.664001,17.913437,17.526155,17.654156,18.376207,20.394669,21.668104,17.417847,21.914259,22.905437,19.505232,14.139078,12.560411,8.94359,10.108719,12.373334,12.744206,8.897642,16.357744,23.302567,23.67672,19.90236,22.872618,27.293541,34.930874,46.05703,55.896618,54.623184,54.258877,58.381134,60.0878,56.782772,50.146465,41.951183,39.666874,44.41272,51.328003,49.57867,38.898876,36.148514,33.975796,30.536207,29.48595,27.657848,25.396515,25.252104,24.897642,17.106052,16.659693,14.257232,12.652308,11.782565,8.763078,7.430565,9.961026,8.513641,3.8531284,5.346462,5.6943593,4.8640003,4.6539493,4.857436,3.2820516,2.6486156,3.4691284,6.931693,9.659078,3.7054362,7.259898,7.3682055,4.706462,1.9265642,3.6726158,7.4010262,5.668103,4.886975,7.2369237,10.656821,9.15036,9.26195,8.3593855,6.810257,7.9917955,8.474257,4.7524104,2.6354873,3.31159,3.3378465,4.529231,4.4701543,3.698872,2.7175386,2.0217438,2.7044106,2.9604106,2.1234872,0.8992821,1.3554872,1.1027694,0.9944616,1.1257436,1.4342566,1.7165129,1.8116925,1.3226668,1.0075898,0.96492314,0.6235898,0.46933338,0.6301539,0.64000005,0.43323082,0.3446154,0.45292312,0.37743592,0.34133336,0.35446155,0.2231795,0.18379489,0.23958977,0.39384618,0.5284103,0.40369233,0.20348719,0.14769232,0.13456412,0.1148718,0.06564103,0.059076928,0.11158975,0.12471796,0.08861539,0.072205134,0.098461546,0.15097436,0.13784617,0.09189744,0.17723078,0.67938465,0.5316923,0.42338464,0.60389745,0.9124103,0.77128214,0.77456415,0.61374366,0.3446154,0.38728207,0.3249231,0.27569234,0.24615386,0.256,0.35446155,0.42338464,0.4397949,0.5218462,0.6268718,0.5481026,0.42338464,0.3446154,0.3314872,0.30851284,0.12471796,0.029538464,0.01969231,0.01969231,0.0032820515,0.0,0.11158975,0.108307704,0.08533334,0.09189744,0.101743594,0.06235898,0.03938462,0.036102567,0.049230773,0.06564103,0.08205129,0.055794876,0.01969231,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.052512825,0.059076928,0.032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.02297436,0.068923086,0.17394873,0.15753847,0.16410258,0.17723078,0.0,0.0,0.03938462,0.06564103,0.10502565,0.27569234,0.5415385,0.4660513,0.36430773,0.3314872,0.21989745,0.08205129,0.032820515,0.016410258,0.009846155,0.01969231,0.0032820515,0.0,0.0032820515,0.0032820515,0.0,0.0,0.006564103,0.006564103,0.0032820515,0.0,0.006564103,0.04266667,0.072205134,0.10502565,0.19364104,0.052512825,0.009846155,0.029538464,0.08205129,0.17066668,0.10502565,0.14441027,0.108307704,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.03938462,0.08205129,0.11158975,0.13128206,0.14441027,0.17394873,0.24615386,0.3249231,0.37743592,0.44964105,0.6695385,1.0043077,1.1946667,1.2996924,1.332513,1.2603078,1.142154,0.92553854,0.65312827,0.38400003,0.17066668,0.128,0.09189744,0.068923086,0.08205129,0.15425642,0.21661541,0.30851284,0.49230772,0.7811283,1.1158975,1.0896411,0.67938465,0.28225642,0.0951795,0.098461546,0.21333335,0.38728207,0.52512825,0.6268718,0.761436,0.8369231,0.77456415,0.702359,0.6432821,0.50543594,0.54482055,0.636718,0.702359,0.7122052,0.6826667,0.67282057,0.58420515,0.47917953,0.43323082,0.5316923,0.571077,0.49230772,0.37415388,0.28882053,0.2986667,0.3511795,0.512,0.60061544,0.58420515,0.57764107,0.69251287,0.77456415,0.81394875,0.79425645,0.69251287,0.5481026,0.46933338,0.44307697,0.46276927,0.512,0.5152821,0.46933338,0.44307697,0.4594872,0.48902568,0.58092314,0.69907695,0.8041026,0.9616411,1.3128207,1.5819489,2.0742567,2.3466668,2.2416413,1.9068719,1.5622566,1.3850257,1.3686155,1.4244103,1.3686155,1.1027694,0.90584624,0.75487185,0.69907695,0.86646163,0.8730257,0.8598975,0.9189744,0.9878975,0.8336411,0.6826667,0.69907695,0.7515898,0.7384616,0.58420515,0.49887183,0.48574364,0.48246157,0.45292312,0.4135385,0.44964105,0.4201026,0.39384618,0.39712822,0.4004103,0.41025645,0.46933338,0.5349744,0.5874872,0.6170257,0.5546667,0.4135385,0.36102566,0.4135385,0.42994875,0.4266667,0.47589746,0.508718,0.48574364,0.36758977,0.33805132,0.3314872,0.318359,0.2986667,0.29210258,0.33476925,0.3249231,0.2986667,0.27569234,0.28225642,0.30194873,0.33476925,0.41682056,0.5349744,0.6465641,0.7089231,0.7220513,0.78769237,0.892718,0.90256417,0.8598975,0.88943595,0.8041026,0.6235898,0.5546667,0.76800007,0.93866676,1.0469744,1.086359,1.0502565,1.1585642,1.3357949,1.4473847,1.4473847,1.3850257,0.009846155,0.02297436,0.02297436,0.032820515,0.04594872,0.04594872,0.059076928,0.036102567,0.009846155,0.0032820515,0.009846155,0.0032820515,0.0,0.0032820515,0.03938462,0.15753847,0.128,0.06564103,0.02297436,0.013128206,0.0,0.016410258,0.049230773,0.118153855,0.256,0.508718,0.8960001,1.2931283,1.8609232,2.5042052,2.8750772,1.9298463,1.3259488,1.2012309,1.339077,1.1913847,0.92225647,1.014154,1.6344616,2.9210258,4.9887185,9.143796,18.582975,25.961027,28.704823,29.023182,28.314259,30.057028,34.215385,40.415184,47.94749,44.580105,36.83118,29.96513,27.520002,31.304207,31.573336,28.21908,24.835283,23.23036,23.42072,21.126566,20.28308,21.195488,22.390156,20.611284,20.883694,22.898874,23.5159,22.321232,21.605745,21.241438,21.924105,24.277336,27.598772,29.88308,35.99754,47.586464,61.16103,71.51919,71.74236,79.20247,85.44165,79.08431,60.77703,43.204926,41.137234,39.696415,41.64267,45.200413,44.061543,33.923286,26.594463,22.849644,21.924105,21.507284,25.261951,27.720207,27.667694,25.77395,24.582565,20.8279,19.91877,19.840002,19.108105,16.761436,17.024002,15.694771,14.674052,14.710155,15.376411,14.729847,14.457437,13.6697445,12.268309,10.932513,9.501539,7.2960005,5.402257,4.2502565,3.620103,4.141949,4.7556925,5.139693,5.467898,6.413129,6.8594875,8.12636,9.288206,10.217027,11.588924,12.714667,13.35795,13.574565,13.5778475,13.74195,12.488206,11.628308,11.270565,11.562668,12.694975,14.227694,14.979283,16.416822,17.88718,16.626873,16.180513,15.186052,13.571283,11.552821,9.619693,8.303591,6.5411286,5.681231,6.1472826,7.4141545,11.172104,13.840411,14.614976,16.443079,26.016823,16.278976,14.106257,15.842463,16.04595,7.4765134,14.536206,24.644924,25.337439,17.381744,14.792206,17.217642,35.698875,39.282875,27.181952,28.773746,25.212719,22.912003,25.80349,29.072412,19.170464,24.887796,33.920002,40.786053,43.421543,43.17539,54.242466,41.67549,25.701746,16.059078,12.002462,12.1928215,12.754052,11.936821,9.882257,8.595693,13.098668,14.326155,11.099898,6.4722056,7.6996927,11.657847,16.866463,18.756924,16.689232,13.945437,7.2303596,10.909539,14.139078,13.564719,13.348104,20.640821,22.06195,18.277744,12.258463,9.271795,16.265848,21.083899,19.377232,14.024206,15.104001,18.58954,17.696821,17.88718,22.485334,32.68267,59.4478,61.138058,50.878365,39.460106,35.33785,33.214363,32.006565,25.225847,13.889642,6.514872,8.792616,13.764924,18.189129,19.8039,17.32595,17.345642,16.896002,18.753643,21.635284,20.20431,22.57395,26.59118,24.874668,18.41231,16.534975,11.749744,12.672001,15.133539,15.396104,10.167795,12.721231,17.526155,18.41559,15.248411,13.932309,16.89272,24.44472,38.862774,53.812515,54.36062,53.234875,54.324516,50.740517,42.837337,38.20308,34.829132,34.0119,39.538876,48.374157,50.642056,45.538464,42.207184,37.86831,33.473644,33.70339,30.263798,27.858053,29.558157,32.338055,27.090054,23.443693,16.869745,11.9860525,9.819899,7.8080006,6.166975,5.297231,4.1747694,4.2141542,9.281642,9.4916935,7.066257,5.8847184,5.98318,3.564308,3.245949,3.4264617,6.6560006,9.770667,3.889231,6.432821,7.6110773,5.7140517,2.6847181,4.135385,8.608821,5.3858466,2.993231,4.5587697,7.8112826,8.152616,10.584617,11.18195,9.032206,6.2523084,8.185436,5.146257,2.5993848,2.2678976,2.1530259,2.868513,2.8521028,2.7470772,2.4057438,0.892718,2.7995899,3.6496413,2.865231,1.4178462,1.8543591,1.6738462,1.4145643,1.529436,1.8937438,1.8412309,2.3762052,1.8445129,1.276718,1.1290257,1.2832822,0.7811283,0.60389745,0.51856416,0.4660513,0.58420515,0.6465641,0.48902568,0.33476925,0.25928208,0.18707694,0.2100513,0.2100513,0.26256412,0.3249231,0.26256412,0.1148718,0.08861539,0.101743594,0.0951795,0.06564103,0.07876924,0.13128206,0.12471796,0.068923086,0.072205134,0.10502565,0.14112821,0.13128206,0.0951795,0.128,0.4660513,0.39056414,0.34133336,0.4660513,0.6301539,0.52512825,0.45620516,0.33476925,0.22646156,0.33805132,0.35774362,0.3052308,0.23302566,0.190359,0.21333335,0.318359,0.33805132,0.3511795,0.41025645,0.53825647,0.52512825,0.38728207,0.3249231,0.36758977,0.3511795,0.13456412,0.032820515,0.013128206,0.029538464,0.029538464,0.07548718,0.049230773,0.03938462,0.059076928,0.06564103,0.04594872,0.059076928,0.049230773,0.02297436,0.049230773,0.101743594,0.08205129,0.03938462,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.009846155,0.02297436,0.01969231,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.08861539,0.16738462,0.29210258,0.33805132,0.0,0.0,0.0,0.0,0.0032820515,0.01969231,0.18707694,0.3117949,0.35774362,0.30851284,0.17066668,0.068923086,0.026256412,0.013128206,0.009846155,0.01969231,0.009846155,0.0032820515,0.0,0.0032820515,0.013128206,0.013128206,0.009846155,0.006564103,0.0,0.0,0.006564103,0.029538464,0.049230773,0.06235898,0.108307704,0.02297436,0.0,0.009846155,0.032820515,0.06564103,0.04594872,0.049230773,0.036102567,0.006564103,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.07876924,0.098461546,0.101743594,0.10502565,0.12471796,0.17394873,0.24943592,0.29538465,0.34133336,0.5152821,0.7975385,1.0404103,1.1979488,1.2471796,1.204513,1.1815386,1.0601027,0.8369231,0.5349744,0.20020515,0.14441027,0.128,0.11158975,0.108307704,0.18051283,0.23958977,0.32164106,0.48246157,0.7450257,1.0732309,1.0043077,0.8533334,0.5513847,0.20020515,0.055794876,0.13456412,0.32164106,0.48902568,0.5973334,0.6892308,0.73517954,0.7220513,0.71548724,0.7122052,0.65969235,0.60389745,0.6071795,0.6268718,0.6301539,0.5874872,0.63343596,0.61374366,0.58092314,0.57764107,0.6465641,0.6826667,0.5677949,0.4397949,0.34789747,0.26912823,0.27897438,0.380718,0.45620516,0.48574364,0.5218462,0.6662565,0.761436,0.8402052,0.8763078,0.8041026,0.574359,0.4660513,0.4397949,0.4594872,0.51856416,0.5415385,0.48246157,0.43651286,0.446359,0.50543594,0.6662565,0.72861546,0.764718,0.8763078,1.1913847,1.4867693,1.910154,2.1267693,2.0676925,1.9068719,1.7690258,1.595077,1.6114873,1.7526156,1.6410258,1.2274873,0.95835906,0.82379496,0.8172308,0.93866676,0.9485129,0.88943595,0.8795898,0.892718,0.761436,0.7089231,0.6629744,0.6432821,0.61374366,0.49887183,0.4397949,0.44307697,0.43651286,0.40369233,0.35446155,0.3446154,0.318359,0.29538465,0.28882053,0.28882053,0.2986667,0.34789747,0.39056414,0.42994875,0.50543594,0.39712822,0.29210258,0.27569234,0.34133336,0.380718,0.38728207,0.40369233,0.46933338,0.50543594,0.3117949,0.29538465,0.26912823,0.256,0.26584616,0.3052308,0.3314872,0.29210258,0.256,0.25271797,0.25928208,0.27241027,0.35774362,0.48902568,0.60061544,0.58092314,0.5513847,0.60061544,0.69579494,0.75487185,0.65312827,0.7220513,0.84348726,0.81394875,0.6662565,0.6662565,0.7811283,0.8566154,0.90584624,0.9156924,0.8533334,1.0075898,1.1881026,1.3522053,1.4178462,1.2931283,0.0,0.01969231,0.016410258,0.006564103,0.0,0.0,0.0,0.009846155,0.016410258,0.02297436,0.02297436,0.0032820515,0.0,0.0,0.02297436,0.098461546,0.03938462,0.009846155,0.0032820515,0.006564103,0.0032820515,0.01969231,0.0951795,0.22646156,0.43651286,0.761436,1.1716924,1.5491283,2.0709746,2.7241027,3.3017437,2.28759,1.7296412,1.5819489,1.5688206,1.1815386,1.0469744,1.3423591,1.9593848,2.9210258,4.3749747,8.553026,18.353231,25.24554,26.650259,25.947899,27.776003,31.730875,37.458054,44.478363,52.17149,45.75836,37.24144,30.158772,27.3559,31.015387,31.763695,29.390772,28.33395,29.653336,31.002258,26.289232,22.770874,20.873848,19.820309,17.6279,18.369642,19.584002,19.734976,18.894772,18.753643,18.159592,19.922052,23.798155,28.658875,32.49231,36.736004,44.40944,55.91303,68.178055,74.68636,69.77313,58.804516,47.60944,39.909748,37.32349,38.505028,36.545643,34.566566,33.122463,30.217848,25.51795,22.554258,21.825644,23.089233,25.399797,27.670977,26.824207,23.857233,20.548925,19.43631,17.739489,17.903591,17.503181,16.118155,15.327181,16.528412,15.734155,14.989129,15.084309,15.530668,13.99795,12.790154,11.82195,10.880001,9.6525135,7.640616,5.687795,4.128821,3.3017437,3.5249233,3.6627696,4.332308,5.1626673,6.1046157,7.433847,8.070564,9.324308,10.768411,12.097642,13.108514,13.571283,13.380924,12.71795,11.96636,11.697231,10.121847,9.350565,9.025641,9.140513,10.036513,11.122872,11.828514,13.978257,16.485744,15.363283,15.747283,14.6182575,11.792411,8.6580515,8.15918,7.640616,6.3573337,8.257642,12.47836,13.351386,15.284514,16.725334,14.76595,11.631591,14.6871805,15.78995,19.761232,25.261951,25.842875,9.944616,16.420103,34.86195,34.34667,16.200207,14.007796,13.971693,26.561644,28.386463,19.689028,24.375797,15.094155,12.511181,17.14872,23.417439,19.600412,21.786259,27.592207,29.630362,27.214771,26.371284,28.822977,24.497232,17.224207,10.138257,5.677949,8.251078,9.485129,7.9261546,5.5532312,7.752206,11.815386,13.275898,9.147078,2.7470772,3.7087183,14.500104,17.870771,17.096207,14.191591,9.941334,7.460103,11.956513,14.674052,13.289026,11.900719,12.652308,12.658873,13.617231,13.74195,7.768616,9.77395,18.192411,22.38359,22.30154,28.49149,34.29744,30.63795,24.359386,20.808207,23.840822,41.53108,51.42975,48.433235,36.60472,29.170874,29.462976,26.98831,20.844309,12.320822,4.900103,5.21518,11.152411,17.821539,21.421951,19.242668,19.27877,17.345642,18.858667,23.108925,23.250053,22.262156,29.010054,30.080002,23.699694,19.761232,16.938667,17.798565,19.600412,19.347694,13.801026,12.819694,11.989334,12.186257,13.095386,13.1872835,10.9686165,15.579899,29.994669,48.28226,55.620926,61.229954,62.821747,55.240208,42.223595,36.41436,37.284107,36.739285,41.114258,51.915493,65.80842,75.053955,68.31262,55.94257,47.01539,49.32267,43.346054,37.2119,35.25908,37.136414,37.828926,32.256004,20.696617,11.851488,8.539898,7.6603084,6.51159,5.5138464,4.1846156,4.4340515,10.5780525,10.541949,7.4174366,6.2588725,6.701949,2.9505644,5.425231,5.7009234,7.834257,10.069334,4.844308,3.6594875,5.786257,6.0717955,4.2436924,4.893539,8.234667,5.691077,3.114667,3.0424619,4.663795,6.409847,9.065026,11.638155,11.54954,4.640821,5.3727183,4.4373336,3.3050258,2.4188719,1.1618463,2.1792822,2.3171284,2.034872,1.5064616,0.63343596,2.5862565,3.5938463,3.2886157,2.409026,2.802872,2.2219489,1.9823592,2.5665643,3.2131286,1.9364104,2.4582565,2.428718,2.0742567,1.8182565,2.2646155,1.5655385,1.1093334,0.8041026,0.702359,0.98461545,0.77128214,0.508718,0.33476925,0.26256412,0.21989745,0.29538465,0.3117949,0.30194873,0.28225642,0.25271797,0.072205134,0.01969231,0.029538464,0.049230773,0.04266667,0.07876924,0.12143591,0.118153855,0.08205129,0.08533334,0.108307704,0.118153855,0.118153855,0.1148718,0.1148718,0.28225642,0.28225642,0.3117949,0.40697438,0.41682056,0.24615386,0.15097436,0.15097436,0.24287182,0.39056414,0.45620516,0.4004103,0.3117949,0.2231795,0.118153855,0.22646156,0.3708718,0.4004103,0.38400003,0.5940513,0.62030774,0.4004103,0.256,0.32164106,0.56451285,0.27241027,0.08533334,0.029538464,0.068923086,0.108307704,0.12471796,0.06235898,0.01969231,0.026256412,0.03938462,0.029538464,0.08205129,0.07548718,0.016410258,0.026256412,0.07548718,0.072205134,0.04594872,0.01969231,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.0032820515,0.016410258,0.016410258,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.118153855,0.3052308,0.39384618,0.08205129,0.03938462,0.009846155,0.013128206,0.029538464,0.02297436,0.036102567,0.17066668,0.19692309,0.11158975,0.12143591,0.08533334,0.03938462,0.009846155,0.0,0.0,0.009846155,0.0032820515,0.0,0.006564103,0.026256412,0.026256412,0.009846155,0.0,0.0,0.0,0.0032820515,0.0,0.0032820515,0.013128206,0.013128206,0.0032820515,0.0032820515,0.009846155,0.029538464,0.055794876,0.20020515,0.13784617,0.049230773,0.01969231,0.03938462,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07876924,0.0951795,0.08861539,0.08861539,0.098461546,0.118153855,0.15753847,0.19692309,0.25271797,0.36430773,0.47917953,0.67938465,0.955077,1.2077949,1.2537436,1.270154,1.1815386,1.0043077,0.7318975,0.3708718,0.2100513,0.17394873,0.15753847,0.14112821,0.17394873,0.23302566,0.31507695,0.47589746,0.73517954,1.0929232,1.0305642,1.0469744,0.8369231,0.40697438,0.06564103,0.0951795,0.2100513,0.3446154,0.46276927,0.5481026,0.64000005,0.702359,0.69907695,0.6662565,0.7253334,0.6859488,0.636718,0.5973334,0.57764107,0.5513847,0.5677949,0.60061544,0.6432821,0.67938465,0.702359,0.827077,0.6662565,0.5284103,0.48902568,0.39056414,0.318359,0.4201026,0.5152821,0.5415385,0.54482055,0.6498462,0.764718,0.86646163,0.9353847,0.95835906,0.7515898,0.60061544,0.50543594,0.47589746,0.5284103,0.56123084,0.53825647,0.512,0.5152821,0.58092314,0.81066674,0.79097444,0.74830776,0.81066674,1.0043077,1.3128207,1.7165129,1.9659488,1.9922053,1.9364104,1.9068719,1.723077,1.6475899,1.7066668,1.6672822,1.463795,1.2504616,1.1126155,1.0469744,0.955077,0.88287187,0.8041026,0.76800007,0.75487185,0.67938465,0.74830776,0.6071795,0.512,0.5218462,0.49887183,0.446359,0.41025645,0.380718,0.34133336,0.2855385,0.23302566,0.22646156,0.2231795,0.21989745,0.26256412,0.28882053,0.3249231,0.32164106,0.30194873,0.3708718,0.27569234,0.21989745,0.25271797,0.33476925,0.34789747,0.3446154,0.3511795,0.39712822,0.4266667,0.30851284,0.29210258,0.27897438,0.26584616,0.26584616,0.28225642,0.3117949,0.29538465,0.26584616,0.24615386,0.2231795,0.24615386,0.4004103,0.5677949,0.6268718,0.4660513,0.44964105,0.5907693,0.761436,0.81066674,0.58092314,0.6465641,0.8467693,0.94523084,0.8960001,0.8467693,0.8041026,0.7089231,0.7056411,0.79097444,0.78769237,0.8960001,0.9911796,1.0765129,1.1388719,1.1684103,0.0,0.049230773,0.02297436,0.0,0.0,0.0,0.0,0.009846155,0.052512825,0.108307704,0.108307704,0.02297436,0.0,0.006564103,0.013128206,0.0,0.0,0.0,0.013128206,0.026256412,0.016410258,0.0032820515,0.06564103,0.18707694,0.41025645,0.82379496,1.3489232,1.8379488,2.2514873,2.5337439,2.5928206,1.7624617,1.719795,2.038154,2.2547693,1.8773335,1.8412309,1.7591796,1.6475899,2.03159,3.9351797,8.123077,18.087385,24.247797,24.654772,25.009233,29.794464,36.10913,41.363697,45.728825,52.12554,46.752823,38.61662,31.7079,28.596516,30.441029,31.504414,30.71672,32.9879,37.789543,39.168003,30.63795,25.993849,23.93272,22.728207,20.263386,20.65395,20.624413,19.324718,17.335796,16.679386,16.640001,18.645334,22.642874,27.864618,32.820515,36.31262,42.164516,51.83016,64.99447,79.60616,68.864006,51.347694,38.78072,34.661747,34.271183,33.14872,29.581131,27.444515,27.690668,28.35036,23.834259,22.163694,21.999592,22.629745,23.972105,23.653746,20.965746,18.665028,18.497643,21.195488,18.619078,18.021746,17.972515,17.841232,17.792002,15.753847,15.471591,15.980309,16.311796,15.51754,13.810873,12.750771,11.877745,10.482873,7.6143594,6.294975,5.0871797,4.378257,3.9647183,3.0358977,2.9013336,3.4002054,4.4734364,5.9569235,7.568411,9.193027,10.450052,11.23118,11.385437,10.725744,10.262975,9.340718,8.083693,6.6428723,5.2053337,5.7764106,7.768616,8.805744,8.891078,10.390975,13.088821,13.29559,12.931283,12.898462,13.092104,11.98277,9.53436,6.7216415,4.59159,4.2896414,5.412103,5.976616,12.297847,20.148514,14.7561035,9.921641,11.378873,11.999181,11.136001,14.601848,22.403284,31.566772,31.77354,22.688822,13.961847,13.033027,30.37867,28.895182,9.370257,10.466462,10.725744,19.99754,21.687796,15.330462,16.587488,10.509129,9.83959,14.8250265,19.662771,12.498053,15.75713,21.451488,23.555285,21.559797,20.46359,28.921438,26.22031,17.558975,8.316719,4.0434875,9.147078,9.55077,6.8496413,7.240206,21.543386,20.14195,21.392412,14.70359,2.7175386,1.3292309,16.951796,18.743795,17.394873,15.192616,6.012718,8.684308,13.154463,16.955078,18.018463,14.647796,19.091694,17.161848,16.899282,18.15631,12.603078,10.906258,10.043077,13.2562065,18.983387,20.873848,18.215385,14.739694,12.199386,11.437949,12.389745,28.235489,43.201645,46.21457,36.04349,21.287386,18.100513,17.02072,17.112617,16.059078,10.161232,4.9493337,6.9710774,14.339283,22.439386,23.939283,29.06585,25.38667,22.183386,23.141745,26.351591,21.458054,26.79795,30.086567,28.317541,27.75631,30.733131,30.194874,29.141336,26.7159,18.218668,13.078976,11.933539,12.950975,14.578873,15.51754,13.699283,15.360002,22.068514,33.992207,49.89703,69.645134,70.8398,60.65888,46.887386,37.90113,34.008617,34.527184,49.06011,78.72329,116.16165,141.53847,124.53088,95.26811,73.85929,70.35734,60.724518,51.570877,43.54954,37.097027,32.41026,25.928207,17.450668,11.424822,8.979693,7.90318,6.6592827,7.2631803,5.687795,2.8389745,4.5489235,9.258667,7.8080006,5.2644105,3.9154875,3.2820516,6.672411,7.706257,9.701744,11.250873,6.2096415,4.4406157,8.63836,9.317744,5.293949,3.7087183,7.3321033,7.269744,5.802667,4.161641,2.5042052,4.9821544,5.681231,6.806975,7.706257,4.896821,2.993231,2.809436,2.9440002,2.3958976,0.56451285,1.1979488,2.4746668,3.255795,2.7831798,0.67282057,0.7089231,1.339077,2.3762052,3.4231799,3.876103,1.7033848,2.0939488,4.322462,5.8518977,2.349949,2.3368206,3.2853336,4.4701543,4.850872,3.0818465,2.9111798,3.0687182,2.5009232,1.3259488,0.8402052,0.5940513,0.52512825,0.446359,0.318359,0.24287182,0.37743592,0.40369233,0.40369233,0.42338464,0.47261542,0.108307704,0.016410258,0.059076928,0.1148718,0.09189744,0.07876924,0.13128206,0.13784617,0.08533334,0.06235898,0.072205134,0.0951795,0.12471796,0.16410258,0.21333335,0.16410258,0.16082053,0.19692309,0.24615386,0.25928208,0.18707694,0.15097436,0.17394873,0.28225642,0.48902568,0.47589746,0.28882053,0.23630771,0.3249231,0.28882053,0.28882053,0.4004103,0.5284103,0.6301539,0.7187693,0.75487185,0.54482055,0.2986667,0.18707694,0.32164106,0.2231795,0.108307704,0.026256412,0.04594872,0.2297436,0.18051283,0.08533334,0.01969231,0.0032820515,0.016410258,0.016410258,0.02297436,0.02297436,0.016410258,0.016410258,0.016410258,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.009846155,0.0,0.0,0.0,0.0,0.006564103,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13456412,0.3511795,0.4135385,0.19364104,0.055794876,0.06235898,0.14441027,0.108307704,0.032820515,0.04266667,0.06235898,0.08533334,0.18379489,0.14769232,0.06564103,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.016410258,0.006564103,0.0,0.0,0.0,0.013128206,0.006564103,0.0,0.0,0.0,0.0,0.009846155,0.026256412,0.06564103,0.15097436,0.88615394,0.636718,0.21661541,0.026256412,0.07548718,0.016410258,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.055794876,0.07876924,0.06235898,0.06235898,0.12143591,0.15425642,0.16082053,0.16738462,0.2297436,0.31507695,0.46276927,0.69579494,0.9485129,1.083077,1.2537436,1.1782565,1.0371283,0.90584624,0.74830776,0.39384618,0.20348719,0.108307704,0.06564103,0.07548718,0.12471796,0.21989745,0.38400003,0.5907693,0.761436,0.78769237,0.81066674,0.79425645,0.6301539,0.15097436,0.09189744,0.15097436,0.31507695,0.47589746,0.4266667,0.5874872,0.7187693,0.69907695,0.60389745,0.702359,0.702359,0.636718,0.571077,0.5415385,0.56451285,0.5415385,0.54482055,0.60389745,0.6892308,0.702359,0.6892308,0.60389745,0.5481026,0.5481026,0.5481026,0.39056414,0.39712822,0.5316923,0.6892308,0.702359,0.60389745,0.6892308,0.83035904,0.9944616,1.2504616,1.2504616,1.0404103,0.7844103,0.60061544,0.56451285,0.5874872,0.5874872,0.5677949,0.5546667,0.58092314,0.71548724,0.7581539,0.8369231,0.9911796,1.1749744,1.1979488,1.3161026,1.5458462,1.8379488,2.044718,1.7624617,1.4276924,1.2012309,1.1520001,1.2504616,1.1651284,1.2077949,1.2077949,1.1257436,1.0535386,1.1257436,0.9616411,0.75487185,0.6301539,0.65641034,0.7056411,0.5874872,0.5021539,0.508718,0.5349744,0.47261542,0.4201026,0.38400003,0.34789747,0.27569234,0.24943592,0.24287182,0.21989745,0.17723078,0.15097436,0.190359,0.27241027,0.29538465,0.26256412,0.27569234,0.22646156,0.23958977,0.30851284,0.38400003,0.39712822,0.38400003,0.380718,0.35774362,0.30851284,0.25928208,0.28225642,0.3446154,0.380718,0.380718,0.380718,0.3314872,0.33805132,0.3708718,0.3708718,0.25928208,0.3314872,0.54482055,0.71548724,0.73517954,0.56451285,0.47917953,0.4955898,0.5316923,0.51856416,0.39712822,0.48246157,0.6859488,0.88943595,1.017436,1.0535386,0.9419488,0.7778462,0.7220513,0.8008206,0.88615394,0.98133343,1.024,1.0075898,0.99774367,1.1454359,0.013128206,0.20676924,0.108307704,0.013128206,0.013128206,0.013128206,0.0032820515,0.009846155,0.032820515,0.059076928,0.068923086,0.013128206,0.006564103,0.009846155,0.0032820515,0.013128206,0.098461546,0.049230773,0.006564103,0.02297436,0.03938462,0.016410258,0.026256412,0.07876924,0.26912823,0.761436,1.591795,2.294154,2.737231,2.8816411,2.7766156,2.2383592,2.2350771,2.4648206,2.8422565,3.4888208,3.948308,3.2525132,2.5173335,2.5271797,3.7284105,8.119796,13.193847,16.633438,18.865232,23.056412,29.88308,34.18585,37.51713,41.554054,48.095184,45.95857,40.23467,33.027283,27.398565,27.365746,26.308926,25.488413,28.360207,32.76144,30.916925,23.995079,21.31036,20.795078,20.900105,20.581745,20.289642,18.681437,16.695797,15.172924,14.834873,16.22318,19.062155,22.767591,26.660105,29.96513,32.879593,35.183594,39.686565,47.524105,58.17108,57.57375,49.35549,39.282875,31.799797,30.01108,27.85477,26.7159,26.624002,26.049643,21.907694,19.557745,19.856411,21.832207,24.267488,25.718155,23.778463,21.865026,20.279797,19.173744,18.520617,16.482462,16.305231,16.90913,17.539284,17.742771,19.111385,18.796309,18.248207,18.267899,18.996513,17.736206,14.257232,10.971898,8.723693,6.7840004,5.435077,4.352,3.8531284,3.7415388,3.2918978,3.4921029,4.1452312,5.297231,6.885744,8.753231,9.908514,9.435898,8.260923,6.9710774,5.832206,4.841026,4.0008206,3.5347695,3.4297438,3.446154,3.95159,5.3858466,7.2861543,9.31118,11.234463,10.962052,11.116308,11.444513,11.234463,9.321027,8.786052,8.641642,8.996103,9.278359,8.231385,10.144821,14.683899,21.796104,24.152617,7.174565,5.0477953,8.342975,15.829334,23.968822,26.919386,21.526976,27.943386,32.76472,27.966362,10.8996935,13.193847,30.119387,27.001438,6.38359,8.0377445,9.770667,15.845745,18.294155,15.783386,13.633642,10.541949,9.419488,12.901745,16.804104,10.115283,9.724719,12.937847,16.508718,17.979078,15.688207,18.855387,17.234053,12.386462,7.0498466,5.142975,7.9294367,7.7423596,8.2215395,11.638155,18.884924,17.306257,20.847591,16.800821,6.5345645,5.5138464,19.14749,21.809233,19.600412,15.16636,7.6964107,11.237744,11.98277,11.904001,12.071385,12.645744,27.90072,20.319181,16.823795,22.104616,18.62236,13.830565,12.22236,11.592206,10.807796,9.777231,7.030154,6.5345645,8.185436,11.273847,14.503386,28.46195,35.413338,38.383595,37.156105,28.255182,13.633642,10.889847,16.820515,23.962257,20.585028,8.060719,4.9920006,9.094564,16.918976,23.880207,35.968002,33.700104,28.035284,25.301334,27.19508,22.974361,24.379078,25.898668,26.850464,31.40595,34.628925,32.01313,31.153233,32.797543,30.851284,23.174566,19.495386,17.076513,15.025232,14.28677,13.003489,17.772308,25.48513,34.195694,43.109745,52.04021,50.008617,43.900723,38.649437,37.24472,38.232616,45.771492,57.75754,78.50339,118.75119,137.52124,120.55632,96.50544,79.66524,69.979904,61.774773,54.47549,45.059284,34.051285,25.524515,18.7799,14.621539,12.514462,11.37559,9.586872,8.500513,7.1647186,5.904411,4.9460516,4.4373336,8.083693,6.764308,4.821334,3.764513,2.281026,5.146257,5.605744,6.114462,6.695385,4.965744,8.838565,16.01641,17.027283,10.9915905,5.6352825,7.4830775,6.7577443,5.832206,4.969026,2.294154,3.8071797,4.670359,5.3037953,5.32677,3.5544617,2.1792822,3.3444104,8.28718,13.10195,8.743385,2.484513,2.7602053,5.362872,6.4295387,2.4549747,0.86974365,0.8598975,3.5183592,9.216001,17.608206,9.088,4.384821,3.3017437,3.8465643,2.228513,1.3456411,2.553436,4.2502565,5.0609236,3.8400004,2.740513,2.3236926,2.428718,2.6387694,2.2678976,1.5753847,0.79097444,0.45620516,0.53825647,0.4266667,0.39712822,0.39384618,0.3446154,0.26256412,0.25271797,0.08205129,0.026256412,0.03938462,0.07548718,0.07876924,0.14441027,0.2297436,0.27241027,0.22646156,0.08533334,0.068923086,0.059076928,0.12143591,0.2231795,0.26256412,0.29210258,0.26584616,0.21661541,0.17066668,0.11158975,0.08861539,0.07876924,0.08205129,0.13128206,0.28225642,0.32820517,0.27897438,0.22646156,0.190359,0.14441027,0.14441027,0.25928208,0.40369233,0.44964105,0.23958977,0.38400003,0.44964105,0.33476925,0.12143591,0.101743594,0.16082053,0.21333335,0.16082053,0.03938462,0.04594872,0.06564103,0.118153855,0.12471796,0.08205129,0.06564103,0.016410258,0.0032820515,0.0032820515,0.0032820515,0.0032820515,0.0032820515,0.0,0.0032820515,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.0032820515,0.0,0.006564103,0.013128206,0.0,0.0,0.052512825,0.20348719,0.35446155,0.256,0.108307704,0.029538464,0.0032820515,0.0,0.0,0.0,0.0,0.006564103,0.013128206,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.026256412,0.108307704,0.27897438,0.23302566,0.08861539,0.06235898,0.18051283,0.28882053,0.20676924,0.20020515,0.16410258,0.118153855,0.20676924,0.21989745,0.23630771,0.18379489,0.068923086,0.0,0.029538464,0.029538464,0.013128206,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.006564103,0.0032820515,0.013128206,0.013128206,0.006564103,0.006564103,0.013128206,0.029538464,0.20676924,0.3249231,0.2297436,0.016410258,0.016410258,0.0032820515,0.0,0.0,0.0032820515,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03938462,0.068923086,0.068923086,0.049230773,0.072205134,0.0951795,0.10502565,0.11158975,0.14441027,0.190359,0.30851284,0.4955898,0.71548724,0.88943595,1.0601027,1.086359,1.0272821,0.9419488,0.88287187,0.6465641,0.37415388,0.190359,0.11158975,0.07548718,0.10502565,0.18707694,0.2986667,0.42338464,0.5546667,0.84348726,0.97805136,0.8566154,0.54482055,0.27569234,0.1148718,0.11158975,0.21333335,0.34789747,0.4135385,0.52512825,0.6498462,0.6465641,0.5513847,0.5907693,0.65969235,0.71548724,0.6892308,0.6301539,0.7220513,0.72861546,0.62030774,0.56451285,0.60061544,0.65312827,0.65969235,0.69579494,0.8336411,0.9944616,0.97805136,0.5940513,0.47589746,0.54482055,0.636718,0.5316923,0.56123084,0.62030774,0.75487185,0.93866676,1.0666667,1.0568206,0.97805136,0.8763078,0.7811283,0.6859488,0.6235898,0.5973334,0.58092314,0.5513847,0.51856416,0.50543594,0.512,0.6071795,0.81066674,1.1027694,1.017436,1.0502565,1.1749744,1.4211283,1.8740515,1.8281027,1.5130258,1.1815386,1.0404103,1.276718,1.2012309,1.1585642,1.1520001,1.1618463,1.1388719,1.1323078,1.0666667,0.86317956,0.61374366,0.571077,0.5907693,0.5316923,0.4955898,0.48902568,0.43651286,0.42338464,0.4135385,0.36758977,0.28882053,0.22646156,0.20020515,0.2100513,0.21333335,0.21989745,0.26256412,0.318359,0.3249231,0.28225642,0.21989745,0.20020515,0.17066668,0.21333335,0.29210258,0.36430773,0.39712822,0.37415388,0.3249231,0.2855385,0.27569234,0.29538465,0.30194873,0.32820517,0.37743592,0.42994875,0.42994875,0.3314872,0.3117949,0.3314872,0.3511795,0.32164106,0.39384618,0.48574364,0.512,0.48246157,0.5152821,0.5284103,0.5316923,0.54482055,0.56123084,0.5677949,0.47589746,0.6301539,0.80738467,0.892718,0.86974365,0.7778462,0.7515898,0.764718,0.81066674,0.88615394,0.8960001,0.98133343,1.0075898,0.94523084,0.88943595,0.006564103,0.098461546,0.06235898,0.016410258,0.006564103,0.016410258,0.009846155,0.02297436,0.036102567,0.04594872,0.07876924,0.12471796,0.08533334,0.029538464,0.009846155,0.04266667,0.101743594,0.04594872,0.0032820515,0.009846155,0.01969231,0.009846155,0.006564103,0.03938462,0.19364104,0.6104616,1.4769232,2.2908719,2.8750772,3.05559,2.6683078,2.2022567,2.1956925,2.3630772,2.8717952,4.338872,5.028103,5.146257,4.457026,3.5807183,3.9975388,7.532308,11.385437,15.261539,19.429745,24.720411,31.002258,33.1159,35.311592,40.037746,47.95077,51.14421,42.95221,31.786669,23.660309,22.193232,21.293951,21.044514,22.393438,23.732515,20.90995,18.241642,18.231796,18.379488,18.116924,18.819284,18.28431,16.646564,15.382976,14.92677,14.683899,16.292105,19.203283,22.46236,25.284925,27.073643,27.785849,28.786875,31.058054,34.691284,38.869335,39.67344,37.175797,33.014156,29.233232,28.278156,27.316515,26.532104,26.12513,25.124104,21.366156,20.260103,20.949335,22.482054,23.545437,22.482054,20.696617,19.662771,18.500925,17.152,16.387283,15.537232,15.642258,15.652103,15.363283,15.40595,16.551386,16.787693,17.529438,19.094976,20.719591,16.699078,12.603078,9.360411,7.276308,6.0258465,5.3825645,4.3716927,3.4560003,2.8455386,2.487795,3.170462,3.6135387,4.2305646,5.097026,5.937231,6.0816417,5.5696416,4.7983594,4.2207184,4.325744,3.82359,4.266667,4.2469745,3.7218463,4.0041027,4.397949,7.0892315,9.281642,10.174359,10.985026,10.443488,10.28595,10.20718,9.724719,8.211693,16.873028,16.548103,15.497848,17.35877,21.126566,18.418873,22.777437,26.115284,22.321232,7.2664623,7.506052,12.097642,18.22195,25.557335,36.28636,27.910566,36.00739,44.32739,39.73908,12.245335,12.540719,27.526566,24.641644,5.6254363,6.5345645,9.242257,11.444513,12.416001,12.1928215,11.585642,9.9282055,8.260923,8.868103,10.164514,6.701949,5.586052,7.1581545,10.561642,13.922462,14.329437,12.219078,10.473026,8.763078,7.39118,7.2664623,7.131898,5.970052,7.7423596,12.530872,16.52513,19.06872,22.078362,19.456001,11.769437,6.2490263,15.993437,21.014977,19.96472,14.299898,8.274052,10.026668,10.305642,10.509129,11.897437,15.596309,34.212105,26.128412,22.324514,28.199387,23.578259,16.07877,13.174155,11.9860525,10.834052,9.238976,4.027077,3.3444104,5.280821,9.019077,14.828309,31.03508,38.839798,44.04185,46.257233,38.925133,18.816002,10.492719,13.732103,22.885746,26.883284,15.560206,10.5780525,9.83959,13.4629755,23.7719,34.002052,30.825027,25.606565,24.523489,28.576822,25.051899,24.86154,25.967592,27.858053,31.540516,34.904617,35.810463,38.324516,41.120823,37.490875,30.592003,24.933746,20.94277,18.930874,19.104822,20.292925,26.86031,33.6279,38.258873,41.265232,39.62749,34.067696,30.82831,32.712208,39.102364,48.08534,51.46913,50.678158,55.988518,86.49847,97.109344,89.885544,82.4517,77.512215,62.85457,60.18298,56.32657,46.247387,31.317335,19.298464,16.193642,15.097437,15.442053,15.734155,13.571283,9.964309,7.568411,9.012513,11.365745,6.121026,8.418462,5.4449234,3.7743592,4.3060517,2.2580514,12.806565,11.881026,7.499488,4.2141542,3.1081028,9.931488,16.472616,15.425642,8.690872,7.4010262,6.688821,6.180103,6.918565,7.325539,3.2229745,2.8750772,3.6069746,6.0980515,7.709539,2.5042052,1.6935385,2.9013336,10.95877,20.486567,15.894976,5.179077,2.8389745,6.1341543,9.304616,3.5478978,1.5163078,0.8795898,2.7766156,9.511385,24.576002,22.377028,12.911591,5.8289237,4.0041027,3.5249233,2.1267693,2.7798977,4.604718,6.0324106,4.8147697,2.7175386,2.477949,3.2886157,3.8432825,2.359795,1.3193847,0.92553854,0.6432821,0.32820517,0.23630771,0.21333335,0.2100513,0.17723078,0.118153855,0.1148718,0.052512825,0.01969231,0.016410258,0.04594872,0.0951795,0.128,0.24287182,0.34133336,0.33476925,0.16410258,0.11158975,0.098461546,0.15425642,0.256,0.32820517,0.38728207,0.30851284,0.21661541,0.15097436,0.08533334,0.08205129,0.06235898,0.06564103,0.13128206,0.30194873,0.43651286,0.40369233,0.27897438,0.14441027,0.08861539,0.118153855,0.17723078,0.25928208,0.28225642,0.11158975,0.16738462,0.3249231,0.32164106,0.14112821,0.036102567,0.068923086,0.16082053,0.16410258,0.06564103,0.0,0.013128206,0.17066668,0.508718,0.7975385,0.56123084,0.25928208,0.07876924,0.009846155,0.006564103,0.0,0.0,0.0,0.006564103,0.016410258,0.026256412,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.0032820515,0.0,0.0032820515,0.0032820515,0.0,0.0,0.026256412,0.14441027,0.28225642,0.21989745,0.190359,0.128,0.068923086,0.032820515,0.01969231,0.055794876,0.026256412,0.0032820515,0.006564103,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01969231,0.098461546,0.16410258,0.072205134,0.049230773,0.128,0.13456412,0.27569234,0.51856416,0.5874872,0.4201026,0.16738462,0.20020515,0.34789747,0.36102566,0.20020515,0.055794876,0.055794876,0.072205134,0.059076928,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.009846155,0.0,0.006564103,0.006564103,0.006564103,0.02297436,0.04266667,0.036102567,0.029538464,0.1148718,0.1148718,0.029538464,0.01969231,0.0032820515,0.0,0.0,0.0,0.006564103,0.009846155,0.009846155,0.016410258,0.02297436,0.0,0.0,0.0,0.0,0.006564103,0.036102567,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.04266667,0.06235898,0.036102567,0.032820515,0.04594872,0.055794876,0.059076928,0.07548718,0.098461546,0.18707694,0.35446155,0.55794877,0.7122052,0.80738467,0.9124103,0.9714873,0.9616411,0.88943595,0.7187693,0.47917953,0.27241027,0.14112821,0.07548718,0.072205134,0.11158975,0.17723078,0.27569234,0.4201026,0.761436,1.2635899,1.3718976,1.0043077,0.58092314,0.21989745,0.098461546,0.1148718,0.190359,0.26584616,0.47261542,0.6432821,0.6235898,0.47589746,0.46276927,0.512,0.6170257,0.6859488,0.69907695,0.69907695,0.7122052,0.6826667,0.67610264,0.7089231,0.7417436,0.761436,0.7811283,0.85005134,0.955077,1.0108719,0.61374366,0.45292312,0.5218462,0.6662565,0.5513847,0.6859488,0.73517954,0.83035904,1.0075898,1.2242053,1.0666667,1.079795,1.1027694,1.0633847,0.98133343,0.78769237,0.6465641,0.5677949,0.5284103,0.4955898,0.4594872,0.44964105,0.49230772,0.6071795,0.80738467,0.82379496,0.88615394,1.0010257,1.1979488,1.5195899,1.5688206,1.4998976,1.2635899,1.0305642,1.1815386,1.0994873,1.0404103,1.086359,1.2077949,1.270154,1.0699488,0.9616411,0.86646163,0.761436,0.67610264,0.6465641,0.53825647,0.46276927,0.446359,0.42994875,0.42994875,0.39712822,0.3314872,0.256,0.2231795,0.20676924,0.19692309,0.2100513,0.24287182,0.28225642,0.3117949,0.3314872,0.3117949,0.256,0.20020515,0.21333335,0.26584616,0.3314872,0.37743592,0.3708718,0.3314872,0.26584616,0.2231795,0.21989745,0.24943592,0.26584616,0.29210258,0.33476925,0.37743592,0.37743592,0.2986667,0.28882053,0.31507695,0.3446154,0.36430773,0.42338464,0.44964105,0.43323082,0.41025645,0.45620516,0.5152821,0.5284103,0.5284103,0.56451285,0.67282057,0.636718,0.67938465,0.73517954,0.7778462,0.81394875,0.67938465,0.65969235,0.7187693,0.8336411,0.9944616,0.92553854,0.88615394,0.84348726,0.7811283,0.71548724,0.0,0.0,0.009846155,0.013128206,0.016410258,0.052512825,0.17066668,0.18379489,0.118153855,0.04266667,0.06235898,0.13128206,0.08861539,0.026256412,0.006564103,0.036102567,0.052512825,0.02297436,0.0032820515,0.0032820515,0.0,0.0,0.0,0.01969231,0.1148718,0.3708718,1.0010257,1.8674873,2.7011285,3.0752823,2.4057438,1.8838975,1.7755898,1.9954873,2.7208207,4.4077954,5.0674877,5.7698464,5.293949,4.2896414,5.297231,7.3091288,9.865847,13.686155,18.986668,25.488413,29.856823,29.75508,32.141132,39.96226,52.141953,57.49498,46.11939,30.887386,20.161642,17.792002,17.952822,18.340103,18.248207,17.194668,14.900514,15.176207,15.816206,15.849027,15.760411,17.506462,16.873028,15.868719,15.471591,15.606155,15.14995,16.774565,18.983387,21.16595,22.78072,23.35508,23.223797,24.595694,26.387693,27.569233,27.16554,27.214771,27.457644,27.82195,28.114054,27.989336,27.69395,25.659079,23.673437,22.232616,20.565334,20.834463,21.943796,22.767591,22.528002,20.804924,20.099283,18.891489,17.545847,16.836924,17.93641,17.329231,16.804104,16.009848,15.209026,15.29436,16.019693,17.430975,21.014977,24.769644,23.19754,16.042667,11.723488,8.746667,6.413129,4.824616,4.4832826,3.6758976,2.789744,2.1956925,2.2416413,2.6683078,2.8947694,3.2656412,3.5380516,2.8914874,2.7273848,2.5862565,2.4943593,2.917744,4.7524104,4.1189747,5.1364107,5.7403083,5.4449234,5.32677,5.868308,8.4512825,10.118565,10.292514,10.791386,9.6065645,9.117539,8.887795,9.993847,15.035078,31.583181,29.571285,25.494976,25.580309,25.790361,18.136618,19.373951,20.768822,17.145437,6.875898,10.811078,19.712002,27.083488,33.345642,45.863388,35.13108,38.14072,42.96862,37.766567,10.765129,9.521232,18.983387,17.476925,5.356308,5.0215387,7.722667,8.395488,8.356103,8.717129,10.371283,8.749949,6.442667,4.9920006,4.4898467,3.5511796,3.0752823,4.027077,6.4032826,9.527796,12.028719,9.330873,7.456821,6.76759,6.918565,6.8562055,5.76,4.2994876,5.8781543,10.341744,13.98154,16.725334,19.40677,19.446156,15.225437,6.091488,11.85477,17.64759,17.77559,12.49477,7.9983597,9.521232,9.508103,10.686359,13.699283,17.112617,28.560413,24.484104,24.339695,29.413746,22.816822,15.133539,11.053949,9.856001,10.033232,9.281642,3.6463592,2.986667,3.7874875,5.4514875,10.325335,23.46995,35.08185,46.63139,53.549953,45.236515,22.92513,11.158976,9.55077,14.818462,20.775387,16.843489,15.61272,12.087796,9.078155,17.207796,26.499285,24.07713,20.345438,20.785233,25.941336,23.968822,24.12636,26.210464,29.144617,30.98585,33.2439,35.51836,38.85949,41.396515,38.334362,31.957336,25.078156,20.345438,19.016207,20.965746,24.274054,28.99036,33.398155,36.4078,37.599182,30.680618,24.336412,22.042257,24.690874,30.601849,38.501747,37.7239,35.183594,38.44267,55.70954,58.49272,60.770466,68.020515,72.56616,53.57621,53.395695,51.876106,42.37457,26.482874,14.020925,16.708925,16.354464,16.246155,18.054565,21.799387,13.249642,9.347282,10.820924,13.702565,9.314463,7.830975,4.164923,2.9997952,4.092718,2.2580514,13.896206,12.343796,7.6143594,4.4996924,2.550154,7.125334,11.168821,10.075898,6.4000006,9.842873,9.412924,6.5083084,6.7610264,8.933744,4.926359,3.1081028,4.2601027,7.0367184,8.1755905,2.5107694,2.3663592,2.2482052,7.972103,16.502155,15.970463,6.298257,2.6518977,4.824616,8.316719,4.325744,2.7831798,2.28759,2.733949,6.75118,19.712002,23.538874,14.641232,6.1013336,3.4166157,4.4767184,3.0720003,3.5446157,6.1472826,8.454565,5.3760004,2.7306669,3.2131286,4.4045134,4.7228723,3.4330258,1.4309745,0.9288206,0.636718,0.17723078,0.0951795,0.18051283,0.16410258,0.108307704,0.06564103,0.06564103,0.04266667,0.01969231,0.006564103,0.02297436,0.07548718,0.08205129,0.22646156,0.38400003,0.44307697,0.3052308,0.24287182,0.18707694,0.2231795,0.3249231,0.37743592,0.40369233,0.35774362,0.25928208,0.15097436,0.108307704,0.1148718,0.08861539,0.08205129,0.14441027,0.31507695,0.64000005,0.61374366,0.446359,0.26584616,0.13128206,0.13128206,0.15425642,0.19364104,0.21661541,0.16738462,0.0951795,0.23630771,0.34133336,0.28225642,0.08533334,0.049230773,0.101743594,0.14769232,0.128,0.013128206,0.0032820515,0.128,0.5316923,1.0108719,1.020718,0.86317956,0.4266667,0.12143591,0.049230773,0.006564103,0.0,0.0,0.0032820515,0.016410258,0.03938462,0.026256412,0.009846155,0.0,0.0,0.006564103,0.006564103,0.0032820515,0.0,0.0,0.006564103,0.0,0.0,0.0,0.0032820515,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.04594872,0.1148718,0.108307704,0.15425642,0.16082053,0.14441027,0.1148718,0.08533334,0.14769232,0.13456412,0.072205134,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0951795,0.0951795,0.098461546,0.108307704,0.049230773,0.190359,0.4594872,0.62030774,0.52512825,0.118153855,0.13456412,0.34133336,0.6301539,0.77128214,0.38400003,0.13456412,0.08533334,0.06235898,0.013128206,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0,0.01969231,0.026256412,0.009846155,0.0,0.0,0.036102567,0.08533334,0.11158975,0.055794876,0.02297436,0.04594872,0.068923086,0.059076928,0.01969231,0.0032820515,0.0,0.0,0.0,0.0,0.006564103,0.009846155,0.01969231,0.026256412,0.0,0.01969231,0.009846155,0.0,0.006564103,0.036102567,0.006564103,0.0,0.009846155,0.01969231,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.036102567,0.036102567,0.029538464,0.026256412,0.02297436,0.026256412,0.03938462,0.04594872,0.10502565,0.2100513,0.3446154,0.4594872,0.5481026,0.73517954,0.8960001,0.94523084,0.827077,0.7450257,0.58420515,0.37415388,0.17723078,0.08861539,0.059076928,0.059076928,0.08861539,0.16738462,0.34133336,0.6432821,1.2898463,1.7394873,1.6640002,0.97805136,0.49887183,0.19692309,0.08861539,0.13784617,0.25271797,0.446359,0.60389745,0.60061544,0.49230772,0.51856416,0.5152821,0.5940513,0.6892308,0.7318975,0.6432821,0.636718,0.67938465,0.74830776,0.80738467,0.81394875,0.892718,0.84348726,0.81394875,0.8566154,0.9189744,0.62030774,0.508718,0.5874872,0.7253334,0.65641034,0.702359,0.764718,0.9124103,1.142154,1.3686155,1.2668719,1.3292309,1.3883078,1.3620514,1.2570257,1.0732309,0.8533334,0.6695385,0.5481026,0.46933338,0.44964105,0.4397949,0.4594872,0.51856416,0.6268718,0.65969235,0.7318975,0.8533334,1.014154,1.1585642,1.2471796,1.3718976,1.3062565,1.1191796,1.1881026,1.0436924,0.9682052,1.0305642,1.1881026,1.2865642,1.0929232,1.0371283,0.9944616,0.9321026,0.8960001,0.7975385,0.6104616,0.4594872,0.40369233,0.4135385,0.40697438,0.35774362,0.29538465,0.24615386,0.2297436,0.22646156,0.22646156,0.25271797,0.29538465,0.3052308,0.33805132,0.3511795,0.3249231,0.26584616,0.20676924,0.25928208,0.2986667,0.3314872,0.3511795,0.3314872,0.30851284,0.23958977,0.18379489,0.16738462,0.17066668,0.19692309,0.26584616,0.3249231,0.35446155,0.35446155,0.3314872,0.34133336,0.35774362,0.3708718,0.39384618,0.39712822,0.380718,0.35774362,0.3446154,0.35446155,0.42338464,0.4660513,0.49230772,0.54482055,0.69907695,0.78769237,0.73517954,0.6465641,0.62030774,0.72861546,0.65641034,0.62030774,0.6859488,0.8467693,1.0305642,0.98461545,0.86317956,0.7056411,0.57764107,0.5546667,0.0032820515,0.0,0.0,0.0032820515,0.029538464,0.108307704,0.3249231,0.3314872,0.20020515,0.049230773,0.029538464,0.06564103,0.03938462,0.009846155,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.0,0.0,0.0,0.006564103,0.03938462,0.13128206,0.4004103,1.2012309,2.1989746,2.7634873,1.9692309,1.3718976,1.3981539,1.910154,2.8488207,4.240411,5.0018463,5.3202057,4.8114877,4.417641,6.416411,7.6734366,9.084719,11.926975,16.879591,24.021336,26.010258,24.566156,28.757336,41.088,57.504826,59.854774,46.565746,30.106258,18.58954,15.793232,16.436514,16.886156,16.154257,14.5952835,13.915898,14.569027,13.88636,13.640206,14.674052,16.922258,15.783386,15.353437,15.570052,15.947489,15.563488,17.897026,19.108105,19.685745,19.958155,20.096,20.742565,22.636309,24.336412,24.864822,23.702976,23.75549,24.6679,26.22359,27.621746,27.490463,26.912823,23.939283,21.074053,19.51836,19.170464,20.263386,21.710772,22.130873,21.530258,21.316925,21.891283,19.826874,17.903591,17.818258,20.164925,19.419899,18.60595,18.097233,18.22195,19.239386,21.458054,24.320002,28.632618,31.087593,24.25108,16.406975,11.9171295,8.763078,5.9569235,3.5347695,2.8882053,2.3860514,2.0250258,1.9659488,2.5304618,2.2744617,2.3368206,2.806154,3.0194874,1.5655385,1.9429746,2.2646155,2.3302567,2.7602053,4.9920006,4.1682053,4.7261543,5.8420515,6.678975,6.380308,7.397744,8.280616,8.87795,9.465437,10.742155,9.179898,9.321027,9.590155,12.826258,26.272823,41.934772,37.796104,32.288822,29.682875,20.069746,9.895386,8.0377445,11.464206,13.925745,5.970052,11.444513,24.152617,34.917747,41.537643,48.77785,36.58831,29.906054,27.02113,22.239182,5.865026,5.1232824,7.9130263,7.975385,4.7458467,3.3345644,5.0018463,6.5444107,6.9710774,7.0498466,9.291488,7.325539,4.585026,2.5600002,1.7427694,1.6246156,1.9593848,2.7437952,3.8334363,5.35959,7.7259493,7.9917955,6.4722056,5.225026,4.7261543,3.8564105,3.9154875,2.9505644,3.6562054,6.567385,10.069334,9.6754875,13.387488,16.738462,15.586463,6.117744,8.736821,12.868924,13.249642,9.639385,6.8004107,9.265231,8.710565,9.997129,13.528616,15.27795,14.260514,15.209026,19.797335,23.762053,16.889437,11.487181,7.4010262,5.973334,6.62318,6.8266673,3.7152824,3.6660516,3.2295387,2.1858463,3.5380516,8.467693,20.919796,38.22277,51.045746,43.414978,23.348515,15.058052,10.66995,7.768616,9.409642,15.153232,21.300514,18.500925,9.744411,10.364718,20.916515,20.575182,18.504206,19.012924,21.563078,19.77436,20.050053,23.296001,27.789131,29.184002,30.25395,30.946465,31.465029,31.911386,32.301952,26.50913,19.99754,15.53395,14.690463,17.85436,21.576206,25.508104,31.159798,36.453747,35.73826,26.574772,20.6999,17.542566,16.055796,14.7331295,14.523078,14.299898,20.450462,32.594055,43.572517,39.394466,44.44554,56.835285,64.49231,45.206978,43.14585,41.449028,33.447388,20.227283,10.610872,18.507488,16.961643,14.083283,15.927796,26.479591,16.57436,11.818667,10.35159,10.699488,11.772718,6.6428723,3.95159,3.4855387,3.9548721,2.9669745,8.211693,6.5739493,6.626462,8.454565,3.6594875,3.4724104,5.2348723,5.723898,5.9503593,11.145847,13.354668,7.2303596,5.5236926,9.055181,6.695385,4.7360005,6.2752824,6.8627696,5.297231,3.629949,4.7983594,2.477949,2.044718,5.179077,9.869129,5.920821,2.674872,2.5009232,4.594872,4.9427695,4.204308,5.4449234,5.402257,4.7228723,7.9491286,13.259488,10.092308,5.0871797,2.5993848,4.716308,3.7021542,4.325744,7.433847,10.04636,5.366154,2.8947694,4.1911798,5.293949,4.969026,4.709744,2.356513,1.2931283,0.7778462,0.43651286,0.27241027,0.37743592,0.30194873,0.18051283,0.101743594,0.098461546,0.059076928,0.026256412,0.009846155,0.009846155,0.026256412,0.03938462,0.18707694,0.37743592,0.50543594,0.45620516,0.39056414,0.25928208,0.256,0.36430773,0.37415388,0.36102566,0.40697438,0.3314872,0.16410258,0.15097436,0.19364104,0.16410258,0.118153855,0.1148718,0.21333335,0.6498462,0.65641034,0.52512825,0.380718,0.18051283,0.13456412,0.16410258,0.19692309,0.21661541,0.26912823,0.13128206,0.19692309,0.3708718,0.46276927,0.17723078,0.0951795,0.11158975,0.190359,0.2231795,0.04594872,0.016410258,0.01969231,0.18707694,0.574359,1.142154,1.3817437,0.81394875,0.29538465,0.12471796,0.052512825,0.013128206,0.0,0.0,0.0032820515,0.02297436,0.026256412,0.013128206,0.0032820515,0.0032820515,0.013128206,0.013128206,0.006564103,0.0032820515,0.0032820515,0.013128206,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.03938462,0.04594872,0.108307704,0.17066668,0.19692309,0.16738462,0.21333335,0.24943592,0.16738462,0.016410258,0.0,0.0,0.0,0.01969231,0.04266667,0.02297436,0.006564103,0.0,0.0,0.0,0.0,0.059076928,0.12471796,0.14441027,0.118153855,0.098461546,0.049230773,0.101743594,0.25928208,0.36430773,0.108307704,0.072205134,0.23302566,0.76800007,1.270154,0.7515898,0.33805132,0.20348719,0.13128206,0.04594872,0.009846155,0.0032820515,0.009846155,0.009846155,0.0,0.0,0.0,0.029538464,0.03938462,0.02297436,0.0032820515,0.0032820515,0.06235898,0.12471796,0.13456412,0.03938462,0.02297436,0.072205134,0.11158975,0.0951795,0.029538464,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.013128206,0.013128206,0.04266667,0.01969231,0.0,0.0,0.0,0.0,0.0,0.01969231,0.03938462,0.0,0.0,0.0,0.0032820515,0.009846155,0.0,0.0,0.006564103,0.006564103,0.009846155,0.052512825,0.04594872,0.029538464,0.016410258,0.016410258,0.026256412,0.026256412,0.049230773,0.07876924,0.118153855,0.190359,0.318359,0.54482055,0.7450257,0.83035904,0.7515898,0.78769237,0.7089231,0.50543594,0.25928208,0.13456412,0.08205129,0.055794876,0.049230773,0.101743594,0.27897438,0.5415385,1.014154,1.6672822,2.0545642,1.3161026,0.82379496,0.36758977,0.13456412,0.15753847,0.31507695,0.38728207,0.5021539,0.56123084,0.58420515,0.7187693,0.6465641,0.6826667,0.7384616,0.7515898,0.67610264,0.6071795,0.64000005,0.7187693,0.78769237,0.8041026,0.93866676,0.8533334,0.7778462,0.79097444,0.78769237,0.6662565,0.6826667,0.7515898,0.79425645,0.7581539,0.6235898,0.7056411,0.92553854,1.1716924,1.3062565,1.3981539,1.4605129,1.4736412,1.4145643,1.2668719,1.2406155,1.0896411,0.8730257,0.65641034,0.51856416,0.48902568,0.4660513,0.48902568,0.5513847,0.61374366,0.56123084,0.57764107,0.67938465,0.81394875,0.88943595,0.98461545,1.1388719,1.214359,1.2209232,1.3292309,1.1158975,1.017436,1.0469744,1.142154,1.1749744,1.1388719,1.2274873,1.1946667,1.0568206,1.1060513,0.95835906,0.7253334,0.5218462,0.40369233,0.3708718,0.36102566,0.32164106,0.28225642,0.25271797,0.23302566,0.23958977,0.26256412,0.3052308,0.34789747,0.3446154,0.4266667,0.4201026,0.34133336,0.24287182,0.20020515,0.27569234,0.29210258,0.2855385,0.27569234,0.28225642,0.29210258,0.24615386,0.18707694,0.14441027,0.1148718,0.13784617,0.23630771,0.318359,0.3511795,0.35774362,0.40369233,0.42338464,0.41682056,0.39384618,0.4004103,0.34133336,0.28882053,0.25928208,0.25271797,0.26256412,0.3511795,0.42994875,0.47917953,0.52512825,0.6432821,0.79425645,0.7220513,0.56123084,0.4594872,0.57764107,0.64000005,0.6268718,0.67938465,0.81394875,0.92225647,0.9747693,0.88943595,0.6662565,0.42338464,0.40369233,0.016410258,0.0032820515,0.0,0.0,0.02297436,0.108307704,0.032820515,0.02297436,0.049230773,0.07876924,0.09189744,0.21333335,0.14441027,0.04594872,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.032820515,0.04594872,0.16738462,0.6104616,1.2832822,1.7362052,1.1749744,0.6268718,1.7427694,2.9636924,3.826872,4.97559,6.7183595,5.85518,4.7524104,4.388103,4.3651285,8.123077,12.744206,16.479181,19.15077,22.14072,21.88472,21.62872,29.252926,44.150158,57.235695,52.719593,38.61662,26.09231,19.541334,16.587488,15.55036,14.769232,13.400617,12.340514,14.221129,14.158771,13.036308,13.459693,15.176207,15.090873,12.22236,11.769437,12.813129,14.427898,15.684924,20.178053,21.064207,20.191181,19.423182,20.644104,21.24472,21.336617,21.809233,22.90872,24.277336,24.34954,25.091284,25.38995,24.999386,24.536617,24.684309,24.408617,24.211695,23.919592,22.675694,21.648413,21.510565,20.65067,19.144207,18.753643,20.158361,18.474669,16.315079,14.864411,13.90277,15.415796,17.880617,20.329027,22.806976,26.38113,32.777847,36.64739,33.024002,23.650463,16.997746,13.725539,9.8592825,6.9809237,5.2414365,3.387077,2.5435898,2.2055387,1.8937438,1.5786668,1.6640002,1.847795,1.5360001,1.6869745,2.2383592,2.0906668,2.8947694,4.4242053,4.637539,3.3575387,2.2580514,3.9417439,4.309334,4.71959,5.6352825,6.636308,8.310155,8.644924,8.408616,8.484103,9.888822,12.524308,16.019693,16.856617,18.14318,29.617233,30.631388,25.071592,23.22708,24.388926,16.846771,6.994052,6.7938466,14.106257,20.775387,12.632616,8.861539,14.25395,18.809437,21.06749,28.1239,25.521233,20.066463,16.659693,13.814155,3.6332312,2.8980515,4.775385,5.412103,3.8596926,2.0906668,2.0775387,3.9975388,5.671385,6.413129,7.0334363,6.229334,3.8662567,1.8510771,1.0994873,1.5261539,2.0250258,1.785436,1.7657437,2.4188719,3.6627696,3.4789746,2.5632823,1.7263591,1.4178462,1.7099489,2.7831798,2.2908719,2.665026,3.767795,2.9144619,5.4416413,10.807796,14.500104,13.430155,5.937231,6.2785645,7.709539,7.525744,5.579488,4.273231,3.8564105,4.7524104,5.6320004,7.2927184,12.665437,7.4404106,8.073847,11.608616,14.290052,11.565949,8.625232,7.138462,6.4590774,6.0947695,5.691077,5.47118,3.9614363,2.3696413,1.6705642,2.609231,3.9154875,8.342975,19.538054,32.57436,33.96595,25.580309,31.209028,28.163284,15.766975,15.366566,27.582361,38.163696,38.915283,30.421335,22.048822,28.800003,27.237745,27.139284,29.105232,24.566156,16.30195,12.461949,14.628103,20.164925,22.20308,25.449028,27.808823,25.360413,19.51836,17.030565,16.101746,13.003489,11.208206,12.0549755,14.739694,16.754873,32.74831,52.77867,63.812927,49.726364,31.796515,21.618874,16.712206,14.112822,10.377847,11.329642,14.624822,17.499899,24.628515,48.12472,37.041233,35.09498,41.193027,47.46503,39.2599,35.45272,30.930054,24.234669,16.33477,10.633847,19.413334,16.59077,11.204924,8.536616,10.085744,14.17518,12.724514,9.833026,8.234667,9.3078985,7.9294367,6.5312824,6.3343596,7.020308,6.7150774,11.109744,7.939283,11.139283,17.207796,5.2348723,5.674667,7.788308,6.2818465,2.9801028,6.8365135,9.435898,6.3606157,5.8157954,8.477539,7.4765134,7.2927184,7.1844106,5.211898,2.8947694,5.2020516,9.340718,5.0018463,1.6147693,2.6190772,5.464616,7.207385,3.9187696,2.0644104,3.4789746,5.3694363,4.699898,10.19077,12.228924,8.546462,4.2272825,10.94236,13.341539,10.535385,5.533539,5.2644105,4.640821,4.4865646,4.955898,5.549949,5.097026,3.5347695,5.0576415,5.668103,4.197744,2.3040001,3.3772311,2.9965131,2.100513,1.2964103,0.86974365,0.6268718,0.41025645,0.24287182,0.15753847,0.18379489,0.08533334,0.02297436,0.013128206,0.026256412,0.016410258,0.026256412,0.0951795,0.23958977,0.41682056,0.5021539,0.380718,0.21333335,0.14112821,0.19364104,0.28882053,0.31507695,0.39384618,0.35774362,0.22646156,0.21333335,0.3708718,0.32164106,0.19364104,0.07876924,0.029538464,0.055794876,0.068923086,0.07548718,0.068923086,0.04594872,0.108307704,0.15097436,0.14441027,0.14769232,0.3052308,0.20676924,0.16410258,0.3052308,0.46933338,0.21333335,0.09189744,0.18051283,0.3249231,0.36430773,0.108307704,0.059076928,0.01969231,0.08533334,0.33476925,0.82379496,0.81066674,0.5973334,0.36758977,0.2231795,0.19692309,0.052512825,0.006564103,0.0,0.0,0.0,0.013128206,0.02297436,0.01969231,0.0,0.0,0.013128206,0.016410258,0.009846155,0.0,0.0,0.049230773,0.02297436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.052512825,0.068923086,0.11158975,0.16738462,0.16738462,0.15425642,0.16082053,0.118153855,0.036102567,0.0,0.0,0.0,0.098461546,0.21989745,0.12143591,0.036102567,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.098461546,0.15753847,0.21333335,0.23958977,0.16738462,0.04594872,0.12471796,0.2100513,0.27569234,0.45620516,0.7384616,0.75487185,0.5415385,0.2297436,0.04594872,0.009846155,0.009846155,0.009846155,0.0,0.0,0.0,0.0,0.006564103,0.016410258,0.016410258,0.016410258,0.016410258,0.009846155,0.0032820515,0.016410258,0.026256412,0.049230773,0.09189744,0.14112821,0.15097436,0.029538464,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.02297436,0.06235898,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02297436,0.049230773,0.0,0.0,0.036102567,0.036102567,0.016410258,0.07548718,0.052512825,0.036102567,0.02297436,0.016410258,0.016410258,0.016410258,0.016410258,0.03938462,0.07876924,0.09189744,0.15097436,0.25928208,0.380718,0.51856416,0.702359,0.8369231,0.8336411,0.67282057,0.4266667,0.24287182,0.12143591,0.06564103,0.04594872,0.068923086,0.16738462,0.4594872,0.7450257,1.1782565,1.5721027,1.3883078,0.8402052,0.4266667,0.16410258,0.04594872,0.04594872,0.16738462,0.35446155,0.4955898,0.5973334,0.79425645,0.6235898,0.69907695,0.7844103,0.81066674,0.88615394,0.67610264,0.6629744,0.6629744,0.6465641,0.7318975,0.76800007,0.761436,0.636718,0.48246157,0.51856416,0.6892308,0.8598975,0.9353847,0.892718,0.79425645,0.7581539,0.81066674,0.8369231,0.84348726,0.97805136,0.93866676,0.95835906,0.90256417,0.7778462,0.7187693,0.827077,0.98133343,0.9944616,0.8730257,0.82379496,0.7253334,0.6301539,0.5874872,0.5874872,0.56451285,0.5415385,0.5152821,0.54482055,0.6301539,0.7187693,0.75487185,0.8369231,0.96492314,1.1585642,1.463795,1.3193847,1.2438976,1.2406155,1.2242053,1.0535386,0.9189744,1.014154,1.1093334,1.1290257,1.1290257,1.0305642,0.8336411,0.6432821,0.50543594,0.39712822,0.39712822,0.3511795,0.29538465,0.256,0.24287182,0.23302566,0.2297436,0.24615386,0.28225642,0.32164106,0.49230772,0.5349744,0.43651286,0.27569234,0.21333335,0.2855385,0.3052308,0.26256412,0.19692309,0.19692309,0.19692309,0.23630771,0.23958977,0.20020515,0.15097436,0.16410258,0.15753847,0.17723078,0.2231795,0.25928208,0.3446154,0.37415388,0.35774362,0.3249231,0.3511795,0.30194873,0.25271797,0.2231795,0.23958977,0.33476925,0.54482055,0.61374366,0.5874872,0.5349744,0.5349744,0.54482055,0.5940513,0.5513847,0.44307697,0.44307697,0.4660513,0.54482055,0.636718,0.702359,0.702359,0.77456415,0.8041026,0.6629744,0.4135385,0.3052308,0.0032820515,0.0,0.0,0.0,0.0032820515,0.02297436,0.016410258,0.009846155,0.01969231,0.055794876,0.1148718,0.101743594,0.06235898,0.032820515,0.02297436,0.013128206,0.0032820515,0.029538464,0.049230773,0.03938462,0.0,0.0,0.0,0.013128206,0.029538464,0.02297436,0.08533334,0.3446154,0.83035904,1.3029745,1.2603078,0.88615394,1.7329233,3.2951798,4.709744,4.7556925,4.965744,5.684513,6.373744,6.925129,7.6242056,9.478565,12.251899,15.363283,18.189129,20.066463,18.218668,16.882874,22.85949,35.764515,48.019695,45.31857,33.496616,24.136208,20.857437,19.30831,16.689232,15.425642,14.060308,13.10195,15.002257,14.588719,13.8765135,14.375385,15.343591,13.784616,11.464206,11.684103,14.089848,17.289848,18.858667,20.089437,20.437334,20.736002,21.07077,20.778667,20.25354,20.345438,21.241438,23.066257,25.888823,25.189745,25.540926,25.70831,25.3079,24.805746,24.054155,24.021336,23.991796,23.5159,22.419695,23.463387,23.243488,22.048822,20.246977,18.264616,19.738258,20.17477,20.841026,21.894566,22.396719,22.94154,25.819899,28.442259,30.644516,34.671593,37.894566,34.671593,27.549541,19.856411,15.704617,12.599796,9.527796,6.9710774,4.962462,3.1081028,2.4418464,1.8904617,1.4276924,1.2570257,1.8084104,2.1792822,2.3171284,5.402257,8.832001,4.2141542,3.4855387,3.2032824,2.6945643,2.1169233,2.4549747,3.131077,4.850872,5.9667697,6.669129,8.969847,9.888822,12.2847185,14.326155,14.162052,9.911796,11.191795,14.408206,15.579899,14.788924,16.167385,16.768002,18.356514,17.952822,16.715488,19.93518,13.804309,10.180923,12.498053,17.621334,15.845745,9.055181,8.802463,9.938052,11.264001,15.524104,17.631182,14.194873,11.050668,9.091283,4.240411,2.5042052,2.5829747,3.2525132,3.3903592,1.9922053,1.6475899,3.4198978,4.07959,3.4822567,4.5456414,3.6693337,2.2580514,1.7033848,1.9429746,1.4539489,1.4244103,1.083077,0.8730257,1.1454359,2.1366155,2.540308,1.8576412,1.0962052,0.827077,1.2077949,1.529436,1.6640002,1.8018463,1.8149745,1.2537436,3.1671798,6.4295387,8.211693,7.0826674,3.006359,2.428718,2.861949,2.8455386,2.0939488,1.4900514,1.3095386,1.5524104,2.3335385,4.394667,9.101129,4.7655387,4.141949,5.9963083,8.162462,7.5388722,5.4941545,4.8705645,4.781949,4.6112823,3.9942567,3.373949,3.18359,2.6157951,2.5961027,5.7829747,8.982975,8.333129,11.08677,18.04472,23.56513,30.628105,29.033028,20.292925,10.581334,10.7158985,12.370052,18.20554,22.268719,21.85518,17.545847,18.340103,18.976822,23.666874,33.430977,46.1358,37.842052,26.105438,19.27877,18.914463,19.771078,20.696617,25.38667,25.56718,19.544617,12.219078,12.179693,13.407181,18.560001,26.942362,34.487797,48.00657,68.31918,79.27467,78.27693,76.28801,47.35344,37.67467,31.908106,23.322258,13.804309,11.195078,13.817437,16.643284,20.752413,33.332516,39.492928,37.792824,35.328003,32.82708,24.661335,21.782976,19.452719,16.981335,14.221129,11.588924,17.122463,19.121233,15.491283,9.334154,8.950154,9.622975,9.002667,9.819899,10.8537445,6.928411,6.925129,6.8299494,7.8080006,9.107693,8.080411,12.836103,9.957745,10.246565,13.545027,8.736821,5.474462,7.7718983,12.826258,14.723283,4.4307694,7.958975,8.2215395,8.1066675,7.5585647,3.5577438,4.4406157,4.089436,3.564308,3.8301542,5.7632823,6.7971287,4.1058464,2.0939488,2.3204105,3.4855387,8.618668,8.887795,6.2851286,3.3476925,3.1507695,1.8642052,3.1573336,4.1058464,4.2896414,5.789539,16.154257,16.846771,11.437949,5.106872,4.6539493,3.945026,4.089436,5.5991797,7.3485136,6.5739493,4.3651285,3.3903592,3.255795,3.2689233,2.4516926,2.7733335,1.9035898,0.9714873,0.5316923,0.56451285,0.4266667,0.28882053,0.17394873,0.108307704,0.13456412,0.0951795,0.049230773,0.02297436,0.016410258,0.016410258,0.026256412,0.0951795,0.20676924,0.34789747,0.49230772,0.48574364,0.3708718,0.32164106,0.43651286,0.72861546,0.35446155,0.36102566,0.40697438,0.33805132,0.190359,0.32820517,0.23630771,0.12471796,0.07876924,0.029538464,0.016410258,0.23958977,0.5349744,0.61374366,0.068923086,0.052512825,0.08205129,0.118153855,0.13784617,0.15753847,0.101743594,0.059076928,0.12143591,0.25928208,0.33476925,0.20348719,0.20348719,0.32820517,0.47917953,0.43651286,0.21333335,0.08533334,0.052512825,0.12471796,0.3117949,0.36758977,0.4135385,0.4201026,0.36102566,0.2100513,0.12143591,0.055794876,0.013128206,0.0,0.0,0.0032820515,0.0032820515,0.0032820515,0.0,0.0,0.0032820515,0.016410258,0.02297436,0.009846155,0.0,0.009846155,0.013128206,0.006564103,0.0,0.0,0.01969231,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.029538464,0.04594872,0.06564103,0.08533334,0.0951795,0.072205134,0.08205129,0.068923086,0.026256412,0.0,0.0,0.0,0.03938462,0.101743594,0.108307704,0.052512825,0.04594872,0.029538464,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.02297436,0.04266667,0.108307704,0.16738462,0.20348719,0.2297436,0.12471796,0.072205134,0.07876924,0.17066668,0.3708718,0.7811283,0.6892308,0.4004103,0.18379489,0.26584616,0.072205134,0.026256412,0.029538464,0.029538464,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0032820515,0.0032820515,0.0032820515,0.0,0.0032820515,0.006564103,0.009846155,0.06235898,0.13784617,0.14112821,0.029538464,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.02297436,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.0,0.0,0.006564103,0.013128206,0.016410258,0.03938462,0.026256412,0.01969231,0.016410258,0.016410258,0.016410258,0.006564103,0.009846155,0.016410258,0.026256412,0.06564103,0.03938462,0.11158975,0.20348719,0.3052308,0.45620516,0.571077,0.6662565,0.67282057,0.56451285,0.34133336,0.20020515,0.101743594,0.052512825,0.055794876,0.0951795,0.28882053,0.5349744,0.8598975,1.2274873,1.522872,1.5885129,0.9419488,0.34789747,0.101743594,0.032820515,0.08861539,0.23302566,0.44964105,0.65641034,0.7450257,0.69907695,0.77128214,0.761436,0.6892308,0.81066674,0.63343596,0.5677949,0.5677949,0.6104616,0.69579494,0.702359,0.7089231,0.7122052,0.71548724,0.71548724,0.9616411,1.3423591,1.9528207,2.2547693,1.0633847,0.77128214,0.8008206,0.9911796,1.1749744,1.1716924,1.3292309,1.3456411,1.3161026,1.2242053,0.9485129,1.0305642,1.0601027,0.98461545,0.8402052,0.7515898,0.69251287,0.6104616,0.53825647,0.49230772,0.4660513,0.5218462,0.5316923,0.52512825,0.5349744,0.58420515,0.60061544,0.73517954,0.88287187,0.99774367,1.0994873,1.1093334,1.1782565,1.2406155,1.2373334,1.1257436,0.9419488,0.84348726,0.827077,0.84348726,0.77456415,0.7056411,0.64000005,0.60389745,0.56123084,0.43323082,0.37415388,0.31507695,0.26584616,0.2297436,0.20676924,0.27241027,0.28882053,0.32164106,0.380718,0.41682056,0.4135385,0.4201026,0.41025645,0.36758977,0.2855385,0.30194873,0.2986667,0.27897438,0.24615386,0.19692309,0.18707694,0.17066668,0.15425642,0.14112821,0.14112821,0.17066668,0.19364104,0.21661541,0.24287182,0.25928208,0.3052308,0.3052308,0.30194873,0.30851284,0.30194873,0.28225642,0.26256412,0.26584616,0.3052308,0.38400003,0.41682056,0.39712822,0.3708718,0.35446155,0.37415388,0.43651286,0.5546667,0.6301539,0.5907693,0.40697438,0.39056414,0.4397949,0.5021539,0.56451285,0.65312827,0.77456415,0.8730257,0.7581539,0.48246157,0.34133336,0.0,0.0,0.0,0.006564103,0.013128206,0.0,0.0032820515,0.013128206,0.02297436,0.03938462,0.07548718,0.049230773,0.036102567,0.10502565,0.17394873,0.016410258,0.009846155,0.036102567,0.049230773,0.032820515,0.0,0.006564103,0.013128206,0.026256412,0.036102567,0.016410258,0.026256412,0.17723078,0.56123084,1.079795,1.4375386,1.2603078,1.3817437,2.0020514,2.861949,3.2164104,3.639795,4.529231,5.658257,7.00718,8.795898,10.7158985,12.202667,14.011078,16.118155,17.72636,15.645539,15.271386,20.545643,30.785643,40.68103,37.776413,29.892925,23.926155,21.632002,19.623386,18.159592,17.64759,17.34236,17.368616,18.68472,19.643078,19.958155,21.195488,22.291695,19.528206,15.937642,15.95077,17.975796,20.397951,21.586054,21.48759,21.444925,21.504002,21.231592,19.731693,19.98113,20.73272,22.098053,23.958977,25.951181,25.353848,25.088001,23.456821,21.241438,21.704206,22.075079,23.305847,23.574976,22.344208,20.368412,22.41313,23.6439,23.135181,21.284103,19.826874,20.342155,21.825644,23.59467,24.740105,24.136208,25.951181,28.921438,31.27467,32.9879,35.800617,35.30831,31.415798,25.271797,18.84554,14.913642,12.406155,9.032206,6.012718,4.0303593,3.239385,3.318154,3.0752823,2.9472823,3.5052311,5.481026,5.405539,7.0104623,8.73354,8.579283,4.132103,2.9997952,2.6157951,2.681436,3.062154,3.7940516,4.916513,6.38359,7.240206,8.064001,10.952206,12.445539,13.988104,15.228719,15.911386,15.8884115,17.220924,16.764719,15.734155,15.576616,17.96595,15.881847,16.41354,13.942155,10.55836,16.055796,15.812924,11.290257,9.915077,13.056001,16.01641,7.5552826,4.854154,4.516103,5.218462,7.716103,10.289231,8.700719,6.2884107,4.4340515,2.546872,1.5885129,2.0250258,3.4822567,5.0576415,5.3202057,4.2240005,3.8531284,2.9144619,1.9298463,3.2361028,3.4198978,1.8281027,1.0075898,1.3161026,0.90256417,0.7811283,0.636718,0.47261542,0.47917953,1.0043077,1.5688206,1.4933335,1.0469744,0.6465641,0.8369231,0.8960001,1.5360001,1.6738462,1.1224617,0.58420515,1.5360001,3.131077,3.8498464,3.0916924,1.1946667,0.85005134,1.142154,1.3062565,1.0338463,0.48246157,0.6104616,1.3062565,3.1934361,5.5171285,6.1407185,3.623385,2.4746668,2.7667694,3.889231,4.5522056,3.9286156,3.7251284,3.4002054,3.0752823,3.515077,2.605949,2.8192823,2.8192823,2.737231,4.1682053,9.55077,8.759795,8.864821,12.836103,19.538054,26.558361,22.665848,16.833643,14.221129,16.144411,9.80677,10.200616,14.605129,19.321438,19.649643,17.585232,17.063385,22.347488,34.55344,51.656208,78.94975,78.57231,72.50708,63.104004,33.089645,22.422976,25.688618,29.604105,26.902977,16.33477,13.361232,16.879591,24.713848,33.854362,40.44472,57.57703,71.97539,72.749954,69.805954,93.86339,55.479797,43.346054,36.68677,27.474054,20.43077,13.289026,12.550565,12.737642,13.062565,17.430975,28.255182,27.720207,25.521233,24.329847,19.784206,17.890463,16.682669,15.645539,14.375385,12.603078,16.843489,21.251284,18.087385,10.06277,10.325335,10.594462,13.197129,12.544001,8.5891285,6.8266673,9.357129,9.639385,9.760821,9.718155,7.387898,16.7319,11.07036,7.7259493,10.581334,10.108719,5.4580517,7.9327188,12.727796,13.653335,3.1343591,6.439385,7.0104623,6.409847,5.149539,2.678154,4.9329233,5.1232824,5.3792825,5.9536414,5.228308,4.896821,3.5938463,2.8192823,2.7470772,2.1956925,6.1768208,8.356103,7.328821,4.132103,2.2088206,1.2537436,2.858667,4.699898,5.540103,5.228308,10.312206,9.846154,7.1023593,4.8016415,5.106872,3.9351797,4.460308,6.5345645,8.257642,5.989744,4.2896414,3.9286156,5.0477953,6.11118,3.9056413,2.4451284,1.273436,0.60389745,0.39384618,0.34133336,0.42338464,0.49230772,0.36758977,0.11158975,0.049230773,0.03938462,0.026256412,0.01969231,0.016410258,0.016410258,0.036102567,0.10502565,0.17394873,0.2231795,0.24943592,0.38400003,0.33476925,0.29210258,0.380718,0.6662565,0.3511795,0.3708718,0.446359,0.40697438,0.20020515,0.23958977,0.15753847,0.08861539,0.07548718,0.03938462,0.016410258,0.7318975,1.3029745,1.1684103,0.0951795,0.04266667,0.04594872,0.08861539,0.128,0.0951795,0.10502565,0.055794876,0.055794876,0.14441027,0.3117949,0.27241027,0.18379489,0.17066668,0.256,0.36430773,0.26912823,0.14769232,0.06564103,0.049230773,0.09189744,0.14441027,0.27569234,0.39384618,0.39712822,0.18707694,0.16410258,0.12471796,0.06235898,0.0032820515,0.01969231,0.009846155,0.0032820515,0.0032820515,0.006564103,0.0,0.0,0.013128206,0.02297436,0.02297436,0.01969231,0.0032820515,0.0032820515,0.006564103,0.006564103,0.0,0.016410258,0.013128206,0.006564103,0.0,0.0,0.0,0.006564103,0.006564103,0.0,0.0,0.009846155,0.016410258,0.02297436,0.04266667,0.08533334,0.118153855,0.13128206,0.12143591,0.108307704,0.118153855,0.04594872,0.009846155,0.009846155,0.032820515,0.068923086,0.049230773,0.108307704,0.09189744,0.0,0.0,0.0,0.026256412,0.026256412,0.0032820515,0.013128206,0.013128206,0.03938462,0.068923086,0.11158975,0.190359,0.13456412,0.71548724,0.69251287,0.08533334,0.17723078,0.40369233,0.48574364,0.43323082,0.34133336,0.39384618,0.31507695,0.17066668,0.09189744,0.0951795,0.072205134,0.036102567,0.03938462,0.029538464,0.006564103,0.0,0.0,0.0,0.013128206,0.04594872,0.08205129,0.10502565,0.04266667,0.07548718,0.17723078,0.108307704,0.029538464,0.0032820515,0.006564103,0.016410258,0.009846155,0.0032820515,0.0,0.0,0.0,0.006564103,0.02297436,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.02297436,0.016410258,0.009846155,0.009846155,0.016410258,0.016410258,0.0032820515,0.0032820515,0.0032820515,0.0032820515,0.02297436,0.0032820515,0.052512825,0.101743594,0.14441027,0.23302566,0.3708718,0.55794877,0.6498462,0.5973334,0.4397949,0.30851284,0.190359,0.101743594,0.055794876,0.059076928,0.19364104,0.38400003,0.65969235,1.0305642,1.5195899,1.5261539,1.0601027,0.56123084,0.24287182,0.08533334,0.07876924,0.15097436,0.34133336,0.6104616,0.8336411,0.7844103,0.76800007,0.72861546,0.67938465,0.7122052,0.5907693,0.5415385,0.5546667,0.61374366,0.6695385,0.6695385,0.63343596,0.63343596,0.6826667,0.7450257,0.86646163,1.083077,1.5425643,2.034872,1.9889232,1.5195899,1.1520001,1.0568206,1.1946667,1.339077,1.3193847,1.4998976,1.5885129,1.4408206,1.0436924,0.98461545,0.9682052,1.0075898,1.0338463,0.90584624,0.7844103,0.6892308,0.5874872,0.48574364,0.43323082,0.48574364,0.4660513,0.446359,0.45620516,0.4955898,0.5218462,0.6301539,0.7450257,0.84348726,0.9419488,0.9419488,1.0108719,1.0962052,1.1388719,1.0699488,0.9353847,0.8598975,0.77128214,0.6432821,0.5218462,0.52512825,0.5218462,0.5021539,0.4660513,0.40697438,0.3708718,0.2855385,0.23302566,0.2231795,0.20676924,0.22646156,0.25271797,0.318359,0.4201026,0.5152821,0.512,0.54482055,0.5415385,0.4660513,0.36102566,0.3446154,0.3117949,0.27241027,0.23630771,0.190359,0.20020515,0.18379489,0.15425642,0.12471796,0.128,0.14441027,0.17066668,0.21333335,0.256,0.25928208,0.26584616,0.24943592,0.256,0.28225642,0.26256412,0.23630771,0.25928208,0.31507695,0.39056414,0.46933338,0.45620516,0.36758977,0.3117949,0.3314872,0.4004103,0.43651286,0.49887183,0.571077,0.58420515,0.43323082,0.3708718,0.4135385,0.47589746,0.51856416,0.5481026,0.6170257,0.7220513,0.7220513,0.5940513,0.43323082,0.0,0.0,0.0,0.006564103,0.013128206,0.0,0.0,0.009846155,0.01969231,0.02297436,0.032820515,0.068923086,0.04266667,0.09189744,0.16738462,0.026256412,0.032820515,0.04594872,0.04266667,0.026256412,0.006564103,0.013128206,0.02297436,0.052512825,0.08205129,0.08205129,0.026256412,0.118153855,0.4004103,0.8336411,1.3029745,1.3423591,1.0010257,0.98133343,1.4441026,2.03159,2.6584618,3.3312824,4.3618464,6.121026,9.051898,10.857026,11.881026,13.11836,14.6642065,15.727591,14.421334,15.035078,19.081848,25.967592,32.978054,30.834875,27.319798,24.22154,21.897848,19.288616,19.393642,19.695591,20.053335,20.693335,22.199797,23.857233,25.849438,27.959797,28.744207,25.550772,21.691078,20.473438,20.8279,21.825644,22.695387,21.129848,20.489847,19.86954,18.960411,18.070976,20.299488,21.589334,22.826668,24.119797,24.799181,24.336412,23.046566,20.233849,17.46708,18.566566,20.401232,22.160412,22.439386,21.13313,19.416616,21.471182,23.341951,23.092514,21.287386,20.985437,21.569643,23.312412,25.51795,26.719181,24.681028,27.759592,30.447592,32.292107,33.18154,33.345642,30.037336,27.346054,23.785027,19.232822,14.933334,12.747488,9.304616,6.882462,6.1374364,6.1308722,6.7971287,7.0531287,7.0957956,7.709539,10.266257,10.249847,12.25518,10.5780525,5.5204105,3.4067695,3.1671798,3.2065644,3.3903592,3.9122055,5.3202057,6.5936418,6.8332314,6.550975,6.8627696,9.452309,15.189335,16.311796,14.841437,14.309745,19.764515,23.617643,18.871796,14.217847,14.979283,23.115488,18.576412,16.367592,11.58236,7.056411,13.338258,16.656412,11.943385,7.6603084,7.8802056,12.304411,5.651693,2.678154,1.7690258,2.0676925,3.501949,5.858462,5.2381544,3.570872,2.0151796,0.97805136,0.9517949,1.6475899,2.9538465,4.4406157,5.356308,4.6145644,3.3050258,1.8543591,1.2307693,2.930872,3.8728209,1.8576412,0.5874872,0.9944616,1.2570257,2.0775387,1.6869745,0.827077,0.17394873,0.3314872,0.7515898,1.3686155,1.2865642,0.7056411,0.9156924,0.64000005,1.2865642,1.4769232,0.9124103,0.35774362,0.7089231,1.214359,1.401436,1.1290257,0.5874872,0.6662565,1.2406155,1.5721027,1.3850257,0.88943595,1.6902566,2.412308,3.8334363,5.0576415,3.5216413,3.0326157,2.034872,1.3686155,1.5064616,2.550154,3.5971284,3.1770258,2.3138463,1.8970258,2.6847181,2.4451284,2.6223593,2.9210258,3.0293336,2.6420515,7.0137444,7.817847,8.218257,10.358154,15.350155,17.493334,15.186052,14.073437,15.793232,17.956104,14.139078,11.881026,13.932309,17.975796,16.617027,14.746258,15.858873,21.274258,31.251696,44.993645,108.75078,126.54278,125.72883,110.92021,63.954056,36.463593,33.283283,39.217236,42.37785,34.212105,24.070566,22.30154,26.351591,33.073235,38.76103,50.79303,57.885544,54.367184,52.21744,81.073235,48.72862,36.164925,31.031797,27.32636,25.399797,13.636924,10.469745,9.4916935,8.441437,9.189744,16.019693,15.783386,15.304206,16.36431,15.714462,16.42995,16.210052,19.03918,21.546669,13.013334,15.95077,19.672617,17.11918,10.820924,12.898462,12.107488,14.8939495,13.302155,7.9852314,8.195283,10.9686165,10.358154,9.386667,8.674462,6.449231,13.344822,8.569437,6.5706673,10.473026,12.06154,7.7357955,7.5191803,9.048616,9.189744,4.06318,7.3682055,8.326565,7.312411,5.366154,4.1747694,5.1922054,5.907693,6.422975,6.426257,5.1659493,4.7917953,4.017231,3.6069746,3.2918978,1.7723079,3.56759,6.0160003,7.4732313,6.774154,3.2164104,2.6256413,5.366154,7.3682055,6.889026,4.532513,5.4449234,4.965744,4.7327185,5.1954875,5.618872,4.6802053,5.0477953,6.0652313,6.4557953,4.3290257,4.46359,5.110154,6.1341543,6.377026,3.6693337,1.6968206,0.90912825,0.827077,0.90584624,0.54482055,1.0338463,0.8402052,0.42338464,0.08861539,0.0,0.009846155,0.016410258,0.02297436,0.02297436,0.02297436,0.029538464,0.09189744,0.13784617,0.14441027,0.10502565,0.23958977,0.23302566,0.20020515,0.24943592,0.48246157,0.3708718,0.4004103,0.4201026,0.36430773,0.23302566,0.17723078,0.118153855,0.07548718,0.052512825,0.026256412,0.016410258,0.6695385,1.142154,0.9747693,0.08205129,0.04594872,0.036102567,0.055794876,0.08861539,0.0951795,0.18707694,0.15753847,0.1148718,0.13128206,0.23958977,0.4660513,0.26584616,0.07876924,0.07548718,0.16738462,0.23630771,0.18051283,0.101743594,0.049230773,0.01969231,0.03938462,0.128,0.24287182,0.30194873,0.17394873,0.14112821,0.1148718,0.06564103,0.01969231,0.072205134,0.0951795,0.059076928,0.02297436,0.016410258,0.02297436,0.029538464,0.026256412,0.036102567,0.06564103,0.1148718,0.049230773,0.01969231,0.009846155,0.006564103,0.0,0.013128206,0.013128206,0.006564103,0.0,0.0,0.0032820515,0.006564103,0.006564103,0.0,0.0,0.0,0.0,0.0032820515,0.02297436,0.07876924,0.13784617,0.17394873,0.16410258,0.13128206,0.15097436,0.08205129,0.032820515,0.006564103,0.013128206,0.06564103,0.03938462,0.108307704,0.128,0.07548718,0.055794876,0.009846155,0.026256412,0.026256412,0.0,0.0,0.0,0.0,0.006564103,0.032820515,0.09189744,0.08205129,0.7089231,0.7417436,0.15097436,0.08533334,0.108307704,0.2231795,0.29538465,0.3052308,0.37415388,0.48246157,0.25928208,0.09189744,0.09189744,0.072205134,0.06235898,0.128,0.14112821,0.072205134,0.006564103,0.0,0.0,0.013128206,0.04594872,0.08205129,0.108307704,0.04594872,0.055794876,0.12471796,0.072205134,0.032820515,0.013128206,0.013128206,0.026256412,0.026256412,0.006564103,0.0,0.0,0.0,0.0,0.02297436,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.01969231,0.013128206,0.009846155,0.016410258,0.016410258,0.0032820515,0.0032820515,0.006564103,0.0032820515,0.0,0.0032820515,0.02297436,0.036102567,0.049230773,0.09189744,0.19692309,0.3708718,0.5021539,0.53825647,0.48902568,0.39056414,0.29538465,0.18707694,0.08205129,0.04594872,0.12471796,0.256,0.5021539,0.88943595,1.3981539,1.4539489,1.1881026,0.81394875,0.46276927,0.20676924,0.13784617,0.14112821,0.256,0.4660513,0.7187693,0.761436,0.761436,0.7581539,0.7450257,0.67282057,0.61374366,0.5940513,0.60389745,0.6301539,0.6695385,0.65312827,0.6104616,0.5874872,0.6170257,0.7318975,0.7122052,0.6629744,0.7975385,1.3981539,2.7963078,2.03159,1.4178462,1.0994873,1.1027694,1.3259488,1.2996924,1.3653334,1.5031796,1.5458462,1.1848207,0.92553854,0.8992821,1.0272821,1.1848207,1.1946667,1.020718,0.86317956,0.7089231,0.571077,0.48902568,0.51856416,0.46276927,0.43323082,0.4660513,0.512,0.5152821,0.571077,0.64000005,0.7122052,0.7975385,0.8369231,0.8992821,0.9682052,1.0338463,1.083077,0.955077,0.8763078,0.74830776,0.56123084,0.39384618,0.39712822,0.4135385,0.4201026,0.41025645,0.39384618,0.38728207,0.3117949,0.27241027,0.28225642,0.24943592,0.20020515,0.21989745,0.30194873,0.41682056,0.49230772,0.5349744,0.61374366,0.6170257,0.53825647,0.4397949,0.43323082,0.37415388,0.30194873,0.24943592,0.22646156,0.21661541,0.190359,0.15753847,0.13456412,0.128,0.13456412,0.17723078,0.23302566,0.27569234,0.26584616,0.26256412,0.21989745,0.20676924,0.23302566,0.23302566,0.2231795,0.27569234,0.34789747,0.41682056,0.46276927,0.45620516,0.37743592,0.3249231,0.33805132,0.38728207,0.4135385,0.46933338,0.5152821,0.512,0.43323082,0.34789747,0.3511795,0.38400003,0.4135385,0.4266667,0.48246157,0.5415385,0.5940513,0.5907693,0.46933338,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.052512825,0.03938462,0.013128206,0.0032820515,0.013128206,0.101743594,0.052512825,0.009846155,0.026256412,0.055794876,0.055794876,0.06235898,0.049230773,0.029538464,0.03938462,0.02297436,0.02297436,0.059076928,0.12143591,0.15425642,0.055794876,0.12471796,0.28882053,0.5546667,1.0075898,1.1749744,0.827077,0.8467693,1.3423591,1.6475899,1.9922053,2.5895386,3.761231,5.8420515,9.16677,9.954462,10.893129,12.356924,13.98154,14.674052,14.322873,14.795488,16.889437,20.555489,24.874668,24.336412,24.57272,23.657028,21.316925,18.934155,19.5479,20.23713,20.384823,20.657232,22.99077,24.106668,27.181952,29.630362,29.945438,27.687387,24.159182,21.313643,19.93518,19.99754,20.683489,18.12677,17.332514,16.8599,16.57436,17.64759,21.077335,22.22277,22.951385,23.840822,24.198566,22.872618,20.568617,18.120207,16.692514,17.75918,19.879387,20.886976,20.906668,20.46359,20.46031,22.029129,24.06072,24.057438,22.340925,22.032412,23.138464,24.201847,25.984001,27.339489,25.238976,28.547285,30.61826,31.753849,31.61272,29.210258,25.59672,24.280617,22.738052,19.892515,16.131283,14.454155,11.385437,10.459898,11.74318,11.82195,10.824206,11.346052,11.772718,11.785847,12.3766165,12.501334,13.433437,9.488411,2.8422565,3.5249233,5.8125134,7.0859494,5.8518977,3.8137438,5.874872,6.6625648,6.688821,6.6067696,6.9382567,8.044309,19.15077,19.551182,14.628103,11.152411,17.27672,23.46995,16.918976,10.157949,11.23118,23.702976,18.136618,14.7331295,9.429334,5.2053337,12.091078,15.786668,11.395283,5.8223596,3.5446157,6.6002054,3.9351797,1.847795,0.8467693,0.96492314,1.7624617,3.9318976,3.5938463,2.7273848,1.972513,0.6301539,0.7187693,1.0469744,1.4769232,1.8642052,2.041436,2.4451284,2.1891284,1.3981539,0.96492314,2.5665643,3.3772311,1.5721027,0.53825647,1.2077949,2.0611284,3.9023592,3.045744,1.339077,0.108307704,0.13128206,0.380718,1.4802053,1.6278975,0.9124103,1.3128207,0.6268718,0.90584624,1.083077,0.78769237,0.35446155,0.56123084,0.5218462,0.46933338,0.56123084,0.88615394,1.086359,1.8018463,2.1070771,1.9823592,2.3269746,3.82359,3.8564105,3.4034874,2.7995899,1.7362052,2.8455386,2.1234872,1.0502565,0.6071795,1.276718,3.5216413,2.9604106,1.8576412,1.339077,1.3817437,2.0676925,2.0775387,2.6912823,3.7448208,3.636513,4.7983594,6.048821,6.692103,7.250052,9.462154,9.248821,10.371283,12.199386,13.692719,13.420309,18.14318,16.617027,15.474873,14.982565,9.019077,8.743385,13.019898,20.197744,29.764925,42.371284,116.79508,145.24391,147.85313,132.3717,94.175186,54.596928,46.194874,53.533543,62.477135,60.192825,43.152412,30.713438,26.029951,28.70154,34.773335,37.376003,38.915283,36.66708,34.89149,44.82298,30.155489,20.76554,19.459284,24.362669,28.92472,12.534155,8.425026,9.084719,10.079181,10.033232,9.878975,8.786052,8.067283,8.726975,11.464206,14.467283,14.792206,22.33108,29.801027,12.763899,14.549335,17.696821,16.626873,12.911591,15.274668,12.560411,12.550565,11.858052,10.410667,11.457642,12.583385,9.521232,7.450257,7.6668725,7.581539,5.979898,4.4012313,6.7610264,12.035283,14.25395,10.256411,6.619898,5.4875903,6.3606157,6.124308,9.580308,10.630565,9.494975,7.430565,6.7249236,4.713026,6.0356927,6.9152827,6.2129235,5.425231,5.8190775,4.9526157,4.1583595,3.5905645,2.2121027,2.3040001,4.4307694,8.080411,10.167795,5.037949,4.2174363,6.747898,7.762052,6.0685134,4.1517954,5.3136415,5.356308,5.4153852,5.756718,5.756718,5.901129,5.7107697,4.7360005,3.4034874,3.006359,4.9427695,5.61559,4.972308,3.4166157,1.8346668,0.9616411,0.8205129,1.1618463,1.4441026,0.83035904,1.5688206,0.955077,0.26912823,0.029538464,0.0032820515,0.026256412,0.029538464,0.026256412,0.026256412,0.032820515,0.01969231,0.052512825,0.09189744,0.12471796,0.18051283,0.18707694,0.16082053,0.13456412,0.17066668,0.37743592,0.37415388,0.39384618,0.34789747,0.26256412,0.27569234,0.26584616,0.17723078,0.09189744,0.03938462,0.009846155,0.02297436,0.12143591,0.21989745,0.2297436,0.055794876,0.055794876,0.049230773,0.032820515,0.032820515,0.108307704,0.25928208,0.26584616,0.2100513,0.16410258,0.18051283,0.61374366,0.36430773,0.108307704,0.06564103,0.029538464,0.13456412,0.14441027,0.11158975,0.06235898,0.009846155,0.0032820515,0.0,0.049230773,0.128,0.14769232,0.068923086,0.032820515,0.01969231,0.03938462,0.14441027,0.21333335,0.16082053,0.09189744,0.06235898,0.072205134,0.07876924,0.055794876,0.059076928,0.118153855,0.2231795,0.11158975,0.052512825,0.02297436,0.006564103,0.0032820515,0.009846155,0.0032820515,0.0,0.0,0.0,0.009846155,0.0032820515,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0,0.009846155,0.052512825,0.08205129,0.14441027,0.14112821,0.07876924,0.068923086,0.08205129,0.052512825,0.01969231,0.01969231,0.072205134,0.02297436,0.04266667,0.101743594,0.14769232,0.108307704,0.026256412,0.0032820515,0.0,0.009846155,0.04266667,0.01969231,0.009846155,0.0032820515,0.0,0.0,0.013128206,0.029538464,0.13456412,0.24615386,0.101743594,0.04594872,0.02297436,0.029538464,0.08205129,0.23630771,0.42994875,0.22646156,0.049230773,0.029538464,0.0,0.055794876,0.18707694,0.27241027,0.2297436,0.026256412,0.009846155,0.0032820515,0.0,0.0,0.0,0.009846155,0.0032820515,0.01969231,0.06564103,0.15097436,0.15425642,0.20348719,0.18379489,0.09189744,0.052512825,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01969231,0.026256412,0.02297436,0.016410258,0.016410258,0.0032820515,0.006564103,0.013128206,0.013128206,0.0032820515,0.009846155,0.0032820515,0.0,0.006564103,0.036102567,0.055794876,0.13456412,0.27241027,0.41682056,0.47917953,0.41682056,0.380718,0.28882053,0.14769232,0.055794876,0.07548718,0.14441027,0.35774362,0.7318975,1.1979488,1.5130258,1.3587693,1.0404103,0.7187693,0.38728207,0.24615386,0.20020515,0.2231795,0.30194873,0.44964105,0.6498462,0.74830776,0.8041026,0.8172308,0.7417436,0.6892308,0.6629744,0.6432821,0.636718,0.65969235,0.63343596,0.63343596,0.61374366,0.6104616,0.72861546,0.67282057,0.42994875,0.34133336,0.90256417,2.7667694,1.8018463,1.3095386,1.1093334,1.0994873,1.2537436,1.3751796,1.1158975,1.1618463,1.4802053,1.3226668,0.9156924,0.8533334,0.92553854,1.0633847,1.3226668,1.2242053,0.9878975,0.8008206,0.7056411,0.5907693,0.62030774,0.55794877,0.508718,0.512,0.5513847,0.51856416,0.53825647,0.58092314,0.6170257,0.62030774,0.7450257,0.8402052,0.90584624,0.98461545,1.142154,1.0043077,0.8566154,0.7089231,0.5546667,0.3708718,0.3117949,0.32820517,0.39056414,0.44307697,0.4135385,0.39712822,0.36102566,0.34789747,0.3511795,0.30194873,0.24615386,0.24615386,0.3249231,0.42994875,0.42994875,0.47589746,0.55794877,0.5973334,0.56451285,0.49230772,0.48902568,0.4135385,0.32820517,0.27569234,0.28225642,0.23302566,0.17723078,0.15425642,0.16082053,0.15097436,0.17066668,0.23958977,0.30194873,0.3249231,0.2855385,0.30194873,0.2231795,0.17723078,0.190359,0.21661541,0.25271797,0.30851284,0.35446155,0.37743592,0.3708718,0.37743592,0.36758977,0.35774362,0.34789747,0.318359,0.3446154,0.43651286,0.46276927,0.4135385,0.39056414,0.3446154,0.28225642,0.256,0.28225642,0.34133336,0.4201026,0.41682056,0.42994875,0.4594872,0.42994875,0.0,0.0,0.0,0.0,0.013128206,0.06235898,0.26912823,0.19364104,0.06564103,0.0,0.0,0.013128206,0.016410258,0.04594872,0.09189744,0.09189744,0.055794876,0.06564103,0.052512825,0.03938462,0.13784617,0.052512825,0.013128206,0.006564103,0.02297436,0.04594872,0.032820515,0.0951795,0.18707694,0.45620516,1.2504616,1.2635899,0.9911796,0.9419488,1.1716924,1.2832822,1.6344616,2.3729234,4.650667,7.837539,9.521232,9.117539,9.163487,10.374565,12.658873,15.136822,14.660924,13.561437,14.027489,16.269129,18.54031,17.207796,19.72513,20.768822,19.203283,18.067694,17.529438,18.346668,17.920002,16.8599,18.996513,19.606976,20.62113,22.098053,23.637335,24.369232,18.14318,14.683899,13.522053,13.686155,13.686155,13.945437,15.097437,17.155283,19.636515,21.589334,22.176823,22.160412,23.08595,25.186464,27.359182,22.94154,20.644104,19.685745,19.685745,20.676924,20.54236,20.178053,20.115694,20.76554,22.400002,23.899899,28.626053,31.110567,29.587694,26.000412,24.891079,23.752207,22.787283,22.294975,22.675694,25.347284,26.601028,26.692924,25.721437,23.620924,24.01149,25.409643,23.840822,19.941746,18.950565,19.59713,16.400412,15.734155,18.084105,18.034874,9.6754875,9.724719,12.1238985,12.1928215,6.6395903,5.0149746,4.644103,3.6496413,2.878359,5.904411,12.849232,17.920002,13.334975,3.3247182,4.1058464,4.824616,9.015796,14.818462,19.016207,17.027283,27.208208,21.743591,13.778052,9.462154,7.9491286,9.964309,7.512616,4.896821,6.308103,15.793232,10.518975,7.4174366,4.1878977,1.8609232,4.7917953,8.477539,6.3343596,3.2984617,2.156308,3.5249233,2.3040001,1.2307693,0.8402052,1.1027694,1.4178462,1.332513,1.6771283,2.228513,2.3991797,1.2504616,0.33476925,0.8566154,1.8149745,2.3958976,1.9692309,2.176,3.3444104,2.8488207,0.8336411,0.19692309,0.24615386,0.14112821,0.24287182,0.62030774,1.024,1.4506668,1.079795,0.56123084,0.27897438,0.3511795,0.86317956,1.9331284,2.0151796,1.2406155,1.4342566,0.8369231,1.0075898,1.0371283,0.7450257,0.67282057,0.6826667,0.44964105,0.25271797,0.43323082,1.3718976,1.3981539,1.404718,1.1651284,1.522872,4.378257,5.5991797,5.1922054,4.588308,3.9220517,2.028308,3.761231,2.3827693,0.85005134,0.34789747,0.27569234,2.0808206,3.0720003,2.7142565,1.4933335,0.9321026,0.5415385,0.37743592,1.7165129,4.457026,7.141744,8.362667,6.3606157,4.059898,3.3936412,5.3103595,9.32759,12.701539,15.287796,15.589745,10.758565,13.138052,13.413745,11.690667,9.494975,9.750975,9.199591,9.521232,20.552206,43.78913,72.402054,113.06339,128.50545,125.30544,109.29888,85.55652,54.564106,55.886772,69.07078,79.442055,78.12267,63.86544,45.30544,32.213337,28.655592,32.99118,31.465029,26.614157,23.532309,22.764309,20.312616,13.328411,8.900924,11.040821,20.808207,36.28636,14.546052,8.461129,12.153437,17.480206,14.037334,11.316514,9.426052,7.069539,6.5936418,13.991385,13.479385,12.3536415,17.030565,22.518156,12.435693,15.501129,25.265232,26.581335,18.838976,15.944206,13.761642,13.515489,12.442257,12.081232,18.294155,20.102566,12.770463,8.310155,10.240001,13.610668,10.692924,5.1954875,5.2480006,10.738873,13.289026,6.820103,6.163693,6.377026,5.796103,6.0258465,8.260923,5.2480006,3.7251284,5.677949,8.362667,6.0652313,9.081436,11.529847,10.112,4.1189747,5.5007186,4.97559,4.059898,3.5052311,3.31159,1.723077,5.034667,9.6065645,11.152411,4.7458467,2.7437952,3.0687182,3.8432825,3.9417439,2.989949,5.395693,4.670359,4.1124105,4.8147697,5.6451287,6.951385,6.738052,5.366154,3.8498464,3.8596926,4.6539493,4.338872,3.3805132,2.284308,1.6016412,1.785436,1.2176411,0.827077,0.7187693,0.18379489,0.20676924,0.25928208,0.17394873,0.0032820515,0.016410258,0.03938462,0.026256412,0.009846155,0.009846155,0.04594872,0.02297436,0.016410258,0.016410258,0.0951795,0.4135385,0.3511795,0.19692309,0.13128206,0.20676924,0.36758977,0.19692309,0.26256412,0.3052308,0.27569234,0.33476925,0.67610264,0.40697438,0.15097436,0.108307704,0.04594872,0.068923086,0.11158975,0.11158975,0.07876924,0.09189744,0.10502565,0.068923086,0.032820515,0.02297436,0.06235898,0.17066668,0.190359,0.16410258,0.14441027,0.16738462,0.18051283,0.16410258,0.14769232,0.1148718,0.029538464,0.006564103,0.009846155,0.016410258,0.02297436,0.04594872,0.02297436,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.032820515,0.16738462,0.21661541,0.24615386,0.25271797,0.21989745,0.12143591,0.098461546,0.08205129,0.08205129,0.101743594,0.13784617,0.11158975,0.068923086,0.04594872,0.03938462,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.016410258,0.006564103,0.0,0.0032820515,0.016410258,0.026256412,0.03938462,0.04594872,0.04594872,0.04594872,0.059076928,0.04266667,0.029538464,0.02297436,0.0,0.0,0.0,0.0,0.0,0.0,0.02297436,0.013128206,0.0,0.04266667,0.21333335,0.10502565,0.049230773,0.01969231,0.0,0.0,0.02297436,0.013128206,0.0,0.0032820515,0.016410258,0.026256412,0.029538464,0.055794876,0.08861539,0.07548718,0.12471796,0.118153855,0.08861539,0.049230773,0.0,0.036102567,0.04594872,0.27241027,0.5021539,0.07548718,0.03938462,0.013128206,0.0,0.0,0.0,0.0,0.0,0.09189744,0.2986667,0.58092314,0.64000005,0.9321026,0.85005134,0.380718,0.07548718,0.016410258,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.04594872,0.052512825,0.016410258,0.016410258,0.0032820515,0.0,0.006564103,0.016410258,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.04594872,0.13784617,0.27241027,0.44307697,0.380718,0.40369233,0.37743592,0.26256412,0.09189744,0.055794876,0.101743594,0.23630771,0.5021539,0.9911796,1.1979488,1.214359,1.1158975,0.92553854,0.5940513,0.37415388,0.26584616,0.2297436,0.27897438,0.47261542,0.5940513,0.65312827,0.7089231,0.79097444,0.8992821,0.72861546,0.6235898,0.5874872,0.5874872,0.5481026,0.574359,0.5973334,0.5973334,0.6071795,0.7187693,0.7778462,0.49230772,0.28882053,0.48574364,1.2668719,0.7778462,0.7187693,0.9878975,1.3653334,1.5097437,1.3751796,1.142154,0.98133343,0.9911796,1.1749744,0.8566154,0.64000005,0.4955898,0.49230772,0.80738467,1.0043077,0.76800007,0.6892308,0.81066674,0.64000005,0.6892308,0.6826667,0.58092314,0.42994875,0.380718,0.40697438,0.44964105,0.5152821,0.571077,0.5349744,0.5349744,0.65312827,0.84348726,1.0075898,1.0075898,1.0075898,0.90584624,0.72861546,0.5284103,0.380718,0.3314872,0.33805132,0.40697438,0.47589746,0.4266667,0.34133336,0.33805132,0.3249231,0.28882053,0.28882053,0.3511795,0.36758977,0.446359,0.57764107,0.6268718,0.56451285,0.5677949,0.5874872,0.56451285,0.44307697,0.3314872,0.26912823,0.23302566,0.2231795,0.25928208,0.24615386,0.20676924,0.19692309,0.21333335,0.21333335,0.24943592,0.3314872,0.40697438,0.4201026,0.33476925,0.36102566,0.29210258,0.24287182,0.23958977,0.2297436,0.26584616,0.32164106,0.3314872,0.30851284,0.32164106,0.3708718,0.39056414,0.41025645,0.4135385,0.36758977,0.3052308,0.27241027,0.25928208,0.28225642,0.36758977,0.47589746,0.40369233,0.34133336,0.35446155,0.36758977,0.36758977,0.32820517,0.3117949,0.3314872,0.380718,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.190359,0.1148718,0.01969231,0.0,0.0,0.06235898,0.04594872,0.02297436,0.029538464,0.07876924,0.052512825,0.08533334,0.07876924,0.029538464,0.03938462,0.02297436,0.006564103,0.0,0.006564103,0.02297436,0.01969231,0.10502565,0.2986667,0.6104616,1.0305642,1.2570257,1.1651284,1.0765129,1.1060513,1.148718,2.359795,4.069744,5.7009234,6.948103,7.765334,7.506052,7.6931286,9.501539,12.2617445,13.453129,10.866873,10.985026,12.668719,14.670771,15.622565,16.636719,15.803078,15.507693,16.233027,16.551386,15.304206,15.363283,16.150976,17.946259,21.891283,23.817848,23.506054,22.73149,22.317951,22.121027,19.666052,17.778873,16.482462,15.954053,16.518566,16.666258,18.674873,20.329027,21.523693,24.228104,25.38995,26.049643,27.040823,27.602053,25.380104,21.520412,20.178053,19.18031,18.336823,19.442873,20.98872,22.537848,23.913027,24.82872,24.900925,26.072617,28.347078,28.727797,26.791388,24.694157,22.111181,21.891283,22.104616,22.442669,24.237951,26.676516,27.030977,26.318771,25.081438,23.351797,22.278566,20.424206,18.743795,18.31713,20.355284,22.741335,21.287386,20.552206,22.629745,27.142567,20.214155,15.402668,12.015591,9.179898,5.832206,3.6135387,6.485334,8.874667,8.818872,7.9786673,11.096616,14.933334,12.324103,4.6244106,1.6771283,2.5895386,3.8728209,6.1505647,8.503796,8.448001,19.488823,18.806156,12.4685135,6.2030773,5.421949,5.5926156,3.7382567,2.6683078,3.7415388,6.8594875,4.7491283,3.4100516,1.9593848,0.9156924,2.2022567,2.861949,2.2383592,1.4112822,1.014154,1.2176411,0.7975385,0.6629744,0.7122052,0.86646163,1.0765129,1.2274873,1.3522053,1.3718976,1.1355898,0.41025645,0.17723078,0.48246157,0.98133343,1.270154,0.88287187,0.7778462,1.4276924,1.4605129,0.7056411,0.19692309,0.3249231,0.25271797,0.25271797,0.40369233,0.58420515,1.1257436,1.585231,2.0873847,2.166154,0.75487185,0.80738467,1.3915899,1.9593848,2.1267693,1.6672822,0.9714873,0.7220513,0.60061544,0.45292312,0.28225642,0.4201026,0.4594872,0.3511795,0.2297436,0.41025645,1.4309745,1.3915899,1.2012309,1.3915899,2.1103592,5.927385,6.8562055,6.0061545,4.33559,2.6387694,2.4681027,2.3138463,1.9265642,1.2668719,0.48246157,0.84348726,1.8904617,2.103795,1.522872,1.7591796,1.9167181,1.4834872,1.8970258,3.5380516,5.723898,6.87918,4.315898,2.3926156,3.186872,6.518154,7.381334,8.795898,9.7673855,10.010257,9.95118,9.196308,9.668923,10.916103,11.802258,10.505847,10.075898,10.755282,13.702565,23.450258,47.894978,101.5598,127.71447,121.49498,94.664215,75.60862,56.723698,57.133953,64.04923,68.77867,66.737236,63.904827,56.92062,44.626053,31.40267,27.191797,32.84349,31.041643,26.499285,21.910976,17.952822,11.684103,6.9645133,11.142565,20.197744,18.73395,9.783795,6.99077,7.0432825,7.781744,8.214975,8.989539,8.119796,6.8594875,7.204103,11.9171295,10.663385,13.728822,17.867489,18.599386,10.213744,11.989334,23.988514,23.906464,12.71795,14.6871805,22.86277,13.843694,8.4053335,13.942155,24.470976,26.01354,16.692514,9.672206,9.810052,13.6467705,11.227899,5.720616,5.3136415,9.281642,8.004924,5.179077,6.0324106,6.0061545,4.5554876,5.149539,8.533334,4.9394875,5.474462,11.444513,14.355694,8.553026,7.6701546,7.650462,6.173539,2.6322052,6.2162056,5.467898,3.9745643,4.1189747,7.059693,2.0053334,7.2336416,14.214565,15.904821,6.7216415,3.1770258,4.7491283,7.3321033,8.316719,6.6034875,5.346462,4.1878977,3.4855387,3.889231,6.340924,6.954667,5.733744,4.2994876,3.4166157,2.9702566,3.373949,3.1442053,2.8980515,2.8750772,2.9440002,1.9265642,1.1618463,1.0043077,1.2800001,1.270154,0.33805132,0.13456412,0.09189744,0.0,0.0032820515,0.14441027,0.118153855,0.049230773,0.07548718,0.3249231,0.068923086,0.0032820515,0.006564103,0.029538464,0.0951795,0.190359,0.16410258,0.13456412,0.190359,0.37743592,0.51856416,0.38728207,0.26912823,0.24943592,0.21333335,0.3117949,0.18379489,0.15097436,0.24615386,0.20348719,0.11158975,0.14769232,0.5874872,0.9714873,0.10502565,0.10502565,0.108307704,0.068923086,0.013128206,0.013128206,0.08205129,0.1148718,0.108307704,0.10502565,0.16738462,0.18051283,0.2231795,0.29210258,0.3052308,0.10502565,0.049230773,0.016410258,0.0032820515,0.0032820515,0.009846155,0.013128206,0.01969231,0.013128206,0.0,0.0,0.0,0.0,0.0,0.013128206,0.059076928,0.08861539,0.15097436,0.21989745,0.25271797,0.19692309,0.24943592,0.2100513,0.13456412,0.08205129,0.08861539,0.055794876,0.029538464,0.016410258,0.009846155,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.03938462,0.08861539,0.13456412,0.14441027,0.108307704,0.052512825,0.026256412,0.01969231,0.026256412,0.036102567,0.04594872,0.068923086,0.055794876,0.029538464,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.013128206,0.04266667,0.16410258,0.17066668,0.12471796,0.059076928,0.013128206,0.013128206,0.06564103,0.09189744,0.08205129,0.06235898,0.06564103,0.04594872,0.029538464,0.032820515,0.052512825,0.03938462,0.03938462,0.036102567,0.029538464,0.02297436,0.013128206,0.009846155,0.016410258,0.06235898,0.101743594,0.016410258,0.026256412,0.01969231,0.006564103,0.0032820515,0.013128206,0.0032820515,0.0,0.01969231,0.068923086,0.16410258,0.20676924,0.49230772,0.5973334,0.43323082,0.23630771,0.37743592,0.16738462,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.009846155,0.016410258,0.06564103,0.013128206,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.06564103,0.16082053,0.23630771,0.37743592,0.40697438,0.36758977,0.29538465,0.20020515,0.08533334,0.098461546,0.18707694,0.37415388,0.73517954,1.1093334,1.1651284,1.1618463,1.2373334,1.4244103,0.8041026,0.43323082,0.2986667,0.3446154,0.4594872,0.54482055,0.62030774,0.764718,0.88943595,0.764718,0.54482055,0.47917953,0.508718,0.57764107,0.5973334,0.61374366,0.65641034,0.67610264,0.65641034,0.62030774,0.6695385,0.57764107,0.43651286,0.3511795,0.44964105,0.4004103,0.508718,0.80738467,1.2373334,1.657436,1.522872,1.2964103,1.1158975,1.0502565,1.0765129,0.96492314,0.9321026,0.8402052,0.6826667,0.60061544,0.8467693,0.86317956,0.8960001,1.0043077,1.0666667,1.0305642,0.9485129,0.81066674,0.6465641,0.5415385,0.4660513,0.4201026,0.4135385,0.42994875,0.4135385,0.46933338,0.5513847,0.63343596,0.7089231,0.78769237,0.78769237,0.7450257,0.6662565,0.5513847,0.39384618,0.31507695,0.2855385,0.32164106,0.40697438,0.47589746,0.4201026,0.42338464,0.41682056,0.3708718,0.30194873,0.31507695,0.35446155,0.39384618,0.45292312,0.5874872,0.6170257,0.5677949,0.5481026,0.5513847,0.4660513,0.33805132,0.3117949,0.29538465,0.25928208,0.24615386,0.20676924,0.16738462,0.14769232,0.16738462,0.22646156,0.3314872,0.36430773,0.39712822,0.43651286,0.41025645,0.35446155,0.3117949,0.2986667,0.29538465,0.25271797,0.25928208,0.30194873,0.32164106,0.32820517,0.3708718,0.40697438,0.38400003,0.3708718,0.43323082,0.5973334,0.4594872,0.3249231,0.24943592,0.23302566,0.23302566,0.32164106,0.36758977,0.39056414,0.38400003,0.318359,0.28882053,0.25271797,0.26256412,0.3446154,0.49230772,0.0,0.0,0.0,0.0,0.0,0.0,0.14769232,0.07876924,0.0032820515,0.016410258,0.08205129,0.068923086,0.032820515,0.009846155,0.026256412,0.0951795,0.08533334,0.08861539,0.13456412,0.18379489,0.14441027,0.03938462,0.013128206,0.006564103,0.0,0.006564103,0.013128206,0.101743594,0.23630771,0.39056414,0.53825647,0.7515898,0.8566154,0.95835906,1.1126155,1.3423591,2.7995899,4.647385,5.868308,6.2588725,6.409847,6.373744,7.5388722,10.535385,13.984821,14.513232,10.427077,9.672206,11.011283,12.954257,13.728822,13.571283,12.435693,12.737642,14.240822,14.060308,13.538463,15.852309,19.38708,23.007181,26.04636,27.615181,26.535387,24.904207,23.968822,24.14277,22.790565,20.427488,17.972515,16.722052,18.353231,19.478975,22.777437,25.380104,26.896412,29.410463,31.097439,30.099695,27.733335,24.950155,22.33436,20.434053,20.158361,19.498669,19.052309,22.019283,23.315695,24.103386,25.163488,26.354874,26.607592,27.776003,28.534157,27.720207,25.744411,24.615387,24.086977,23.666874,23.5159,23.670156,24.024618,25.173336,24.526772,23.318975,21.671387,18.615797,16.22318,14.060308,13.584412,15.031796,17.411283,16.905848,15.238565,17.824821,24.22154,28.137028,27.529848,22.30154,16.101746,11.562668,10.289231,14.506668,16.528412,13.929027,9.357129,10.522257,9.124104,8.530052,8.080411,6.5444107,2.1202054,1.6213335,1.7362052,2.5731285,3.6036925,3.6660516,8.277334,10.230155,7.8145647,3.31159,3.006359,2.6322052,1.7952822,1.4408206,1.7887181,2.3335385,1.7263591,1.5556924,1.1027694,0.5973334,1.2373334,0.9189744,0.6629744,0.52512825,0.45292312,0.29210258,0.20348719,0.49887183,0.7581539,0.78769237,0.5973334,0.93866676,1.083077,1.2373334,1.5425643,2.0841026,2.1103592,1.4211283,0.95835906,1.1224617,1.7920002,1.1552821,1.1684103,1.1355898,0.8533334,0.6104616,0.63343596,0.508718,0.34133336,0.3117949,0.67282057,1.5130258,2.3072822,3.2164104,3.69559,2.5304618,1.8084104,1.654154,1.8018463,1.9232821,1.6147693,1.0699488,0.6432821,0.446359,0.37743592,0.14769232,0.23630771,0.3249231,0.318359,0.22646156,0.15097436,0.9124103,1.8379488,2.5698464,2.7766156,2.1464617,5.47118,5.87159,4.9460516,3.6529233,2.297436,1.9068719,2.7700515,2.9440002,1.9856411,0.955077,0.65641034,1.4342566,1.6443079,1.2373334,1.7493335,2.172718,2.1464617,2.3040001,3.0358977,4.4832826,5.72718,4.141949,3.3575387,4.516103,6.2523084,5.5565133,5.618872,5.674667,5.664821,6.245744,6.47877,6.5247183,8.054154,10.463181,10.889847,17.503181,12.603078,9.032206,14.099693,29.607388,88.19529,130.94073,127.829346,89.46873,67.09498,52.916515,50.04144,51.77108,53.950363,54.97108,53.3399,51.57744,45.748516,35.67262,24.917336,28.813131,27.395285,21.648413,14.736411,11.989334,12.6063595,13.042872,13.197129,12.937847,12.091078,10.522257,9.964309,9.140513,7.788308,6.6494365,7.1548724,6.9152827,7.13518,8.208411,9.7214365,7.4469748,16.387283,19.856411,14.647796,11.024411,9.905231,13.948719,14.247386,10.975181,13.384206,25.521233,13.978257,6.491898,11.497026,18.133335,23.601233,16.521847,8.513641,6.47877,12.586668,10.8767185,7.0531287,6.242462,8.4972315,8.79918,5.0576415,6.373744,6.8955903,5.211898,4.352,8.349539,4.8016415,5.2315903,11.894155,17.80513,7.817847,4.5390773,4.128821,3.945026,2.5600002,5.865026,4.788513,3.4756925,4.07959,6.76759,2.5764105,9.754257,18.520617,20.345438,7.9491286,4.342154,5.943795,7.9130263,8.086975,6.9677954,5.681231,5.405539,4.5522056,3.6660516,5.4153852,6.055385,5.1856413,4.0467696,3.1671798,2.3696413,2.4713848,2.349949,2.1530259,2.048,2.1989746,1.8937438,1.3620514,1.1158975,1.214359,1.2832822,0.43651286,0.16738462,0.098461546,0.059076928,0.108307704,0.27241027,0.14769232,0.06235898,0.14769232,0.34133336,0.10502565,0.01969231,0.01969231,0.04594872,0.016410258,0.098461546,0.13456412,0.16082053,0.20676924,0.30851284,0.5349744,0.47589746,0.4135385,0.4266667,0.36758977,0.32164106,0.15097436,0.08205129,0.16410258,0.24287182,0.15753847,0.18379489,0.5415385,0.8533334,0.17066668,0.128,0.118153855,0.098461546,0.052512825,0.01969231,0.072205134,0.1148718,0.1148718,0.10502565,0.18707694,0.30851284,0.29538465,0.26584616,0.23958977,0.13128206,0.08533334,0.036102567,0.006564103,0.0,0.0,0.0032820515,0.009846155,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.02297436,0.03938462,0.08533334,0.13456412,0.16738462,0.17723078,0.24287182,0.19692309,0.12143591,0.07876924,0.08533334,0.06235898,0.032820515,0.009846155,0.0,0.006564103,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.01969231,0.049230773,0.21333335,0.3511795,0.36430773,0.22646156,0.101743594,0.036102567,0.016410258,0.01969231,0.01969231,0.036102567,0.032820515,0.016410258,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.016410258,0.029538464,0.07876924,0.08533334,0.08205129,0.06564103,0.049230773,0.07876924,0.15425642,0.16082053,0.13128206,0.12471796,0.20348719,0.36430773,0.18707694,0.036102567,0.029538464,0.03938462,0.48902568,0.24943592,0.013128206,0.006564103,0.016410258,0.009846155,0.006564103,0.006564103,0.009846155,0.01969231,0.04266667,0.029538464,0.01969231,0.026256412,0.02297436,0.0032820515,0.006564103,0.006564103,0.006564103,0.032820515,0.03938462,0.15097436,0.21661541,0.28225642,0.5940513,0.51856416,0.2100513,0.01969231,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.029538464,0.006564103,0.0,0.0032820515,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01969231,0.06564103,0.13784617,0.25271797,0.33805132,0.36102566,0.32164106,0.24615386,0.128,0.09189744,0.12143591,0.24615386,0.5152821,0.79097444,0.9288206,1.020718,1.2012309,1.6410258,1.1191796,0.6071795,0.32164106,0.318359,0.4660513,0.5415385,0.6235898,0.6826667,0.6859488,0.61374366,0.48246157,0.42338464,0.44307697,0.5218462,0.60061544,0.57764107,0.6268718,0.67282057,0.6695385,0.60389745,0.6170257,0.571077,0.49887183,0.42994875,0.36430773,0.38728207,0.48574364,0.7450257,1.1126155,1.4112822,1.4867693,1.2340513,1.0404103,1.014154,0.97805136,1.0436924,1.0469744,1.0502565,1.0469744,0.97805136,0.92225647,0.9288206,1.1126155,1.3718976,1.4211283,1.1913847,1.1027694,1.0633847,0.9944616,0.827077,0.5907693,0.46276927,0.4135385,0.39384618,0.3446154,0.40369233,0.47261542,0.51856416,0.54482055,0.60389745,0.6268718,0.6301539,0.6104616,0.54482055,0.4135385,0.36758977,0.34133336,0.35446155,0.40369233,0.48902568,0.4397949,0.42994875,0.4004103,0.33805132,0.25928208,0.3117949,0.40369233,0.48246157,0.5415385,0.5973334,0.6104616,0.55794877,0.5349744,0.52512825,0.41025645,0.34789747,0.36102566,0.34133336,0.27569234,0.24287182,0.23302566,0.20676924,0.17723078,0.18051283,0.27569234,0.3446154,0.36102566,0.380718,0.41682056,0.4266667,0.36102566,0.37743592,0.4135385,0.42338464,0.36102566,0.36758977,0.38400003,0.39384618,0.39056414,0.3708718,0.41025645,0.38400003,0.3708718,0.42338464,0.5546667,0.45620516,0.3708718,0.3052308,0.25271797,0.19692309,0.23302566,0.29210258,0.32820517,0.3314872,0.3052308,0.29210258,0.26912823,0.28882053,0.36758977,0.508718,0.0,0.0,0.0,0.0,0.0,0.0,0.08205129,0.03938462,0.0032820515,0.026256412,0.11158975,0.118153855,0.049230773,0.02297436,0.068923086,0.11158975,0.07876924,0.059076928,0.108307704,0.19692309,0.20348719,0.06235898,0.02297436,0.01969231,0.01969231,0.02297436,0.072205134,0.14441027,0.17723078,0.17066668,0.19692309,0.46276927,0.7056411,0.9288206,1.1782565,1.5425643,2.802872,4.0303593,4.969026,5.4449234,5.3760004,5.930667,8.454565,11.894155,14.621539,14.427898,10.118565,8.677744,9.892103,12.465232,14.040616,12.793437,11.720206,12.100924,13.692719,14.736411,17.365335,22.547693,27.241028,29.93231,30.63795,31.366566,29.479387,26.801233,24.615387,23.660309,23.030155,21.704206,20.453745,20.217438,22.081642,23.716105,27.720207,30.67077,31.586464,31.924515,31.415798,28.14031,24.14277,21.257847,21.113438,21.35631,22.101336,21.743591,21.428514,25.03877,25.668924,25.928207,26.7159,27.782566,27.743181,28.143593,27.789131,26.79795,25.88554,26.377848,25.028925,24.241232,23.538874,22.672413,21.59918,22.360617,20.260103,18.566566,17.54913,14.477129,12.143591,10.771693,10.939077,12.301129,13.564719,12.150155,10.469745,15.543797,23.978668,21.973335,22.921848,20.847591,16.833643,13.315283,14.099693,23.335386,28.09436,23.942566,15.530668,16.594053,13.4859495,8.933744,7.4371285,8.4512825,6.409847,3.006359,1.6836925,1.4539489,1.5458462,1.4145643,1.5031796,3.3280003,3.2918978,1.4276924,1.4080001,1.1027694,0.86646163,0.7384616,0.67938465,0.56451285,0.5021539,0.96492314,0.9419488,0.53825647,0.9616411,0.58420515,0.3117949,0.26912823,0.32820517,0.09189744,0.052512825,0.58420515,1.020718,1.0535386,0.7318975,1.017436,0.9944616,1.024,1.4276924,2.487795,3.442872,2.5600002,1.8543591,2.2678976,3.6890259,2.3926156,1.7755898,1.5064616,1.3357949,1.1060513,1.1552821,1.0108719,0.7384616,0.5546667,0.827077,1.7033848,2.3236926,3.1540515,3.9187696,3.5872824,2.7175386,2.2416413,1.9495386,1.7887181,1.847795,1.4080001,0.8763078,0.7187693,0.7581539,0.17066668,0.14441027,0.20020515,0.2986667,0.3511795,0.23630771,0.79425645,2.3663592,3.508513,3.5314875,2.5107694,3.761231,4.082872,3.5413337,2.484513,1.5589745,1.6771283,3.0752823,3.639795,2.7667694,1.3686155,0.8566154,1.0929232,1.1585642,0.97805136,1.332513,1.5392822,1.847795,2.7109745,3.8498464,4.2338467,5.175795,5.1922054,5.5958977,6.0980515,4.788513,3.9417439,4.325744,4.0008206,3.0162053,3.3936412,5.4153852,5.546667,6.0947695,8.093539,11.290257,20.614565,12.688411,6.76759,10.673231,20.79836,70.57724,116.864006,122.35488,90.28596,64.4398,51.51508,44.58667,42.942364,45.810875,52.34544,47.20903,45.157745,43.986053,39.161438,23.817848,26.292515,25.212719,18.763489,10.069334,7.1680007,12.360206,15.90154,13.46954,8.119796,10.308924,11.227899,11.490462,11.083488,9.750975,6.99077,6.925129,6.314667,6.0947695,6.4722056,6.944821,11.657847,16.472616,16.09518,11.789129,11.382154,8.769642,7.4797955,8.677744,11.779283,14.427898,21.888002,12.320822,5.333334,7.174565,10.748719,18.520617,15.632411,8.444718,3.8367183,9.199591,10.125129,9.028924,8.36595,8.868103,9.554052,4.7458467,7.8047185,9.9282055,8.218257,5.674667,8.402052,4.8672824,4.95918,10.236719,13.915898,5.0477953,2.8389745,3.7284105,4.8738465,4.1714873,5.4186673,3.945026,2.878359,3.7120004,6.298257,4.1124105,8.661334,15.783386,18.793028,8.461129,5.612308,5.8289237,6.6133337,6.8955903,7.066257,6.6428723,6.7183595,5.586052,3.8104618,4.2272825,5.106872,4.322462,3.2984617,2.6683078,2.2678976,2.281026,2.2055387,1.9922053,1.7985642,1.9922053,1.8707694,1.5163078,1.211077,1.0765129,1.0666667,0.65969235,0.34133336,0.16082053,0.11158975,0.13456412,0.24943592,0.12143591,0.06235898,0.15097436,0.24287182,0.0951795,0.032820515,0.04594872,0.072205134,0.009846155,0.08205129,0.18051283,0.23302566,0.24615386,0.29538465,0.55794877,0.508718,0.4201026,0.40697438,0.4397949,0.33805132,0.15425642,0.049230773,0.07548718,0.17723078,0.16082053,0.2297436,0.4004103,0.5152821,0.22646156,0.14441027,0.11158975,0.128,0.14112821,0.04266667,0.08533334,0.14112821,0.18379489,0.20348719,0.21661541,0.34789747,0.2855385,0.18379489,0.118153855,0.0951795,0.072205134,0.04266667,0.016410258,0.0,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.016410258,0.03938462,0.055794876,0.072205134,0.108307704,0.14112821,0.118153855,0.08205129,0.06235898,0.072205134,0.06564103,0.03938462,0.013128206,0.0,0.0,0.013128206,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.006564103,0.009846155,0.15425642,0.3117949,0.39712822,0.36102566,0.3249231,0.20348719,0.0951795,0.032820515,0.0,0.006564103,0.009846155,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.016410258,0.02297436,0.029538464,0.01969231,0.032820515,0.055794876,0.09189744,0.17066668,0.26256412,0.22646156,0.15753847,0.15425642,0.31507695,0.47261542,0.3117949,0.256,0.32164106,0.11158975,0.5481026,0.27897438,0.01969231,0.006564103,0.009846155,0.009846155,0.006564103,0.009846155,0.032820515,0.10502565,0.16738462,0.108307704,0.049230773,0.032820515,0.02297436,0.0032820515,0.009846155,0.013128206,0.006564103,0.009846155,0.0032820515,0.0032820515,0.009846155,0.11158975,0.49230772,0.35774362,0.15097436,0.032820515,0.02297436,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.06564103,0.13456412,0.24287182,0.3249231,0.33476925,0.27241027,0.17723078,0.098461546,0.07876924,0.15097436,0.3446154,0.5415385,0.6892308,0.8172308,1.020718,1.4539489,1.1946667,0.7384616,0.39712822,0.30851284,0.44964105,0.5218462,0.58092314,0.5677949,0.5021539,0.5021539,0.46276927,0.40369233,0.41025645,0.56123084,0.9189744,0.6662565,0.61374366,0.64000005,0.65641034,0.6301539,0.67610264,0.62030774,0.53825647,0.47917953,0.44307697,0.54482055,0.67938465,0.8566154,1.0469744,1.1848207,1.2570257,1.0601027,0.8960001,0.86646163,0.88287187,1.017436,0.99774367,1.0371283,1.142154,1.0896411,1.017436,1.1355898,1.404718,1.6082052,1.3554872,1.2635899,1.2504616,1.2668719,1.2307693,1.017436,0.8336411,0.65641034,0.5218462,0.42338464,0.3249231,0.34133336,0.38400003,0.4135385,0.4201026,0.446359,0.47261542,0.512,0.5677949,0.60389745,0.53825647,0.48902568,0.4594872,0.446359,0.446359,0.48246157,0.44307697,0.4135385,0.36430773,0.30194873,0.27241027,0.3117949,0.39384618,0.49230772,0.56451285,0.5677949,0.61374366,0.5907693,0.5513847,0.50543594,0.4266667,0.44964105,0.47589746,0.4266667,0.31507695,0.24287182,0.23630771,0.2297436,0.21333335,0.20348719,0.27569234,0.34133336,0.37415388,0.38400003,0.37743592,0.3708718,0.35446155,0.39384618,0.4397949,0.46276927,0.43323082,0.43651286,0.41682056,0.40697438,0.40369233,0.3708718,0.39056414,0.39056414,0.4135385,0.4660513,0.52512825,0.49887183,0.48246157,0.41682056,0.30194873,0.20348719,0.20348719,0.23958977,0.26256412,0.26584616,0.26256412,0.28225642,0.29538465,0.3314872,0.4004103,0.49887183,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.026256412,0.07876924,0.16082053,0.098461546,0.07548718,0.12471796,0.098461546,0.032820515,0.04266667,0.055794876,0.07548718,0.18051283,0.14112821,0.0951795,0.098461546,0.14112821,0.14112821,0.24615386,0.256,0.19364104,0.12143591,0.16082053,0.56123084,0.8336411,0.9911796,1.1323078,1.4473847,2.2219489,2.8160002,3.761231,4.772103,4.7622566,6.196513,9.524513,12.081232,12.754052,11.972924,8.644924,7.9524107,9.872411,13.220103,15.658668,15.136822,14.224411,15.159796,18.697847,24.113234,28.964106,33.22421,35.01621,34.307285,32.912415,32.006565,29.778053,27.008001,24.218258,21.661541,23.095797,24.25108,25.232412,26.177643,27.264002,28.281439,31.455181,32.994465,31.793234,29.443285,26.207182,21.96349,19.334566,19.56759,22.54113,22.948105,24.323284,24.677746,24.536617,26.93908,26.407387,26.574772,27.103182,27.359182,26.397541,25.993849,25.225847,25.219284,26.12513,27.14913,22.596926,22.475489,22.564104,21.398975,20.309336,20.12554,16.321642,13.856822,13.5778475,12.20595,10.640411,10.095591,10.039796,10.138257,10.262975,12.849232,12.964104,17.686975,23.673437,17.171694,15.179488,14.854566,13.594257,11.844924,13.111795,20.992002,29.433437,29.371078,22.321232,20.394669,19.56431,14.857847,10.804514,9.6754875,11.467488,5.5663595,2.7733335,1.529436,0.9156924,0.6498462,0.65641034,0.7811283,0.7450257,0.574359,0.636718,0.77128214,0.71548724,0.636718,0.5940513,0.5546667,0.41025645,0.9156924,0.96492314,0.574359,0.8763078,0.56123084,0.3249231,0.3446154,0.44964105,0.12143591,0.032820515,0.67610264,1.4244103,1.8281027,1.5885129,1.8642052,1.6902566,1.2340513,0.9944616,1.8018463,4.059898,3.7284105,3.2853336,3.9614363,5.733744,3.757949,2.605949,2.1431797,1.9692309,1.4145643,2.2416413,1.975795,1.4834872,1.1913847,1.086359,1.5327181,1.9265642,2.4451284,2.9735386,3.0949745,2.8521028,2.6912823,2.3302567,1.9889232,2.3762052,2.0053334,1.3357949,1.1257436,1.1552821,0.21989745,0.118153855,0.16410258,0.3314872,0.48246157,0.3708718,1.1027694,2.8192823,3.7842054,3.3805132,2.1202054,1.6968206,2.878359,3.05559,1.8773335,1.2373334,1.7558975,2.8849232,3.5741541,3.2525132,1.8346668,1.1126155,0.7318975,0.7417436,1.083077,1.5885129,0.9517949,1.0535386,3.0687182,5.6976414,5.1954875,5.149539,5.9995904,6.567385,5.756718,2.556718,2.3368206,3.8137438,3.5380516,1.7296412,2.284308,5.618872,6.3277955,5.7665644,6.232616,10.971898,16.987898,11.349334,6.9842057,9.80677,18.697847,47.829338,81.94298,97.578674,88.15919,63.980312,53.251286,44.672005,41.524517,45.42031,56.306877,48.863182,44.44554,43.139286,39.33867,21.737028,24.359386,24.12636,18.54031,9.862565,5.093744,10.020103,12.560411,11.224616,8.231385,9.494975,9.403078,9.334154,9.816616,9.931488,7.322257,7.138462,5.586052,3.7054362,3.0752823,5.8092313,18.159592,12.389745,7.79159,9.898667,10.489437,7.893334,7.3616414,9.025641,12.898462,18.865232,14.831591,9.38995,5.3005133,4.4406157,7.788308,13.817437,15.159796,10.295795,3.5905645,5.297231,10.197334,11.848206,11.286975,9.754257,8.694155,4.44718,8.63836,12.038565,11.158976,8.267488,8.214975,4.650667,5.1298466,8.792616,6.3343596,2.6847181,3.8104618,5.868308,6.5903597,5.277539,4.516103,3.0358977,2.2186668,3.511795,8.421744,6.0816417,4.673641,8.644924,14.759386,12.074668,7.755488,5.366154,5.5958977,7.4765134,8.39877,7.1876926,6.521436,5.4843082,4.096,3.308308,4.128821,2.989949,2.0020514,1.9823592,2.484513,2.537026,2.3302567,2.297436,2.5304618,2.7864618,2.038154,1.6869745,1.3850257,1.0633847,0.9353847,0.8467693,0.47917953,0.20348719,0.12143591,0.07548718,0.13128206,0.101743594,0.08533334,0.1148718,0.15425642,0.049230773,0.032820515,0.068923086,0.0951795,0.013128206,0.09189744,0.23630771,0.3117949,0.32164106,0.40697438,0.6662565,0.52512825,0.2986667,0.19692309,0.34133336,0.28225642,0.16410258,0.09189744,0.08205129,0.072205134,0.1148718,0.22646156,0.32164106,0.32820517,0.21333335,0.14441027,0.10502565,0.15425642,0.20676924,0.052512825,0.08205129,0.15097436,0.256,0.32164106,0.2231795,0.23630771,0.18379489,0.108307704,0.04594872,0.026256412,0.026256412,0.032820515,0.02297436,0.0032820515,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.013128206,0.016410258,0.036102567,0.026256412,0.03938462,0.04266667,0.032820515,0.03938462,0.04266667,0.036102567,0.01969231,0.0032820515,0.0,0.009846155,0.013128206,0.006564103,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.013128206,0.02297436,0.049230773,0.0951795,0.18051283,0.33476925,0.571077,0.5316923,0.36430773,0.17723078,0.036102567,0.006564103,0.0,0.009846155,0.026256412,0.04594872,0.009846155,0.0,0.0,0.0,0.0,0.0,0.013128206,0.026256412,0.03938462,0.049230773,0.03938462,0.029538464,0.049230773,0.11158975,0.2231795,0.3117949,0.25271797,0.16410258,0.15425642,0.33805132,0.37415388,0.4201026,0.636718,0.8041026,0.33476925,0.256,0.15425642,0.108307704,0.0951795,0.0,0.0,0.006564103,0.013128206,0.04266667,0.17066668,0.28882053,0.256,0.14441027,0.03938462,0.059076928,0.03938462,0.026256412,0.016410258,0.016410258,0.01969231,0.013128206,0.013128206,0.013128206,0.016410258,0.02297436,0.059076928,0.055794876,0.049230773,0.04266667,0.026256412,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.068923086,0.15425642,0.24615386,0.30851284,0.28225642,0.22646156,0.13784617,0.07876924,0.098461546,0.21333335,0.42994875,0.54482055,0.6662565,0.8467693,1.1191796,1.0994873,0.9124103,0.6826667,0.5021539,0.40697438,0.47917953,0.51856416,0.5218462,0.49887183,0.4594872,0.42338464,0.36758977,0.38400003,0.6071795,1.1979488,0.79097444,0.65969235,0.636718,0.64000005,0.65641034,0.7811283,0.73517954,0.60389745,0.47589746,0.43651286,0.6498462,0.9124103,1.086359,1.142154,1.1749744,0.99774367,0.9189744,0.85005134,0.80738467,0.9189744,0.97805136,0.90584624,0.90584624,0.9616411,0.85005134,0.98461545,1.2406155,1.4834872,1.5097437,1.0404103,1.270154,1.3522053,1.3915899,1.3751796,1.1684103,1.1126155,0.92553854,0.71548724,0.53825647,0.39056414,0.3249231,0.31507695,0.31507695,0.30851284,0.32164106,0.3511795,0.39384618,0.512,0.65641034,0.67610264,0.62030774,0.55794877,0.508718,0.47917953,0.45620516,0.43651286,0.4004103,0.3446154,0.30194873,0.33805132,0.3446154,0.36430773,0.41682056,0.47917953,0.5021539,0.61374366,0.63343596,0.571077,0.49230772,0.51856416,0.5677949,0.58420515,0.5284103,0.4135385,0.28882053,0.2231795,0.21333335,0.21661541,0.21333335,0.2297436,0.33476925,0.4135385,0.4266667,0.38400003,0.31507695,0.3446154,0.36102566,0.3708718,0.39712822,0.4397949,0.43651286,0.38728207,0.36430773,0.37415388,0.37743592,0.36758977,0.4004103,0.45620516,0.5152821,0.54482055,0.5907693,0.60389745,0.51856416,0.35774362,0.23302566,0.21661541,0.2297436,0.23630771,0.2231795,0.19692309,0.24615386,0.28882053,0.36430773,0.4660513,0.54482055,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01969231,0.09189744,0.01969231,0.118153855,0.18707694,0.13456412,0.0,0.013128206,0.15097436,0.19692309,0.14441027,0.2297436,0.42338464,0.3249231,0.3446154,0.50543594,0.45620516,0.5907693,0.44307697,0.26584616,0.2100513,0.32164106,0.6629744,0.8402052,0.79097444,0.65312827,0.761436,0.92225647,2.2711797,3.9417439,5.077334,4.821334,6.9710774,9.173334,9.67877,8.736821,8.592411,6.6494365,8.333129,11.264001,13.912617,15.609437,17.490053,18.966976,25.37354,37.00513,49.09949,47.57662,40.677746,33.686977,29.423592,28.212515,23.049849,22.547693,24.500515,26.689644,26.886566,32.88944,34.310566,32.47262,29.863386,30.119387,29.633644,29.574566,27.572515,24.109951,22.521437,23.095797,21.333336,20.46359,21.91754,25.360413,20.857437,21.96349,24.73354,26.912823,27.940105,24.119797,22.09149,20.54236,19.134361,18.5239,19.817028,20.480001,22.78072,24.841848,20.630976,17.8839,20.93949,24.864822,27.060514,27.267284,20.736002,15.724309,11.881026,9.449026,9.278359,6.616616,6.6560006,6.76759,6.370462,6.941539,17.670565,22.468925,24.201847,25.718155,29.830566,30.611694,21.53354,12.714667,7.9950776,4.9460516,3.626667,3.7185643,5.989744,8.628513,7.250052,11.546257,13.489232,12.1698475,9.4916935,10.161232,5.8420515,4.0369234,2.9013336,1.6508719,0.56451285,0.7844103,0.6301539,0.36102566,0.13784617,0.016410258,1.1749744,1.6738462,1.7362052,1.6902566,1.9823592,1.0568206,0.8598975,0.8172308,0.75487185,0.8992821,0.30194873,0.28882053,0.508718,0.574359,0.06235898,0.013128206,0.4201026,1.782154,3.249231,2.6387694,3.7251284,4.279795,3.6824617,2.8389745,4.1813335,6.439385,5.7140517,4.381539,4.391385,7.24677,4.6966157,3.1343591,2.5304618,2.3040001,1.3259488,4.585026,3.7448208,2.4320002,2.100513,2.0151796,1.5622566,2.6289232,2.9538465,2.1070771,1.4966155,1.9954873,2.5600002,2.3958976,1.9003079,2.6715899,2.6223593,1.7755898,0.94523084,0.45292312,0.12143591,0.098461546,0.20020515,0.35446155,0.44307697,0.32164106,0.955077,3.255795,4.6834874,3.9023592,0.7778462,1.5360001,3.1803079,3.8990772,3.3017437,2.412308,2.5074873,2.1858463,2.1103592,2.4582565,2.8849232,1.4309745,0.6826667,0.7811283,1.8937438,4.2272825,2.0545642,1.2537436,3.5052311,7.1089234,6.987488,5.2545643,4.2896414,2.5632823,0.43323082,0.15425642,0.26256412,0.7384616,0.8730257,0.6826667,0.9156924,5.87159,6.498462,5.5204105,5.3431797,8.041026,12.642463,11.651283,9.6065645,9.849437,14.50995,20.60472,40.418465,60.478363,68.608,53.970055,51.200005,48.12472,44.71467,44.02872,52.230568,49.972515,47.090874,42.39754,33.48021,16.708925,14.244103,13.863386,12.576821,9.170052,4.2272825,7.4732313,8.267488,8.723693,9.127385,7.9195905,5.5991797,4.9099493,6.5903597,8.602257,6.1505647,4.3552823,2.7437952,1.7132308,3.308308,11.23118,8.861539,4.781949,4.2502565,7.5946674,10.20718,6.363898,6.820103,7.8637953,11.687386,26.397541,9.931488,7.817847,8.52677,7.8112826,8.726975,9.911796,14.007796,12.12718,5.5532312,5.737026,13.049437,16.049232,13.8765135,9.38995,9.170052,6.2884107,4.893539,6.2162056,8.779488,8.375795,6.117744,3.1638978,4.7228723,8.982975,7.141744,4.417641,6.7774363,6.619898,2.9210258,1.2373334,1.4441026,1.2668719,1.2537436,4.138667,14.831591,6.738052,3.1573336,9.110975,20.949335,26.38113,12.928001,7.269744,8.172308,11.657847,10.985026,4.9788723,3.2032824,3.7842054,4.417641,2.3794873,2.284308,1.6640002,1.3522053,1.6771283,2.4713848,2.3860514,1.7165129,1.9889232,3.0194874,2.8849232,2.5665643,2.3236926,1.7591796,1.0075898,0.702359,0.50543594,0.23958977,0.072205134,0.06564103,0.13784617,0.2231795,0.20676924,0.17066668,0.15425642,0.16738462,0.032820515,0.0,0.06235898,0.13456412,0.06235898,0.013128206,0.118153855,0.30194873,0.49230772,0.6268718,0.69907695,0.6170257,0.40369233,0.19692309,0.24287182,0.37743592,0.26584616,0.17394873,0.15753847,0.06235898,0.072205134,0.07548718,0.17394873,0.27569234,0.09189744,0.128,0.14769232,0.14769232,0.11158975,0.016410258,0.026256412,0.11158975,0.2100513,0.24615386,0.13784617,0.06564103,0.04594872,0.032820515,0.016410258,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.02297436,0.026256412,0.016410258,0.026256412,0.029538464,0.02297436,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.108307704,0.16410258,0.128,0.055794876,0.09189744,0.54482055,0.92225647,0.96492314,0.6465641,0.18379489,0.036102567,0.0,0.04266667,0.13128206,0.2297436,0.04594872,0.0,0.0,0.0,0.0,0.0,0.026256412,0.052512825,0.072205134,0.12143591,0.12143591,0.08533334,0.06235898,0.07548718,0.13784617,0.18707694,0.17066668,0.14112821,0.15425642,0.28882053,0.55794877,0.7450257,0.8730257,0.92225647,0.82379496,0.6301539,0.42338464,0.40697438,0.4266667,0.0,0.0,0.0,0.0,0.0,0.0,0.098461546,0.40697438,0.4004103,0.13128206,0.2297436,0.19364104,0.09189744,0.02297436,0.029538464,0.09189744,0.06564103,0.02297436,0.006564103,0.02297436,0.04594872,0.04594872,0.055794876,0.07876924,0.11158975,0.13784617,0.026256412,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08205129,0.15097436,0.18379489,0.24287182,0.26912823,0.21989745,0.128,0.055794876,0.09189744,0.2855385,0.508718,0.6629744,0.764718,0.9616411,1.1093334,1.3259488,1.4080001,1.1520001,0.380718,0.45620516,0.53825647,0.63343596,0.6695385,0.47261542,0.3249231,0.28225642,0.2986667,0.3446154,0.380718,0.5874872,0.7417436,0.761436,0.67938465,0.65641034,0.7417436,0.7811283,0.7384616,0.6071795,0.4135385,0.44964105,0.81394875,1.2668719,1.5425643,1.3587693,1.0666667,1.0010257,1.086359,1.2373334,1.3587693,1.1749744,1.020718,0.9353847,0.92553854,0.9616411,0.75487185,0.5907693,0.6826667,0.97805136,1.1749744,1.1979488,1.214359,1.4145643,1.6935385,1.6311796,1.204513,1.0338463,0.9419488,0.8172308,0.6104616,0.4266667,0.3446154,0.28882053,0.24615386,0.25928208,0.3708718,0.3511795,0.3708718,0.46933338,0.58092314,0.6301539,0.512,0.4201026,0.40697438,0.380718,0.380718,0.380718,0.3511795,0.31507695,0.3511795,0.47261542,0.4955898,0.48246157,0.47917953,0.5021539,0.5152821,0.5546667,0.53825647,0.48246157,0.51856416,0.46933338,0.47589746,0.54482055,0.5940513,0.47261542,0.28882053,0.20676924,0.190359,0.20348719,0.2297436,0.3249231,0.4135385,0.512,0.55794877,0.4135385,0.37415388,0.35774362,0.3446154,0.35446155,0.4266667,0.46276927,0.41682056,0.38728207,0.39056414,0.36758977,0.36758977,0.38400003,0.40369233,0.41025645,0.39712822,0.54482055,0.5349744,0.47261542,0.40369233,0.3052308,0.23302566,0.2231795,0.2297436,0.2231795,0.19692309,0.23630771,0.26256412,0.39712822,0.6170257,0.761436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.01969231,0.013128206,0.029538464,0.036102567,0.026256412,0.0,0.013128206,0.108307704,0.190359,0.2231795,0.23958977,0.30851284,0.38400003,0.49230772,0.574359,0.50543594,0.7384616,0.56123084,0.36102566,0.3052308,0.35774362,0.7384616,0.5874872,0.40697438,0.41025645,0.5316923,1.3817437,2.5895386,4.204308,5.543385,5.1987696,6.235898,7.2237954,7.77518,7.9327188,8.188719,8.766359,11.723488,14.884104,17.391592,19.721848,23.6439,31.438772,49.762466,71.56513,76.11406,57.50154,40.72698,29.177439,24.30031,25.600002,23.719387,26.453335,31.330463,35.042465,33.440823,34.750362,33.125748,30.529644,28.980515,30.585438,31.891695,32.869747,30.664207,26.026669,23.328823,25.85272,24.726976,24.152617,25.839592,29.010054,28.343798,28.432413,28.133745,27.254156,26.57149,24.421745,21.208616,18.83241,18.113642,18.793028,19.843283,21.746874,24.264208,24.454565,16.699078,14.979283,14.162052,14.953027,16.239592,15.110565,11.099898,8.444718,7.8670774,9.042052,10.607591,9.265231,8.667898,7.860513,6.3310776,4.013949,10.975181,15.619284,17.821539,18.884924,21.543386,24.999386,21.270975,20.998566,23.588104,17.184822,13.213539,12.104206,11.241027,11.339488,16.46277,12.3536415,7.3025646,4.33559,4.578462,7.269744,4.6769233,2.5074873,1.5721027,1.6804104,1.6377437,1.0371283,0.81066674,0.52512825,0.14441027,0.0032820515,0.55794877,1.7493335,2.425436,2.2777438,1.8379488,0.67610264,0.38400003,0.44307697,0.5546667,0.6301539,0.18051283,0.17394873,0.2986667,0.32164106,0.12143591,0.02297436,0.18051283,0.7778462,1.6180514,2.0906668,3.1573336,3.8465643,3.7415388,3.1967182,3.3378465,5.4514875,5.156103,4.3027697,4.1846156,5.5269747,4.7228723,3.5249233,2.7109745,2.4057438,2.0709746,2.1956925,2.1366155,1.9495386,1.8313848,2.1366155,2.0742567,2.5304618,3.4789746,4.0533338,2.5435898,2.176,1.9593848,1.6377437,1.5491283,2.6223593,2.8947694,2.553436,1.8576412,1.0699488,0.47589746,0.24615386,0.23958977,0.33476925,0.47261542,0.6629744,1.2471796,3.1573336,4.4832826,4.4734364,3.5249233,2.8849232,3.639795,4.6211286,4.772103,3.117949,4.9460516,4.1222568,3.05559,3.1934361,5.0576415,3.2918978,1.5885129,1.270154,2.858667,6.0685134,2.9604106,3.2000003,4.896821,6.3212314,5.914257,4.5128207,2.7306669,1.394872,1.0075898,1.7526156,1.8806155,1.6508719,2.4549747,4.97559,9.189744,7.0859494,3.8596926,2.674872,3.7940516,4.588308,6.1341543,6.882462,7.020308,8.093539,13.010053,22.498463,42.912823,56.3758,55.122055,41.521233,37.07077,38.95139,39.49621,37.779694,39.647182,37.96349,36.391388,33.621334,28.205952,18.550156,12.63918,10.381129,9.531077,9.353847,10.610872,11.641437,9.947898,8.349539,7.5520005,6.1505647,5.549949,5.21518,6.951385,9.4916935,8.493949,6.482052,5.3103595,4.906667,5.474462,7.4699492,4.342154,3.4100516,4.086154,7.3649235,15.835898,7.752206,4.338872,4.7524104,13.354668,39.712822,14.546052,12.645744,18.881643,20.325745,6.262154,4.4307694,9.754257,11.145847,6.951385,4.969026,9.731283,12.967385,12.209231,8.641642,7.0957956,5.717334,3.7874875,5.113436,9.386667,12.196103,6.0324106,4.204308,5.1298466,6.173539,3.636513,3.8367183,7.7456417,8.674462,6.2687182,6.49518,8.129642,12.301129,13.275898,11.533129,13.768207,8.274052,4.6244106,9.117539,18.898052,21.976618,13.249642,9.216001,8.73354,10.118565,11.155693,6.567385,3.8038976,2.681436,2.3893335,1.5031796,1.6672822,1.6114873,1.6672822,2.0644104,2.934154,2.665026,2.2482052,2.409026,3.6758976,6.373744,4.699898,3.2656412,2.294154,1.7263591,1.214359,0.77456415,0.31507695,0.06564103,0.055794876,0.101743594,0.128,0.17066668,0.16738462,0.12471796,0.108307704,0.03938462,0.02297436,0.032820515,0.049230773,0.072205134,0.072205134,0.052512825,0.068923086,0.17066668,0.380718,0.88287187,0.6662565,0.32164106,0.17723078,0.3052308,0.3314872,0.2297436,0.16082053,0.14769232,0.06235898,0.032820515,0.04266667,0.15097436,0.27241027,0.17723078,0.0951795,0.098461546,0.1148718,0.101743594,0.06564103,0.055794876,0.06564103,0.12143591,0.17394873,0.06564103,0.029538464,0.02297436,0.013128206,0.0032820515,0.0032820515,0.0,0.006564103,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.016410258,0.016410258,0.016410258,0.01969231,0.016410258,0.013128206,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.032820515,0.08861539,0.09189744,0.04266667,0.029538464,0.40369233,0.7417436,0.94523084,0.88615394,0.40369233,0.19692309,0.059076928,0.013128206,0.03938462,0.068923086,0.013128206,0.0,0.0,0.0,0.0,0.0,0.04266667,0.09189744,0.118153855,0.108307704,0.108307704,0.101743594,0.128,0.18051283,0.2231795,0.23302566,0.20020515,0.19364104,0.23958977,0.3249231,0.3117949,0.3314872,0.42994875,0.56451285,0.60389745,0.6629744,0.49230772,0.30194873,0.16738462,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.01969231,0.22646156,0.26584616,0.14112821,0.2297436,0.318359,0.21989745,0.14441027,0.128,0.04266667,0.055794876,0.052512825,0.04594872,0.036102567,0.02297436,0.02297436,0.23630771,0.25928208,0.07548718,0.03938462,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.029538464,0.03938462,0.055794876,0.098461546,0.15753847,0.17394873,0.20348719,0.17066668,0.08533334,0.04266667,0.14112821,0.33805132,0.5349744,0.7122052,0.9353847,1.083077,1.1946667,1.0732309,0.7417436,0.42994875,0.4660513,0.55794877,0.6432821,0.65969235,0.58420515,0.4955898,0.39712822,0.33805132,0.30851284,0.24615386,0.4660513,0.67938465,0.79425645,0.81066674,0.81394875,0.73517954,0.7253334,0.7253334,0.6662565,0.4594872,0.41025645,0.5546667,0.9353847,1.3850257,1.5524104,1.2012309,1.0732309,1.079795,1.204513,1.4933335,1.719795,1.6213335,1.4112822,1.214359,1.0962052,0.8402052,0.8041026,0.7844103,0.7417436,0.8205129,1.2373334,1.2471796,1.2471796,1.4769232,2.0118976,1.7099489,1.3456411,1.083077,0.892718,0.53825647,0.3446154,0.26584616,0.256,0.26584616,0.24615386,0.23958977,0.21333335,0.2231795,0.28882053,0.41025645,0.5152821,0.508718,0.47589746,0.43651286,0.3314872,0.30194873,0.3117949,0.3249231,0.3314872,0.33805132,0.4135385,0.4201026,0.4004103,0.37743592,0.380718,0.4135385,0.44307697,0.48246157,0.5349744,0.5907693,0.54482055,0.55794877,0.67610264,0.8008206,0.6695385,0.4955898,0.44307697,0.36758977,0.26256412,0.27897438,0.33476925,0.39384618,0.446359,0.48574364,0.48574364,0.4397949,0.4266667,0.4135385,0.38728207,0.35446155,0.36102566,0.3511795,0.3446154,0.34133336,0.318359,0.36758977,0.5152821,0.63343596,0.65969235,0.58092314,0.69579494,0.69579494,0.6235898,0.51856416,0.40369233,0.26256412,0.21989745,0.24615386,0.2986667,0.3314872,0.37743592,0.3446154,0.31507695,0.35446155,0.48246157,0.01969231,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0032820515,0.006564103,0.01969231,0.049230773,0.101743594,0.03938462,0.04594872,0.07548718,0.108307704,0.14441027,0.2231795,0.38728207,0.50543594,0.52512825,0.48246157,0.7089231,0.67282057,0.508718,0.34789747,0.3117949,0.48902568,0.3314872,0.2100513,0.26912823,0.4266667,1.7165129,2.6420515,3.7743592,4.9362054,5.1954875,5.4153852,5.664821,6.0947695,6.8004107,7.821129,10.033232,14.089848,18.980104,24.06072,29.062567,36.079594,54.37703,79.75713,96.08206,75.30995,49.83467,33.7559,25.3079,23.007181,25.652515,27.697233,31.015387,33.99549,35.091694,32.836926,35.492104,35.11467,32.42995,29.686155,30.683899,31.24513,30.191591,27.64472,24.832003,24.050873,26.640411,28.3799,30.020926,31.392822,31.396105,28.868925,27.181952,25.15036,22.90872,21.90113,21.40554,20.214155,19.337847,19.34113,20.33231,19.206566,17.732924,17.224207,17.092924,14.864411,11.592206,10.013539,10.387693,12.081232,13.561437,10.157949,7.1909747,9.494975,15.274668,16.065641,15.780104,15.232001,13.5778475,11.700514,12.20595,9.970873,10.994873,11.825232,12.534155,16.695797,21.225027,18.904617,16.321642,15.688207,14.864411,17.80513,17.900309,14.815181,11.218052,12.754052,10.860309,6.9645133,4.2863593,3.8662567,4.568616,2.8389745,1.7263591,2.0020514,2.9768207,2.4943593,1.5688206,1.2438976,0.78769237,0.16410258,0.009846155,0.39712822,1.3686155,1.9429746,1.8904617,1.7362052,0.8598975,0.40697438,0.32820517,0.5021539,0.74830776,0.38400003,0.37743592,0.508718,0.5546667,0.30194873,0.25928208,0.26584616,0.48574364,0.8598975,1.1191796,1.8904617,2.5009232,2.4976413,2.0906668,2.166154,3.0785644,2.9801028,2.8717952,3.3017437,4.3552823,4.1878977,3.4625645,2.7733335,2.3958976,2.3138463,2.2678976,2.3072822,1.9626669,1.6344616,2.5862565,2.3696413,2.28759,2.989949,3.8367183,2.9078977,2.038154,1.3817437,1.0272821,1.1126155,1.847795,2.3926156,2.5796926,2.284308,1.6475899,1.0666667,0.90584624,0.6465641,0.47917953,0.5677949,1.0765129,1.6147693,3.1606157,4.70318,5.6254363,5.720616,3.817026,3.4166157,3.9089234,4.2535386,2.9768207,3.7973337,3.2196925,2.1333334,1.5491283,2.5698464,2.169436,1.9692309,1.9692309,2.7208207,5.3234878,2.9669745,4.0008206,5.402257,5.6287184,4.601436,4.772103,4.204308,3.1967182,2.481231,3.2328207,3.131077,3.5446157,4.092718,4.7917953,6.0783596,5.2348723,3.6036925,4.352,6.672411,5.7829747,4.0008206,3.8367183,4.1124105,5.169231,8.854975,17.946259,33.83467,45.443287,46.916927,37.609028,27.69395,32.580925,38.65272,38.288414,29.863386,26.866875,25.137232,24.018053,22.17354,17.56554,11.85477,8.868103,8.3823595,9.577026,11.044104,10.84718,7.8802056,5.2348723,4.027077,3.3805132,3.4166157,5.5893335,8.392206,9.947898,8.018052,6.76759,4.900103,9.941334,16.042667,3.9942567,2.8947694,3.7284105,4.594872,6.9152827,15.43877,7.6570263,3.2328207,4.194462,13.190565,33.47036,12.681848,10.30236,14.8709755,16.170668,5.2512827,3.4494362,7.5585647,9.53436,7.3058467,4.7950773,5.835488,8.953437,10.43036,9.29477,7.2894363,6.12759,4.5128207,5.943795,9.45559,9.619693,4.772103,6.229334,7.9097443,6.5706673,1.8084104,3.0391798,6.4754877,8.283898,7.4436927,5.7698464,6.941539,11.372309,11.323078,7.3780518,8.4512825,7.059693,5.0018463,6.803693,11.510155,12.688411,8.4283085,8.608821,9.504821,9.317744,8.198565,5.7764106,3.2787695,1.8248206,1.6672822,2.1530259,1.913436,1.9495386,2.3105643,3.0424619,4.1682053,4.0041027,4.056616,4.1583595,4.4865646,5.5630774,3.8071797,2.8324106,2.1989746,1.7362052,1.5261539,1.0404103,0.4135385,0.06564103,0.06235898,0.128,0.08205129,0.108307704,0.15753847,0.16410258,0.036102567,0.016410258,0.029538464,0.08533334,0.14769232,0.12143591,0.06235898,0.01969231,0.0032820515,0.036102567,0.13784617,0.4397949,0.32820517,0.15097436,0.09189744,0.17394873,0.2100513,0.2297436,0.2231795,0.18707694,0.1148718,0.04266667,0.06564103,0.3249231,0.761436,1.1126155,0.30194873,0.09189744,0.08861539,0.101743594,0.15753847,0.118153855,0.068923086,0.06564103,0.08205129,0.036102567,0.026256412,0.01969231,0.013128206,0.006564103,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.006564103,0.006564103,0.006564103,0.006564103,0.006564103,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.032820515,0.04266667,0.02297436,0.006564103,0.17066668,0.35446155,0.5513847,0.63343596,0.36758977,0.21333335,0.08533334,0.01969231,0.006564103,0.013128206,0.0032820515,0.0,0.0032820515,0.006564103,0.0,0.0,0.01969231,0.04266667,0.06564103,0.068923086,0.055794876,0.055794876,0.09189744,0.14769232,0.20676924,0.2297436,0.22646156,0.27241027,0.3708718,0.446359,0.33805132,0.20676924,0.17394873,0.24615386,0.3117949,0.37415388,0.26584616,0.13128206,0.052512825,0.032820515,0.02297436,0.013128206,0.006564103,0.0,0.0,0.0,0.07876924,0.17723078,0.21989745,0.09189744,0.18379489,0.14112821,0.08533334,0.06235898,0.013128206,0.02297436,0.02297436,0.02297436,0.016410258,0.006564103,0.07876924,0.21333335,0.19692309,0.04594872,0.032820515,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.009846155,0.013128206,0.052512825,0.16410258,0.118153855,0.16410258,0.17723078,0.12471796,0.059076928,0.07876924,0.21989745,0.40369233,0.60061544,0.8467693,0.9517949,1.0108719,0.93866676,0.7450257,0.5349744,0.43323082,0.48246157,0.64000005,0.78769237,0.7384616,0.5546667,0.38400003,0.27897438,0.23630771,0.19692309,0.38728207,0.49887183,0.5940513,0.7056411,0.827077,0.74830776,0.71548724,0.73517954,0.7417436,0.5907693,0.52512825,0.55794877,0.761436,1.1060513,1.463795,1.332513,1.2996924,1.3883078,1.5753847,1.8084104,2.0939488,2.2219489,2.1169233,1.8543591,1.6508719,1.273436,1.0765129,0.9419488,0.83035904,0.8041026,1.142154,1.2438976,1.2209232,1.2209232,1.4375386,1.3883078,1.3095386,1.1815386,1.024,0.8763078,0.7253334,0.4397949,0.27569234,0.27897438,0.28882053,0.23958977,0.18051283,0.15753847,0.18051283,0.23958977,0.30851284,0.33476925,0.33476925,0.3117949,0.24615386,0.22646156,0.23302566,0.26584616,0.3052308,0.3249231,0.3511795,0.36430773,0.3708718,0.3708718,0.37743592,0.40697438,0.43323082,0.4594872,0.48574364,0.51856416,0.49230772,0.508718,0.6071795,0.73517954,0.7187693,0.53825647,0.54482055,0.49230772,0.3708718,0.39056414,0.446359,0.48574364,0.5316923,0.5677949,0.5316923,0.4397949,0.4201026,0.42338464,0.41025645,0.36430773,0.33476925,0.32164106,0.32164106,0.33476925,0.36102566,0.38400003,0.45620516,0.54482055,0.5973334,0.5513847,0.6695385,0.7089231,0.65969235,0.5415385,0.4266667,0.3117949,0.29210258,0.3117949,0.35446155,0.4397949,0.5481026,0.45620516,0.33476925,0.3052308,0.4201026,0.04266667,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.01969231,0.049230773,0.108307704,0.03938462,0.013128206,0.01969231,0.04594872,0.08861539,0.23630771,0.37743592,0.42994875,0.40697438,0.4266667,0.57764107,0.6432821,0.51856416,0.27241027,0.17066668,0.19364104,0.14112821,0.128,0.20348719,0.34133336,1.6640002,2.556718,3.4198978,4.2601027,4.6933336,4.414359,4.342154,4.7655387,5.76,7.181129,10.377847,15.126975,21.589334,29.650053,38.908722,49.48021,67.90565,85.648415,89.29478,60.576824,37.586056,25.560617,21.346462,22.170258,25.64595,29.630362,33.391594,35.649643,36.240414,36.12554,37.428516,35.862976,32.718773,30.063593,30.736412,30.401644,28.291285,27.224617,28.5079,31.93108,32.055798,33.792004,35.13436,34.46154,30.549335,26.312206,23.742361,21.211899,18.786463,18.20554,18.858667,19.216412,18.898052,18.153027,17.857643,14.857847,12.153437,10.883283,11.122872,11.867898,8.900924,7.9786673,8.3134365,9.527796,11.657847,8.65477,6.2851286,9.7673855,16.459488,15.835898,15.012104,13.351386,11.611898,11.264001,14.477129,11.21477,10.640411,8.960001,7.6143594,13.29559,17.673847,15.973744,10.939077,6.9710774,10.098872,15.409232,16.41354,14.132514,10.496001,8.310155,8.083693,6.0061545,4.0533338,3.0096412,2.481231,1.657436,1.4966155,2.5764105,3.879385,2.7864618,1.9068719,1.5360001,1.1027694,0.48574364,0.016410258,0.5513847,1.4211283,1.7427694,1.4834872,1.4572309,1.3423591,0.8172308,0.5940513,0.80738467,1.0272821,0.93866676,1.083077,1.0601027,0.7844103,0.49230772,0.5415385,0.45292312,0.45292312,0.571077,0.6268718,1.1651284,1.3423591,1.2373334,1.1027694,1.3784616,1.5327181,1.5491283,2.0086155,2.8947694,3.5905645,3.4855387,3.3345644,3.0884104,2.934154,3.2951798,3.436308,3.0687182,2.359795,1.9692309,3.0391798,2.28759,1.8116925,2.0184617,2.546872,2.2547693,1.3489232,0.764718,0.63343596,0.9124103,1.3850257,1.7526156,2.169436,2.2153847,1.8412309,1.3554872,1.2635899,1.1323078,1.0535386,1.0962052,1.3029745,1.9462565,2.6223593,4.2305646,6.2752824,6.8397956,4.818052,3.564308,3.2295387,3.3444104,2.8225644,3.4297438,2.8258464,1.6705642,0.6432821,0.43323082,0.77128214,1.5360001,1.7329233,1.8576412,3.892513,2.7044106,4.128821,5.3858466,5.330052,4.460308,5.1232824,5.156103,4.3651285,3.511795,4.312616,4.4274874,5.3858466,5.651693,4.637539,2.6912823,4.571898,5.723898,6.882462,7.5421543,5.940513,4.0467696,4.378257,3.9286156,2.9046156,4.709744,11.552821,20.758976,29.42031,34.609234,33.368618,22.255592,24.237951,30.33272,32.17067,22.019283,21.16595,20.059898,18.153027,15.875283,14.611693,10.758565,7.8736415,7.3780518,8.5661545,8.595693,7.145026,4.4077954,2.4057438,1.9167181,2.484513,2.3138463,5.543385,8.418462,8.756514,5.9470773,5.6352825,4.637539,9.9282055,15.714462,3.4198978,3.4330258,4.7950773,6.925129,9.616411,13.052719,6.242462,2.7241027,4.663795,12.393026,24.375797,9.787078,7.24677,10.31877,12.71795,8.297027,5.395693,6.8660517,8.73354,8.5661545,5.4843082,4.4307694,6.4065647,9.002667,10.023385,7.4929237,6.7117953,6.173539,7.0990777,8.169026,5.536821,3.1277952,7.680001,10.010257,6.954667,1.3686155,2.5698464,5.2611284,7.686565,8.605539,7.282872,8.214975,8.697436,8.224821,6.928411,5.58277,4.4964104,4.4373336,5.4383593,7.1548724,8.881231,6.941539,7.788308,8.507077,7.8736415,6.3540516,4.394667,2.4648206,1.5524104,1.8904617,2.9801028,2.4385643,2.4746668,3.121231,4.132103,5.0051284,5.113436,5.1331286,4.9985647,4.670359,4.1091285,2.7766156,2.3827693,2.0184617,1.5064616,1.3850257,1.0666667,0.4660513,0.08861539,0.072205134,0.17723078,0.06564103,0.059076928,0.101743594,0.118153855,0.0,0.0,0.016410258,0.098461546,0.18379489,0.1148718,0.029538464,0.0032820515,0.0,0.009846155,0.04594872,0.10502565,0.08205129,0.049230773,0.049230773,0.101743594,0.13128206,0.18707694,0.20020515,0.17066668,0.15097436,0.059076928,0.08861539,0.5546667,1.4080001,2.225231,0.6301539,0.13128206,0.06235898,0.08205129,0.17723078,0.16410258,0.1148718,0.06564103,0.036102567,0.029538464,0.03938462,0.032820515,0.026256412,0.02297436,0.006564103,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.009846155,0.006564103,0.0,0.02297436,0.07548718,0.17723078,0.256,0.190359,0.15753847,0.108307704,0.06564103,0.032820515,0.02297436,0.0032820515,0.0032820515,0.016410258,0.029538464,0.013128206,0.0032820515,0.0,0.009846155,0.029538464,0.06564103,0.07876924,0.098461546,0.15753847,0.26256412,0.39056414,0.39712822,0.38728207,0.4266667,0.5152821,0.5677949,0.44964105,0.21333335,0.068923086,0.06564103,0.09189744,0.10502565,0.059076928,0.026256412,0.055794876,0.16738462,0.17066668,0.15425642,0.21661541,0.27897438,0.10502565,0.118153855,0.055794876,0.08533334,0.16082053,0.0,0.04266667,0.03938462,0.016410258,0.0,0.0,0.0,0.0032820515,0.009846155,0.016410258,0.013128206,0.08205129,0.12471796,0.128,0.11158975,0.11158975,0.02297436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02297436,0.108307704,0.068923086,0.10502565,0.14441027,0.14112821,0.08861539,0.055794876,0.128,0.28225642,0.48246157,0.6826667,0.83035904,0.9485129,0.93866676,0.8008206,0.6432821,0.44964105,0.45620516,0.6301539,0.8598975,0.9353847,0.62030774,0.39712822,0.26912823,0.2100513,0.18379489,0.28225642,0.32820517,0.40697438,0.5415385,0.7220513,0.7384616,0.7220513,0.7515898,0.79097444,0.69579494,0.6301539,0.6465641,0.76800007,1.0043077,1.3718976,1.4178462,1.4342566,1.5753847,1.7920002,1.8412309,2.0709746,2.412308,2.5304618,2.4024618,2.3171284,1.8346668,1.4276924,1.1552821,1.0108719,0.9353847,1.1158975,1.2668719,1.2537436,1.1027694,0.9911796,0.9714873,1.1060513,1.2340513,1.3029745,1.3653334,1.2471796,0.75487185,0.380718,0.28225642,0.28882053,0.24943592,0.17066668,0.12471796,0.128,0.13456412,0.16082053,0.17394873,0.18051283,0.17723078,0.16738462,0.16082053,0.16738462,0.19364104,0.23630771,0.27241027,0.29538465,0.3249231,0.34789747,0.36430773,0.36758977,0.40369233,0.43323082,0.44307697,0.4397949,0.45292312,0.4594872,0.45292312,0.49230772,0.57764107,0.6432821,0.5677949,0.6498462,0.65312827,0.53825647,0.47589746,0.48246157,0.49887183,0.54482055,0.5907693,0.54482055,0.47589746,0.45620516,0.4594872,0.44964105,0.3708718,0.3446154,0.3446154,0.33805132,0.33476925,0.39712822,0.39056414,0.380718,0.41025645,0.46933338,0.4660513,0.571077,0.6498462,0.636718,0.53825647,0.4397949,0.39384618,0.3708718,0.36430773,0.4004103,0.5316923,0.64000005,0.5513847,0.4201026,0.3511795,0.41025645,0.049230773,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.016410258,0.013128206,0.036102567,0.07548718,0.08861539,0.26584616,0.318359,0.30851284,0.2986667,0.36758977,0.45292312,0.49230772,0.36430773,0.12471796,0.016410258,0.016410258,0.049230773,0.0951795,0.15753847,0.24287182,1.3095386,2.3335385,3.3509746,4.1911798,4.4996924,3.8367183,3.629949,4.092718,5.1626673,6.5345645,10.276103,15.688207,22.790565,31.619284,42.22031,53.730465,61.781338,63.612724,57.442467,42.466465,28.261745,20.578463,18.586258,20.65395,24.356104,28.389746,32.784412,36.52267,39.446976,42.24985,38.87918,34.6519,32.26913,32.390568,33.61149,34.195694,32.81395,33.94626,38.531284,43.96308,39.384617,37.832207,36.36185,32.82708,25.882257,21.881437,19.557745,17.54913,15.849027,15.82277,16.83036,17.293129,16.374155,14.201437,11.894155,9.252103,8.854975,9.019077,8.726975,7.6307697,6.9677954,6.816821,6.7150774,6.5739493,6.672411,5.1200004,5.110154,8.188719,12.009027,10.338462,7.975385,4.7360005,3.373949,4.8836927,8.503796,12.632616,13.062565,8.996103,4.673641,9.366975,12.337232,11.940104,8.973129,6.675693,10.755282,10.94236,11.034257,11.244308,10.860309,8.214975,5.3398976,3.0818465,1.7033848,1.3981539,2.284308,1.9626669,1.8084104,2.609231,3.5807183,2.3827693,2.0151796,1.7657437,1.654154,1.3226668,0.03938462,0.67938465,1.6836925,1.847795,1.2471796,1.2537436,1.9003079,1.4080001,1.1224617,1.3193847,1.2209232,1.4572309,1.7690258,1.5327181,0.8730257,0.65641034,0.69579494,0.55794877,0.42994875,0.4397949,0.64000005,1.0305642,0.7056411,0.5218462,0.75487185,1.1093334,1.4473847,1.6377437,2.349949,3.2918978,3.2196925,2.9768207,3.4133337,3.7185643,3.8629746,4.588308,4.348718,3.5249233,2.789744,2.6190772,3.2787695,2.0742567,1.3587693,1.2340513,1.4572309,1.4342566,0.69579494,0.4955898,0.7811283,1.2668719,1.401436,1.332513,1.6049232,1.7690258,1.6213335,1.214359,1.0765129,1.5163078,2.3040001,2.7470772,1.7066668,2.3958976,1.782154,3.0194874,5.930667,7.000616,6.6395903,5.1364107,3.7284105,3.0982566,3.3542566,4.7425647,4.9132314,3.8531284,2.0873847,0.65641034,0.64000005,1.0601027,0.9944616,0.9911796,3.0785644,2.8750772,3.9942567,4.906667,5.0084105,4.647385,5.146257,5.149539,4.644103,4.33559,5.668103,6.2916927,6.875898,6.872616,5.7632823,3.0523078,5.7435904,8.080411,7.8506675,5.5269747,4.2469745,4.8607183,6.8529234,5.602462,2.0184617,2.550154,8.490667,11.372309,13.863386,17.857643,24.467693,19.685745,16.04595,16.689232,19.39036,16.571077,21.579489,20.808207,15.973744,10.962052,11.825232,9.357129,6.7938466,5.927385,6.3376417,5.408821,3.0851285,1.6475899,1.3095386,2.0217438,3.4691284,2.6190772,4.768821,6.4000006,6.0947695,4.5456414,4.023795,5.2020516,5.549949,4.7228723,4.571898,4.7983594,6.5739493,10.404103,13.4400015,9.478565,4.141949,2.934154,6.2162056,12.678565,19.344412,8.963283,7.256616,10.745437,14.49354,12.117334,8.054154,6.8562055,8.425026,10.023385,6.2752824,5.028103,5.756718,8.556309,10.84718,7.3682055,7.2270775,7.64718,7.653744,6.4623594,3.4724104,1.9331284,6.7249236,8.756514,5.756718,2.294154,3.4822567,5.605744,7.7259493,9.616411,11.762873,13.705847,10.35159,11.218052,14.27036,5.8945646,3.4100516,6.889026,9.386667,9.383386,10.807796,9.90195,8.516924,7.6964107,7.506052,7.0104623,3.8695388,2.3926156,2.2777438,2.986667,3.748103,3.570872,3.5971284,4.2174363,5.0510774,4.955898,5.9503593,5.477744,4.772103,4.2535386,3.5052311,2.6256413,2.3860514,1.9922053,1.3456411,1.0371283,0.9616411,0.48902568,0.128,0.072205134,0.19692309,0.06235898,0.032820515,0.02297436,0.0,0.0,0.0,0.0032820515,0.055794876,0.12143591,0.06564103,0.013128206,0.0,0.0,0.016410258,0.07876924,0.07876924,0.059076928,0.052512825,0.08205129,0.15097436,0.19364104,0.16082053,0.1148718,0.098461546,0.14769232,0.07548718,0.08861539,0.6170257,1.6443079,2.6912823,1.0075898,0.27897438,0.059076928,0.052512825,0.12143591,0.2231795,0.20020515,0.1148718,0.03938462,0.029538464,0.052512825,0.052512825,0.04594872,0.036102567,0.016410258,0.006564103,0.0032820515,0.006564103,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.08533334,0.12471796,0.16738462,0.18379489,0.10502565,0.01969231,0.006564103,0.032820515,0.06235898,0.06235898,0.02297436,0.016410258,0.04266667,0.098461546,0.17723078,0.22646156,0.22646156,0.3052308,0.512,0.82379496,0.761436,0.6662565,0.6071795,0.5907693,0.58092314,0.46276927,0.21333335,0.049230773,0.01969231,0.0032820515,0.0032820515,0.0,0.013128206,0.08533334,0.28225642,0.3117949,0.30194873,0.446359,0.5940513,0.23958977,0.28882053,0.18051283,0.068923086,0.016410258,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.02297436,0.032820515,0.02297436,0.013128206,0.04594872,0.12143591,0.19692309,0.18707694,0.03938462,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01969231,0.03938462,0.08533334,0.13456412,0.12143591,0.049230773,0.06235898,0.17723078,0.35774362,0.49887183,0.7187693,0.96492314,0.96492314,0.7581539,0.69579494,0.53825647,0.5284103,0.6235898,0.7975385,1.0404103,0.7318975,0.512,0.36102566,0.25928208,0.18379489,0.16738462,0.23302566,0.32164106,0.4266667,0.574359,0.73517954,0.75487185,0.7778462,0.81394875,0.7417436,0.67282057,0.7384616,0.8992821,1.1224617,1.3686155,1.3915899,1.332513,1.4244103,1.6180514,1.585231,1.7526156,2.1989746,2.5107694,2.609231,2.737231,2.4516926,1.9954873,1.5556924,1.2504616,1.0994873,1.1749744,1.2800001,1.2898463,1.1815386,1.0305642,0.8008206,0.8763078,1.1618463,1.4933335,1.6410258,1.6771283,1.1881026,0.67610264,0.37743592,0.27241027,0.2297436,0.15097436,0.108307704,0.108307704,0.108307704,0.1148718,0.108307704,0.101743594,0.101743594,0.108307704,0.108307704,0.118153855,0.128,0.14769232,0.18379489,0.24615386,0.28882053,0.31507695,0.3249231,0.31507695,0.36430773,0.40369233,0.4266667,0.4397949,0.45620516,0.48574364,0.44307697,0.41682056,0.446359,0.5284103,0.574359,0.7384616,0.81394875,0.7220513,0.49887183,0.44307697,0.4201026,0.4397949,0.48246157,0.49887183,0.52512825,0.5316923,0.52512825,0.49230772,0.36430773,0.37415388,0.4004103,0.38728207,0.3511795,0.39384618,0.38728207,0.36102566,0.36430773,0.38728207,0.37743592,0.45620516,0.55794877,0.574359,0.50543594,0.446359,0.46933338,0.4201026,0.40697438,0.48246157,0.63343596,0.6432821,0.60061544,0.5218462,0.42994875,0.380718,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.026256412,0.013128206,0.0,0.0032820515,0.016410258,0.06564103,0.0951795,0.18707694,0.3052308,0.3052308,0.48902568,0.37743592,0.20020515,0.07548718,0.016410258,0.016410258,0.032820515,0.026256412,0.036102567,0.18379489,1.0633847,1.8215386,3.2131286,5.07077,6.3179493,5.0116925,4.44718,4.5489235,5.3005133,6.7282057,10.745437,17.7559,24.677746,29.170874,29.650053,33.923286,35.40349,35.718567,34.264618,28.182976,23.860516,21.90113,20.36513,19.557745,22.048822,27.076925,30.431181,33.923286,37.254566,38.02585,34.169437,34.47467,38.29498,43.14585,44.708107,49.588516,48.292107,48.213337,49.870773,46.903797,36.614567,32.735184,30.385233,26.17436,18.20554,14.116103,11.976206,11.175385,11.099898,11.122872,11.625027,12.507898,12.662155,11.464206,8.805744,10.341744,11.825232,9.957745,5.8945646,5.2480006,4.7228723,4.5554876,4.4406157,4.266667,4.1189747,5.8781543,8.109949,10.7848215,12.452104,10.253129,7.860513,5.8157954,4.010667,3.5347695,6.6822567,13.51877,13.203693,8.743385,3.8498464,2.9440002,2.8127182,4.2240005,6.373744,10.607591,20.447182,16.259283,13.236514,12.832822,13.453129,10.436924,4.2601027,1.975795,1.3653334,2.176,6.117744,4.1156926,2.8488207,2.3269746,2.1267693,1.3587693,2.297436,2.487795,2.8521028,2.7864618,0.13784617,0.25928208,0.8205129,0.827077,0.62030774,1.8773335,2.3663592,1.8642052,1.529436,1.5261539,1.0371283,1.148718,1.1848207,1.1520001,1.0469744,0.8402052,0.54482055,0.46276927,0.3708718,0.26256412,0.33476925,0.33476925,0.16082053,0.19364104,0.508718,0.8992821,1.8642052,2.4155898,3.239385,4.0008206,3.3411283,2.9636924,3.8465643,4.4045134,4.2207184,4.073026,3.6594875,3.0687182,2.674872,2.6912823,3.2032824,2.3630772,1.5392822,1.4342566,2.0086155,2.4713848,1.4703591,1.4211283,2.0578463,2.487795,1.204513,1.204513,1.1126155,1.1749744,1.276718,0.94523084,0.65312827,1.7427694,4.44718,6.5280004,3.2820516,3.367385,1.7952822,2.0939488,4.706462,6.987488,10.308924,9.196308,6.242462,4.023795,5.110154,5.172513,10.049642,10.738873,5.976616,2.2416413,2.156308,2.4024618,1.7788719,1.1749744,3.5544617,4.240411,3.9351797,3.7251284,3.5249233,2.0611284,4.893539,6.8627696,7.1122055,6.764308,8.92718,9.366975,8.457847,7.3485136,6.1768208,4.089436,5.7731285,6.3868723,6.1078978,5.346462,4.7622566,5.8223596,6.088206,4.348718,2.1234872,3.6627696,14.513232,13.472821,8.15918,5.3760004,11.126155,18.668308,17.010874,13.899488,13.275898,15.287796,25.042053,19.938463,12.809847,10.249847,12.619488,8.772923,5.8814363,4.59159,4.210872,2.6847181,1.719795,1.4703591,1.8313848,2.6026669,3.495385,1.9692309,3.1540515,3.56759,3.5216413,7.1089234,3.373949,4.84759,5.044513,2.8389745,2.4713848,5.756718,9.9282055,12.550565,10.9686165,2.2908719,2.4582565,4.890257,10.489437,16.292105,15.488001,10.935796,11.424822,13.341539,13.177437,7.5388722,8.562873,6.449231,6.5345645,8.300308,5.3727183,3.5905645,5.4514875,9.898667,13.115078,8.513641,8.01477,7.5946674,7.387898,7.0137444,5.586052,2.03159,1.2537436,1.8346668,3.0391798,4.821334,7.3353853,8.237949,7.837539,8.050873,12.419283,16.571077,18.258053,21.943796,22.28513,4.135385,8.077128,20.122257,24.100105,16.932104,8.621949,11.0375395,11.989334,12.977232,13.026463,8.681026,5.3366156,4.2535386,4.5095387,5.175795,5.3103595,6.5805135,6.3277955,6.0061545,5.7140517,4.210872,7.716103,7.1089234,5.398975,4.066462,3.0654361,2.4681027,2.412308,2.0578463,1.3915899,1.2209232,1.1848207,0.5874872,0.13128206,0.049230773,0.12143591,0.036102567,0.006564103,0.0,0.0,0.0,0.0,0.009846155,0.06564103,0.12471796,0.07548718,0.016410258,0.0,0.0,0.006564103,0.029538464,0.029538464,0.03938462,0.08205129,0.15097436,0.19692309,0.4660513,0.36102566,0.17066668,0.072205134,0.12143591,0.108307704,0.068923086,0.20348719,0.6662565,1.5556924,1.3850257,0.6465641,0.13456412,0.072205134,0.12143591,0.39056414,0.34789747,0.17723078,0.029538464,0.029538464,0.04266667,0.055794876,0.049230773,0.026256412,0.016410258,0.016410258,0.016410258,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.026256412,0.10502565,0.35446155,0.58092314,0.27569234,0.055794876,0.0,0.02297436,0.08533334,0.18379489,0.098461546,0.08533334,0.16410258,0.3249231,0.51856416,0.46933338,0.29210258,0.26912823,0.58092314,1.3128207,1.142154,0.8960001,0.67282057,0.4955898,0.33476925,0.190359,0.07876924,0.01969231,0.0032820515,0.016410258,0.016410258,0.006564103,0.0,0.0032820515,0.016410258,0.06564103,0.0951795,0.13784617,0.18051283,0.16738462,0.25271797,0.4135385,0.3446154,0.08533334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01969231,0.055794876,0.08861539,0.07548718,0.026256412,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.055794876,0.14769232,0.18379489,0.06235898,0.03938462,0.08861539,0.20348719,0.4135385,0.49887183,0.8041026,0.8763078,0.6826667,0.6104616,0.65969235,0.67282057,0.63343596,0.6268718,0.80738467,0.86974365,0.72861546,0.5415385,0.36758977,0.18379489,0.15753847,0.19692309,0.28225642,0.39056414,0.48902568,0.8533334,0.88287187,0.85005134,0.85005134,0.7778462,0.72861546,0.8369231,1.0371283,1.2471796,1.3587693,1.1749744,0.955077,0.92553854,1.1454359,1.5097437,1.5721027,1.9987694,2.3171284,2.409026,2.5173335,3.190154,3.0358977,2.412308,1.6968206,1.2832822,1.1716924,1.1815386,1.3029745,1.3981539,1.1913847,0.81066674,0.73517954,0.8467693,1.0436924,1.2504616,1.8609232,1.7952822,1.3357949,0.77128214,0.380718,0.2231795,0.13784617,0.108307704,0.108307704,0.108307704,0.0951795,0.08205129,0.07548718,0.072205134,0.06235898,0.06235898,0.06235898,0.072205134,0.098461546,0.12143591,0.19692309,0.23958977,0.27241027,0.28882053,0.28882053,0.30194873,0.3511795,0.41682056,0.48246157,0.51856416,0.50543594,0.44964105,0.39384618,0.39384618,0.5021539,0.39384618,0.61374366,0.827077,0.8172308,0.48902568,0.49887183,0.4135385,0.33805132,0.3249231,0.3511795,0.44964105,0.5284103,0.5349744,0.47261542,0.4135385,0.4135385,0.42994875,0.42994875,0.40697438,0.380718,0.39384618,0.39712822,0.37743592,0.32820517,0.24287182,0.34133336,0.44964105,0.43651286,0.34789747,0.39712822,0.46933338,0.42338464,0.48574364,0.67282057,0.79425645,0.63343596,0.60389745,0.5907693,0.5284103,0.380718,0.036102567,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.02297436,0.036102567,0.026256412,0.029538464,0.013128206,0.0,0.0032820515,0.016410258,0.026256412,0.08205129,0.17394873,0.25271797,0.23302566,0.25928208,0.24287182,0.19692309,0.13456412,0.06564103,0.055794876,0.032820515,0.016410258,0.02297436,0.072205134,0.35774362,1.3128207,2.605949,3.8367183,4.535795,5.0149746,5.7829747,6.445949,7.1844106,8.779488,11.283693,14.683899,18.73395,23.151592,27.621746,31.123695,31.149952,29.938873,28.852514,28.3799,25.022362,24.244514,24.07713,24.4119,26.981745,33.270157,36.39467,38.902157,40.776207,39.46667,36.545643,38.508312,39.574978,39.61436,44.146873,49.683697,51.757954,51.44944,48.62031,41.911797,34.865234,28.343798,21.96677,16.416822,13.456411,10.8307705,9.672206,9.527796,10.289231,12.199386,10.315488,9.4916935,8.881231,7.9097443,6.2523084,5.927385,7.8506675,7.2631803,4.3585644,4.2962055,4.076308,4.135385,3.9712822,3.5938463,3.5347695,4.900103,5.61559,5.976616,5.970052,5.287385,3.8301542,5.602462,8.04759,9.051898,6.928411,6.157129,6.629744,6.409847,5.097026,3.8104618,14.339283,9.783795,3.9023592,4.2436924,12.160001,17.686975,12.744206,7.529026,5.5663595,3.6758976,1.8740515,1.0699488,0.6826667,0.7844103,2.0906668,1.9922053,1.7558975,1.7657437,1.8018463,1.0535386,0.8992821,1.8838975,3.6660516,4.8607183,3.0424619,1.7493335,1.7526156,1.5556924,0.8763078,0.62030774,0.8533334,0.8533334,1.2570257,1.9922053,2.294154,1.975795,1.2012309,0.90256417,1.1388719,1.1093334,0.9517949,0.6695385,0.56123084,0.7253334,1.0305642,0.6104616,0.23630771,0.3314872,0.8172308,1.1191796,1.4900514,1.9889232,2.4352822,2.7569232,2.986667,2.3663592,3.3444104,4.772103,5.4153852,3.9384618,3.4166157,2.6486156,2.7831798,3.8301542,4.644103,2.7175386,2.0053334,2.15959,2.5731285,2.3630772,1.2537436,1.6180514,2.5271797,2.8488207,1.2537436,1.1749744,2.2580514,3.4560003,3.698872,1.8740515,1.0535386,1.270154,3.2918978,6.439385,8.602257,3.3476925,1.9790771,1.9167181,2.169436,3.3378465,7.5979495,7.680001,5.9667697,4.194462,3.4625645,3.2328207,4.841026,6.0061545,5.989744,5.6254363,8.4283085,8.362667,5.832206,3.5807183,6.705231,8.756514,7.1876926,4.926359,3.3575387,2.353231,5.4383593,7.525744,8.2445135,8.103385,8.487385,10.518975,10.223591,10.345026,11.559385,12.448821,12.76718,9.245539,6.875898,6.678975,5.7140517,6.012718,8.073847,6.5870776,3.0752823,5.8847184,11.1294365,8.54318,4.309334,3.2196925,8.644924,13.679591,18.04472,18.566566,14.736411,8.73354,17.893745,16.213335,10.873437,6.744616,6.370462,5.5893335,8.438154,8.349539,4.97559,4.161641,3.764513,3.3411283,3.56759,4.0434875,3.2754874,3.114667,3.314872,6.7938466,10.243283,4.1583595,2.3729234,4.352,5.1364107,3.817026,3.508513,5.602462,13.568001,15.872002,10.742155,6.193231,6.298257,6.426257,11.234463,16.338053,8.3364105,7.1614366,8.211693,10.463181,11.001437,4.9985647,8.933744,8.096821,6.5936418,5.9470773,5.077334,2.740513,4.4832826,9.672206,14.483693,11.933539,7.643898,7.325539,7.9458466,7.568411,5.32677,2.986667,2.8422565,2.674872,2.2711797,3.4166157,6.744616,6.941539,8.086975,11.74318,16.97477,36.44718,34.454975,29.43672,23.840822,4.135385,11.23118,28.320822,32.105026,20.70318,13.650052,12.268309,10.440206,12.189539,15.00554,9.829744,7.3649235,9.642668,10.532104,8.474257,6.4689236,7.525744,6.232616,5.648411,6.5345645,7.3485136,8.041026,6.3343596,4.273231,3.131077,3.4100516,1.9692309,1.3817437,1.3784616,1.5589745,1.3686155,1.2635899,0.7450257,0.27241027,0.06235898,0.08533334,0.049230773,0.016410258,0.0,0.0,0.0,0.0,0.016410258,0.04266667,0.06235898,0.052512825,0.049230773,0.049230773,0.029538464,0.06564103,0.33476925,1.2537436,0.8172308,0.24615386,0.068923086,0.13784617,0.2986667,0.28882053,0.18707694,0.098461546,0.15753847,0.16738462,0.118153855,0.108307704,0.2986667,0.8960001,1.3718976,1.2471796,0.8369231,0.38728207,0.08533334,0.20676924,0.35446155,0.37415388,0.27241027,0.21333335,0.18707694,0.16082053,0.128,0.09189744,0.052512825,0.02297436,0.006564103,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.006564103,0.013128206,0.009846155,0.0032820515,0.006564103,0.01969231,0.118153855,0.26912823,0.33476925,0.06564103,0.0,0.0032820515,0.098461546,0.45292312,0.32820517,0.2231795,0.16738462,0.15097436,0.14112821,0.20020515,0.16738462,0.18051283,0.33476925,0.67610264,0.65312827,0.4955898,0.37743592,0.32164106,0.20020515,0.10502565,0.1148718,0.08533334,0.009846155,0.052512825,0.09189744,0.098461546,0.09189744,0.068923086,0.0032820515,0.013128206,0.01969231,0.032820515,0.04594872,0.032820515,0.049230773,0.08861539,0.08533334,0.03938462,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.032820515,0.03938462,0.118153855,0.068923086,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016410258,0.055794876,0.12143591,0.068923086,0.049230773,0.068923086,0.13456412,0.25271797,0.39712822,0.61374366,0.73517954,0.7417436,0.7581539,0.78769237,0.80738467,0.8205129,0.8369231,0.892718,0.955077,0.8205129,0.60389745,0.40369233,0.318359,0.21333335,0.190359,0.21333335,0.3249231,0.6465641,0.8172308,0.8172308,0.83035904,0.8992821,0.9124103,0.8730257,0.85005134,0.9189744,1.0633847,1.1618463,1.1552821,1.214359,1.2996924,1.4178462,1.6082052,1.9331284,2.0151796,2.1267693,2.3072822,2.359795,2.6880002,2.9472823,2.8291285,2.3072822,1.6475899,1.6935385,1.4998976,1.3653334,1.3587693,1.3357949,0.93866676,0.702359,0.65641034,0.7811283,1.020718,1.591795,1.7329233,1.8018463,1.6968206,0.8566154,0.4660513,0.24615386,0.15425642,0.12471796,0.108307704,0.08533334,0.07876924,0.06564103,0.052512825,0.049230773,0.049230773,0.055794876,0.059076928,0.059076928,0.072205134,0.118153855,0.16410258,0.20348719,0.23630771,0.26584616,0.30851284,0.34789747,0.38728207,0.41682056,0.43323082,0.4201026,0.38400003,0.35446155,0.34133336,0.3446154,0.4594872,0.5218462,0.56451285,0.6301539,0.76800007,0.702359,0.5349744,0.43323082,0.4135385,0.3511795,0.42994875,0.48246157,0.44964105,0.3708718,0.38728207,0.34789747,0.3511795,0.40369233,0.45620516,0.39384618,0.40697438,0.4004103,0.35774362,0.28225642,0.20676924,0.27569234,0.29538465,0.25271797,0.19364104,0.21333335,0.26584616,0.34133336,0.4397949,0.56123084,0.6826667,0.6235898,0.56451285,0.5284103,0.49230772,0.40697438,0.5021539,0.108307704,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.016410258,0.013128206,0.013128206,0.0032820515,0.009846155,0.036102567,0.068923086,0.14441027,0.2100513,0.23958977,0.22646156,0.18707694,0.22646156,0.30851284,0.29538465,0.19364104,0.18707694,0.055794876,0.013128206,0.006564103,0.009846155,0.01969231,0.072205134,0.7253334,1.654154,2.5764105,3.245949,4.388103,5.586052,6.4754877,7.3616414,9.209436,11.575796,15.366566,18.582975,20.785233,23.095797,26.095592,26.486156,25.800207,25.104412,24.986258,24.01149,24.467693,25.731283,27.319798,28.8919,31.136824,33.65744,34.904617,34.47467,33.106052,34.435284,39.171284,42.824207,45.026466,49.54585,51.459286,49.67385,46.01108,41.216003,34.95385,29.213541,22.761028,16.915693,12.763899,11.142565,9.015796,8.293744,8.4283085,9.255385,11.021129,8.907488,8.182155,7.9786673,7.75877,7.2992826,6.3245134,6.308103,6.1013336,5.290667,4.204308,3.8465643,4.565334,6.0783596,7.719385,8.457847,8.753231,8.093539,6.8627696,6.4754877,9.370257,8.920616,7.177847,7.204103,8.825437,8.664616,8.612103,6.442667,4.818052,4.7917953,5.8125134,14.336001,12.288001,6.1046157,1.8642052,5.297231,10.8996935,11.1064625,8.953437,6.055385,2.605949,1.4145643,0.78769237,0.5284103,0.5415385,0.8467693,1.3029745,1.3554872,1.2668719,1.142154,0.9321026,0.8172308,1.9167181,3.7316926,4.9460516,3.4297438,1.9593848,2.1267693,2.2121027,1.6902566,1.2373334,1.1749744,0.9944616,0.9616411,1.1618463,1.5031796,1.4112822,0.92553854,0.69907695,0.81394875,0.79097444,0.88943595,0.60061544,0.48902568,0.88287187,1.8642052,1.1191796,0.47589746,0.3249231,0.7122052,1.3292309,1.5425643,1.657436,1.9232821,2.3040001,2.4681027,2.3335385,2.9965131,4.2338467,5.356308,5.1954875,3.7842054,3.0096412,3.4002054,4.5554876,5.169231,3.0227695,2.2022567,2.038154,2.0118976,1.7591796,1.024,1.2209232,2.1825643,2.9604106,1.8051283,0.93866676,1.4605129,2.225231,2.3991797,1.4572309,0.96492314,0.79425645,2.409026,4.95918,5.284103,3.062154,3.2131286,2.9407182,1.8740515,2.041436,5.970052,6.2588725,4.565334,2.6847181,2.540308,2.3204105,2.5993848,3.2131286,3.9680004,4.6112823,7.6176414,8.395488,6.567385,4.1025643,5.293949,8.362667,8.172308,6.1440005,3.5840003,1.7132308,5.1626673,7.0925136,7.6668725,7.6931286,8.641642,11.533129,11.697231,12.530872,15.891693,22.111181,20.89354,13.121642,7.7325134,6.885744,5.970052,4.460308,4.4767184,3.442872,2.5961027,6.987488,10.043077,6.87918,3.4822567,3.5872824,8.684308,24.736822,23.512617,16.708925,10.673231,6.409847,10.223591,10.827488,9.363693,7.197539,5.914257,10.016821,12.455385,11.204924,7.1515903,4.092718,3.0949745,2.8947694,3.2853336,4.450462,6.9645133,4.8311796,4.5817437,8.674462,12.566976,4.716308,3.2853336,4.4077954,5.805949,6.1407185,5.0149746,10.952206,13.860104,11.867898,7.5979495,8.169026,8.533334,7.076103,9.432616,12.839386,6.1440005,4.841026,7.076103,9.708308,9.714872,4.2174363,7.312411,9.924924,8.470975,4.8344617,6.3310776,4.0369234,4.082872,7.4174366,11.162257,8.648206,6.055385,6.738052,8.283898,8.231385,4.0467696,3.4592824,4.128821,4.1222568,3.4231799,3.9286156,4.9887185,5.98318,8.251078,11.388719,13.249642,32.12472,33.234055,30.352413,25.301334,7.9261546,19.584002,39.87036,44.389748,30.900515,19.321438,15.553642,14.621539,17.424412,19.93518,13.174155,13.696001,16.528412,15.104001,9.67877,7.3452315,7.24677,5.687795,5.7074876,7.525744,8.536616,7.433847,7.259898,5.8978467,3.69559,3.4658465,1.847795,1.1979488,1.1323078,1.3259488,1.4966155,1.3357949,0.86974365,0.38728207,0.08861539,0.049230773,0.032820515,0.016410258,0.006564103,0.0,0.0,0.0,0.013128206,0.02297436,0.029538464,0.036102567,0.032820515,0.08205129,0.068923086,0.032820515,0.16410258,1.1520001,0.7122052,0.15753847,0.02297436,0.059076928,0.118153855,0.13784617,0.13784617,0.15753847,0.23958977,0.19364104,0.16082053,0.13784617,0.190359,0.45620516,0.9321026,1.3128207,1.270154,0.79425645,0.17723078,0.13128206,0.2100513,0.3117949,0.380718,0.42338464,0.3446154,0.27241027,0.19364104,0.12471796,0.13456412,0.04594872,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.013128206,0.009846155,0.029538464,0.013128206,0.02297436,0.07876924,0.15097436,0.07548718,0.02297436,0.0,0.06564103,0.3249231,0.38400003,0.37743592,0.3446154,0.27241027,0.101743594,0.128,0.14769232,0.20676924,0.32820517,0.5284103,0.45292312,0.3117949,0.23302566,0.24615386,0.3052308,0.256,0.24615386,0.17723078,0.059076928,0.04266667,0.09189744,0.12143591,0.12471796,0.09189744,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0032820515,0.009846155,0.009846155,0.006564103,0.02297436,0.02297436,0.009846155,0.0,0.0,0.013128206,0.016410258,0.02297436,0.029538464,0.04594872,0.029538464,0.02297436,0.02297436,0.029538464,0.02297436,0.15425642,0.25271797,0.17723078,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.02297436,0.06235898,0.052512825,0.04266667,0.055794876,0.101743594,0.17723078,0.2855385,0.46276927,0.62030774,0.7450257,0.8763078,0.8205129,0.85005134,0.9189744,0.9911796,1.0436924,1.0896411,0.9878975,0.86974365,0.72861546,0.43323082,0.25271797,0.20348719,0.2231795,0.318359,0.55794877,0.6498462,0.7253334,0.8369231,0.9419488,0.88287187,0.83035904,0.81066674,0.9189744,1.148718,1.3686155,1.2964103,1.2603078,1.2898463,1.3587693,1.404718,1.6049232,1.6672822,1.6771283,1.7460514,2.0184617,2.1891284,2.5829747,2.7963078,2.6880002,2.3630772,2.1464617,2.0873847,1.913436,1.5819489,1.2537436,0.955077,0.7318975,0.61374366,0.62030774,0.76800007,1.0535386,1.3161026,1.5622566,1.6410258,1.2504616,0.73517954,0.39712822,0.2231795,0.17066668,0.16082053,0.13784617,0.12143591,0.08533334,0.04266667,0.036102567,0.036102567,0.04594872,0.049230773,0.04594872,0.052512825,0.08205129,0.108307704,0.13784617,0.16738462,0.19692309,0.25928208,0.30851284,0.34789747,0.39384618,0.44964105,0.48902568,0.4201026,0.33805132,0.28882053,0.2855385,0.37743592,0.44307697,0.49887183,0.571077,0.6662565,0.7122052,0.64000005,0.60061544,0.5973334,0.48902568,0.43651286,0.42994875,0.40369233,0.36430773,0.3708718,0.39056414,0.40369233,0.43323082,0.46933338,0.46933338,0.5349744,0.512,0.4397949,0.34133336,0.25271797,0.26256412,0.24287182,0.19692309,0.15097436,0.14112821,0.15097436,0.23630771,0.35774362,0.47917953,0.56451285,0.636718,0.61374366,0.5349744,0.46933338,0.47589746,1.6213335,0.36430773,0.01969231,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.02297436,0.055794876,0.068923086,0.16738462,0.20676924,0.190359,0.14769232,0.13784617,0.23958977,0.3446154,0.36102566,0.27897438,0.18051283,0.03938462,0.006564103,0.006564103,0.0032820515,0.0,0.032820515,0.36102566,0.9616411,1.6705642,2.166154,3.4231799,4.6080003,5.405539,6.0258465,7.1909747,9.83959,13.863386,16.443079,16.978052,17.096207,19.623386,21.385847,21.904411,21.622156,21.897848,23.519182,24.582565,26.003695,27.621746,28.196104,27.559387,29.377644,31.097439,31.947489,32.938667,37.041233,42.725746,47.412518,49.79857,49.85108,47.379696,42.292515,37.060925,32.68923,28.708105,22.938257,17.522873,13.095386,10.079181,8.687591,7.4174366,7.030154,8.585847,10.8996935,10.555078,8.362667,7.765334,7.578257,7.680001,9.009232,7.2861543,5.9995904,6.189949,6.7807183,4.565334,3.767795,4.266667,6.0225644,8.208411,9.216001,8.910769,7.6701546,6.160411,6.009436,9.787078,11.303386,7.6734366,5.937231,7.762052,9.4457445,10.033232,6.76759,4.2568207,4.414359,6.449231,13.223386,14.053744,9.061745,2.4057438,2.2514873,4.6112823,7.584821,8.723693,7.0793853,3.2361028,1.785436,0.9124103,0.574359,0.60389745,0.7056411,0.90912825,0.90912825,0.7581539,0.6498462,0.92553854,1.1388719,2.0742567,3.498667,4.562052,3.7710772,2.7241027,2.6912823,2.605949,2.1464617,1.7165129,1.5097437,1.1552821,0.72861546,0.48574364,0.8467693,1.017436,0.8566154,0.69579494,0.8008206,1.3587693,1.142154,0.6465641,0.5513847,1.0633847,1.913436,1.3259488,0.7253334,0.43651286,0.5907693,1.1060513,1.3029745,1.6607181,1.9823592,2.2153847,2.4451284,2.1891284,2.6847181,3.6594875,5.044513,7.003898,5.0084105,3.8006158,4.2830772,5.605744,5.1626673,3.1245131,2.4352822,2.2055387,2.03159,1.9954873,1.5064616,1.1060513,2.0020514,3.3969233,2.4910772,1.1552821,0.9419488,0.9682052,0.98461545,1.3751796,1.0699488,0.79097444,1.7952822,3.121231,1.5786668,2.4746668,3.629949,3.2328207,2.0841026,3.6168208,6.5345645,6.2752824,4.6966157,3.948308,6.4689236,4.890257,3.2886157,2.487795,2.6420515,3.2328207,4.84759,5.536821,4.6900516,3.121231,3.0687182,5.835488,7.2336416,6.6100516,4.332308,1.7657437,4.6145644,5.723898,5.9536414,6.6494365,9.632821,12.087796,11.441232,10.994873,13.5318985,21.32677,20.09272,12.153437,6.882462,6.2916927,5.028103,3.006359,1.7723079,1.332513,2.681436,7.8014364,8.536616,5.927385,4.6802053,6.1046157,8.136206,27.90072,21.024822,10.601027,6.445949,5.113436,4.57518,7.1647186,9.045334,8.320001,5.034667,9.442462,10.768411,9.475283,6.4032826,2.7864618,1.7887181,1.8149745,2.353231,3.5872824,6.38359,5.943795,6.8496413,9.869129,11.930258,6.1407185,4.2141542,4.023795,5.182359,6.810257,7.5454364,16.28554,13.787898,8.576,6.163693,9.07159,8.864821,6.9021544,7.958975,11.257437,10.456616,5.179077,7.1187696,10.43036,10.843898,5.681231,6.311385,10.781539,9.435898,3.692308,6.045539,6.6560006,7.076103,7.571693,7.4436927,5.034667,5.4416413,7.24677,8.78277,8.267488,3.8400004,2.934154,3.9220517,4.59159,4.4307694,4.6244106,3.6036925,5.435077,8.073847,9.685334,8.641642,22.28513,26.925951,27.421541,24.38236,14.152206,34.89149,62.759388,75.66441,68.174774,51.538055,42.610874,37.9799,36.07303,32.256004,18.802874,18.6519,19.492104,16.06236,9.7903595,8.786052,7.4141545,5.651693,5.989744,7.8506675,7.571693,6.810257,7.3649235,6.2720003,3.7415388,3.1606157,1.9035898,1.4539489,1.2570257,1.1290257,1.270154,1.5491283,1.0896411,0.50543594,0.13456412,0.029538464,0.013128206,0.009846155,0.006564103,0.0,0.0,0.0032820515,0.013128206,0.016410258,0.016410258,0.01969231,0.016410258,0.08205129,0.108307704,0.07548718,0.06564103,0.54482055,0.30851284,0.04266667,0.0032820515,0.009846155,0.016410258,0.032820515,0.08861539,0.18379489,0.28882053,0.21333335,0.18707694,0.17394873,0.18379489,0.2855385,0.48574364,0.96492314,1.2077949,0.96492314,0.24943592,0.10502565,0.11158975,0.23630771,0.39056414,0.42338464,0.41682056,0.45620516,0.3708718,0.190359,0.14769232,0.072205134,0.036102567,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.016410258,0.036102567,0.016410258,0.0032820515,0.009846155,0.02297436,0.08861539,0.04266667,0.0,0.02297436,0.118153855,0.30194873,0.46933338,0.5874872,0.5874872,0.36430773,0.4594872,0.4660513,0.49230772,0.5513847,0.57764107,0.47589746,0.35774362,0.2855385,0.2986667,0.39712822,0.3708718,0.33805132,0.24287182,0.1148718,0.049230773,0.06235898,0.08861539,0.101743594,0.08533334,0.006564103,0.0,0.0,0.0032820515,0.006564103,0.006564103,0.0,0.0,0.0,0.0,0.0,0.032820515,0.026256412,0.009846155,0.0,0.0,0.006564103,0.013128206,0.02297436,0.029538464,0.04594872,0.036102567,0.03938462,0.03938462,0.029538464,0.016410258,0.098461546,0.21661541,0.17394873,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.02297436,0.032820515,0.032820515,0.04594872,0.08533334,0.14112821,0.20348719,0.33805132,0.49887183,0.69579494,0.9747693,0.9189744,0.9353847,0.9878975,1.0601027,1.1520001,1.2471796,1.2176411,1.1454359,0.9944616,0.5874872,0.36758977,0.27569234,0.256,0.29538465,0.41682056,0.5218462,0.7089231,0.92553854,1.0633847,0.9321026,0.86974365,0.88287187,1.0108719,1.214359,1.3883078,1.270154,1.3357949,1.5261539,1.7165129,1.719795,1.6738462,1.654154,1.5753847,1.5031796,1.6640002,1.8445129,2.231795,2.5140514,2.6223593,2.740513,2.3696413,2.422154,2.3630772,2.0250258,1.6147693,1.1093334,0.77456415,0.571077,0.4955898,0.56123084,0.67282057,0.9517949,1.2209232,1.3850257,1.4408206,1.0305642,0.60061544,0.32820517,0.23630771,0.2231795,0.18379489,0.16082053,0.1148718,0.059076928,0.036102567,0.036102567,0.04266667,0.049230773,0.055794876,0.06564103,0.06564103,0.072205134,0.08533334,0.10502565,0.128,0.18051283,0.24943592,0.31507695,0.37415388,0.43651286,0.47589746,0.40369233,0.31507695,0.25928208,0.256,0.28882053,0.3446154,0.41682056,0.47589746,0.4955898,0.60389745,0.702359,0.764718,0.7778462,0.7318975,0.6170257,0.49887183,0.39712822,0.32820517,0.3117949,0.4004103,0.46276927,0.508718,0.5513847,0.58092314,0.65641034,0.62030774,0.5218462,0.4135385,0.31507695,0.27897438,0.24287182,0.190359,0.13456412,0.108307704,0.098461546,0.14441027,0.23958977,0.34789747,0.42338464,0.5349744,0.56451285,0.5218462,0.46933338,0.49887183,2.550154,0.6432821,0.068923086,0.0032820515,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01969231,0.04266667,0.049230773,0.013128206,0.06564103,0.06235898,0.03938462,0.03938462,0.09189744,0.20020515,0.3117949,0.36102566,0.29538465,0.052512825,0.02297436,0.013128206,0.013128206,0.013128206,0.0,0.08205129,0.256,0.65641034,1.1618463,1.3686155,2.609231,3.7349746,4.4964104,4.9526157,5.4613338,8.057437,10.794667,12.340514,12.665437,13.02318,14.831591,17.165129,18.31713,18.602669,20.36513,23.40759,24.339695,24.802464,25.393232,25.665644,25.45231,27.401848,31.130259,35.862976,40.438156,44.5079,47.980312,49.65744,48.24944,42.368004,37.53026,32.817234,28.970669,26.112001,23.742361,17.352207,12.911591,9.521232,7.0400004,6.058667,5.930667,6.2194877,9.475283,13.279181,10.256411,7.9819493,7.1909747,6.678975,6.695385,8.920616,7.194257,6.226052,6.8233852,7.578257,4.8607183,4.086154,4.4800005,5.5926156,6.616616,6.3934364,6.0258465,6.5444107,6.6494365,6.1997952,6.1997952,8.083693,6.380308,6.294975,8.267488,7.962257,6.7840004,5.0904617,4.017231,4.066462,5.1265645,14.224411,15.02195,10.28595,4.5095387,3.9023592,2.9144619,3.5478978,4.7261543,5.113436,3.114667,1.9790771,1.086359,0.6498462,0.6170257,0.6892308,0.5152821,0.48902568,0.5874872,0.83035904,1.2504616,1.5819489,2.3401027,3.5971284,5.0051284,5.792821,4.8114877,3.764513,2.7831798,1.9659488,1.3554872,1.276718,0.9911796,0.6498462,0.5481026,1.1093334,1.273436,1.0568206,0.8402052,1.0962052,2.422154,1.7427694,1.1716924,1.1224617,1.4145643,1.2800001,1.1191796,0.8763078,0.702359,0.636718,0.5973334,0.8730257,2.044718,2.6190772,2.4713848,2.861949,1.9889232,2.412308,3.318154,4.821334,7.939283,6.616616,4.906667,5.3924108,7.066257,5.3136415,3.3345644,2.934154,2.9046156,2.8324106,3.0851285,2.556718,1.5753847,2.3072822,4.023795,3.0982566,1.8149745,1.404718,1.0666667,0.86974365,1.7624617,1.401436,1.2242053,1.5425643,1.8576412,0.84348726,2.1398976,3.5774362,3.186872,2.4549747,6.3277955,8.119796,7.4075904,6.373744,7.145026,11.782565,8.195283,4.6834874,2.917744,3.0523078,3.69559,3.7087183,3.186872,2.5042052,2.0053334,2.0020514,3.3608208,5.3070774,6.193231,5.3366156,3.0227695,4.1222568,4.056616,4.0992823,5.5597954,9.787078,10.850462,9.45559,7.3058467,6.7544622,10.794667,10.9226675,7.6734366,5.9634876,6.012718,3.31159,2.412308,2.0873847,2.5042052,4.20759,8.113232,6.8627696,6.0849237,7.318975,9.16677,7.315693,17.801847,11.283693,5.5729237,5.723898,4.0041027,1.9495386,5.651693,9.360411,9.265231,3.5052311,3.4855387,4.4734364,4.4110775,2.9046156,1.2373334,1.0535386,1.0929232,1.5163078,2.103795,2.2678976,7.6734366,8.910769,9.176616,9.045334,6.4590774,4.276513,3.7021542,4.5587697,7.072821,11.88759,16.827078,12.616206,8.316719,7.650462,8.992821,8.093539,6.5312824,7.637334,12.087796,17.877335,7.50277,7.3583593,10.906258,12.727796,8.530052,7.1614366,10.965334,9.609847,3.515077,3.8695388,9.005949,11.424822,9.714872,5.7042055,4.4800005,6.6527185,8.720411,9.29477,7.8014364,4.466872,2.0545642,3.1409233,4.417641,4.706462,4.969026,3.5216413,5.2053337,7.7357955,9.091283,7.4896417,17.539284,22.393438,22.852924,21.169233,21.034668,51.6759,86.87262,109.88965,112.34134,94.23098,79.52739,69.10688,60.150158,47.980312,26.059488,20.98872,19.081848,15.074463,9.777231,10.066052,8.136206,6.442667,6.7905645,8.021334,5.98318,6.554257,6.193231,5.0215387,3.6135387,3.0227695,2.1333334,1.8904617,1.6410258,1.2274873,1.0010257,1.9429746,1.3915899,0.60061544,0.16410258,0.026256412,0.006564103,0.0,0.0,0.0,0.0032820515,0.016410258,0.016410258,0.013128206,0.013128206,0.013128206,0.016410258,0.059076928,0.12471796,0.17066668,0.14112821,0.03938462,0.0032820515,0.0,0.0032820515,0.013128206,0.02297436,0.01969231,0.055794876,0.14112821,0.25271797,0.21661541,0.18707694,0.17394873,0.2100513,0.33476925,0.26584616,0.47917953,0.7417436,0.77128214,0.24615386,0.101743594,0.1148718,0.25928208,0.41025645,0.3446154,0.45620516,0.65312827,0.6104616,0.33476925,0.15425642,0.13456412,0.09189744,0.052512825,0.029538464,0.032820515,0.02297436,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.013128206,0.013128206,0.0032820515,0.006564103,0.016410258,0.02297436,0.08205129,0.03938462,0.0,0.0,0.0,0.14769232,0.40369233,0.67938465,0.83035904,0.67610264,0.86646163,0.8763078,0.8467693,0.7975385,0.6170257,0.5677949,0.5284103,0.508718,0.4955898,0.45620516,0.40697438,0.35446155,0.26584616,0.15425642,0.09189744,0.06564103,0.072205134,0.08861539,0.08205129,0.016410258,0.0032820515,0.0,0.0032820515,0.013128206,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.01969231,0.013128206,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.032820515,0.032820515,0.013128206,0.013128206,0.0032820515,0.0032820515,0.006564103,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.02297436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.013128206,0.02297436,0.036102567,0.06564103,0.1148718,0.17066668,0.24615386,0.36758977,0.58420515,0.96492314,1.0436924,1.0601027,1.0469744,1.0568206,1.1651284,1.3981539,1.4473847,1.339077,1.1093334,0.78769237,0.571077,0.39056414,0.27897438,0.25928208,0.34789747,0.45620516,0.6826667,0.9517949,1.1552821,1.1290257,1.0436924,1.0502565,1.0994873,1.1454359,1.1585642,1.1881026,1.5327181,1.913436,2.1530259,2.1924105,2.0676925,1.9922053,1.9167181,1.7952822,1.5753847,1.7952822,2.034872,2.1300514,2.1825643,2.5698464,2.4385643,2.487795,2.4910772,2.3762052,2.1891284,1.3883078,0.8598975,0.55794877,0.43323082,0.43651286,0.5481026,0.74830776,0.9944616,1.2176411,1.3423591,1.270154,0.8598975,0.49887183,0.32820517,0.28225642,0.2231795,0.21333335,0.18707694,0.13128206,0.06564103,0.055794876,0.055794876,0.055794876,0.068923086,0.098461546,0.068923086,0.06235898,0.06235898,0.06564103,0.08533334,0.10502565,0.18707694,0.27569234,0.3446154,0.38400003,0.39056414,0.33805132,0.2986667,0.27897438,0.23958977,0.25271797,0.256,0.28225642,0.33476925,0.38400003,0.44964105,0.6892308,0.85005134,0.892718,0.9911796,0.94523084,0.72861546,0.47589746,0.29210258,0.24615386,0.34133336,0.43651286,0.54482055,0.6432821,0.6629744,0.7056411,0.6826667,0.5973334,0.47261542,0.3708718,0.3249231,0.2986667,0.2297436,0.13784617,0.10502565,0.08533334,0.098461546,0.13128206,0.19364104,0.28882053,0.34789747,0.41025645,0.45292312,0.46276927,0.44307697,1.404718,0.5973334,0.17723078,0.01969231,0.0,0.0,0.0,0.009846155,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.055794876,0.072205134,0.036102567,0.0,0.02297436,0.02297436,0.009846155,0.01969231,0.09189744,0.055794876,0.38400003,0.3708718,0.016410258,0.016410258,0.016410258,0.006564103,0.006564103,0.013128206,0.0,0.072205134,0.19364104,0.39384618,0.73517954,1.2964103,2.6157951,3.9712822,5.5072823,7.499488,10.345026,11.992617,13.321847,14.102976,14.815181,16.646564,17.19795,16.49231,16.584206,17.851078,18.996513,20.683489,21.231592,21.274258,21.454771,22.42954,23.762053,28.248617,33.14544,37.973335,44.54072,47.89826,46.28349,42.804516,38.583797,32.76144,29.623796,27.392002,25.317745,22.6199,18.49436,11.779283,7.9327188,6.373744,6.117744,5.7534366,5.605744,7.3550773,9.321027,9.596719,6.058667,5.421949,5.172513,5.654975,6.186667,5.0510774,7.066257,6.7905645,6.875898,7.1187696,4.4701543,5.58277,9.265231,13.092104,14.50995,10.84718,9.93477,17.010874,21.208616,18.297438,10.679795,5.297231,4.7589746,7.899898,10.256411,4.0434875,2.4451284,2.2744617,2.3729234,2.4648206,3.1737437,13.354668,12.760616,8.694155,6.514872,9.626257,5.2709746,2.4681027,1.1323078,0.9419488,1.3587693,1.0896411,0.85005134,0.7581539,0.7384616,0.51856416,0.67610264,0.9747693,1.529436,2.166154,2.412308,2.5074873,3.1934361,4.8082056,7.3550773,10.466462,7.9163084,5.2742567,3.0326157,1.4998976,0.79425645,1.1355898,0.94523084,0.83035904,1.0732309,1.6475899,1.5753847,1.1618463,0.85005134,0.9714873,1.7394873,1.9462565,2.4943593,2.5435898,1.913436,1.083077,0.827077,0.8730257,0.9353847,0.84348726,0.5481026,1.1848207,2.6880002,3.5807183,3.4494362,2.9604106,2.5435898,2.2777438,2.8882053,4.3749747,6.012718,7.4043083,6.452513,6.885744,8.388924,6.6067696,4.4340515,3.8367183,3.4691284,3.121231,3.7087183,3.170462,2.3401027,2.7503593,3.9647183,3.5872824,2.2416413,2.0184617,1.7920002,1.3128207,1.1913847,1.3259488,1.5491283,1.8609232,2.0151796,1.5261539,3.2229745,5.5958977,5.546667,4.056616,6.180103,7.2894363,7.6964107,6.994052,6.1308722,7.4010262,4.2994876,2.353231,2.5731285,4.5390773,6.3934364,6.2588725,5.100308,3.9351797,3.1113849,2.3204105,2.5271797,3.9417439,5.3891287,5.927385,4.850872,3.764513,3.2098465,3.498667,4.4767184,5.540103,5.477744,7.200821,7.5191803,5.7403083,3.6791797,4.568616,8.224821,10.06277,7.936001,2.1530259,2.3466668,3.2098465,5.0543594,6.941539,6.698667,8.247795,10.7158985,11.237744,9.95118,9.964309,7.6570263,8.070564,10.020103,10.486155,4.578462,1.8182565,3.764513,8.418462,11.625027,7.0957956,4.007385,2.934154,2.1989746,1.3456411,1.1126155,1.2242053,1.020718,0.86317956,1.5360001,4.2568207,13.6697445,8.4512825,3.5544617,3.9089234,4.4110775,3.5905645,5.4482055,8.408616,12.438975,19.042463,8.569437,5.858462,7.683283,9.8592825,7.24677,8.12636,7.138462,7.2369237,10.883283,20.050053,9.245539,6.738052,8.3364105,10.545232,10.545232,9.701744,12.209231,11.972924,7.5552826,2.1989746,8.740103,10.230155,8.556309,6.432821,7.384616,9.216001,9.45559,9.153642,7.8112826,3.3575387,2.612513,4.844308,5.8814363,5.139693,5.61559,5.0642056,5.0477953,7.8736415,11.808822,11.076924,20.404514,21.00513,18.326975,18.107079,26.38113,57.206158,83.96144,100.23714,102.334366,89.31119,76.73437,71.7358,66.28431,54.682262,33.552414,23.93272,21.842052,17.624617,10.564924,8.881231,7.9786673,7.768616,8.910769,9.892103,7.0334363,6.5083084,5.3727183,5.4153852,6.0225644,4.1813335,2.7175386,2.4057438,2.1530259,1.7099489,1.6475899,2.4549747,1.6114873,0.60389745,0.11158975,0.016410258,0.0032820515,0.0,0.0,0.0032820515,0.016410258,0.026256412,0.02297436,0.009846155,0.013128206,0.06235898,0.036102567,0.049230773,0.07876924,0.09189744,0.029538464,0.006564103,0.0,0.0,0.013128206,0.06235898,0.12143591,0.06564103,0.016410258,0.032820515,0.108307704,0.16738462,0.14769232,0.16410258,0.27569234,0.45620516,0.3117949,0.28225642,0.29538465,0.28225642,0.19692309,0.101743594,0.15097436,0.36430773,0.6268718,0.6859488,0.6629744,0.6826667,0.6662565,0.571077,0.4135385,0.30194873,0.17394873,0.118153855,0.14441027,0.16738462,0.108307704,0.04594872,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.006564103,0.0,0.0,0.0,0.0,0.0,0.013128206,0.02297436,0.0,0.0,0.0,0.006564103,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.04594872,0.26584616,0.5546667,0.58092314,0.4955898,0.65641034,0.73517954,0.64000005,0.51856416,0.46933338,0.61374366,0.7778462,0.8369231,0.702359,0.54482055,0.38400003,0.256,0.17723078,0.15097436,0.17723078,0.2100513,0.21661541,0.16082053,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.016410258,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.055794876,0.108307704,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.016410258,0.029538464,0.09189744,0.16410258,0.20020515,0.24943592,0.37743592,0.67282057,0.97805136,1.1093334,1.0896411,1.020718,1.0666667,1.4966155,1.5556924,1.4408206,1.2504616,1.0075898,0.81066674,0.48902568,0.29210258,0.2986667,0.39712822,0.36102566,0.37743592,0.56123084,0.92225647,1.3718976,1.1913847,1.1093334,1.0272821,0.9878975,1.1585642,1.5885129,1.7755898,1.6049232,1.2635899,1.2504616,1.5556924,2.034872,2.297436,2.2580514,2.1366155,2.15959,1.9659488,1.7591796,1.7394873,2.1070771,2.678154,2.740513,2.4549747,2.0545642,1.847795,1.5031796,1.0994873,0.761436,0.54482055,0.4135385,0.43651286,0.49887183,0.69251287,0.9288206,0.9156924,1.2832822,1.1454359,0.79097444,0.46276927,0.36758977,0.32820517,0.36758977,0.38400003,0.32164106,0.13784617,0.101743594,0.09189744,0.07876924,0.072205134,0.12143591,0.12143591,0.0951795,0.068923086,0.06235898,0.06235898,0.06235898,0.1148718,0.20020515,0.2986667,0.39712822,0.46933338,0.37743592,0.34133336,0.37415388,0.28882053,0.25271797,0.23630771,0.24615386,0.27569234,0.27569234,0.3117949,0.5481026,0.76800007,0.9189744,1.1126155,1.2242053,1.0666667,0.761436,0.45620516,0.32164106,0.24615386,0.26584616,0.37415388,0.5284103,0.6268718,0.6498462,0.74830776,0.7220513,0.5677949,0.45620516,0.4201026,0.4397949,0.3708718,0.22646156,0.15097436,0.1148718,0.108307704,0.11158975,0.14441027,0.2297436,0.27897438,0.30851284,0.3446154,0.3708718,0.32164106,1.024,0.56123084,0.2100513,0.055794876,0.049230773,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.013128206,0.006564103,0.0,0.032820515,0.01969231,0.0032820515,0.006564103,0.029538464,0.032820515,0.0951795,0.08533334,0.016410258,0.026256412,0.016410258,0.006564103,0.006564103,0.013128206,0.0,0.013128206,0.11158975,0.22646156,0.38728207,0.7220513,1.522872,3.2098465,5.5171285,8.274052,11.418258,14.982565,17.555695,18.95713,18.87836,16.89272,15.048206,14.001232,13.883078,14.54277,15.543797,17.32595,18.786463,20.896822,23.670156,26.14154,30.8119,35.410053,39.522465,42.98831,45.89621,42.57477,38.006157,33.414566,29.535181,26.633848,25.38995,24.503798,20.630976,14.086565,8.825437,7.640616,8.057437,8.182155,7.381334,6.301539,5.658257,6.7905645,7.975385,8.484103,8.595693,6.701949,4.8836927,4.673641,6.6592827,10.496001,10.020103,9.196308,7.6701546,6.1308722,6.314667,10.587898,12.432411,11.057232,7.936001,6.820103,4.9788723,5.7796926,7.318975,8.093539,7.020308,3.5610259,2.930872,5.2414365,7.4797955,3.4822567,1.4539489,1.2176411,1.9528207,3.4330258,6.055385,7.650462,7.062975,5.172513,3.3772311,3.6102567,2.484513,1.332513,0.6498462,0.5481026,0.74830776,0.81066674,0.6104616,0.5284103,0.6498462,0.761436,1.2537436,1.719795,2.3040001,2.6289232,1.8018463,2.2482052,3.2918978,4.8114877,7.017026,10.443488,8.283898,5.85518,3.9351797,2.8356924,2.3794873,2.0578463,1.4966155,0.9944616,0.80738467,1.148718,1.0633847,1.2373334,1.4473847,1.6672822,2.0578463,2.294154,2.356513,2.484513,2.3335385,0.98461545,0.90584624,1.6311796,2.0873847,1.7296412,0.5481026,0.84348726,2.3630772,3.6660516,4.1583595,4.1189747,4.056616,4.2207184,3.8498464,3.367385,4.388103,4.2272825,4.394667,6.0356927,8.12636,7.4863596,4.7556925,4.9329233,5.0576415,4.2436924,3.7087183,3.629949,2.7536411,3.436308,4.9394875,3.4264617,1.7920002,1.148718,1.9200002,3.3772311,3.6562054,3.564308,3.6693337,3.7316926,3.3411283,1.9167181,4.0434875,7.958975,9.386667,7.860513,6.741334,6.298257,6.491898,6.5280004,6.114462,5.4613338,4.84759,4.089436,4.8836927,6.633026,6.416411,7.131898,6.6560006,5.395693,3.9154875,2.917744,1.6705642,1.5491283,2.2219489,3.4034874,4.8771286,5.2447186,4.086154,3.2984617,3.1967182,2.5107694,2.1956925,6.4656415,9.258667,9.032206,8.756514,11.1983595,12.583385,10.092308,5.346462,4.4340515,5.2447186,8.664616,12.035283,13.46954,11.848206,13.692719,11.096616,7.381334,4.8607183,4.8607183,4.70318,10.259693,12.763899,9.862565,5.61559,3.170462,2.5435898,4.2830772,7.062975,7.680001,5.6385646,4.7589746,3.3411283,1.6443079,1.8707694,1.5327181,1.1290257,2.7831798,5.868308,7.026872,4.5062566,2.6978464,3.639795,5.986462,5.031385,3.9909747,5.9930263,11.851488,17.14872,12.268309,6.3442054,6.941539,8.920616,9.133949,6.4065647,5.789539,4.788513,5.664821,9.419488,15.766975,8.615385,4.6178465,5.2545643,8.457847,8.602257,9.508103,11.69395,11.382154,8.260923,5.481026,9.622975,7.640616,5.658257,7.0793853,12.57354,12.304411,11.293539,10.466462,9.317744,5.907693,2.6453335,3.570872,4.519385,4.772103,7.0432825,9.353847,7.532308,4.8311796,3.2656412,3.6069746,7.318975,8.786052,10.893129,15.261539,22.268719,40.231388,57.22585,64.00657,58.98831,48.24944,46.592003,46.208004,41.373543,32.226463,24.77949,17.864206,14.293334,11.936821,9.970873,8.881231,9.393231,9.626257,9.783795,9.616411,8.438154,6.9743595,6.3934364,6.73477,6.928411,4.7917953,2.7109745,2.553436,2.553436,2.0742567,1.6114873,1.6049232,1.0732309,0.45620516,0.052512825,0.0032820515,0.009846155,0.013128206,0.006564103,0.0,0.0032820515,0.026256412,0.02297436,0.009846155,0.006564103,0.036102567,0.052512825,0.029538464,0.026256412,0.03938462,0.01969231,0.0032820515,0.0,0.0,0.02297436,0.108307704,0.16082053,0.23302566,0.29538465,0.27897438,0.059076928,0.059076928,0.07548718,0.12471796,0.21661541,0.36102566,0.28225642,0.2855385,0.25928208,0.18051283,0.12471796,0.055794876,0.39056414,0.90256417,1.4112822,1.785436,1.3587693,1.2964103,1.3620514,1.2898463,0.7778462,0.73517954,0.8533334,1.1552821,1.3357949,0.764718,0.35446155,0.16738462,0.13128206,0.16738462,0.20676924,0.13784617,0.06235898,0.04266667,0.06564103,0.036102567,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0,0.02297436,0.049230773,0.0,0.0,0.006564103,0.029538464,0.052512825,0.036102567,0.055794876,0.06235898,0.052512825,0.036102567,0.02297436,0.032820515,0.16738462,0.15425642,0.0,0.0,0.0,0.009846155,0.052512825,0.11158975,0.1148718,0.098461546,0.190359,0.29210258,0.36102566,0.38400003,0.37415388,0.41682056,0.4660513,0.49230772,0.4955898,0.5021539,0.47917953,0.4201026,0.318359,0.17723078,0.2297436,0.24287182,0.19364104,0.101743594,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.006564103,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.0032820515,0.0,0.0,0.0032820515,0.013128206,0.02297436,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08205129,0.14112821,0.13128206,0.06235898,0.052512825,0.01969231,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.009846155,0.029538464,0.07548718,0.14769232,0.19692309,0.256,0.45292312,0.78769237,1.1224617,1.1979488,1.0305642,0.9353847,1.0305642,1.1749744,1.3817437,1.5524104,1.4834872,1.0633847,0.65312827,0.40369233,0.3446154,0.3708718,0.33476925,0.39056414,0.52512825,0.7581539,1.142154,1.2504616,1.1749744,1.0371283,0.9747693,1.1355898,1.3292309,1.2668719,1.5261539,2.2482052,3.1540515,2.7963078,2.553436,2.4451284,2.3433847,1.9790771,2.3138463,2.3729234,2.0775387,1.6869745,1.8018463,2.2088206,2.550154,2.6912823,2.540308,2.028308,1.8642052,1.4145643,0.98461545,0.7089231,0.5349744,0.4594872,0.4397949,0.47917953,0.5546667,0.6104616,0.90912825,1.142154,1.0666667,0.7187693,0.4266667,0.4201026,0.36102566,0.28225642,0.19692309,0.101743594,0.11158975,0.1148718,0.0951795,0.072205134,0.12143591,0.14112821,0.14769232,0.13784617,0.118153855,0.108307704,0.09189744,0.0951795,0.118153855,0.16082053,0.23958977,0.4201026,0.47261542,0.42338464,0.33805132,0.30194873,0.23630771,0.23958977,0.24287182,0.2297436,0.24943592,0.3052308,0.41025645,0.55794877,0.73517954,0.9321026,1.1979488,1.2931283,1.0601027,0.67282057,0.636718,0.50543594,0.3708718,0.31507695,0.34789747,0.40697438,0.51856416,0.636718,0.6170257,0.48902568,0.45620516,0.39056414,0.35774362,0.3052308,0.23958977,0.21333335,0.13784617,0.12471796,0.13784617,0.14441027,0.14441027,0.17394873,0.23630771,0.3052308,0.3446154,0.29538465,1.782154,1.1552821,0.512,0.6268718,1.2668719,1.1979488,0.23958977,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.013128206,0.006564103,0.013128206,0.068923086,0.17066668,0.15425642,0.07876924,0.009846155,0.029538464,0.10502565,0.049230773,0.0032820515,0.016410258,0.055794876,0.009846155,0.068923086,0.13128206,0.20020515,0.37743592,0.90912825,1.9922053,3.6036925,5.720616,8.320001,11.707078,15.090873,16.774565,16.160822,13.7386675,12.711386,12.097642,12.058257,12.688411,14.020925,15.78995,18.04472,21.80595,26.640411,30.647797,35.19344,39.502773,42.61744,44.00903,43.598774,38.495182,33.686977,30.06031,28.022156,27.480618,26.73231,24.592413,20.496412,15.195899,10.738873,10.706052,11.0375395,10.686359,9.856001,9.990565,12.826258,12.619488,10.131693,7.315693,7.3091288,5.737026,4.637539,6.1013336,9.734565,12.642463,9.590155,8.523488,8.933744,10.9456415,15.317334,13.584412,11.175385,9.104411,8.39877,10.06277,8.103385,6.196513,5.602462,6.1505647,6.2490263,3.9975388,2.9538465,3.2131286,3.6693337,2.0151796,0.77128214,0.9321026,1.7952822,3.1015387,5.0084105,4.634257,4.900103,4.1485133,2.3926156,1.3193847,1.2931283,0.90256417,0.65641034,0.63343596,0.4955898,0.48574364,0.44964105,0.44307697,0.5284103,0.761436,1.3686155,1.6738462,1.9922053,2.2416413,1.9495386,1.8149745,2.03159,2.8882053,4.4701543,6.6560006,6.380308,4.9788723,3.570872,2.5895386,1.7985642,1.4703591,1.0043077,0.6859488,0.65969235,0.93866676,1.1782565,1.2996924,1.4309745,1.6640002,2.0808206,2.2219489,2.2613335,2.5337439,2.5862565,1.1520001,1.020718,1.5097437,1.7427694,1.3456411,0.4397949,0.7056411,1.6311796,2.6026669,3.3247182,3.82359,4.6244106,5.612308,5.3760004,4.4865646,5.4843082,4.069744,3.5544617,4.5423594,6.038975,5.47118,4.0467696,4.8836927,6.3277955,7.3583593,7.581539,5.4941545,4.1714873,4.325744,5.1298466,4.2305646,2.5632823,1.273436,1.2996924,2.5665643,3.9712822,3.9253337,4.650667,6.294975,7.3058467,4.4307694,4.2469745,6.744616,8.825437,8.789334,6.3310776,6.1472826,4.9493337,4.7589746,5.8125134,6.567385,6.117744,5.353026,5.2480006,5.8092313,6.0685134,7.4699492,6.8365135,5.356308,4.07959,3.8990772,2.2383592,1.401436,1.3981539,2.1103592,3.308308,5.028103,4.6276927,3.639795,2.7208207,1.6278975,1.6377437,4.781949,7.499488,8.234667,7.4174366,10.233437,11.073642,8.772923,5.2315903,5.425231,7.643898,11.657847,14.700309,15.579899,14.677335,15.684924,9.7673855,4.414359,2.5600002,2.5961027,4.821334,9.67877,11.608616,9.639385,7.4043083,6.2523084,4.384821,3.442872,3.8728209,4.9362054,4.8738465,3.8367183,2.5304618,1.6278975,1.7493335,1.9429746,2.2383592,3.882667,6.311385,7.1614366,3.6496413,2.1989746,2.9440002,4.381539,3.3476925,2.7536411,5.3136415,10.8767185,14.592001,6.885744,5.2709746,6.997334,7.8670774,6.564103,4.647385,4.706462,4.460308,5.7403083,8.15918,9.117539,6.432821,4.4077954,4.059898,5.2611284,6.7183595,7.5191803,8.618668,8.730257,8.690872,11.447796,13.718975,9.987283,7.817847,9.7214365,13.157744,10.8996935,9.170052,7.250052,5.3366156,4.522667,2.3072822,4.709744,5.333334,3.7349746,5.431795,8.641642,7.512616,4.706462,2.4516926,2.537026,4.4832826,5.546667,7.9983597,12.49477,18.064411,27.477335,38.508312,41.288208,35.748104,31.606155,32.82708,31.471592,27.64472,22.68554,19.177027,14.178463,11.372309,11.044104,11.733335,10.236719,12.199386,11.365745,9.865847,8.933744,8.881231,8.267488,7.3616414,6.554257,5.7632823,4.4045134,2.6683078,2.349949,2.0742567,1.4966155,1.3095386,1.2176411,0.83035904,0.3708718,0.049230773,0.06564103,0.026256412,0.009846155,0.0032820515,0.0,0.0,0.016410258,0.016410258,0.009846155,0.0032820515,0.02297436,0.04594872,0.032820515,0.04594872,0.08861539,0.098461546,0.128,0.08861539,0.06564103,0.098461546,0.15753847,0.40369233,0.58092314,0.69907695,0.6826667,0.37415388,0.098461546,0.052512825,0.11158975,0.24615386,0.51856416,0.52512825,0.5677949,0.6268718,0.6071795,0.35446155,0.15425642,0.37743592,0.73517954,1.0469744,1.2274873,0.9517949,1.1093334,1.4080001,1.5163078,1.079795,0.6301539,0.65641034,0.9517949,1.1191796,0.55794877,0.26912823,0.11158975,0.06564103,0.09189744,0.15097436,0.07876924,0.032820515,0.049230773,0.09189744,0.06564103,0.049230773,0.055794876,0.03938462,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.02297436,0.0,0.0,0.009846155,0.026256412,0.04266667,0.04594872,0.08533334,0.17066668,0.23958977,0.24943592,0.18707694,0.118153855,0.15425642,0.20676924,0.21333335,0.14769232,0.029538464,0.0,0.0,0.009846155,0.055794876,0.055794876,0.07876924,0.13784617,0.24615386,0.42338464,0.45292312,0.42338464,0.34133336,0.24615386,0.2231795,0.27241027,0.49887183,0.6301539,0.57764107,0.4201026,0.35774362,0.27897438,0.17066668,0.059076928,0.009846155,0.009846155,0.13456412,0.43323082,0.61374366,0.072205134,0.013128206,0.0032820515,0.0032820515,0.0,0.0,0.013128206,0.006564103,0.0,0.0032820515,0.009846155,0.0032820515,0.0,0.0,0.0,0.006564103,0.0,0.0,0.0,0.0,0.006564103,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.42338464,0.90584624,1.0010257,0.6662565,0.25928208,0.072205134,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.029538464,0.07548718,0.12143591,0.190359,0.3249231,0.5907693,0.8992821,1.0896411,1.1191796,1.0666667,1.0272821,1.083077,1.211077,1.3522053,1.401436,1.1093334,0.8336411,0.5677949,0.36430773,0.34789747,0.38400003,0.39712822,0.4135385,0.5316923,0.892718,1.0666667,1.2012309,1.1782565,1.0896411,1.211077,1.1782565,1.6344616,3.259077,6.0192823,9.160206,5.7501545,3.6758976,2.678154,2.3204105,2.0020514,2.1530259,2.7044106,2.793026,2.3171284,1.9265642,2.0217438,2.0808206,2.3138463,2.5632823,2.2777438,2.044718,1.6213335,1.2635899,1.0272821,0.79425645,0.65312827,0.5316923,0.46276927,0.44307697,0.45292312,0.56451285,0.827077,1.0305642,0.99774367,0.5973334,0.4594872,0.3708718,0.28882053,0.20020515,0.128,0.13128206,0.14112821,0.12143591,0.08533334,0.10502565,0.13456412,0.16410258,0.18051283,0.190359,0.2231795,0.21989745,0.18051283,0.15097436,0.15097436,0.190359,0.31507695,0.37415388,0.35774362,0.318359,0.36102566,0.3314872,0.29538465,0.25928208,0.2297436,0.22646156,0.23630771,0.28882053,0.4201026,0.6170257,0.8205129,0.9124103,1.2012309,1.2242053,0.9517949,0.77128214,0.6170257,0.47589746,0.380718,0.34789747,0.36102566,0.42994875,0.508718,0.51856416,0.47589746,0.5316923,0.47917953,0.41682056,0.33805132,0.26584616,0.24615386,0.19692309,0.17723078,0.17723078,0.17394873,0.15097436,0.16738462,0.20348719,0.24615386,0.26912823,0.23630771,1.6902566,1.1355898,0.5415385,1.2274873,2.674872,2.5173335,0.5021539,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.006564103,0.01969231,0.0951795,0.20348719,0.21661541,0.13456412,0.036102567,0.055794876,0.10502565,0.049230773,0.009846155,0.029538464,0.055794876,0.029538464,0.07548718,0.10502565,0.1148718,0.190359,0.4955898,0.92553854,1.6114873,2.6420515,4.0402055,6.2720003,9.028924,10.752001,10.932513,10.102155,10.115283,10.036513,10.394258,11.487181,13.403898,15.609437,18.980104,23.56513,29.010054,34.566566,39.401028,42.305645,43.165543,42.033234,39.161438,34.888206,32.338055,31.0679,30.690464,30.86113,27.316515,22.275284,17.913437,15.100719,13.37436,14.647796,14.628103,13.239796,11.772718,12.852514,16.305231,15.186052,11.178667,6.8299494,5.540103,5.333334,5.041231,6.2720003,8.530052,9.206155,6.678975,5.8125134,6.810257,9.8363085,15.00554,14.122667,9.931488,8.257642,10.322052,12.73436,11.001437,9.124104,7.857231,7.0892315,5.87159,4.394667,3.2820516,2.2711797,1.3751796,0.892718,0.42994875,0.82379496,1.6147693,2.3926156,2.809436,2.550154,3.0654361,2.9243078,1.847795,0.71548724,0.85005134,0.74830776,0.6301539,0.5415385,0.35446155,0.2986667,0.33476925,0.37415388,0.4397949,0.6695385,1.0601027,1.2406155,1.4080001,1.6246156,1.8149745,1.6508719,1.719795,2.2153847,2.9538465,3.370667,3.4231799,2.8816411,2.2350771,1.6640002,1.0404103,1.3095386,0.9485129,0.61374366,0.6268718,1.0010257,1.2242053,1.1454359,1.148718,1.3718976,1.7263591,1.8445129,2.0250258,2.3204105,2.3958976,1.5491283,1.339077,1.7001027,1.7362052,1.214359,0.56123084,0.8041026,1.1257436,1.5589745,2.0644104,2.5238976,3.5282054,4.6276927,4.9985647,5.07077,6.5083084,5.208616,3.8990772,3.7743592,4.4832826,4.1222568,3.4789746,4.076308,6.1505647,8.884514,10.407386,7.3616414,5.5138464,5.1922054,5.681231,5.218462,4.519385,3.006359,1.8182565,1.7887181,3.4198978,3.9680004,4.663795,6.669129,8.648206,6.7938466,4.965744,5.0018463,6.2096415,7.3583593,6.705231,7.3747697,4.824616,3.5446157,4.7917953,6.5870776,6.12759,5.3136415,4.6966157,4.6080003,5.1626673,6.747898,6.180103,5.028103,4.31918,4.5456414,3.255795,2.1497438,1.6016412,1.6640002,2.0873847,4.417641,4.5062566,3.6036925,2.556718,1.7788719,1.8904617,3.0096412,4.588308,5.546667,4.2896414,6.1505647,7.3058467,6.987488,6.0652313,7.062975,9.419488,10.962052,11.277129,10.768411,10.637129,10.9226675,6.3540516,2.733949,2.028308,2.3827693,5.477744,9.051898,9.7903595,7.8506675,6.885744,6.498462,5.0904617,3.308308,1.9987694,2.2121027,2.7273848,1.9495386,1.3029745,1.2668719,1.3587693,2.0775387,3.058872,4.338872,5.668103,6.521436,4.9854364,3.7021542,3.2229745,3.245949,2.6026669,2.2186668,4.066462,7.3353853,9.235693,4.9854364,5.3169236,6.2916927,6.3934364,5.4908724,4.818052,4.893539,5.2578464,7.755488,10.020103,5.481026,6.6560006,6.5411286,4.95918,3.4658465,5.349744,6.038975,6.5444107,7.1548724,9.304616,15.596309,19.72513,14.381949,10.44677,11.008,11.34277,7.39118,5.8256416,4.6834874,3.629949,3.948308,2.802872,5.8190775,6.1997952,3.4888208,3.564308,7.322257,8.461129,8.146052,6.8627696,4.414359,4.890257,4.6900516,6.8594875,11.526565,15.90154,19.984411,25.90195,28.320822,26.804514,25.813335,23.217232,21.320208,19.968002,18.30072,14.759386,12.3076935,12.186257,12.35036,11.769437,10.417232,13.843694,13.147899,10.952206,9.242257,9.373539,9.544206,8.710565,7.273026,5.61559,4.1058464,2.6486156,2.0053334,1.529436,1.148718,1.3751796,1.4178462,0.8402052,0.29210258,0.06235898,0.08205129,0.02297436,0.006564103,0.0032820515,0.0,0.0,0.006564103,0.009846155,0.006564103,0.0032820515,0.02297436,0.07548718,0.072205134,0.072205134,0.0951795,0.1148718,0.16082053,0.1148718,0.0951795,0.12471796,0.1148718,0.3446154,0.74830776,1.2898463,1.5031796,0.49887183,0.15753847,0.055794876,0.15097436,0.40369233,0.7811283,0.6629744,0.7220513,0.8533334,0.8730257,0.49887183,0.33476925,0.45292312,0.61374366,0.67610264,0.5973334,0.4594872,0.69579494,0.98461545,1.0896411,0.8730257,0.36102566,0.3117949,0.508718,0.6432821,0.33805132,0.9485129,0.47589746,0.036102567,0.013128206,0.068923086,0.013128206,0.0,0.026256412,0.059076928,0.04594872,0.04594872,0.055794876,0.03938462,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.02297436,0.013128206,0.0032820515,0.006564103,0.02297436,0.06235898,0.13784617,0.18051283,0.27241027,0.36102566,0.40369233,0.36430773,0.256,0.18379489,0.21989745,0.318359,0.34133336,0.14112821,0.059076928,0.032820515,0.036102567,0.055794876,0.10502565,0.12143591,0.14441027,0.21989745,0.39384618,0.45620516,0.46933338,0.35774362,0.17723078,0.11158975,0.20676924,0.5415385,0.7220513,0.6498462,0.54482055,0.4266667,0.28225642,0.19692309,0.15425642,0.02297436,0.19364104,0.47917953,1.079795,1.4802053,0.4397949,0.18707694,0.07548718,0.052512825,0.059076928,0.02297436,0.032820515,0.032820515,0.04266667,0.06564103,0.08861539,0.1148718,0.11158975,0.08533334,0.04266667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.9288206,1.9167181,1.9889232,1.1651284,0.4594872,0.09189744,0.02297436,0.02297436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.01969231,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.009846155,0.02297436,0.059076928,0.12143591,0.20676924,0.38728207,0.6301539,0.90584624,1.142154,1.2373334,1.1126155,1.142154,1.1651284,1.1716924,1.2832822,1.0994873,0.9124103,0.6662565,0.4135385,0.3249231,0.36430773,0.3708718,0.3708718,0.4397949,0.702359,0.8533334,1.1158975,1.2176411,1.1782565,1.3095386,1.3817437,2.1464617,3.9581542,6.6100516,9.334154,5.4383593,3.1803079,2.1497438,1.8773335,1.847795,1.7558975,2.3991797,2.7995899,2.5961027,2.0611284,1.9298463,1.7985642,1.975795,2.3302567,2.284308,2.0118976,1.7263591,1.4408206,1.1815386,1.0010257,0.8598975,0.65312827,0.5021539,0.4397949,0.39712822,0.39056414,0.5415385,0.7811283,0.9517949,0.7811283,0.508718,0.40697438,0.33805132,0.256,0.190359,0.14441027,0.14441027,0.14112821,0.12471796,0.13456412,0.17066668,0.21333335,0.23630771,0.24287182,0.28882053,0.28882053,0.24943592,0.21661541,0.20348719,0.20020515,0.24943592,0.27569234,0.28225642,0.28882053,0.33476925,0.3314872,0.29210258,0.26584616,0.25928208,0.21989745,0.190359,0.2297436,0.33805132,0.508718,0.7187693,0.69907695,0.99774367,1.1716924,1.0633847,0.81394875,0.7450257,0.6301539,0.4955898,0.39056414,0.37743592,0.39712822,0.43651286,0.45292312,0.44964105,0.48902568,0.46276927,0.4135385,0.35446155,0.2986667,0.26584616,0.23958977,0.2100513,0.18379489,0.17066668,0.16082053,0.17066668,0.16082053,0.16410258,0.17723078,0.16082053,0.7056411,0.4955898,0.30194873,1.3784616,3.062154,2.7995899,0.56123084,0.0,0.0,0.0,0.0,0.009846155,0.013128206,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.013128206,0.009846155,0.016410258,0.08533334,0.190359,0.28225642,0.26256412,0.15753847,0.108307704,0.032820515,0.0032820515,0.02297436,0.052512825,0.02297436,0.072205134,0.12471796,0.1148718,0.068923086,0.098461546,0.21661541,0.34133336,0.512,0.73517954,0.9714873,1.9659488,3.121231,4.6802053,6.3442054,7.2664623,7.529026,7.8473854,8.871386,10.824206,13.528616,16.38072,20.834463,25.947899,31.655388,38.79385,43.91385,43.634876,41.232414,38.094772,33.70995,31.671797,32.07549,32.659695,32.482464,31.921234,26.164515,21.35631,18.556719,17.680412,17.509745,19.216412,18.169437,15.520822,13.170873,13.7386675,14.296617,12.619488,9.757539,6.8365135,5.080616,6.3179493,6.052103,4.965744,3.757949,3.1343591,3.8465643,3.6430771,3.0654361,3.1671798,5.5138464,11.460924,9.915077,8.487385,9.705027,11.0145645,9.997129,9.537642,8.815591,7.2960005,4.71959,3.692308,2.865231,1.9167181,0.9419488,0.47589746,0.30851284,0.6465641,1.5655385,2.3794873,1.6278975,1.0699488,1.0994873,1.273436,1.2012309,0.56451285,0.6465641,0.6301539,0.45620516,0.26256412,0.4135385,0.4397949,0.37415388,0.380718,0.51856416,0.7450257,0.67282057,0.8402052,1.0633847,1.2209232,1.2406155,1.7920002,2.553436,3.0129232,2.8750772,2.0676925,1.0305642,0.86646163,0.9288206,0.9189744,0.90256417,1.9003079,1.5589745,0.92553854,0.69251287,1.214359,1.1520001,1.0404103,1.0732309,1.2209232,1.2406155,1.467077,1.7690258,1.9561027,1.9922053,2.0053334,1.8182565,2.281026,2.3663592,1.8642052,1.394872,1.214359,0.99774367,0.9747693,1.1191796,1.1290257,1.529436,1.9692309,2.7503593,4.0336413,5.8518977,5.9536414,4.778667,3.9581542,4.1156926,4.8705645,4.056616,3.69559,5.1954875,8.090257,10.056206,7.683283,5.7665644,5.5105643,6.3474874,5.940513,6.3442054,5.408821,3.7120004,2.3794873,3.0720003,4.2272825,4.2601027,5.034667,6.816821,8.2904625,6.5837955,4.6178465,3.882667,4.8771286,7.1023593,9.209436,6.5280004,4.20759,4.204308,5.290667,5.3366156,4.7491283,4.240411,4.0533338,3.9548721,5.218462,5.156103,4.713026,4.5456414,4.9952826,4.7261543,3.5380516,2.5271797,2.0939488,1.9331284,4.010667,4.073026,3.4297438,2.7798977,2.2055387,1.8904617,1.719795,2.2580514,2.930872,2.038154,2.605949,4.6080003,6.2096415,7.0531287,8.27077,9.019077,7.204103,4.8016415,3.2032824,3.2131286,3.249231,3.0096412,2.7175386,2.6617439,3.2065644,5.1167183,8.625232,8.484103,4.9854364,3.9712822,3.5840003,3.6430771,2.7044106,1.0994873,0.90256417,0.65641034,0.5349744,0.6104616,0.8467693,1.1158975,1.7920002,3.0194874,4.1025643,4.850872,5.546667,5.7764106,5.2480006,4.634257,4.2929235,4.2469745,3.4724104,3.6168208,4.2469745,5.037949,5.76,5.5269747,5.0609236,5.353026,6.308103,6.7577443,5.8978467,6.3343596,10.371283,13.748514,5.661539,8.786052,9.324308,6.8266673,3.5741541,4.59159,5.330052,5.6418467,6.38359,8.795898,14.513232,21.028105,15.455181,10.161232,9.140513,8.004924,3.882667,3.7120004,4.9526157,5.72718,4.8114877,3.7743592,6.3868723,7.017026,4.6145644,2.6978464,7.387898,10.630565,12.035283,10.742155,5.4416413,4.345436,3.4855387,6.5837955,12.544001,15.461744,16.006565,17.792002,21.75672,25.531078,23.463387,15.044924,14.332719,15.254975,14.283488,10.44677,11.565949,15.274668,14.943181,10.860309,10.210463,14.230975,14.611693,12.76718,10.499283,9.984001,10.194052,10.226872,9.189744,6.957949,4.1682053,2.789744,1.8904617,1.585231,1.7427694,1.9790771,1.785436,0.86646163,0.20348719,0.068923086,0.03938462,0.009846155,0.02297436,0.026256412,0.016410258,0.0032820515,0.0032820515,0.009846155,0.02297436,0.04266667,0.06235898,0.14441027,0.14441027,0.10502565,0.072205134,0.08533334,0.09189744,0.06564103,0.06235898,0.072205134,0.013128206,0.016410258,0.58420515,1.5885129,2.1070771,0.41025645,0.21333335,0.098461546,0.24943592,0.636718,0.98461545,0.67938465,0.82379496,0.9911796,0.9288206,0.5415385,0.49230772,0.60389745,0.77128214,0.86646163,0.73517954,0.48246157,0.5316923,0.53825647,0.4135385,0.318359,0.18051283,0.20348719,0.32820517,0.44307697,0.37415388,1.8412309,0.98133343,0.10502565,0.026256412,0.06564103,0.026256412,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01969231,0.04594872,0.032820515,0.013128206,0.0032820515,0.02297436,0.10502565,0.29538465,0.35446155,0.35774362,0.35774362,0.37415388,0.4004103,0.36430773,0.27897438,0.2297436,0.28225642,0.4660513,0.32164106,0.21661541,0.16082053,0.12471796,0.059076928,0.12471796,0.16082053,0.18379489,0.22646156,0.32820517,0.35774362,0.43651286,0.39384618,0.23958977,0.16410258,0.32820517,0.7417436,0.93866676,0.81394875,0.60061544,0.44964105,0.26584616,0.2297436,0.27241027,0.049230773,0.42338464,0.80738467,1.4769232,1.9298463,0.88615394,0.6268718,0.49230772,0.45292312,0.4201026,0.25271797,0.2297436,0.20676924,0.21989745,0.26256412,0.27569234,0.33476925,0.3052308,0.21333335,0.098461546,0.0,0.0,0.0,0.0,0.006564103,0.029538464,0.04594872,0.01969231,0.0,0.0,0.0,0.0,0.0,0.0,0.032820515,0.16082053,1.2603078,2.3236926,2.2646155,1.2340513,0.6104616,0.19692309,0.1148718,0.0951795,0.03938462,0.026256412,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.026256412,0.055794876,0.016410258,0.013128206,0.006564103,0.0032820515,0.0032820515,0.013128206,0.0032820515,0.0032820515,0.0032820515,0.0,0.0,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.009846155,0.026256412,0.049230773,0.0951795,0.20348719,0.40697438,0.69251287,1.0075898,1.276718,1.142154,1.2176411,1.2307693,1.1684103,1.270154,1.079795,0.90912825,0.7089231,0.48246157,0.28882053,0.26584616,0.31507695,0.4135385,0.5284103,0.6170257,0.702359,0.95835906,1.1290257,1.1782565,1.2832822,1.7165129,2.2613335,2.8553848,3.3247182,3.3903592,2.6978464,1.6147693,1.0666667,1.2077949,1.4276924,1.2832822,1.6213335,2.0053334,2.156308,1.9561027,1.8313848,1.7493335,1.8412309,2.03159,2.0545642,1.8576412,1.7920002,1.5721027,1.2274873,1.0929232,1.017436,0.8041026,0.61374366,0.4955898,0.40697438,0.38728207,0.41025645,0.47917953,0.6104616,0.8369231,0.5907693,0.46276927,0.3708718,0.28225642,0.2231795,0.14112821,0.13128206,0.14769232,0.17066668,0.19692309,0.24287182,0.3052308,0.3249231,0.3117949,0.34133336,0.3117949,0.2986667,0.28225642,0.256,0.23630771,0.24615386,0.25271797,0.25271797,0.24615386,0.23630771,0.2231795,0.21661541,0.24287182,0.27569234,0.22646156,0.19692309,0.2297436,0.29210258,0.39384618,0.58420515,0.6268718,0.79097444,0.9419488,0.9714873,0.7975385,0.8402052,0.77128214,0.6104616,0.44307697,0.40697438,0.40697438,0.42994875,0.42338464,0.38400003,0.3249231,0.33476925,0.33476925,0.33476925,0.32164106,0.26584616,0.24943592,0.21333335,0.17394873,0.15097436,0.15753847,0.15753847,0.12143591,0.101743594,0.101743594,0.101743594,0.7187693,0.44964105,0.3446154,0.61374366,1.0043077,0.80738467,0.16082053,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.049230773,0.068923086,0.04594872,0.02297436,0.12143591,0.49887183,0.7056411,0.67938465,0.46276927,0.18379489,0.08533334,0.02297436,0.02297436,0.072205134,0.12143591,0.15753847,0.19692309,0.128,0.013128206,0.06235898,0.21989745,0.2855385,0.38400003,0.58092314,0.88615394,1.276718,1.7591796,2.937436,4.4340515,4.896821,5.58277,6.3212314,8.155898,11.293539,15.090873,17.77559,22.147284,28.950977,37.671387,46.50667,47.205746,41.33744,36.214157,33.257027,27.986053,29.462976,30.116104,28.960823,26.63713,25.38995,27.66113,34.829132,40.772926,41.58031,35.55118,30.267078,22.593643,17.539284,15.911386,14.313026,14.020925,10.843898,7.755488,6.2162056,6.180103,7.53559,6.9677954,5.4153852,3.7185643,2.609231,5.293949,6.1505647,5.1167183,3.4264617,3.5872824,4.562052,9.081436,8.726975,4.1550775,5.080616,6.045539,6.5050263,6.1538467,4.916513,2.9768207,1.975795,1.1552821,0.7056411,0.52512825,0.24287182,0.14769232,0.47917953,2.2678976,4.276513,3.006359,1.2964103,1.2832822,1.4342566,1.0896411,0.44307697,0.5152821,0.49887183,0.39384618,0.43651286,1.083077,1.1323078,0.81394875,0.69907695,0.9517949,1.3423591,0.892718,0.92553854,1.1618463,1.2898463,0.9616411,1.8510771,2.605949,2.5337439,1.8018463,1.4342566,1.2274873,1.3226668,1.3587693,1.2077949,0.97805136,1.9659488,1.8182565,1.2012309,0.81066674,1.3718976,1.5425643,1.7329233,1.7952822,1.6311796,1.1913847,1.6049232,1.9003079,2.048,2.103795,2.2121027,2.2121027,2.231795,2.4024618,2.8225644,3.5544617,2.0644104,0.90584624,0.55794877,0.8598975,1.0075898,0.8598975,0.8795898,1.1651284,1.8510771,3.0818465,4.6572313,4.9493337,4.1682053,3.882667,7.020308,6.6034875,5.720616,5.940513,7.076103,7.1876926,4.7458467,3.9975388,4.4734364,5.5138464,6.2720003,5.4547696,5.9995904,5.579488,4.1091285,3.767795,4.2207184,4.3716927,4.644103,5.973334,9.780514,8.766359,6.298257,4.1878977,3.43959,4.2568207,9.580308,9.107693,7.506052,6.803693,6.377026,6.6461544,6.0356927,4.8640003,3.6496413,3.1113849,3.9187696,4.1550775,3.8071797,3.8498464,6.23918,7.6209235,6.4000006,4.916513,3.8728209,2.3335385,3.7021542,4.3552823,4.5062566,4.0369234,2.487795,1.3883078,1.1684103,1.6377437,2.100513,1.3423591,2.4155898,6.0258465,8.51036,8.109949,4.97559,3.436308,2.858667,3.1113849,3.7251284,3.9220517,3.6529233,4.4012313,4.716308,4.269949,3.8301542,3.170462,6.193231,6.8266673,3.9811285,1.5425643,1.4178462,2.1956925,1.8576412,0.52512825,0.4266667,0.56123084,0.7056411,0.8336411,0.98133343,1.2504616,1.1651284,2.2514873,2.917744,2.8947694,3.249231,6.6560006,6.1440005,5.7468724,6.8004107,7.9327188,6.3606157,6.0291286,5.8157954,5.4416413,5.477744,4.023795,3.5347695,4.571898,6.4623594,7.2927184,6.806975,6.9120007,10.610872,13.925745,5.904411,7.857231,8.933744,7.204103,4.056616,4.164923,3.6036925,2.678154,2.737231,4.066462,5.858462,5.7140517,5.3760004,4.7655387,3.8531284,2.6715899,2.1825643,4.9985647,7.269744,6.9120007,3.6168208,3.31159,7.8473854,9.711591,6.8233852,2.5632823,8.434873,11.067078,9.508103,5.100308,1.4506668,1.4867693,3.0785644,8.188719,14.204719,13.961847,11.008,12.852514,18.648617,24.477541,23.332104,15.126975,13.883078,12.455385,8.822155,6.088206,11.142565,18.602669,19.59713,14.65436,13.702565,15.740719,14.841437,12.967385,11.218052,9.826463,9.852718,11.0375395,10.512411,7.64718,4.059898,3.314872,2.5238976,2.7569232,3.5314875,2.8225644,1.3587693,0.48902568,0.12143591,0.06564103,0.016410258,0.016410258,0.068923086,0.101743594,0.07548718,0.016410258,0.016410258,0.052512825,0.118153855,0.18379489,0.18379489,0.20676924,0.21333335,0.19692309,0.17066668,0.18379489,0.108307704,0.06564103,0.032820515,0.013128206,0.0,0.02297436,0.15097436,0.55794877,0.9714873,0.64000005,0.34789747,0.2297436,0.4135385,0.7778462,0.9616411,0.8992821,1.4342566,1.6902566,1.3817437,0.80738467,0.4660513,0.45620516,0.92553854,1.5885129,1.723077,1.1979488,0.9944616,0.7811283,0.46276927,0.18379489,0.23302566,0.380718,0.44964105,0.4135385,0.4135385,0.764718,0.4594872,0.15425642,0.08861539,0.07548718,0.07548718,0.029538464,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.04594872,0.032820515,0.013128206,0.01969231,0.11158975,0.380718,0.5284103,0.47261542,0.32164106,0.16738462,0.108307704,0.27897438,0.256,0.256,0.3314872,0.380718,0.47917953,0.5021539,0.4594872,0.37415388,0.28882053,0.13128206,0.08205129,0.108307704,0.23302566,0.5481026,0.35446155,0.25928208,0.23958977,0.23958977,0.15097436,0.33476925,1.2504616,1.9528207,1.9200002,1.0535386,0.5874872,0.28882053,0.118153855,0.06235898,0.12143591,0.29210258,0.60061544,0.892718,1.0075898,0.761436,1.4211283,1.723077,1.7427694,1.5097437,1.020718,0.9616411,0.7811283,0.67610264,0.6662565,0.58092314,0.54482055,0.4135385,0.23302566,0.06235898,0.0,0.0,0.0,0.0,0.029538464,0.15097436,0.22646156,0.098461546,0.0,0.0,0.0,0.0,0.0,0.0,0.16082053,0.80738467,1.273436,1.1224617,0.80738467,0.6235898,0.7318975,0.52512825,0.35446155,0.24943592,0.19692309,0.13784617,0.026256412,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.029538464,0.07548718,0.07548718,0.06564103,0.032820515,0.016410258,0.02297436,0.06235898,0.013128206,0.009846155,0.009846155,0.0,0.0,0.013128206,0.006564103,0.0,0.0,0.0,0.0,0.009846155,0.016410258,0.02297436,0.04594872,0.108307704,0.23302566,0.40369233,0.65312827,1.0666667,1.1913847,1.1651284,1.1290257,1.1224617,1.0994873,0.97805136,0.955077,0.80738467,0.508718,0.2297436,0.20348719,0.25271797,0.45620516,0.6892308,0.64000005,0.58092314,0.8566154,1.1027694,1.1224617,0.9156924,1.4769232,1.5983591,1.2438976,0.72861546,0.7187693,4.1846156,2.3040001,0.6859488,0.9878975,0.9156924,0.97805136,1.2471796,1.332513,1.273436,1.5425643,1.7001027,1.5556924,1.591795,1.847795,1.9068719,1.8084104,1.9495386,1.9265642,1.6049232,1.1290257,1.142154,1.1257436,0.9747693,0.69907695,0.44307697,0.40697438,0.34133336,0.318359,0.38400003,0.58092314,0.6662565,0.5021539,0.31507695,0.19692309,0.13784617,0.11158975,0.12471796,0.14441027,0.15753847,0.18379489,0.26912823,0.36430773,0.44307697,0.49887183,0.5481026,0.49887183,0.4594872,0.37415388,0.27241027,0.25928208,0.27241027,0.256,0.23302566,0.2100513,0.19692309,0.18707694,0.16410258,0.17723078,0.21333335,0.21333335,0.21333335,0.23302566,0.24943592,0.28882053,0.4135385,0.5349744,0.60061544,0.7220513,0.8336411,0.6859488,0.6629744,0.72861546,0.7122052,0.57764107,0.44307697,0.40697438,0.42338464,0.4004103,0.31507695,0.2297436,0.31507695,0.3708718,0.3708718,0.31507695,0.2297436,0.23958977,0.23630771,0.21661541,0.19692309,0.18379489,0.17066668,0.15097436,0.118153855,0.08861539,0.07548718,0.7778462,0.7253334,0.40369233,0.20348719,0.20020515,0.16082053,0.072205134,0.01969231,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.013128206,0.009846155,0.02297436,0.108307704,0.3511795,0.5349744,0.5907693,0.50543594,0.34133336,0.30194873,0.118153855,0.0032820515,0.013128206,0.02297436,0.09189744,0.128,0.08533334,0.0032820515,0.013128206,0.36758977,0.50543594,0.60061544,0.77128214,1.0568206,1.3784616,2.1366155,2.865231,3.4330258,4.0434875,5.546667,8.6580515,11.969642,14.647796,16.433231,20.690052,29.732105,41.81662,52.75898,55.94257,47.1959,38.514874,33.217644,31.130259,28.583387,29.229952,28.399591,27.579079,27.792412,29.61395,34.783184,42.06277,53.149544,62.736416,58.512413,40.12308,28.6359,21.474463,16.393847,11.493745,10.614155,8.425026,6.774154,6.265436,6.2785645,6.042257,4.818052,3.8334363,3.2984617,2.4024618,3.4756925,5.6254363,6.294975,5.796103,7.3321033,3.7120004,3.170462,2.7569232,1.8576412,2.1989746,3.114667,3.2853336,2.806154,1.9200002,1.0338463,0.64000005,0.5284103,0.47261542,0.380718,0.3052308,0.3052308,0.39056414,2.9505644,6.265436,4.5062566,1.4605129,1.5195899,2.2482052,2.228513,1.0535386,0.46276927,0.35774362,0.7384616,1.5458462,2.681436,1.4998976,1.2274873,1.0043077,0.62030774,0.512,0.84348726,1.204513,1.3292309,1.1290257,0.69251287,1.3193847,1.8412309,1.8346668,1.394872,1.1158975,1.5524104,1.7526156,1.4834872,0.9288206,0.65969235,1.276718,1.3817437,1.214359,1.086359,1.3850257,1.401436,1.5885129,1.657436,1.7001027,2.1792822,3.1015387,2.5271797,1.8543591,1.7329233,2.0676925,1.9692309,1.6114873,1.4211283,1.7723079,2.9801028,3.3280003,2.1136413,1.4211283,1.8116925,2.349949,1.3161026,0.96492314,1.1684103,1.7920002,2.6912823,4.0041027,5.3792825,5.405539,4.7425647,6.1407185,6.3901544,5.730462,5.874872,6.7971287,6.770872,4.6145644,3.7973337,4.013949,5.0051284,6.550975,5.970052,5.277539,4.9427695,4.900103,4.5489235,3.8695388,4.2994876,5.106872,5.943795,6.8529234,5.1364107,4.1911798,3.6102567,3.255795,3.242667,4.269949,6.6494365,8.763078,10.016821,10.820924,8.726975,5.8420515,4.7622566,5.2348723,4.1517954,5.3366156,5.756718,4.923077,3.9351797,5.4974365,6.9152827,7.5421543,6.426257,4.3716927,3.9581542,3.0785644,3.8531284,4.7950773,4.84759,3.367385,1.7591796,1.5655385,2.0118976,2.281026,1.5130258,3.5347695,5.6451287,6.6461544,5.986462,3.7776413,2.678154,3.1507695,3.7087183,3.3247182,1.4309745,1.2603078,1.5195899,2.0118976,2.231795,1.3522053,0.955077,3.0391798,3.9253337,2.6683078,1.0666667,1.1684103,2.0512822,1.7920002,0.53825647,0.48902568,0.7187693,1.7591796,2.225231,1.7952822,1.214359,1.8707694,2.7273848,2.7273848,1.972513,1.7132308,3.2328207,4.2863593,7.686565,11.733335,10.194052,5.356308,4.2469745,4.194462,4.089436,4.378257,3.698872,4.4242053,5.5171285,6.432821,7.1483083,7.968821,8.27077,11.162257,13.443283,5.5893335,7.0137444,6.6822567,6.183385,6.3376417,7.181129,5.8190775,8.388924,11.88759,13.308719,9.655796,4.2568207,3.3575387,3.6069746,3.387077,2.8160002,3.7054362,6.413129,8.684308,8.349539,3.3345644,4.84759,11.72677,12.501334,6.124308,1.9889232,11.592206,14.670771,11.050668,4.2568207,1.5360001,1.7001027,6.186667,9.494975,8.953437,4.7458467,5.464616,9.242257,13.860104,18.20554,22.291695,15.58318,11.437949,9.206155,8.385642,8.63836,10.187488,16.961643,21.11672,20.361847,17.975796,15.258258,13.653335,13.042872,12.875488,12.156719,13.423591,13.2562065,11.808822,9.278359,5.914257,4.164923,3.6332312,4.0992823,4.4996924,2.934154,1.654154,0.6104616,0.12143591,0.0951795,0.026256412,0.036102567,0.08861539,0.101743594,0.072205134,0.03938462,0.049230773,0.08205129,0.128,0.18051283,0.21989745,0.128,0.08861539,0.10502565,0.14441027,0.14769232,0.11158975,0.068923086,0.032820515,0.013128206,0.0,0.08205129,0.15753847,0.29210258,0.49230772,0.6892308,0.39712822,0.32164106,0.37743592,0.45620516,0.42338464,0.85005134,1.1618463,1.404718,1.4802053,1.1520001,0.88615394,0.49887183,0.4397949,0.7515898,1.0535386,1.083077,1.1290257,0.96492314,0.6235898,0.39056414,0.55794877,0.9485129,1.6443079,1.9790771,0.5349744,0.3708718,0.20676924,0.08205129,0.026256412,0.052512825,0.06235898,0.026256412,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.032820515,0.0951795,0.13128206,0.098461546,0.059076928,0.055794876,0.12143591,0.27241027,0.3314872,0.61374366,0.5973334,0.2855385,0.20348719,0.25928208,0.25271797,0.23302566,0.26584616,0.44307697,0.44307697,0.5218462,0.67610264,0.77128214,0.55794877,0.30194873,0.19364104,0.17394873,0.19692309,0.21989745,0.09189744,0.101743594,0.20348719,0.29538465,0.23958977,0.5481026,1.2176411,1.6443079,1.6016412,1.2242053,0.6235898,0.37743592,0.22646156,0.13784617,0.318359,0.8598975,0.93866676,1.1585642,1.5688206,1.6672822,1.6508719,1.6607181,2.0250258,2.5337439,2.425436,1.595077,1.339077,1.3751796,1.5097437,1.6311796,1.3193847,0.9485129,0.58420515,0.318359,0.26912823,0.15097436,0.12143591,0.118153855,0.12471796,0.190359,0.18379489,0.21333335,0.22646156,0.20348719,0.14769232,0.128,0.1148718,0.108307704,0.15097436,0.30851284,0.44964105,0.38728207,0.52512825,0.94523084,1.4145643,1.276718,0.86646163,0.55794877,0.4594872,0.41682056,0.32820517,0.23958977,0.16082053,0.101743594,0.072205134,0.013128206,0.0,0.0,0.0,0.0,0.0,0.029538464,0.049230773,0.049230773,0.049230773,0.059076928,0.068923086,0.055794876,0.029538464,0.03938462,0.026256412,0.013128206,0.006564103,0.013128206,0.013128206,0.04266667,0.02297436,0.0032820515,0.0032820515,0.013128206,0.0032820515,0.009846155,0.006564103,0.0,0.0,0.0,0.0032820515,0.006564103,0.01969231,0.032820515,0.04594872,0.09189744,0.20348719,0.41025645,0.7253334,1.1224617,1.1651284,1.0699488,1.014154,1.148718,1.1126155,0.98133343,0.8369231,0.6662565,0.37415388,0.25271797,0.22646156,0.3117949,0.4660513,0.60389745,0.56123084,0.764718,0.9124103,0.8992821,0.83035904,1.3029745,1.6836925,1.4309745,0.7089231,0.37415388,1.0305642,0.60061544,0.256,0.4135385,0.7187693,0.5677949,0.86646163,1.1618463,1.3883078,1.8707694,2.2350771,1.972513,1.6311796,1.5458462,1.8707694,1.7920002,2.0118976,2.100513,1.8215386,1.1290257,1.1027694,1.1520001,1.1552821,1.017436,0.6629744,0.4004103,0.3249231,0.30851284,0.318359,0.39712822,0.48246157,0.4660513,0.37415388,0.24615386,0.13784617,0.11158975,0.13128206,0.15425642,0.16738462,0.17066668,0.21661541,0.27241027,0.34789747,0.44307697,0.5481026,0.51856416,0.574359,0.58420515,0.512,0.39384618,0.32820517,0.27897438,0.24287182,0.21333335,0.16082053,0.16082053,0.14769232,0.15097436,0.16082053,0.14112821,0.13128206,0.15425642,0.18707694,0.2297436,0.31507695,0.40697438,0.4594872,0.5218462,0.57764107,0.5284103,0.49230772,0.5218462,0.60061544,0.6465641,0.5021539,0.39712822,0.39384618,0.37743592,0.318359,0.23958977,0.2986667,0.38400003,0.39056414,0.3117949,0.26584616,0.25928208,0.24615386,0.2297436,0.2100513,0.20676924,0.19692309,0.19692309,0.17394873,0.12471796,0.06564103,1.0404103,1.0272821,0.58092314,0.27569234,0.20348719,0.0,0.01969231,0.009846155,0.0,0.0,0.0,0.0,0.0,0.049230773,0.0951795,0.0,0.006564103,0.0032820515,0.0,0.0,0.0,0.029538464,0.049230773,0.032820515,0.009846155,0.04266667,0.20676924,0.34789747,0.39712822,0.3249231,0.15097436,0.14441027,0.055794876,0.006564103,0.03938462,0.118153855,0.052512825,0.06564103,0.06564103,0.029538464,0.0,0.256,0.47917953,0.7318975,1.0436924,1.4276924,2.0644104,3.2196925,4.5423594,5.8190775,6.9710774,9.419488,13.016617,16.52513,20.04677,25.025642,34.743797,46.093132,54.104618,55.975388,51.081852,39.25662,32.43323,29.587694,29.062567,28.596516,28.836105,27.214771,25.813335,25.947899,28.163284,31.875284,35.075283,41.613132,48.879593,47.842464,36.178055,30.391798,24.67118,17.234053,10.322052,8.651488,7.351795,6.485334,5.986462,5.651693,7.4404106,6.189949,5.8223596,6.7249236,5.737026,5.618872,7.8408213,7.8080006,5.7796926,6.8594875,3.8301542,2.1858463,1.5556924,1.4178462,1.086359,1.273436,1.2274873,0.96492314,0.61374366,0.42994875,0.3249231,0.36102566,0.32820517,0.2231795,0.26584616,0.28225642,0.24943592,1.7755898,3.8596926,2.8947694,1.3981539,1.5458462,1.8248206,1.4998976,0.62030774,0.39712822,0.5940513,0.94523084,1.3062565,1.6278975,1.024,1.214359,1.0666667,0.47589746,0.36102566,1.0666667,1.6278975,1.7887181,1.6344616,1.595077,0.955077,1.3522053,1.529436,1.2012309,1.0568206,1.2438976,1.1158975,0.7975385,0.5940513,1.0108719,1.3226668,0.9878975,0.65641034,0.6859488,1.1224617,1.2307693,1.6705642,2.0906668,2.3040001,2.281026,3.6594875,2.540308,1.5458462,1.7460514,2.6420515,2.0808206,1.6180514,1.4867693,2.3433847,5.2545643,2.7634873,1.9626669,1.9593848,2.097231,1.9364104,1.3653334,1.1290257,1.4375386,2.284308,3.446154,4.8082056,6.2884107,6.918565,6.8660517,7.4207187,8.487385,8.989539,8.598975,7.7981544,7.8670774,8.687591,7.1581545,5.3070774,4.4438977,5.156103,5.4449234,4.637539,4.194462,4.46359,4.673641,5.179077,6.921847,8.116513,7.7948723,5.7796926,6.0717955,5.7829747,4.4996924,3.121231,3.8596926,4.7917953,5.668103,6.948103,8.828718,11.227899,8.723693,5.8420515,4.9460516,5.668103,4.9329233,4.9526157,5.2414365,4.6211286,3.442872,3.5905645,6.2194877,8.162462,7.0400004,3.948308,3.4756925,3.2065644,3.5840003,4.709744,5.8190775,5.2611284,3.3378465,3.058872,3.0129232,2.5993848,2.0512822,3.826872,5.139693,5.5236926,4.7622566,2.8914874,2.3433847,2.7011285,2.678154,1.910154,0.96492314,0.71548724,0.6235898,0.79425645,1.0010257,0.67610264,0.3052308,1.4998976,2.2711797,1.8937438,0.9288206,0.7056411,1.7887181,1.8871796,0.8205129,0.512,0.57764107,1.8773335,2.8521028,2.8488207,2.1202054,2.0250258,2.0053334,1.7066668,1.2340513,1.1618463,1.6180514,3.3936412,7.3747697,10.791386,7.197539,4.5456414,5.5926156,5.579488,3.889231,4.023795,5.1232824,7.397744,8.772923,8.339693,6.3507695,8.605539,8.881231,9.718155,9.783795,3.8596926,4.1878977,4.516103,6.2194877,8.815591,9.96759,6.514872,9.465437,15.415796,19.085129,13.305437,5.287385,4.601436,6.554257,7.9294367,6.9645133,6.232616,7.653744,8.749949,7.709539,3.383795,9.275078,21.425232,20.168207,6.626462,2.7076926,11.972924,14.043899,9.544206,2.678154,1.1979488,1.1749744,5.586052,8.480822,7.3550773,3.1376412,5.218462,7.3485136,11.339488,17.575386,24.999386,23.446976,15.914668,9.419488,7.3419495,9.432616,9.803488,14.020925,18.41231,20.315899,18.090668,14.381949,15.835898,16.73518,15.360002,13.978257,15.346873,14.785643,12.550565,9.4457445,6.8266673,6.2588725,5.661539,5.0543594,4.2469745,2.8225644,1.4276924,0.512,0.118153855,0.0951795,0.10502565,0.101743594,0.09189744,0.08861539,0.0951795,0.09189744,0.10502565,0.101743594,0.11158975,0.16410258,0.30194873,0.19364104,0.128,0.16738462,0.256,0.2100513,0.13456412,0.16738462,0.19692309,0.16738462,0.08205129,0.06235898,0.10502565,0.13456412,0.18379489,0.380718,0.3314872,0.32164106,0.2855385,0.21333335,0.14441027,0.62030774,0.78769237,0.9517949,1.2176411,1.4834872,1.5031796,1.0043077,0.54482055,0.39056414,0.51856416,0.6662565,0.8795898,0.8369231,0.6301539,0.75487185,0.6859488,1.0666667,1.7920002,2.5140514,2.6322052,1.0666667,0.3052308,0.06235898,0.059076928,0.036102567,0.032820515,0.108307704,0.09189744,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.036102567,0.036102567,0.07548718,0.15425642,0.24287182,0.27241027,0.23630771,0.15097436,0.118153855,0.16082053,0.22646156,0.22646156,0.38400003,0.45620516,0.4266667,0.5316923,0.41025645,0.2986667,0.24287182,0.256,0.30194873,0.32164106,0.3446154,0.38728207,0.4135385,0.31507695,0.15097436,0.14769232,0.20676924,0.27241027,0.34789747,0.4660513,0.56451285,0.5874872,0.48246157,0.2231795,0.40369233,0.574359,0.6629744,0.6465641,0.5513847,0.27569234,0.23958977,0.6071795,1.2504616,1.7296412,1.9922053,1.6508719,1.5261539,1.8182565,2.1103592,2.4352822,2.8980515,3.9056413,5.100308,5.35959,4.1124105,3.2689233,3.1442053,3.5282054,3.6758976,2.8389745,1.7296412,0.96492314,0.764718,0.9485129,1.0075898,0.69907695,0.46933338,0.44307697,0.4266667,0.38728207,0.39056414,0.39056414,0.36758977,0.33805132,0.32164106,0.31507695,0.318359,0.3314872,0.33805132,0.33476925,0.28225642,0.40369233,0.8172308,1.5425643,2.2744617,2.2022567,1.7001027,1.1158975,0.761436,0.58092314,0.4594872,0.36758977,0.27897438,0.19364104,0.08861539,0.06564103,0.055794876,0.036102567,0.0,0.0,0.013128206,0.029538464,0.032820515,0.02297436,0.036102567,0.049230773,0.04266667,0.026256412,0.029538464,0.026256412,0.01969231,0.01969231,0.02297436,0.009846155,0.029538464,0.01969231,0.006564103,0.0,0.006564103,0.009846155,0.006564103,0.006564103,0.006564103,0.0,0.0,0.0,0.0032820515,0.006564103,0.013128206,0.026256412,0.04594872,0.11158975,0.23958977,0.4201026,0.8336411,0.86646163,0.8172308,0.86317956,1.0404103,1.0568206,0.9353847,0.82379496,0.7253334,0.47589746,0.3446154,0.21989745,0.21333335,0.36102566,0.6301539,0.55794877,0.6498462,0.79425645,0.8960001,0.88287187,0.9878975,1.2537436,1.1848207,0.7384616,0.318359,0.23302566,0.15425642,0.13128206,0.2297436,0.54482055,0.32820517,0.47261542,0.8598975,1.4276924,2.162872,2.4320002,2.2482052,2.0151796,1.9692309,2.1924105,1.6935385,1.6049232,1.782154,1.9068719,1.4769232,1.273436,1.2570257,1.2668719,1.1946667,1.0010257,0.7056411,0.4660513,0.33476925,0.30851284,0.3511795,0.43651286,0.39712822,0.2986667,0.19692309,0.14769232,0.12143591,0.128,0.14112821,0.15425642,0.16738462,0.21989745,0.23958977,0.318359,0.4594872,0.60389745,0.6170257,0.67938465,0.72861546,0.6826667,0.46276927,0.37743592,0.32164106,0.26912823,0.21661541,0.16082053,0.14769232,0.12471796,0.11158975,0.118153855,0.12143591,0.101743594,0.108307704,0.13128206,0.16738462,0.22646156,0.26584616,0.32164106,0.4004103,0.46933338,0.4594872,0.42994875,0.4397949,0.48574364,0.5284103,0.49887183,0.44307697,0.41682056,0.37743592,0.318359,0.24287182,0.22646156,0.256,0.26584616,0.24943592,0.256,0.26584616,0.26912823,0.25271797,0.21989745,0.20348719,0.21333335,0.21333335,0.190359,0.13128206,0.052512825,0.92553854,0.92553854,0.5021539,0.23302566,0.20348719,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06564103,0.13456412,0.01969231,0.009846155,0.0032820515,0.0,0.0,0.0,0.029538464,0.068923086,0.055794876,0.009846155,0.049230773,0.118153855,0.18707694,0.20676924,0.15097436,0.0,0.01969231,0.009846155,0.006564103,0.03938462,0.118153855,0.02297436,0.02297436,0.036102567,0.029538464,0.0,0.15425642,0.33476925,0.6235898,1.0568206,1.6049232,2.6847181,4.5554876,6.9710774,9.852718,13.305437,18.566566,23.364925,27.536413,32.42667,40.914055,49.778877,54.13416,52.414364,45.604107,37.20862,28.970669,25.888823,25.819899,27.040823,28.248617,27.887592,25.93149,24.448002,24.359386,25.445745,26.318771,28.01231,31.291079,34.304,32.600616,28.777027,26.95877,22.626463,15.510976,9.577026,7.6242056,6.816821,6.4656415,6.0783596,5.35959,7.765334,8.310155,8.694155,9.206155,8.720411,8.864821,9.563898,7.817847,4.5095387,4.414359,3.1409233,1.9167181,1.2931283,1.1618463,0.7581539,0.508718,0.37743592,0.28882053,0.23630771,0.29538465,0.26584616,0.35774362,0.50543594,0.6301539,0.6695385,0.48574364,0.39712822,0.92225647,1.7329233,1.6278975,2.0184617,2.4549747,2.1464617,1.1881026,0.57764107,0.6826667,0.8402052,0.9353847,0.9124103,0.8041026,0.7811283,1.0108719,0.98461545,0.7515898,0.9156924,1.6278975,1.913436,1.9429746,1.9396925,2.1956925,0.955077,0.9944616,1.2274873,1.1815386,1.0305642,0.83035904,0.6071795,0.57764107,0.83035904,1.3259488,1.1815386,0.60389745,0.33805132,0.6268718,1.1946667,1.142154,1.5786668,1.9626669,1.975795,1.5097437,2.5238976,1.9626669,1.5097437,1.8543591,2.7175386,2.0512822,1.9200002,1.8773335,2.4910772,5.3103595,1.8543591,1.9003079,2.4615386,2.2908719,1.8740515,1.591795,1.4473847,1.8051283,2.6420515,3.5249233,5.277539,6.7117953,7.460103,7.4830775,7.0793853,8.346257,9.750975,9.764103,8.651488,8.470975,10.522257,9.563898,7.0957956,4.772103,4.4077954,5.0510774,4.8344617,4.562052,4.7228723,5.4843082,6.2785645,7.9983597,9.042052,8.802463,7.6668725,10.134975,9.403078,6.7117953,4.201026,4.893539,5.5302567,5.474462,5.733744,6.7183595,8.224821,6.47877,4.7524104,4.4800005,5.5630774,6.377026,4.6867695,4.381539,4.1222568,3.4658465,2.868513,6.3540516,8.090257,6.8266673,3.9745643,3.6102567,3.8498464,3.570872,3.9712822,5.2545643,6.6395903,5.218462,4.138667,3.4527183,3.1507695,3.1442053,3.3903592,4.352,4.788513,4.128821,2.4418464,2.7109745,2.5074873,1.8379488,1.1290257,1.2077949,0.9156924,0.88615394,0.9189744,0.8566154,0.5677949,0.5513847,2.3236926,3.43959,3.006359,1.6836925,1.394872,1.6836925,1.5360001,0.8566154,0.47589746,0.44307697,1.6607181,2.737231,2.9210258,2.097231,2.5074873,2.3991797,2.2121027,2.2121027,2.4976413,2.9604106,5.5893335,7.722667,7.8112826,5.4186673,5.979898,6.698667,5.7140517,3.9187696,4.962462,7.3583593,9.537642,9.6754875,8.592411,9.760821,12.967385,12.868924,10.20718,6.1538467,2.3236926,2.8356924,4.2272825,7.680001,11.989334,13.568001,6.7872825,7.4896417,13.147899,17.604925,11.090053,5.333334,5.3727183,8.254359,10.65354,8.868103,6.7807183,6.514872,7.565129,8.011488,4.5062566,11.687386,25.347284,24.362669,9.764103,4.7524104,9.517949,9.452309,5.730462,1.3029745,0.892718,1.3095386,6.5411286,9.731283,8.192,3.3936412,4.95918,6.180103,10.368001,18.067694,27.073643,29.239798,18.993233,9.498257,6.5936418,8.79918,8.78277,12.701539,17.417847,20.276514,19.104822,15.780104,17.24718,17.88718,16.384,15.717745,16.479181,15.455181,13.078976,10.456616,9.340718,8.231385,6.9809237,5.431795,3.8038976,2.7142565,1.2406155,0.50543594,0.24287182,0.20348719,0.15097436,0.14441027,0.108307704,0.08861539,0.108307704,0.17066668,0.21661541,0.16738462,0.13128206,0.17723078,0.3314872,0.27897438,0.17066668,0.18379489,0.29210258,0.28225642,0.19692309,0.24615386,0.3052308,0.30194873,0.2100513,0.12143591,0.14769232,0.17066668,0.17066668,0.24615386,0.28225642,0.25271797,0.17066668,0.08205129,0.068923086,0.48246157,0.6104616,0.65969235,0.8205129,1.2832822,1.4966155,1.211077,0.79425645,0.46933338,0.3052308,0.55794877,0.7811283,0.8336411,0.80738467,1.0404103,1.211077,1.5261539,1.6804104,1.8215386,2.5600002,1.0502565,0.2855385,0.04266667,0.06564103,0.055794876,0.04266667,0.118153855,0.101743594,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.032820515,0.06564103,0.072205134,0.06235898,0.072205134,0.07876924,0.16410258,0.28225642,0.37743592,0.4135385,0.44307697,0.3511795,0.25928208,0.24287182,0.3117949,0.36102566,0.46933338,0.6301539,0.827077,1.020718,0.6465641,0.3314872,0.18379489,0.17394873,0.13128206,0.15425642,0.3117949,0.3446154,0.20676924,0.06564103,0.013128206,0.08861539,0.19692309,0.29210258,0.36758977,0.5481026,0.65312827,0.61374366,0.4397949,0.2297436,0.4397949,0.46276927,0.56123084,0.7778462,0.955077,1.083077,1.2603078,1.975795,3.0785644,3.7874875,3.6135387,2.6486156,1.8773335,1.7723079,2.2646155,3.308308,4.381539,5.5729237,6.560821,6.6100516,5.5302567,5.3366156,5.533539,5.802667,6.0225644,5.425231,3.4034874,1.7558975,1.2209232,1.4736412,1.5622566,1.2865642,1.1290257,1.1520001,0.9878975,0.90584624,0.8402052,0.76800007,0.7056411,0.6859488,0.6695385,0.6629744,0.6695385,0.6826667,0.67282057,0.6170257,0.5415385,0.5218462,0.7056411,1.3226668,2.8127182,3.3312824,2.9965131,2.176,1.4834872,1.0010257,0.7253334,0.574359,0.47917953,0.38728207,0.256,0.17394873,0.118153855,0.06235898,0.006564103,0.0,0.0032820515,0.009846155,0.013128206,0.006564103,0.013128206,0.02297436,0.029538464,0.032820515,0.036102567,0.032820515,0.029538464,0.029538464,0.029538464,0.02297436,0.016410258,0.016410258,0.013128206,0.009846155,0.006564103,0.009846155,0.0032820515,0.006564103,0.013128206,0.006564103,0.006564103,0.0032820515,0.0,0.0,0.006564103,0.026256412,0.04594872,0.07876924,0.13784617,0.23958977,0.5349744,0.6432821,0.702359,0.79425645,0.9485129,0.9747693,0.9288206,0.827077,0.67610264,0.45292312,0.36430773,0.2297436,0.18051283,0.28225642,0.5415385,0.5513847,0.5973334,0.702359,0.8205129,0.827077,0.7187693,0.892718,0.9321026,0.69251287,0.3052308,0.21333335,0.16410258,0.13456412,0.15753847,0.3052308,0.20676924,0.256,0.5546667,1.1290257,1.9331284,2.2482052,2.425436,2.556718,2.6157951,2.4549747,1.8084104,1.4178462,1.4572309,1.8018463,2.0020514,1.7132308,1.467077,1.332513,1.273436,1.1651284,0.9682052,0.79425645,0.64000005,0.5021539,0.380718,0.4135385,0.3511795,0.24615386,0.16082053,0.15097436,0.13784617,0.13128206,0.13456412,0.14769232,0.16738462,0.21333335,0.2231795,0.2855385,0.42338464,0.5973334,0.6629744,0.75487185,0.8598975,0.8730257,0.60389745,0.47917953,0.39384618,0.3249231,0.25928208,0.18707694,0.14112821,0.11158975,0.098461546,0.10502565,0.10502565,0.098461546,0.0951795,0.098461546,0.118153855,0.15753847,0.19692309,0.256,0.35446155,0.45292312,0.47261542,0.44307697,0.4201026,0.39712822,0.39056414,0.43323082,0.47917953,0.4955898,0.44307697,0.34133336,0.26912823,0.2231795,0.20348719,0.20020515,0.20676924,0.21333335,0.24287182,0.25928208,0.24943592,0.21989745,0.2100513,0.2100513,0.19364104,0.16410258,0.118153855,0.059076928,0.47917953,0.5218462,0.2297436,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.032820515,0.07548718,0.036102567,0.006564103,0.0,0.0,0.0,0.0,0.0,0.04266667,0.04266667,0.01969231,0.098461546,0.09189744,0.101743594,0.1148718,0.098461546,0.016410258,0.052512825,0.02297436,0.0,0.0032820515,0.01969231,0.016410258,0.016410258,0.01969231,0.029538464,0.04594872,0.17066668,0.24615386,0.4397949,0.8533334,1.5261539,3.1409233,5.8420515,9.363693,14.139078,21.303797,30.41149,37.22503,42.36144,47.327183,54.531284,54.705235,47.35344,37.64513,29.049438,23.328823,21.507284,21.546669,23.177849,25.659079,27.782566,26.998156,25.088001,23.972105,23.936003,23.611078,22.465643,25.15036,28.406157,29.236515,24.884514,23.552002,21.07077,16.932104,12.064821,8.818872,7.177847,6.8627696,7.0957956,7.145026,6.3376417,6.6461544,9.609847,10.643693,9.229129,8.904206,9.875693,8.595693,5.805949,2.9210258,2.0184617,1.6410258,0.94523084,0.53825647,0.5349744,0.54482055,0.41025645,0.3117949,0.25271797,0.21989745,0.20020515,0.14441027,0.32820517,0.7811283,1.2603078,1.2537436,0.80738467,0.7581539,1.0305642,1.4375386,1.6836925,2.8750772,3.4527183,2.8816411,1.6082052,1.0765129,1.1323078,0.8795898,0.7581539,0.86317956,0.96492314,0.86646163,0.7220513,0.8566154,1.3161026,1.8707694,2.228513,1.8576412,1.5360001,1.6246156,2.0742567,1.1979488,0.7515898,0.85005134,1.1815386,1.0108719,0.6071795,0.5513847,0.9485129,1.4900514,1.4473847,0.7450257,0.35774362,0.512,1.086359,1.591795,1.1355898,1.2504616,1.2274873,0.8763078,0.52512825,0.67282057,1.1618463,1.595077,1.8674873,2.166154,1.7920002,2.0184617,1.9528207,1.7493335,2.5895386,1.3357949,2.156308,2.6945643,2.3630772,2.356513,1.8609232,1.6968206,1.9462565,2.3762052,2.4418464,4.2371287,5.5926156,6.12759,5.7829747,4.8377438,5.737026,7.4371285,8.549745,8.454565,7.2894363,8.182155,8.874667,7.9425645,5.904411,5.2315903,5.4416413,6.0849237,6.518154,6.747898,7.456821,7.0859494,7.1614366,7.3353853,7.817847,9.383386,12.57354,11.444513,8.54318,6.042257,5.733744,4.893539,5.5729237,5.8814363,5.1987696,4.1780515,3.6824617,3.1934361,3.4855387,4.9788723,7.7357955,5.7107697,4.33559,3.879385,4.017231,3.8465643,7.282872,7.824411,6.6133337,5.1626673,5.35959,4.9460516,4.013949,3.2032824,3.6102567,6.770872,6.442667,4.2994876,3.0326157,3.3509746,3.9844105,2.5764105,3.4297438,4.1878977,3.7776413,2.425436,3.4100516,2.7208207,1.9331284,1.8313848,2.412308,2.2055387,2.2449234,2.4648206,2.3269746,0.8205129,1.4802053,4.824616,6.7971287,5.796103,2.6847181,2.4516926,1.5163078,0.8041026,0.58092314,0.4594872,0.47917953,1.4112822,2.1333334,2.048,1.079795,3.1081028,3.8629746,4.204308,4.535795,4.7655387,6.0324106,8.825437,8.306872,5.1889234,5.733744,7.75877,6.0685134,4.6572313,5.5105643,8.608821,10.331899,9.731283,7.1876926,6.3868723,14.319591,17.732924,16.68595,11.024411,3.9876926,2.2153847,3.9680004,5.805949,9.156924,13.121642,14.460719,6.2720003,5.3694363,10.039796,14.10954,6.931693,4.2568207,4.493129,6.951385,9.225847,7.1680007,5.5663595,4.4242053,6.6395903,9.846154,6.413129,9.905231,19.538054,20.995283,12.888617,6.744616,6.550975,4.194462,1.8904617,0.8008206,1.0436924,3.3444104,9.885539,12.534155,8.992821,2.7766156,3.245949,5.346462,10.102155,17.503181,26.512413,27.588924,17.204514,8.736821,6.9710774,8.067283,7.8047185,12.960821,18.06113,20.614565,21.110155,19.908924,18.051283,17.14872,18.031591,20.768822,18.323694,16.042667,13.978257,12.501334,12.294565,9.314463,7.328821,5.405539,3.4789746,2.356513,1.1881026,0.636718,0.44964105,0.36758977,0.15097436,0.14112821,0.13456412,0.128,0.15097436,0.27897438,0.36758977,0.27569234,0.20348719,0.23302566,0.3249231,0.32164106,0.18051283,0.13456412,0.2297436,0.3249231,0.28882053,0.27241027,0.2855385,0.3117949,0.30194873,0.24943592,0.28882053,0.3708718,0.45292312,0.48902568,0.35774362,0.190359,0.07548718,0.04594872,0.0951795,0.47261542,0.7515898,0.761436,0.6071795,0.67282057,0.86317956,0.9288206,0.8402052,0.61374366,0.3052308,0.74830776,0.8533334,0.9124103,0.99774367,0.9714873,1.6016412,1.8871796,1.5327181,0.81394875,0.56451285,0.37415388,0.39712822,0.37743592,0.3314872,0.54482055,0.35446155,0.24615386,0.24615386,0.28882053,0.23302566,0.09189744,0.02297436,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.032820515,0.026256412,0.032820515,0.02297436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13784617,0.21333335,0.21989745,0.16738462,0.11158975,0.128,0.256,0.39712822,0.50543594,0.62030774,0.8041026,0.76800007,0.5973334,0.4397949,0.53825647,0.79425645,1.1027694,1.2931283,1.3554872,1.4309745,0.80738467,0.31507695,0.068923086,0.036102567,0.026256412,0.14112821,0.7089231,0.9485129,0.6826667,0.34133336,0.21661541,0.37743592,0.5513847,0.60389745,0.53825647,0.63343596,0.58092314,0.6268718,0.764718,0.7450257,1.0633847,1.1946667,1.5458462,2.156308,2.7109745,3.1737437,3.4888208,4.0533338,4.9460516,5.914257,5.5007186,3.95159,2.5173335,1.9856411,2.665026,4.2929235,5.9930263,7.322257,7.8112826,6.9710774,5.5007186,6.439385,7.574975,7.968821,7.955693,7.6143594,5.113436,2.789744,1.7723079,1.9790771,1.9954873,2.048,2.169436,2.2088206,1.8084104,1.6902566,1.6016412,1.4736412,1.332513,1.2931283,1.2635899,1.2340513,1.2209232,1.214359,1.2012309,1.1224617,1.014154,0.90912825,0.9156924,1.2504616,3.117949,4.1846156,4.2207184,3.4330258,2.4943593,1.6705642,1.1388719,0.8402052,0.69907695,0.6301539,0.48246157,0.33805132,0.21989745,0.128,0.06564103,0.036102567,0.026256412,0.02297436,0.016410258,0.016410258,0.016410258,0.02297436,0.029538464,0.032820515,0.04266667,0.036102567,0.032820515,0.032820515,0.032820515,0.029538464,0.01969231,0.016410258,0.01969231,0.026256412,0.016410258,0.006564103,0.0032820515,0.006564103,0.016410258,0.016410258,0.016410258,0.006564103,0.0032820515,0.0032820515,0.013128206,0.02297436,0.052512825,0.07548718,0.101743594,0.18051283,0.33476925,0.55794877,0.7187693,0.81066674,0.94523084,0.92553854,0.93866676,0.8369231,0.60389745,0.37415388,0.3117949,0.23630771,0.190359,0.21989745,0.35446155,0.508718,0.574359,0.5973334,0.6104616,0.6301539,0.60389745,0.7778462,0.7811283,0.5349744,0.23958977,0.20348719,0.21989745,0.21989745,0.18379489,0.14441027,0.16082053,0.21333335,0.318359,0.5677949,1.148718,1.6738462,2.3630772,2.9111798,3.0523078,2.5435898,2.2121027,1.7001027,1.4506668,1.6475899,2.2121027,2.0545642,1.6902566,1.4473847,1.3620514,1.1881026,1.083077,1.1355898,1.1290257,0.9747693,0.7056411,0.5152821,0.38400003,0.27569234,0.18707694,0.15753847,0.15097436,0.13784617,0.14441027,0.16410258,0.17394873,0.20676924,0.21989745,0.24943592,0.3314872,0.49887183,0.6235898,0.79097444,0.98461545,1.0765129,0.8205129,0.60389745,0.46276927,0.37743592,0.31507695,0.21333335,0.14769232,0.118153855,0.108307704,0.108307704,0.08205129,0.101743594,0.098461546,0.08861539,0.09189744,0.1148718,0.18707694,0.24943592,0.34133336,0.44964105,0.5021539,0.48574364,0.4266667,0.36102566,0.3249231,0.3511795,0.46276927,0.5546667,0.52512825,0.4004103,0.3249231,0.27569234,0.24615386,0.2231795,0.20348719,0.16738462,0.19364104,0.2100513,0.2100513,0.2100513,0.21661541,0.17723078,0.14112821,0.11158975,0.09189744,0.07548718,0.380718,0.45620516,0.26256412,0.072205134,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06235898,0.14112821,0.17723078,0.15097436,0.07548718,0.06564103,0.02297436,0.0,0.01969231,0.09189744,0.07876924,0.08533334,0.10502565,0.14441027,0.2297436,0.26584616,0.45620516,0.6465641,0.892718,1.463795,3.8695388,6.925129,11.155693,17.604925,27.848207,38.416412,45.65662,49.99549,50.868515,46.706875,37.51713,29.879797,24.992823,22.826668,22.15713,21.592617,21.956924,23.689848,26.12185,27.464207,27.795694,26.368002,24.579285,23.233643,22.537848,21.635284,20.886976,20.256823,19.830154,19.80718,21.40554,19.104822,15.284514,11.480617,8.392206,7.1122055,8.372514,9.563898,9.69518,9.412924,7.3386674,9.714872,10.738873,8.562873,5.280821,4.8147697,3.748103,2.5928206,1.7493335,1.4802053,1.1126155,0.6465641,0.28225642,0.10502565,0.09189744,0.16410258,0.14769232,0.15753847,0.20020515,0.15097436,0.1148718,0.18051283,0.4660513,0.85005134,0.9616411,0.6301539,0.8598975,1.1946667,1.4276924,1.5885129,2.172718,1.8510771,1.3751796,1.1027694,0.9911796,1.017436,0.6104616,0.6104616,0.96492314,0.7318975,0.39056414,0.3249231,0.77456415,1.6640002,2.5796926,2.225231,1.3292309,0.64000005,0.7089231,1.8937438,1.270154,0.7384616,0.64000005,0.92553854,1.1454359,0.6432821,0.41025645,0.8598975,1.6672822,1.7394873,0.7253334,0.54482055,0.88287187,1.3850257,1.6771283,1.0929232,0.96492314,0.9288206,0.8041026,0.6104616,0.8172308,0.81394875,1.1257436,1.7165129,1.9823592,1.6311796,1.2668719,1.1618463,1.2373334,1.0535386,1.2242053,1.7427694,1.913436,1.6836925,1.6475899,1.3193847,1.3653334,1.3653334,1.1979488,1.0371283,1.1224617,1.7657437,2.3893335,2.9440002,3.9220517,4.7622566,6.633026,7.680001,6.8233852,3.7218463,4.2371287,5.32677,6.229334,6.7314878,7.171283,6.7577443,8.080411,9.770667,10.738873,10.177642,9.31118,7.9130263,6.557539,5.284103,3.5872824,5.3202057,6.377026,6.7183595,6.564103,6.3934364,5.3202057,5.681231,5.2414365,3.8006158,3.190154,3.8859491,3.7021542,3.1343591,3.4264617,6.5772314,8.467693,5.654975,3.5872824,4.0533338,5.1889234,8.116513,8.546462,7.9852314,7.5552826,7.9950776,6.616616,5.2742567,3.9351797,3.4888208,5.720616,5.979898,4.0467696,2.3269746,1.9462565,2.7766156,1.9823592,2.8291285,3.5380516,3.3903592,2.7306669,3.4034874,2.665026,2.6289232,4.06318,6.3934364,6.380308,5.408821,5.723898,6.193231,2.2744617,3.3247182,6.889026,9.498257,8.4972315,2.0742567,0.9517949,0.571077,0.42338464,0.37415388,0.65641034,0.7056411,1.1388719,1.529436,1.5195899,0.82379496,2.5206156,3.9876926,5.2447186,5.901129,5.156103,7.243488,6.889026,5.362872,3.8432825,3.4034874,4.0500517,4.073026,6.7840004,12.235488,17.227488,14.857847,8.664616,3.9023592,3.698872,9.032206,11.989334,9.091283,5.028103,2.937436,4.4242053,6.157129,7.433847,7.4699492,6.2555904,4.5489235,3.1671798,7.325539,16.177233,22.839796,14.404924,5.2742567,3.3280003,4.4964104,5.802667,5.3858466,6.0225644,6.4623594,8.897642,11.372309,7.781744,4.4734364,7.686565,10.266257,9.258667,5.8912826,7.8047185,4.578462,1.8445129,1.5688206,2.044718,8.379078,12.022155,10.893129,6.0258465,1.5556924,2.5337439,5.037949,9.580308,16.036104,23.666874,17.24718,11.943385,9.334154,9.216001,9.5835905,9.435898,11.779283,14.257232,16.324924,19.242668,25.002668,22.734772,22.002874,26.788105,35.492104,23.013746,18.287592,16.068924,13.650052,10.817642,9.340718,7.79159,5.5204105,2.8455386,1.0371283,0.90256417,0.6859488,0.49887183,0.34789747,0.15097436,0.09189744,0.14112821,0.22646156,0.31507695,0.4135385,0.47261542,0.36102566,0.29210258,0.33805132,0.4135385,0.33805132,0.23958977,0.18379489,0.21661541,0.3511795,0.3511795,0.2855385,0.21333335,0.18051283,0.2297436,0.26584616,0.37415388,0.62030774,0.90256417,0.97805136,0.6104616,0.26256412,0.072205134,0.04594872,0.04594872,0.37415388,1.1158975,1.3850257,0.9878975,0.4266667,0.40369233,0.5349744,0.4135385,0.098461546,0.12143591,0.6235898,0.58420515,0.5349744,0.54482055,0.21333335,0.190359,0.4594872,1.014154,1.5163078,1.2964103,0.9321026,1.6344616,1.8313848,1.5360001,2.3663592,1.4506668,1.0272821,1.1520001,1.4539489,1.1585642,0.46276927,0.1148718,0.0,0.0,0.0,0.0,0.0,0.0,0.032820515,0.16738462,0.13128206,0.16738462,0.118153855,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.34133336,0.4266667,0.3708718,0.27241027,0.19692309,0.2231795,0.38400003,0.53825647,0.7056411,1.083077,1.4605129,1.5655385,1.3095386,0.90256417,0.8533334,1.5130258,2.0808206,2.03159,1.5163078,1.3587693,0.636718,0.2297436,0.052512825,0.016410258,0.016410258,0.6268718,1.7657437,2.281026,1.9889232,1.7099489,1.086359,1.5885129,2.0644104,2.0873847,1.9528207,2.2449234,1.7526156,2.0676925,3.0162053,2.6256413,2.550154,2.2482052,2.487795,3.3936412,4.457026,5.2611284,5.618872,5.586052,5.8157954,7.5388722,7.269744,5.691077,4.1714873,3.56759,4.2272825,5.874872,8.546462,11.54954,13.279181,11.23118,6.3245134,5.5893335,7.77518,10.200616,8.772923,6.1374364,4.4996924,3.3575387,2.7602053,3.31159,3.6758976,3.751385,3.6594875,3.3608208,2.6387694,2.5796926,2.5632823,2.4418464,2.2580514,2.2580514,2.1956925,2.1169233,2.044718,1.9823592,1.9232821,1.8116925,1.6836925,1.5622566,1.6049232,2.1070771,4.352,5.654975,5.58277,4.44718,3.31159,2.5665643,1.847795,1.3062565,0.98133343,0.82379496,0.67610264,0.5874872,0.4955898,0.380718,0.25928208,0.16082053,0.09189744,0.049230773,0.026256412,0.016410258,0.016410258,0.02297436,0.029538464,0.029538464,0.029538464,0.04266667,0.04594872,0.04594872,0.04266667,0.029538464,0.029538464,0.02297436,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.009846155,0.0,0.0,0.0,0.026256412,0.068923086,0.118153855,0.16738462,0.25271797,0.36758977,0.53825647,0.761436,1.0075898,0.8467693,0.8008206,0.77456415,0.69251287,0.47261542,0.30194873,0.21333335,0.190359,0.21989745,0.3052308,0.39056414,0.44964105,0.44307697,0.4135385,0.47261542,0.6695385,0.67282057,0.5316923,0.3249231,0.16738462,0.2297436,0.3249231,0.47261542,0.571077,0.4135385,0.15425642,0.15425642,0.18707694,0.18379489,0.24287182,0.7187693,1.7263591,2.5764105,2.8947694,2.6387694,2.7503593,2.284308,1.9364104,1.785436,1.2964103,1.4802053,1.7001027,1.7723079,1.6508719,1.4178462,1.1881026,1.1191796,1.3587693,1.7427694,1.8149745,1.0601027,0.5677949,0.3117949,0.21989745,0.18379489,0.14769232,0.118153855,0.14441027,0.19692309,0.19692309,0.25928208,0.26584616,0.27241027,0.30194873,0.3511795,0.54482055,0.7975385,1.0601027,1.1979488,0.9911796,0.636718,0.4397949,0.33476925,0.27569234,0.21333335,0.17723078,0.13128206,0.0951795,0.08205129,0.108307704,0.108307704,0.098461546,0.07876924,0.06564103,0.09189744,0.15097436,0.20348719,0.27897438,0.3708718,0.44307697,0.5021539,0.46276927,0.41025645,0.37415388,0.3511795,0.37415388,0.446359,0.4955898,0.48246157,0.39712822,0.26256412,0.20020515,0.190359,0.19364104,0.16738462,0.15425642,0.15097436,0.16410258,0.18051283,0.16738462,0.118153855,0.07876924,0.06235898,0.06564103,0.07548718,0.636718,0.20348719,0.052512825,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.06564103,0.101743594,0.0951795,0.052512825,0.01969231,0.013128206,0.006564103,0.029538464,0.15097436,0.09189744,0.04266667,0.059076928,0.12143591,0.118153855,0.16410258,0.21989745,0.32164106,0.6235898,1.3915899,3.6791797,6.813539,11.552821,18.395899,27.602053,36.289642,41.747696,43.3559,40.67118,33.414566,28.215797,25.62954,24.54318,24.139488,23.876925,24.320002,26.518976,29.295591,31.53395,32.164104,30.628105,26.14154,22.547693,21.18236,20.87713,20.919796,20.483284,19.498669,18.566566,18.950565,19.242668,16.393847,12.465232,8.950154,6.76759,6.5017443,7.6767187,9.590155,10.827488,9.268514,7.5946674,6.0750775,4.5390773,3.1737437,2.546872,3.1474874,2.0512822,1.0404103,0.73517954,0.61374366,1.8871796,2.028308,1.204513,0.16410258,0.24943592,0.3052308,0.18707694,0.108307704,0.13456412,0.16410258,0.17723078,0.21661541,0.32164106,0.5677949,1.0601027,1.4309745,2.1070771,2.2646155,1.7591796,1.1355898,1.0568206,0.9944616,1.0043077,1.0272821,0.9189744,1.1684103,1.339077,1.204513,0.8041026,0.4135385,0.512,1.8740515,2.6617439,2.3663592,1.7985642,1.4244103,0.97805136,0.7187693,0.95835906,2.0742567,1.404718,0.9714873,0.7122052,0.54482055,0.37415388,0.16738462,0.101743594,0.508718,1.2865642,1.8970258,1.4605129,1.3653334,1.5261539,1.6475899,1.2274873,1.3062565,1.3718976,1.4441026,1.4769232,1.3784616,1.3522053,1.5392822,1.5786668,1.3981539,1.2274873,1.086359,0.9911796,0.99774367,1.2603078,2.0053334,0.9944616,1.2603078,1.7493335,1.8543591,1.4145643,1.1257436,1.0043077,1.0338463,1.1191796,1.086359,1.211077,1.5261539,1.9954873,2.6978464,3.8596926,6.987488,8.146052,7.0334363,5.1265645,5.687795,4.9427695,5.1364107,5.7435904,6.4065647,6.951385,6.2063594,5.2053337,5.0642056,6.229334,8.467693,8.100103,7.02359,5.5072823,3.7874875,2.0611284,2.6322052,4.4865646,5.8157954,5.789539,4.57518,4.565334,4.8640003,4.532513,3.5446157,2.7864618,3.7448208,4.010667,3.373949,3.1540515,6.186667,10.761847,8.78277,6.377026,6.055385,6.701949,6.8299494,6.0750775,5.464616,5.428513,5.8092313,4.8114877,4.2535386,3.7284105,3.367385,3.8432825,4.6539493,3.8662567,2.5928206,1.6475899,1.5327181,1.4309745,2.041436,3.1376412,4.066462,3.7185643,3.3378465,2.1300514,3.006359,7.9983597,18.271181,10.932513,5.904411,5.8157954,8.385642,6.409847,2.7241027,4.017231,5.4186673,4.71959,2.3794873,3.767795,2.7766156,1.3587693,0.7187693,1.2898463,1.0666667,1.401436,1.9331284,2.2416413,1.847795,1.8576412,1.9495386,2.733949,3.7185643,3.314872,4.3290257,4.588308,3.6627696,2.8422565,5.149539,4.1550775,5.3366156,8.700719,12.875488,15.104001,8.694155,6.8266673,6.4000006,5.7698464,4.7360005,4.4307694,4.2338467,5.0116925,6.186667,5.7435904,5.3103595,4.775385,5.1200004,6.669129,9.101129,4.2141542,5.467898,11.017847,15.668514,10.86359,6.4590774,4.1747694,4.391385,6.8463597,10.610872,12.885334,10.889847,7.9195905,5.2545643,2.1431797,2.166154,5.6418467,8.073847,7.512616,4.585026,5.9930263,5.221744,3.190154,1.9626669,4.7425647,7.581539,7.282872,5.110154,2.550154,1.3259488,5.8256416,7.243488,8.87795,11.431385,12.987078,10.295795,9.521232,12.5374365,18.599386,24.313438,23.650463,17.575386,13.29559,13.801026,17.860924,22.715078,22.455797,22.078362,24.218258,29.131489,24.625233,21.828924,19.203283,16.154257,13.039591,11.290257,8.746667,5.8814363,3.2656412,1.5753847,1.3128207,0.9419488,0.67282057,0.5284103,0.3249231,0.25271797,0.32820517,0.38400003,0.39056414,0.44964105,0.42338464,0.31507695,0.28225642,0.32820517,0.31507695,0.20348719,0.2100513,0.24615386,0.26256412,0.23958977,0.26912823,0.31507695,0.45292312,0.6071795,0.55794877,0.4004103,0.45292312,0.65969235,1.0535386,1.7690258,1.4244103,0.8763078,0.5284103,0.512,0.6695385,0.44964105,1.0272821,1.8182565,2.176,1.3784616,1.0732309,1.2504616,1.0601027,0.46933338,0.26912823,0.5152821,0.39712822,0.37415388,0.6301539,1.079795,1.0962052,0.6695385,0.76800007,1.5524104,2.3958976,2.3696413,2.4516926,2.422154,2.4943593,3.3050258,3.2196925,3.5183592,3.9581542,4.2436924,4.027077,3.245949,2.3171284,1.4736412,0.8336411,0.40369233,0.08205129,0.0,0.03938462,0.14441027,0.33805132,0.36102566,0.44964105,0.41025645,0.26584616,0.256,0.27569234,0.25271797,0.20676924,0.17066668,0.17066668,0.24943592,0.29210258,0.27897438,0.22646156,0.17394873,0.26584616,0.50543594,0.73517954,0.90912825,1.0699488,1.1651284,1.3522053,1.404718,1.394872,1.7099489,2.425436,2.5107694,1.7690258,0.6892308,0.44307697,0.21989745,0.08861539,0.029538464,0.016410258,0.026256412,0.90256417,1.9462565,2.481231,2.5173335,2.7831798,3.0490258,4.397949,5.425231,5.7501545,6.0061545,5.2447186,4.493129,4.6933336,5.7698464,6.626462,4.650667,3.570872,3.3903592,4.0467696,5.431795,6.6100516,7.2270775,8.51036,10.420513,11.664412,12.097642,11.099898,10.315488,10.049642,9.255385,10.404103,14.70359,19.255796,21.444925,18.944002,14.309745,9.012513,6.6395903,7.276308,7.4797955,5.7796926,5.2315903,5.225026,5.3431797,5.3727183,4.8114877,5.0051284,5.3037953,5.3136415,4.886975,4.2568207,3.9614363,3.882667,3.879385,3.7710772,3.623385,3.4789746,3.4100516,3.4297438,3.498667,3.2984617,3.0260515,2.8914874,3.4297438,5.474462,8.100103,7.5881033,5.8978467,4.33559,3.5446157,2.6617439,2.1300514,1.7723079,1.4933335,1.276718,1.1191796,1.017436,0.92225647,0.8041026,0.6629744,0.4955898,0.35774362,0.23302566,0.12143591,0.052512825,0.02297436,0.016410258,0.02297436,0.029538464,0.029538464,0.04266667,0.04594872,0.04594872,0.04594872,0.04266667,0.032820515,0.029538464,0.026256412,0.029538464,0.03938462,0.029538464,0.01969231,0.009846155,0.006564103,0.016410258,0.016410258,0.029538464,0.029538464,0.009846155,0.0,0.0,0.013128206,0.03938462,0.07876924,0.118153855,0.19364104,0.23958977,0.380718,0.6268718,0.8598975,0.9747693,0.8402052,0.69579494,0.6071795,0.48574364,0.31507695,0.31507695,0.3511795,0.33805132,0.20676924,0.26256412,0.29210258,0.29210258,0.31507695,0.47261542,0.6695385,0.5546667,0.38400003,0.3249231,0.4594872,0.6498462,2.6617439,3.2623591,2.038154,1.401436,0.51856416,0.18707694,0.14112821,0.24287182,0.48902568,0.5349744,0.95835906,1.6935385,2.428718,2.5895386,2.4746668,2.4057438,2.4648206,2.4910772,2.0906668,1.6672822,1.5458462,1.5556924,1.5655385,1.4802053,1.394872,1.3554872,1.394872,1.6213335,2.2416413,2.100513,1.4572309,0.8041026,0.40369233,0.26912823,0.20348719,0.16082053,0.15425642,0.17723078,0.19692309,0.2297436,0.24943592,0.26584616,0.28225642,0.30194873,0.380718,0.5513847,0.76800007,0.9747693,1.0896411,0.8041026,0.6301539,0.42994875,0.2231795,0.20020515,0.13456412,0.10502565,0.09189744,0.098461546,0.13128206,0.14112821,0.13456412,0.12143591,0.118153855,0.15097436,0.20348719,0.25271797,0.3117949,0.36430773,0.3708718,0.4201026,0.40697438,0.38728207,0.36758977,0.31507695,0.2986667,0.3314872,0.3708718,0.40369233,0.446359,0.36102566,0.27569234,0.2297436,0.21333335,0.16738462,0.17394873,0.17066668,0.14441027,0.098461546,0.059076928,0.049230773,0.049230773,0.049230773,0.052512825,0.06564103,0.6301539,0.12471796,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.032820515,0.16410258,0.2231795,0.20676924,0.18379489,0.16738462,0.101743594,0.01969231,0.026256412,0.049230773,0.055794876,0.06564103,0.07548718,0.029538464,0.01969231,0.04594872,0.036102567,0.08533334,0.12471796,0.3249231,0.92553854,2.2350771,4.1780515,6.5444107,9.80677,14.569027,21.592617,28.928001,32.479183,32.741745,30.552618,27.060514,25.747694,26.213745,28.448822,32.518566,38.580517,43.80226,44.73108,41.248825,35.488823,31.839182,28.599796,24.224823,21.185642,20.217438,20.325745,20.010668,19.472412,18.852104,18.356514,18.244925,16.479181,13.650052,10.66995,8.254359,6.931693,6.889026,7.5552826,8.477539,8.756514,7.0531287,6.012718,4.6244106,2.930872,1.4408206,1.1191796,1.394872,0.8402052,0.4397949,0.4201026,0.26912823,1.7558975,1.9659488,1.1881026,0.18707694,0.21661541,0.17723078,0.20020515,0.31507695,0.43651286,0.3708718,0.21661541,0.26256412,0.5677949,1.0436924,1.4309745,1.1520001,1.3653334,1.3686155,1.0568206,0.92225647,0.764718,0.7253334,0.7450257,0.7581539,0.67282057,0.81394875,0.84348726,0.69251287,0.49887183,0.58420515,0.761436,1.2471796,1.401436,1.0929232,0.6859488,0.85005134,0.85005134,0.7581539,0.7450257,1.0962052,1.0929232,1.7591796,1.8379488,1.1158975,0.42994875,0.3708718,0.45620516,0.8467693,1.394872,1.6738462,1.4966155,1.5721027,1.7788719,1.7591796,0.93866676,1.1979488,1.5491283,1.5622566,1.204513,0.83035904,0.95835906,1.2898463,1.4539489,1.332513,1.0732309,0.8795898,0.9156924,1.1585642,1.9298463,3.882667,1.6672822,0.99774367,1.4145643,2.4024618,3.3805132,1.6738462,1.148718,1.2242053,1.6443079,2.4713848,1.8740515,2.2121027,2.7963078,3.2853336,3.6791797,5.218462,5.464616,5.1265645,5.5532312,8.743385,7.0957956,6.2687182,6.6592827,7.975385,9.232411,8.326565,6.76759,5.7435904,5.858462,7.1089234,7.259898,6.521436,5.8420515,5.4514875,4.8836927,4.342154,4.8311796,6.0816417,6.9382567,5.366154,4.7360005,4.709744,4.5587697,4.023795,3.3247182,3.626667,3.3772311,2.9472823,3.2000003,5.4941545,9.291488,8.661334,7.1154876,6.5378466,7.181129,6.774154,5.431795,4.2305646,3.7054362,3.8465643,3.1770258,2.9965131,3.045744,2.9702566,2.3466668,3.2262566,3.6496413,3.570872,2.986667,1.9528207,1.7329233,1.8182565,2.8849232,4.2272825,3.7842054,4.0008206,2.5796926,2.8816411,5.6254363,8.881231,5.3234878,3.1474874,4.312616,7.059693,5.907693,2.5829747,3.2656412,3.5052311,2.156308,1.3489232,4.4242053,4.46359,2.7798977,0.96492314,0.86317956,1.214359,2.15959,3.8432825,5.4613338,5.2545643,3.2196925,2.4681027,2.7273848,3.0916924,2.0118976,3.186872,3.5446157,3.2328207,3.1015387,4.716308,3.6562054,4.2568207,6.11118,8.01477,7.962257,5.228308,9.091283,12.091078,10.617436,4.926359,2.7175386,5.0510774,7.9163084,8.736821,6.36718,6.452513,7.0432825,8.694155,11.063796,12.911591,7.9195905,5.832206,6.9842057,8.730257,5.464616,4.1550775,3.0260515,3.0654361,5.2709746,10.643693,10.929232,7.2172313,3.7251284,2.2416413,2.1136413,5.297231,9.26195,9.665642,6.409847,3.626667,6.2687182,7.128616,5.1200004,2.5304618,5.024821,6.2916927,8.274052,6.73477,2.546872,1.6705642,9.199591,9.780514,9.8363085,11.369026,11.953232,8.093539,8.480822,14.165335,24.12308,35.25908,26.167797,16.81395,11.59877,12.06154,16.876308,17.329231,19.908924,21.83549,22.793848,24.960001,27.14913,26.581335,22.528002,16.682669,13.174155,11.69395,8.851693,5.6418467,3.0654361,2.1398976,1.6278975,1.2077949,1.0601027,1.0436924,0.69579494,0.6301539,0.65312827,0.6826667,0.702359,0.761436,0.49230772,0.4266667,0.47917953,0.5021539,0.28882053,0.118153855,0.17723078,0.30194873,0.36758977,0.26912823,0.35774362,0.5152821,0.83035904,1.142154,1.017436,0.8369231,0.8566154,1.0469744,1.4506668,2.2055387,1.7920002,1.3718976,1.0043077,0.8205129,1.0535386,0.764718,0.96492314,2.156308,3.7842054,4.2174363,3.2295387,3.5380516,3.0687182,1.6213335,0.8467693,0.9911796,0.65969235,0.4660513,0.8533334,2.0939488,4.263385,3.5478978,2.1398976,1.7558975,3.6496413,3.8071797,4.056616,4.450462,5.1922054,6.6428723,6.3540516,6.485334,6.4623594,6.0816417,5.504,5.586052,5.7632823,5.2053337,3.8990772,2.6453335,2.097231,1.5360001,1.0043077,0.636718,0.6826667,0.72861546,0.7253334,0.7253334,0.7417436,0.7515898,0.7384616,0.6268718,0.51856416,0.41025645,0.21333335,0.3708718,0.3511795,0.26256412,0.21989745,0.3249231,0.3314872,0.48574364,0.7384616,0.9517949,0.88615394,0.93866676,1.148718,1.6475899,2.359795,3.0129232,2.484513,1.9035898,1.1224617,0.34789747,0.13128206,0.13456412,0.068923086,0.04594872,0.101743594,0.18707694,0.90584624,1.6607181,1.8674873,1.719795,2.1825643,2.4713848,4.2896414,5.861744,6.8430777,8.320001,8.500513,9.472001,11.907283,14.309745,13.013334,10.601027,8.982975,8.149334,8.687591,11.792411,13.046155,14.736411,16.748308,18.399181,18.44513,17.83795,16.91241,16.62359,16.361027,13.919181,13.170873,16.66954,22.459078,27.382156,27.090054,20.955898,17.660719,14.936617,11.831796,8.684308,6.994052,6.62318,6.8299494,7.1680007,7.509334,7.384616,7.53559,7.9097443,8.39877,8.845129,9.025641,8.333129,7.328821,6.4590774,6.045539,6.124308,6.226052,6.678975,7.3386674,7.5881033,6.62318,5.733744,6.1046157,7.8834877,10.180923,9.107693,7.3091288,5.6385646,4.457026,3.6102567,2.986667,2.6190772,2.3958976,2.2088206,1.9561027,1.723077,1.5524104,1.4145643,1.2865642,1.148718,0.9419488,0.7417436,0.5349744,0.33476925,0.190359,0.101743594,0.04594872,0.02297436,0.02297436,0.02297436,0.032820515,0.04266667,0.049230773,0.055794876,0.055794876,0.04266667,0.03938462,0.03938462,0.03938462,0.036102567,0.032820515,0.026256412,0.01969231,0.009846155,0.016410258,0.016410258,0.029538464,0.036102567,0.029538464,0.009846155,0.016410258,0.016410258,0.026256412,0.052512825,0.08861539,0.17723078,0.32164106,0.380718,0.3708718,0.4955898,0.77128214,0.7778462,0.6826667,0.5973334,0.5874872,0.39712822,0.32820517,0.29210258,0.23302566,0.13784617,0.30194873,0.33805132,0.2855385,0.26256412,0.446359,0.9189744,1.4834872,2.5698464,3.8498464,4.2338467,2.1825643,2.225231,2.3827693,1.9298463,1.3915899,0.6170257,0.26912823,0.16410258,0.20676924,0.37415388,0.40369233,0.5316923,1.2209232,2.1530259,2.231795,2.4910772,2.92759,3.0293336,2.7831798,2.6551797,2.5140514,2.0020514,1.6147693,1.4966155,1.4408206,1.4441026,1.4145643,1.3915899,1.4605129,1.7624617,2.0118976,2.1431797,1.9331284,1.3522053,0.5546667,0.3052308,0.20676924,0.17066668,0.17066668,0.21661541,0.23958977,0.256,0.26584616,0.27569234,0.28225642,0.2986667,0.37743592,0.5021539,0.6826667,0.9321026,0.9189744,0.8369231,0.574359,0.24615386,0.19692309,0.13128206,0.0951795,0.098461546,0.12143591,0.13784617,0.128,0.16410258,0.20020515,0.21333335,0.20348719,0.25271797,0.29538465,0.32820517,0.34789747,0.34133336,0.35446155,0.35446155,0.34789747,0.3249231,0.2855385,0.31507695,0.3314872,0.33805132,0.34133336,0.35774362,0.38728207,0.30851284,0.24943592,0.23958977,0.20348719,0.19364104,0.17723078,0.14441027,0.09189744,0.02297436,0.029538464,0.032820515,0.036102567,0.03938462,0.052512825,0.47589746,0.14769232,0.026256412,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.049230773,0.03938462,0.02297436,0.01969231,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.04266667,0.21333335,0.40369233,0.7515898,0.99774367,0.92225647,0.31507695,0.101743594,0.09189744,0.14769232,0.17394873,0.14112821,0.12471796,0.049230773,0.0,0.0032820515,0.01969231,0.03938462,0.07876924,0.3249231,1.0108719,2.4418464,4.312616,6.042257,7.7390776,10.059488,14.224411,18.953848,21.044514,21.589334,21.779694,22.928411,25.590157,29.505644,35.29518,43.008003,52.10585,57.025646,53.123287,44.435696,35.6759,32.23631,26.394258,22.098053,19.899078,19.777643,21.136412,21.024822,19.715284,18.619078,17.929848,16.656412,13.5778475,11.411694,9.961026,9.163487,9.107693,7.6964107,7.3583593,7.207385,6.669129,5.5072823,4.3552823,3.5577438,2.3926156,1.0436924,0.5940513,0.44307697,0.37415388,0.43323082,0.49230772,0.24287182,1.1191796,1.2635899,0.8369231,0.25271797,0.15097436,0.0951795,0.35774362,0.574359,0.5973334,0.5021539,0.4004103,0.6268718,0.97805136,1.2373334,1.1881026,0.6465641,0.54482055,0.5316923,0.5218462,0.702359,0.6662565,0.8172308,0.84348726,0.69579494,0.60389745,0.58092314,0.38400003,0.24287182,0.3117949,0.6859488,0.7417436,0.48246157,0.3314872,0.38728207,0.42994875,0.58420515,0.636718,0.5677949,0.42338464,0.31507695,0.571077,1.5031796,1.7920002,1.211077,0.6301539,0.6235898,0.8402052,1.2274873,1.5688206,1.4539489,1.5195899,1.5491283,1.7066668,1.7362052,0.9517949,1.0338463,1.4080001,1.5130258,1.2340513,0.8795898,0.81394875,0.9911796,1.1815386,1.2898463,1.3193847,1.6213335,1.3522053,1.3095386,2.2383592,4.8344617,2.8914874,1.4834872,1.5786668,2.9440002,4.1550775,2.6715899,2.4713848,2.9538465,3.9778464,5.865026,6.160411,6.997334,7.213949,6.3934364,4.84759,4.332308,3.9876926,4.768821,7.0400004,10.561642,9.061745,8.254359,8.4512825,9.737847,11.989334,11.815386,10.660104,9.232411,8.054154,7.450257,7.4207187,7.0859494,7.171283,7.683283,7.88677,6.432821,7.1154876,8.484103,9.045334,7.2631803,5.8518977,4.9427695,4.57518,4.562052,4.4996924,4.647385,3.9975388,3.2787695,3.190154,4.394667,7.030154,7.433847,6.941539,6.7183595,7.7423596,8.024616,6.189949,4.1682053,3.186872,3.7349746,3.3969233,3.255795,3.6135387,4.076308,3.5544617,4.2962055,4.818052,4.903385,4.4438977,3.4231799,3.0818465,2.9538465,3.4034874,3.9122055,3.0884104,3.7874875,2.861949,3.0129232,3.6890259,1.0666667,0.9353847,1.6705642,4.128821,6.8693337,6.170257,2.993231,3.515077,3.9122055,2.7864618,1.1946667,3.3247182,3.9581542,2.865231,1.0732309,0.88287187,1.1323078,1.9889232,3.6824617,5.395693,5.2611284,3.495385,2.7995899,2.9702566,3.2656412,2.3696413,3.43959,3.6430771,3.4592824,3.3805132,3.9220517,3.7842054,3.5577438,4.066462,4.8311796,4.066462,4.096,9.363693,13.5089245,12.560411,4.9427695,2.7011285,5.0576415,7.3649235,7.2992826,4.84759,5.4186673,7.1220517,8.858257,10.066052,10.725744,8.077128,7.13518,8.136206,9.104411,5.8190775,3.3903592,4.4045134,5.3694363,5.7435904,7.9524107,5.976616,3.0129232,2.162872,3.501949,4.073026,7.1023593,10.791386,10.939077,7.4108725,4.1452312,7.2631803,8.237949,6.491898,3.620103,3.3936412,5.6254363,10.33518,9.353847,3.8334363,4.2568207,13.636924,14.808617,12.721231,10.791386,10.929232,9.596719,9.334154,14.562463,24.474258,33.056824,20.004105,12.560411,10.722463,13.334975,18.084105,14.706873,18.389336,22.449232,23.80472,22.977642,25.714874,25.678772,22.344208,17.28,14.132514,11.621744,9.603283,7.5388722,5.2578464,2.9702566,2.5337439,2.0644104,1.7723079,1.595077,1.1848207,1.142154,1.083077,1.020718,0.99774367,1.083077,0.7417436,0.63343596,0.6662565,0.6662565,0.380718,0.23630771,0.32820517,0.45292312,0.48574364,0.40369233,0.56451285,0.78769237,1.1224617,1.404718,1.2537436,1.3653334,1.5327181,1.657436,1.8740515,2.5665643,2.7569232,2.2547693,1.5360001,1.0568206,1.2603078,1.1618463,1.0765129,2.100513,4.020513,5.3103595,4.4996924,4.650667,4.0992823,2.7470772,2.0775387,1.654154,1.4605129,1.7460514,2.422154,3.058872,4.7294364,3.7284105,2.8914874,4.279795,9.186462,8.917334,7.8736415,7.768616,9.176616,11.526565,11.053949,10.975181,10.35159,8.786052,6.439385,5.3760004,7.5946674,9.179898,8.78277,7.5946674,7.2861543,6.0685134,4.3060517,2.7142565,2.3630772,1.9954873,1.9692309,2.1333334,2.2613335,2.03159,1.7755898,1.8773335,1.8018463,1.4080001,0.94523084,1.1684103,1.4145643,1.7296412,2.0906668,2.4418464,2.5796926,2.6387694,2.7667694,3.0391798,3.436308,3.4855387,2.7306669,2.3236926,2.5206156,2.6715899,1.6246156,1.2832822,0.90912825,0.44964105,0.54482055,0.6826667,0.49230772,0.39384618,0.65641034,1.394872,1.2635899,1.3686155,1.3653334,1.332513,1.7788719,1.9035898,3.8334363,6.4656415,9.340718,12.63918,15.156514,18.372925,21.72718,23.814566,22.400002,22.416412,22.4919,21.513847,20.096,20.575182,21.00513,24.408617,28.609644,31.232002,29.69272,30.470566,29.922464,29.525335,28.737642,25.01908,22.17354,22.216208,26.49272,32.24944,32.60718,27.201643,25.790361,23.785027,19.190155,12.586668,9.042052,8.178872,8.579283,9.373539,10.233437,10.939077,11.565949,12.524308,13.61395,14.01436,14.171899,13.13477,11.648001,10.640411,11.234463,11.126155,11.07036,11.195078,11.234463,10.518975,8.884514,7.972103,8.687591,10.604308,11.943385,9.426052,7.5454364,6.242462,5.3202057,4.4045134,3.948308,3.5872824,3.3378465,3.131077,2.8291285,2.537026,2.3105643,2.100513,1.8970258,1.7263591,1.4834872,1.2274873,0.95835906,0.6892308,0.43323082,0.26584616,0.14769232,0.07548718,0.04594872,0.052512825,0.04594872,0.03938462,0.04594872,0.055794876,0.06235898,0.049230773,0.04594872,0.04266667,0.03938462,0.036102567,0.032820515,0.029538464,0.026256412,0.02297436,0.02297436,0.016410258,0.01969231,0.029538464,0.03938462,0.04594872,0.03938462,0.029538464,0.026256412,0.036102567,0.07548718,0.17066668,0.3446154,0.3708718,0.24943592,0.23958977,0.4397949,0.67938465,0.80738467,0.77128214,0.6268718,0.446359,0.34133336,0.26584616,0.21333335,0.20348719,0.39384618,0.40697438,0.31507695,0.256,0.4135385,1.0633847,2.3171284,3.82359,4.9952826,5.0084105,2.7076926,1.8182565,1.6213335,1.5360001,1.1093334,0.65969235,0.43323082,0.30851284,0.2297436,0.2231795,0.34789747,0.5218462,1.1093334,1.8904617,2.0644104,2.176,2.6026669,2.7208207,2.5665643,2.8324106,3.1409233,2.8389745,2.412308,2.0644104,1.7394873,1.4966155,1.3981539,1.3915899,1.404718,1.3292309,1.591795,2.0939488,2.3040001,2.0118976,1.3489232,0.92553854,0.48902568,0.2297436,0.18379489,0.2297436,0.24943592,0.256,0.25928208,0.26584616,0.27569234,0.27569234,0.30194873,0.380718,0.5218462,0.7220513,0.80738467,0.7581539,0.5513847,0.2986667,0.2297436,0.16410258,0.118153855,0.11158975,0.12143591,0.108307704,0.108307704,0.15425642,0.20676924,0.23302566,0.21661541,0.25928208,0.29538465,0.31507695,0.31507695,0.3117949,0.2855385,0.27569234,0.28225642,0.28882053,0.27569234,0.3052308,0.3117949,0.30194873,0.28882053,0.28882053,0.35774362,0.3249231,0.28882053,0.27897438,0.26584616,0.24943592,0.21333335,0.16738462,0.11158975,0.03938462,0.032820515,0.029538464,0.029538464,0.029538464,0.04594872,0.318359,0.17066668,0.052512825,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.11158975,0.0951795,0.059076928,0.03938462,0.0,0.07876924,0.14112821,0.13456412,0.06564103,0.0,0.0,0.0,0.0,0.01969231,0.098461546,0.37743592,1.204513,1.8412309,1.7329233,0.49230772,0.190359,0.14769232,0.22646156,0.318359,0.34133336,0.22646156,0.101743594,0.029538464,0.026256412,0.052512825,0.01969231,0.04266667,0.19692309,0.67938465,1.7920002,3.620103,5.2348723,6.2490263,6.997334,8.54318,10.000411,11.378873,13.105232,15.497848,18.770052,24.178873,30.998978,38.862774,46.76267,53.06421,52.749134,44.471798,35.92862,31.471592,32.137848,24.67118,20.09272,18.477951,19.623386,23.03672,24.070566,21.943796,19.419899,17.335796,14.621539,11.257437,9.911796,10.010257,10.925949,11.949949,8.592411,7.5552826,6.951385,6.0750775,5.4153852,4.0992823,3.0818465,1.9495386,0.86646163,0.58420515,0.39712822,0.48902568,0.65641034,0.67610264,0.30851284,0.40369233,0.508718,0.47589746,0.30851284,0.18051283,0.3446154,0.6662565,0.73517954,0.5481026,0.48902568,0.6268718,1.0436924,1.1782565,0.90912825,0.5481026,0.45292312,0.43651286,0.48574364,0.5481026,0.512,0.5218462,0.9189744,1.0568206,0.85005134,0.79097444,0.8402052,0.48246157,0.2297436,0.3249231,0.7450257,0.75487185,0.52512825,0.47261542,0.6662565,0.83035904,0.508718,0.34133336,0.3052308,0.318359,0.23302566,0.22646156,0.4266667,0.6104616,0.7220513,0.8566154,0.8336411,1.0568206,1.3850257,1.6180514,1.4802053,1.7887181,1.6049232,1.5622566,1.654154,1.2471796,1.024,1.3915899,1.7952822,1.9035898,1.6114873,1.0502565,0.9156924,0.98133343,1.1782565,1.6016412,2.989949,2.5862565,2.1267693,2.8553848,5.4974365,4.713026,2.7733335,2.4057438,3.6594875,3.889231,3.7415388,4.1813335,4.9920006,6.314667,8.628513,10.650257,11.818667,11.844924,10.417232,7.207385,6.0324106,5.8289237,7.2631803,9.8592825,12.022155,10.916103,10.420513,10.489437,11.497026,14.234258,15.2155905,15.031796,13.666463,11.631591,9.93477,9.206155,8.979693,9.202872,9.603283,9.665642,7.466667,9.219283,10.79795,10.492719,9.005949,7.273026,5.431795,4.6244106,4.9427695,5.4514875,5.802667,6.009436,5.3366156,4.1091285,3.7185643,5.4449234,6.3967185,6.7282057,6.987488,8.132924,9.222565,7.4371285,5.152821,4.0402055,5.093744,5.106872,4.7228723,4.844308,5.5138464,5.930667,6.298257,6.5805135,6.3179493,5.58277,4.97559,4.585026,4.7458467,4.709744,4.073026,2.7831798,2.9735386,2.9078977,3.6627696,4.342154,2.0742567,1.1684103,2.1924105,5.4941545,9.238976,9.412924,4.1813335,3.8006158,5.4416413,6.1538467,2.858667,1.8215386,1.9331284,1.7427694,1.1651284,1.467077,1.017436,1.2012309,1.7263591,2.231795,2.3138463,2.6978464,2.3827693,2.5173335,3.3575387,4.2601027,4.450462,4.1583595,3.626667,3.259077,3.626667,4.388103,4.076308,4.210872,4.818052,4.4406157,3.7874875,6.380308,9.91836,10.771693,3.9844105,2.934154,3.4231799,3.9056413,3.570872,2.3302567,2.537026,3.8498464,4.4373336,4.1714873,4.6211286,4.84759,7.683283,11.388719,13.243078,9.5606165,5.093744,8.3823595,10.660104,8.697436,4.7983594,2.1136413,1.6016412,3.95159,7.00718,5.7665644,6.052103,8.178872,10.006975,9.980719,7.138462,8.425026,8.018052,6.774154,4.8311796,1.6410258,6.2096415,11.073642,9.668923,4.6276927,7.752206,17.191385,18.464823,13.761642,7.6077952,6.8627696,11.884309,11.185231,13.984821,20.066463,19.761232,10.745437,8.845129,11.378873,16.111591,21.241438,16.787693,18.582975,22.872618,25.869131,23.762053,21.894566,20.470156,19.403488,18.25477,16.239592,12.235488,11.316514,10.9456415,9.048616,4.0041027,3.9220517,3.31159,2.612513,2.0578463,1.6738462,1.6902566,1.522872,1.2931283,1.148718,1.2340513,1.0272821,0.83035904,0.7417436,0.7089231,0.508718,0.47261542,0.58420515,0.6170257,0.5415385,0.5349744,0.72861546,0.94523084,1.276718,1.5589745,1.3522053,1.7394873,2.1431797,2.2153847,2.1956925,2.9078977,3.945026,3.2131286,2.1103592,1.4834872,1.6311796,1.6246156,1.4080001,1.7591796,2.7766156,3.8990772,4.345436,4.906667,5.3727183,5.4514875,4.7556925,2.6190772,2.5698464,3.8465643,5.221744,4.9788723,3.5413337,1.8609232,2.806154,7.4240007,14.933334,14.034052,11.260718,10.482873,12.665437,15.875283,15.911386,16.544823,16.65313,14.680616,8.628513,6.0816417,10.473026,14.55918,15.510976,14.897232,14.395078,12.731078,9.7903595,6.678975,5.6943593,5.152821,5.0084105,5.110154,5.152821,4.670359,3.817026,4.007385,3.95159,3.3411283,2.8521028,3.1474874,4.0434875,5.2053337,6.226052,6.626462,6.8955903,6.816821,6.449231,6.2687182,7.181129,6.925129,4.713026,2.7208207,1.6968206,0.9944616,0.5349744,1.0469744,1.2307693,1.0108719,1.522872,1.9823592,1.7296412,1.529436,1.9823592,3.5314875,2.556718,1.9790771,2.0250258,2.5206156,2.8882053,3.5347695,6.1013336,9.796924,14.122667,18.898052,24.359386,29.77149,32.94195,33.496616,32.896004,34.835693,36.325745,35.20985,31.343592,26.597746,27.421541,32.18708,38.606773,43.506874,42.834053,47.61272,48.397133,47.980312,46.664207,42.292515,37.349747,32.66954,33.046978,36.949337,36.512825,33.680412,31.977028,31.090874,28.662155,20.28636,14.208001,12.593232,13.019898,13.869949,14.326155,15.530668,16.873028,18.395899,19.584002,19.370668,18.471386,17.496616,16.745028,16.918976,19.124514,17.979078,16.961643,15.944206,14.634667,12.603078,11.053949,10.509129,10.781539,11.319796,11.1983595,10.259693,9.114257,7.975385,6.957949,6.058667,5.4974365,5.0215387,4.6539493,4.3585644,4.0303593,3.6660516,3.370667,3.0654361,2.740513,2.477949,2.1792822,1.8642052,1.5524104,1.2274873,0.8533334,0.57764107,0.3708718,0.2231795,0.13128206,0.1148718,0.072205134,0.04594872,0.03938462,0.049230773,0.06235898,0.052512825,0.049230773,0.04266667,0.032820515,0.04266667,0.036102567,0.032820515,0.032820515,0.029538464,0.029538464,0.01969231,0.01969231,0.02297436,0.04266667,0.08533334,0.06235898,0.052512825,0.04266667,0.03938462,0.07876924,0.17066668,0.29538465,0.35446155,0.3117949,0.20676924,0.17723078,0.5546667,0.90256417,0.94523084,0.55794877,0.45292312,0.38400003,0.3314872,0.30851284,0.33805132,0.47261542,0.5152821,0.446359,0.3446154,0.40697438,0.9156924,2.3302567,3.1442053,2.9407182,2.3696413,2.1267693,2.3630772,2.1924105,1.5031796,0.9419488,0.7581539,0.8598975,0.764718,0.4135385,0.18707694,0.32820517,0.6695385,1.1323078,1.6377437,2.1267693,1.7526156,1.7329233,1.8576412,2.0906668,2.550154,3.1081028,3.4691284,3.4724104,3.114667,2.5435898,1.8116925,1.4506668,1.3850257,1.4408206,1.3456411,1.3620514,1.5556924,1.8281027,2.0873847,2.2646155,1.7985642,1.0502565,0.52512825,0.34789747,0.26584616,0.25271797,0.25271797,0.24943592,0.24943592,0.27897438,0.28225642,0.30851284,0.380718,0.48574364,0.5513847,0.5513847,0.48246157,0.40697438,0.35446155,0.30851284,0.22646156,0.18379489,0.15097436,0.108307704,0.06235898,0.08861539,0.10502565,0.13456412,0.18051283,0.20348719,0.24943592,0.27241027,0.28225642,0.28225642,0.26584616,0.21661541,0.18707694,0.20676924,0.25271797,0.256,0.25928208,0.25271797,0.24287182,0.24615386,0.2855385,0.31507695,0.3314872,0.3314872,0.32164106,0.3117949,0.31507695,0.27569234,0.2100513,0.14112821,0.08205129,0.04266667,0.032820515,0.026256412,0.02297436,0.04266667,0.3052308,0.06235898,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.072205134,0.08205129,0.04594872,0.0,0.0,0.39056414,0.7089231,0.67610264,0.32820517,0.0,0.0,0.0,0.0,0.0,0.0,0.08533334,0.4004103,0.72861546,0.77128214,0.13784617,0.101743594,0.036102567,0.108307704,0.28225642,0.3052308,0.26912823,0.21333335,0.14769232,0.08861539,0.07548718,0.016410258,0.0,0.02297436,0.32820517,1.3883078,2.231795,4.0533338,5.3103595,5.7107697,6.2096415,6.7117953,8.146052,10.282667,12.701539,14.8020525,18.901335,23.83754,28.110771,31.054771,32.836926,31.494566,27.828514,24.996105,23.936003,23.361643,20.066463,17.391592,17.079796,19.813745,25.222567,27.26072,25.737848,22.193232,17.929848,14.024206,10.482873,9.048616,10.092308,12.268309,12.511181,9.485129,9.724719,9.065026,6.7840004,5.5991797,6.442667,5.408821,3.1803079,1.0108719,0.7187693,0.571077,0.6071795,0.73517954,0.7220513,0.19692309,0.03938462,0.08205129,0.13128206,0.18051283,0.4135385,1.1946667,0.9485129,0.69251287,0.6826667,0.4266667,0.53825647,0.67610264,0.6629744,0.5973334,0.8533334,0.8172308,0.6892308,0.67282057,0.7450257,0.67282057,0.47589746,0.53825647,0.6826667,0.8402052,1.020718,1.7165129,0.9124103,0.2297436,0.4135385,1.3423591,1.782154,1.214359,0.53825647,0.21989745,0.3052308,0.318359,0.27569234,0.45620516,0.7187693,0.48902568,0.6104616,0.57764107,0.60061544,0.86974365,1.5425643,1.4178462,1.3620514,1.4211283,1.6016412,1.847795,2.1136413,1.9790771,1.7624617,1.6377437,1.6640002,1.3226668,2.481231,3.18359,2.6486156,1.2832822,0.7187693,0.67938465,0.8402052,1.0666667,1.4178462,3.7251284,4.8607183,5.3070774,6.1341543,9.002667,7.5618467,4.417641,3.564308,5.3070774,6.2720003,4.4045134,4.010667,3.8695388,3.8301542,4.8082056,5.4416413,5.3727183,7.460103,10.456616,9.002667,8.832001,9.842873,12.416001,15.622565,17.194668,14.460719,11.874462,12.045129,14.562463,15.990155,16.955078,18.294155,17.897026,15.780104,14.083283,13.22995,12.0549755,11.720206,12.058257,11.58236,8.602257,7.200821,7.5946674,8.992821,9.567181,7.686565,6.193231,5.540103,5.425231,4.7917953,3.9614363,7.499488,9.6295395,8.310155,5.2348723,4.4767184,6.0192823,7.0859494,6.9120007,6.7282057,7.584821,7.8080006,7.0432825,5.8125134,5.5072823,5.861744,5.044513,3.8432825,3.170462,4.073026,3.4756925,5.927385,7.5913854,7.0498466,5.280821,4.2535386,5.0051284,6.189949,6.567385,5.0051284,3.7120004,3.7448208,4.6112823,5.152821,3.5413337,1.4539489,1.6082052,5.9536414,12.370052,14.6642065,6.521436,3.2951798,5.5729237,9.340718,5.9963083,2.225231,1.4112822,1.5130258,1.5031796,1.3587693,1.2964103,1.8576412,2.1103592,2.1431797,3.0818465,3.9844105,2.8488207,1.7132308,2.356513,6.2851286,5.333334,3.761231,2.9046156,3.1113849,3.7218463,3.9318976,4.7622566,4.7655387,3.767795,2.8521028,1.6344616,3.7251284,7.328821,9.284924,5.097026,4.6802053,4.9985647,5.0182567,4.210872,2.5632823,2.612513,2.0118976,2.4385643,3.754667,3.9975388,4.7425647,5.3858466,6.4722056,6.987488,4.348718,6.0816417,10.561642,12.803283,10.338462,3.2361028,1.6836925,2.048,4.667077,7.5388722,6.3179493,5.8912826,5.07077,7.200821,11.58236,13.472821,10.043077,7.4929237,6.045539,5.0215387,2.8389745,8.198565,10.341744,7.50277,3.515077,7.8112826,14.966155,10.850462,5.1626673,2.6880002,3.31159,10.148104,11.720206,12.616206,13.046155,8.835282,6.5411286,10.65354,13.436719,15.14995,24.047592,21.556515,18.563284,19.820309,24.95672,28.471798,23.686565,20.512821,18.884924,18.179283,17.227488,14.785643,13.08554,11.851488,9.849437,4.8836927,4.857436,4.0008206,3.0982566,2.477949,2.0151796,2.15959,1.8051283,1.394872,1.1585642,1.0994873,1.0010257,0.86646163,0.7187693,0.58420515,0.47261542,0.48574364,0.58092314,0.54482055,0.4135385,0.47261542,0.571077,0.69579494,1.4342566,2.3171284,1.8149745,1.7066668,2.0709746,2.284308,2.3827693,3.0654361,3.5544617,3.117949,2.6354873,2.5337439,2.7766156,2.2646155,1.9068719,1.6508719,1.6180514,2.1070771,4.082872,7.6701546,11.69395,13.751796,10.223591,4.535795,3.4330258,5.0871797,7.8112826,10.069334,7.752206,4.6080003,3.698872,5.6418467,8.621949,8.132924,7.499488,8.92718,12.544001,16.387283,17.939693,21.264412,25.744411,26.584618,14.831591,16.73518,22.577232,25.682053,24.579285,22.977642,19.682463,18.336823,15.730873,11.907283,10.161232,11.408411,10.538668,9.537642,9.225847,9.26195,7.3321033,6.2752824,5.87159,5.8912826,6.088206,6.8693337,8.546462,10.354873,11.52,11.277129,10.873437,10.407386,8.805744,6.6428723,6.117744,4.788513,2.550154,1.0994873,0.8008206,0.702359,0.65312827,0.9419488,1.4736412,2.097231,2.609231,3.9778464,4.1714873,4.0500517,4.2994876,5.4482055,5.3136415,4.821334,5.028103,5.8912826,6.2555904,9.196308,14.683899,17.88718,18.996513,23.207386,31.264822,39.12862,45.11508,46.61498,40.083694,35.334568,30.936617,27.913849,25.767387,22.44595,29.745234,33.713234,37.43508,42.883286,50.901337,58.53211,62.060314,63.48144,62.87426,58.39426,50.56985,42.929234,40.15262,42.11857,43.897438,40.723694,39.125336,41.54749,43.552822,33.811695,27.782566,25.760822,24.84513,23.35836,20.844309,21.697643,22.800411,22.98749,22.580515,23.361643,22.18995,22.216208,23.558565,25.62954,27.145847,23.958977,21.12,19.557745,19.035898,18.15631,17.975796,16.738462,15.182771,13.846975,13.075693,11.953232,10.9226675,9.9282055,8.937026,7.9491286,7.1548724,6.619898,6.294975,6.0947695,5.874872,5.2644105,4.7622566,4.348718,3.9680004,3.5413337,3.1606157,2.793026,2.4024618,1.9889232,1.585231,1.1355898,0.77456415,0.48902568,0.27569234,0.15097436,0.07876924,0.052512825,0.04594872,0.049230773,0.06235898,0.06235898,0.06235898,0.049230773,0.029538464,0.029538464,0.04266667,0.04594872,0.03938462,0.029538464,0.029538464,0.029538464,0.029538464,0.036102567,0.049230773,0.06235898,0.08533334,0.08205129,0.08205129,0.09189744,0.09189744,0.20020515,0.4135385,0.508718,0.4397949,0.3052308,0.19692309,0.34133336,0.5481026,0.6432821,0.47261542,0.48574364,0.45292312,0.36758977,0.27897438,0.28882053,0.5218462,0.88287187,0.9189744,0.6268718,0.44307697,0.45620516,1.2077949,1.7952822,1.9331284,1.9692309,2.359795,2.9144619,2.7503593,1.8215386,0.9321026,0.9321026,1.8642052,1.8707694,0.80738467,0.25928208,0.23630771,0.37415388,0.86974365,1.5655385,1.9692309,2.297436,2.1530259,2.0053334,1.9790771,1.8313848,2.4155898,2.937436,3.3969233,3.7185643,3.754667,2.7273848,1.7591796,1.3062565,1.4080001,1.6640002,1.5425643,1.5458462,1.7362052,2.03159,2.228513,1.9462565,1.719795,1.3915899,0.92553854,0.4135385,0.30194873,0.24615386,0.23630771,0.25271797,0.28882053,0.31507695,0.32820517,0.36102566,0.39384618,0.380718,0.4660513,0.47917953,0.45620516,0.42994875,0.44307697,0.3314872,0.29538465,0.24615386,0.15753847,0.06235898,0.049230773,0.055794876,0.09189744,0.15425642,0.2297436,0.30194873,0.3117949,0.29210258,0.26584616,0.2297436,0.18051283,0.15753847,0.15097436,0.15753847,0.18379489,0.24287182,0.26912823,0.24287182,0.21333335,0.27569234,0.3249231,0.3446154,0.3446154,0.3249231,0.27569234,0.2986667,0.31507695,0.28225642,0.20348719,0.108307704,0.059076928,0.036102567,0.029538464,0.029538464,0.029538464,1.1946667,0.23958977,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016410258,0.08533334,0.35446155,0.45620516,0.508718,0.47261542,0.17066668,0.25928208,0.4135385,0.40697438,0.21333335,0.0,0.0,0.0,0.0,0.0,0.0,0.04594872,0.101743594,0.16410258,0.19692309,0.15097436,0.21989745,0.23302566,0.23302566,0.2231795,0.15753847,0.15097436,0.20676924,0.23302566,0.17394873,0.016410258,0.0032820515,0.0,0.032820515,0.17394873,0.5349744,1.404718,3.1474874,4.594872,5.2053337,5.0642056,5.58277,6.764308,8.356103,10.532104,13.909334,17.77559,21.563078,24.07713,25.140514,25.586874,25.504822,24.113234,21.96349,19.534771,17.234053,16.25272,16.406975,17.089642,18.638771,22.317951,23.96554,23.604515,22.25231,20.581745,18.930874,16.738462,13.991385,11.972924,10.758565,9.216001,7.6931286,6.5805135,5.5663595,4.903385,5.428513,5.674667,5.3037953,3.7907696,1.6705642,0.55794877,0.5677949,0.57764107,0.4660513,0.24287182,0.03938462,0.006564103,0.5513847,0.86974365,0.98461545,1.7558975,1.5983591,1.1651284,0.7515898,0.508718,0.4266667,1.211077,1.0043077,0.6268718,0.512,0.7187693,0.5874872,0.5513847,0.81394875,1.1191796,0.7450257,0.73517954,0.761436,0.8008206,0.9944616,1.6443079,3.308308,2.4352822,1.0699488,0.37743592,0.65969235,0.81394875,0.6662565,0.5218462,0.508718,0.574359,0.8992821,0.69251287,0.55794877,0.65312827,0.69579494,1.3456411,1.0338463,1.1224617,1.9331284,2.7602053,1.9659488,1.7165129,1.7362052,1.8773335,2.1530259,2.166154,1.7690258,1.7329233,2.2580514,3.006359,1.9889232,1.5031796,1.8510771,2.6157951,2.6354873,1.2340513,0.8041026,0.9911796,1.3620514,1.394872,2.100513,2.5140514,3.0916924,4.4964104,7.5979495,6.5312824,4.4373336,3.82359,4.7392826,4.7950773,3.7185643,3.3969233,3.3214362,3.3969233,3.95159,4.529231,4.972308,7.02359,9.097847,6.2687182,5.9995904,7.27959,9.511385,12.045129,14.158771,13.824001,11.136001,10.866873,13.39077,14.674052,14.943181,15.750566,15.497848,14.309745,14.060308,14.171899,12.829539,11.785847,11.864616,12.960821,11.680821,11.0605135,10.345026,9.498257,9.212719,8.720411,7.9524107,7.3419495,7.282872,8.123077,4.197744,4.647385,7.2303596,8.825437,5.4153852,4.1222568,5.208616,6.633026,7.381334,7.460103,9.596719,10.233437,9.3078985,7.4141545,5.789539,7.394462,7.003898,5.605744,4.210872,3.8531284,2.4648206,3.0982566,4.082872,4.397949,3.692308,2.28759,2.297436,3.3050258,4.2207184,3.2853336,4.6080003,5.5597954,6.445949,6.961231,6.1997952,3.2065644,1.6311796,3.498667,7.75877,10.31877,5.83877,2.868513,2.5337439,3.7842054,3.3969233,2.0939488,1.3489232,1.3357949,1.7952822,2.028308,3.1113849,4.1058464,3.9876926,3.43959,4.827898,4.128821,2.172718,1.2635899,2.5600002,6.0783596,6.180103,5.149539,4.0008206,3.5347695,4.322462,4.919795,5.8486156,5.730462,4.4996924,3.3903592,5.431795,7.834257,8.43159,6.764308,4.069744,4.6900516,5.346462,5.1659493,4.3749747,4.309334,4.2502565,4.069744,3.7054362,3.6036925,4.706462,3.8104618,2.6978464,2.103795,1.9593848,1.3817437,1.7001027,3.7973337,4.571898,3.3247182,1.7460514,3.6332312,3.9975388,4.916513,8.03118,14.54277,17.027283,9.800206,4.4406157,5.0477953,8.237949,7.433847,7.50277,6.73477,4.821334,2.8488207,4.9493337,7.4699492,7.509334,6.3245134,9.350565,8.838565,5.208616,3.1081028,3.6463592,4.384821,5.9470773,7.8703594,10.115283,10.8767185,6.5772314,6.088206,9.993847,12.635899,13.761642,18.530462,29.59426,25.74113,19.478975,18.28431,24.602259,25.540926,23.013746,19.67918,17.145437,15.970463,16.613745,14.808617,11.812103,8.690872,6.311385,5.904411,5.3792825,4.71959,3.8071797,2.4155898,2.281026,2.1169233,1.8674873,1.5491283,1.2438976,1.0699488,1.017436,0.892718,0.6662565,0.49887183,0.508718,0.56123084,0.6104616,0.73517954,1.1191796,1.079795,1.0896411,1.4736412,2.0217438,2.0118976,1.8313848,2.225231,2.5796926,2.7667694,3.1277952,3.8596926,3.6824617,3.367385,3.1770258,2.8750772,2.1464617,1.8838975,1.7329233,1.4998976,1.1290257,2.1497438,4.7458467,7.936001,9.701744,6.9645133,2.7798977,2.9768207,5.398975,8.677744,12.25518,9.849437,6.521436,4.2896414,4.3060517,6.8627696,8.710565,6.6002054,7.4797955,12.3076935,16.04595,17.578669,20.128822,24.746668,26.164515,12.816411,12.133744,21.041233,26.292515,24.582565,22.564104,21.320208,20.243694,17.746052,14.572309,13.810873,17.391592,18.898052,18.504206,17.079796,16.219898,13.568001,10.768411,9.53436,9.954462,10.482873,10.325335,10.502565,10.709334,10.811078,10.860309,10.154668,10.295795,9.012513,6.314667,4.4701543,3.4822567,2.5173335,2.359795,3.4100516,5.6943593,6.2884107,4.594872,3.3378465,3.2262566,2.937436,4.2568207,7.0990777,8.960001,9.347282,9.780514,9.002667,7.896616,8.493949,10.994873,13.761642,17.194668,22.002874,23.962257,25.156925,33.985645,42.47303,50.64862,55.06626,55.581543,55.378056,48.413544,41.32103,35.314873,31.015387,28.438976,34.215385,37.00185,39.926155,43.716927,46.71672,49.923286,52.07303,55.171288,59.250877,62.385235,62.01108,56.18872,51.817028,52.66708,59.38872,57.173336,55.460106,54.13744,51.597134,44.737644,38.229336,34.031593,30.792208,28.002464,26.006977,24.12636,22.678976,23.243488,26.079182,30.12267,30.12267,30.034054,30.726566,32.452927,34.835693,30.897234,27.181952,25.088001,24.690874,24.74995,25.426054,24.434874,21.3399,17.207796,14.601848,13.039591,12.22236,11.369026,10.368001,9.7673855,9.15036,8.664616,8.254359,7.837539,7.315693,6.803693,6.2030773,5.602462,5.074052,4.6867695,4.348718,3.9876926,3.698872,3.4789746,3.2229745,2.5961027,1.913436,1.3489232,0.92225647,0.50543594,0.29538465,0.18379489,0.15753847,0.15425642,0.049230773,0.059076928,0.06235898,0.052512825,0.04266667,0.04266667,0.036102567,0.03938462,0.03938462,0.029538464,0.029538464,0.029538464,0.02297436,0.01969231,0.02297436,0.036102567,0.072205134,0.098461546,0.10502565,0.08861539,0.07876924,0.2100513,0.32164106,0.4135385,0.4660513,0.4397949,0.25271797,0.2231795,0.35774362,0.52512825,0.47261542,0.4266667,0.4004103,0.36758977,0.30851284,0.20348719,0.7187693,0.9747693,0.90912825,0.69579494,0.74830776,0.8467693,1.719795,2.8717952,3.7218463,3.5905645,3.1245131,3.1409233,3.0162053,2.5206156,1.8346668,1.657436,1.9035898,1.7723079,1.1093334,0.39384618,0.32164106,0.4135385,0.7122052,1.2438976,2.0184617,2.3171284,2.477949,2.5862565,2.6322052,2.5140514,2.231795,2.477949,2.9144619,3.249231,3.2295387,3.629949,2.7667694,1.8248206,1.4080001,1.5163078,1.5031796,1.5360001,1.6607181,1.7624617,1.5688206,1.394872,1.394872,1.401436,1.3357949,1.204513,0.5973334,0.36758977,0.29210258,0.24943592,0.21661541,0.25928208,0.26584616,0.28225642,0.31507695,0.3314872,0.39712822,0.44307697,0.45620516,0.446359,0.41682056,0.36758977,0.3314872,0.2855385,0.2231795,0.14769232,0.1148718,0.101743594,0.13456412,0.20348719,0.26584616,0.318359,0.3249231,0.2986667,0.27569234,0.27897438,0.24943592,0.2231795,0.18379489,0.14112821,0.14769232,0.19692309,0.24287182,0.24615386,0.23958977,0.2986667,0.318359,0.37743592,0.42994875,0.43651286,0.34789747,0.3446154,0.3511795,0.33476925,0.27897438,0.18051283,0.11158975,0.06235898,0.03938462,0.029538464,0.029538464,0.57764107,0.1148718,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.04266667,0.21333335,0.29538465,0.35446155,0.35446155,0.16738462,0.19364104,0.18051283,0.13456412,0.072205134,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.016410258,0.029538464,0.052512825,0.06235898,0.101743594,0.2986667,0.41025645,0.318359,0.049230773,0.049230773,0.08205129,0.101743594,0.07876924,0.0,0.0,0.0,0.059076928,0.16410258,0.2297436,0.98461545,2.678154,4.20759,4.9460516,4.7655387,4.844308,5.717334,7.3649235,9.895386,13.512206,16.121437,18.566566,19.951591,20.663797,22.354053,22.373745,21.3399,19.065437,16.091898,13.679591,14.020925,15.29436,16.577642,17.749334,19.505232,20.614565,21.48431,22.593643,23.732515,24.001642,23.896618,21.930668,18.218668,13.745232,10.377847,9.179898,7.2894363,5.4580517,4.4832826,5.1856413,5.904411,5.602462,4.0992823,1.9790771,0.60061544,0.45292312,0.30194873,0.16082053,0.06235898,0.06564103,0.43651286,1.5392822,1.8215386,1.3292309,1.7066668,1.4473847,1.1585642,0.73517954,0.47261542,1.0601027,1.2635899,0.86646163,0.5940513,0.6695385,0.8041026,1.211077,1.2570257,1.2668719,1.2964103,1.1388719,1.1323078,0.8467693,0.6465641,0.6695385,0.8402052,1.719795,1.9922053,1.6869745,1.0732309,0.6629744,1.1716924,0.955077,0.79097444,1.014154,1.5392822,1.9922053,1.5983591,1.1027694,0.86974365,0.8763078,2.1267693,1.6705642,1.6213335,2.4976413,3.1967182,1.8215386,1.8379488,2.1267693,2.2416413,2.4188719,2.3794873,2.1070771,1.8051283,1.7952822,2.5173335,2.7700515,1.9364104,1.7624617,2.6847181,3.8367183,2.3991797,1.8084104,2.3794873,3.7120004,4.713026,4.056616,3.3476925,2.7700515,2.8291285,4.33559,4.466872,3.5183592,2.9472823,2.9472823,2.4484105,2.2219489,2.4155898,2.7766156,3.170462,3.6004105,4.6900516,6.7872825,7.79159,7.1089234,5.648411,5.9569235,7.6603084,9.895386,11.753027,12.3076935,14.260514,12.340514,10.9456415,11.477334,12.320822,12.688411,12.678565,12.580104,12.681848,13.275898,13.095386,11.651283,10.886565,11.355898,12.251899,12.2847185,14.070155,14.224411,11.871181,8.63836,8.572719,8.503796,8.549745,8.602257,8.326565,5.0674877,3.9417439,5.0871797,6.99077,6.47877,4.896821,5.3169236,7.194257,9.065026,8.549745,9.179898,9.750975,8.736821,6.482052,5.208616,7.1187696,7.177847,5.910975,4.3027697,3.8006158,3.4789746,2.7798977,2.9111798,3.82359,4.2207184,5.435077,5.9569235,5.7501545,4.640821,2.3138463,4.1517954,5.1922054,5.58277,6.2687182,9.009232,7.7325134,4.201026,2.6880002,3.8564105,4.7360005,4.0008206,2.5796926,1.8576412,2.1924105,2.9111798,3.2886157,3.3641028,2.7109745,1.847795,2.2514873,5.3924108,6.62318,5.7665644,4.1550775,4.634257,3.0424619,2.0217438,2.0545642,3.121231,4.699898,5.7764106,5.8420515,5.0642056,4.06318,3.9122055,4.1747694,4.4767184,4.378257,4.194462,4.9985647,9.114257,11.414975,9.977437,6.2129235,4.8672824,6.11118,5.2480006,4.269949,4.4734364,6.4557953,7.9228725,9.196308,8.841846,6.675693,3.7842054,2.1989746,1.2800001,1.0699488,1.3128207,1.463795,1.0108719,1.4966155,2.4713848,3.7842054,5.5663595,6.173539,4.516103,3.511795,5.4547696,12.032001,15.911386,8.779488,2.674872,2.038154,3.7218463,3.6430771,4.4701543,4.2272825,2.7569232,1.719795,4.2174363,8.329846,10.299078,10.233437,12.1238985,8.14277,4.315898,3.3936412,4.7589746,4.453744,3.767795,5.1232824,7.4436927,8.651488,5.654975,6.409847,10.522257,13.046155,14.578873,21.241438,33.060104,29.239798,20.837746,16.088617,20.404514,22.875898,23.168001,22.016,19.794052,16.489027,17.463797,15.90154,12.435693,8.720411,7.4174366,6.675693,5.989744,5.868308,5.677949,3.6430771,2.8127182,2.5632823,2.425436,2.1530259,1.7132308,1.5163078,1.2603078,1.017436,0.81066674,0.60389745,0.5513847,0.65641034,0.75487185,0.9156924,1.4375386,1.3357949,1.148718,1.2242053,1.5360001,1.7132308,1.8674873,2.1267693,2.3630772,2.5206156,2.6026669,3.2722054,3.18359,2.8849232,2.7044106,2.733949,2.231795,2.0644104,1.9593848,1.6771283,1.0404103,1.1848207,2.4155898,4.0434875,5.1659493,4.6834874,2.802872,3.245949,5.2709746,7.9983597,10.404103,7.4896417,6.189949,6.301539,7.3058467,8.346257,11.881026,11.680821,10.289231,9.691898,11.300103,17.096207,19.216412,20.919796,20.499695,11.286975,12.389745,20.20431,24.618668,23.847387,24.457848,27.02113,25.271797,22.396719,20.814772,22.176823,23.322258,24.556309,23.273027,19.777643,17.253744,15.727591,14.431181,15.553642,18.185848,18.320412,15.094155,13.121642,11.497026,10.233437,10.243283,11.638155,13.6467705,13.929027,11.746463,7.975385,7.4830775,6.9382567,6.738052,6.997334,7.5552826,7.7718983,5.989744,4.397949,4.1911798,5.546667,7.0957956,9.603283,12.501334,14.887385,15.53395,14.240822,12.872206,13.725539,17.742771,24.500515,27.218054,28.75077,31.43549,36.775387,45.43344,55.325542,59.795696,59.55939,56.976414,56.064003,54.564106,52.713028,52.40452,54.061954,56.641644,55.138466,52.78195,51.33785,51.19016,51.344414,53.927387,55.158157,56.933746,59.86134,63.248417,69.46134,69.09047,67.531494,69.35303,78.28677,74.8078,70.00616,64.65642,58.098877,48.239594,39.27303,37.093746,35.226257,31.396105,27.546259,24.674463,23.282873,24.953438,28.649029,30.71672,30.614977,31.382977,33.48349,36.181335,37.572926,34.310566,32.292107,31.48472,31.294361,30.552618,27.972925,26.768412,24.362669,20.667078,18.07754,16.436514,15.704617,14.65436,13.292309,12.842668,12.143591,11.552821,10.952206,10.240001,9.314463,8.67118,7.7948723,6.951385,6.3179493,5.9634876,5.684513,5.21518,4.844308,4.6867695,4.667077,3.7152824,3.0326157,2.4451284,1.8674873,1.2898463,0.8992821,0.6695385,0.49230772,0.3446154,0.28225642,0.13456412,0.1148718,0.101743594,0.1148718,0.32164106,0.11158975,0.049230773,0.03938462,0.029538464,0.029538464,0.02297436,0.016410258,0.016410258,0.01969231,0.029538464,0.059076928,0.098461546,0.12143591,0.1148718,0.10502565,0.15097436,0.190359,0.27241027,0.39384618,0.47261542,0.30194873,0.21333335,0.2297436,0.3052308,0.318359,0.33805132,0.32820517,0.32820517,0.318359,0.2297436,0.47917953,0.5677949,0.6235898,0.7220513,0.8960001,1.3062565,3.045744,4.2568207,4.31918,3.879385,2.858667,3.6135387,4.1156926,3.5216413,2.169436,2.2711797,2.100513,1.6640002,1.0305642,0.35446155,0.2986667,0.3249231,0.512,0.8763078,1.3718976,1.8018463,2.2022567,2.4484105,2.5928206,2.8488207,2.993231,2.8980515,2.665026,2.4320002,2.3729234,2.802872,2.7963078,2.5238976,2.284308,2.5042052,1.9593848,1.7362052,1.7493335,1.8182565,1.6508719,1.657436,1.2668719,0.9124103,0.77128214,0.77128214,0.4266667,0.32164106,0.2986667,0.27897438,0.25271797,0.25928208,0.256,0.26912823,0.29538465,0.3117949,0.35774362,0.41025645,0.46276927,0.49230772,0.48574364,0.45620516,0.40369233,0.3511795,0.30194873,0.24943592,0.20020515,0.16082053,0.15425642,0.18379489,0.2297436,0.26256412,0.27241027,0.27241027,0.27569234,0.318359,0.29210258,0.24615386,0.19364104,0.14769232,0.118153855,0.14441027,0.20676924,0.24287182,0.25271797,0.26912823,0.3249231,0.39056414,0.45620516,0.47917953,0.40369233,0.38400003,0.36430773,0.34133336,0.30851284,0.26256412,0.15097436,0.07876924,0.03938462,0.029538464,0.02297436,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.04266667,0.07548718,0.10502565,0.128,0.12471796,0.11158975,0.052512825,0.01969231,0.029538464,0.029538464,0.006564103,0.0,0.0,0.0,0.0,0.0,0.006564103,0.072205134,0.15097436,0.09189744,0.14112821,0.24943592,0.3052308,0.23302566,0.0,0.02297436,0.032820515,0.09189744,0.13784617,0.0,0.0,0.0,0.055794876,0.13784617,0.12471796,0.62030774,2.0086155,3.387077,4.210872,4.3027697,4.2240005,5.277539,7.2336416,9.668923,11.940104,13.315283,14.890668,15.954053,16.78113,18.642054,19.2,18.5239,16.62031,14.313026,13.243078,12.901745,14.070155,15.694771,16.918976,17.106052,17.522873,19.114668,21.366156,23.584822,24.917336,26.12185,25.554052,22.235899,16.869745,11.808822,9.8363085,8.152616,6.6625648,5.435077,4.6966157,4.9493337,4.7228723,3.6857438,2.100513,0.85005134,0.61374366,0.4135385,0.190359,0.01969231,0.101743594,0.56123084,1.4703591,2.0906668,2.1792822,1.9922053,1.8510771,1.1848207,0.62030774,0.55794877,1.1684103,1.014154,0.85005134,0.79425645,0.8008206,0.65312827,1.1815386,1.2537436,1.1290257,1.0338463,1.1618463,1.1257436,0.7778462,0.5152821,0.4397949,0.3446154,0.36102566,1.1126155,1.6804104,1.7033848,1.3817437,2.048,1.8445129,1.585231,1.7427694,2.4418464,2.6026669,2.03159,1.2800001,0.88615394,1.4080001,2.5337439,1.9889232,1.7460514,2.3269746,2.8160002,1.6804104,2.1398976,2.8258464,2.9538465,2.3171284,2.3335385,2.2711797,2.1530259,1.9922053,1.7920002,2.3958976,1.7920002,1.4473847,1.9790771,3.1573336,2.4352822,1.8970258,2.3072822,3.6594875,5.1954875,4.348718,3.5577438,2.7536411,2.1497438,2.225231,2.6715899,2.7142565,2.7175386,2.5435898,1.5491283,1.5885129,2.156308,2.7864618,3.1540515,3.0687182,4.0500517,6.2227697,6.75118,5.7698464,6.380308,6.75118,8.257642,10.699488,12.668719,11.539693,13.584412,12.970668,12.379898,12.416001,11.611898,10.84718,10.121847,10.541949,12.015591,13.233232,12.521027,11.244308,10.545232,10.453334,9.90195,9.796924,11.674257,12.599796,11.385437,8.595693,8.631796,8.825437,9.393231,10.010257,9.796924,6.7183595,4.388103,3.9975388,5.4875903,7.5421543,5.901129,5.3924108,6.816821,9.124104,9.393231,8.684308,9.012513,8.402052,6.701949,5.612308,7.975385,8.27077,7.000616,5.1626673,4.2436924,4.31918,3.8071797,3.6496413,4.571898,7.076103,8.937026,8.146052,6.4754877,4.7261543,2.6978464,4.785231,5.5532312,4.9526157,4.637539,7.9524107,7.899898,4.4734364,2.7076926,3.501949,3.6135387,3.1113849,2.3204105,2.034872,2.409026,2.9735386,4.332308,5.2348723,4.8738465,3.8301542,4.069744,6.2096415,6.11118,4.97559,3.9056413,3.9122055,3.1770258,4.164923,5.668103,6.5411286,5.717334,5.080616,5.2709746,5.661539,5.8125134,5.474462,5.421949,5.0904617,4.388103,4.013949,5.4580517,8.802463,9.908514,8.096821,5.3005133,6.038975,7.2927184,5.9634876,6.170257,8.4512825,9.770667,8.310155,9.18318,9.432616,7.394462,2.7109745,1.2274873,1.2964103,2.4320002,3.7218463,3.820308,2.0578463,2.038154,3.7349746,5.9634876,6.373744,5.100308,3.4002054,2.6157951,3.4560003,6.0028725,8.43159,4.8738465,1.7493335,1.2340513,1.2832822,1.211077,1.7985642,1.8740515,1.3029745,1.0043077,5.0215387,7.181129,8.057437,8.963283,11.972924,10.44677,7.6767187,6.813539,7.3419495,5.074052,4.2240005,5.7435904,8.155898,9.366975,6.6428723,7.460103,10.952206,13.197129,15.940925,26.59118,33.70339,28.580105,20.529232,15.980309,18.474669,18.924309,19.761232,19.961437,19.124514,17.490053,18.628925,17.42113,14.050463,10.236719,9.242257,8.198565,7.650462,7.397744,6.741334,4.4996924,3.7842054,3.7284105,3.3903592,2.6387694,2.169436,2.0873847,1.7099489,1.3686155,1.1782565,1.024,0.84348726,1.0075898,1.1552821,1.2438976,1.5458462,1.4802053,1.270154,1.148718,1.1749744,1.2307693,1.585231,1.9954873,2.422154,2.6420515,2.231795,2.5140514,2.2514873,1.972513,2.0118976,2.5074873,2.8455386,2.858667,2.7536411,2.3991797,1.3226668,2.0020514,2.0217438,2.0808206,2.4188719,2.8160002,3.8695388,5.6287184,7.4240007,8.457847,7.79159,6.87918,8.277334,10.331899,11.542975,10.561642,14.257232,15.681643,14.55918,12.727796,14.12595,18.642054,19.232822,19.994259,19.928617,12.954257,15.182771,22.14072,26.026669,25.826464,27.332926,33.194668,32.784412,31.763695,32.623592,34.658463,32.26913,32.196926,28.435694,21.192207,16.889437,18.074257,18.838976,21.14954,23.70954,21.96349,18.248207,16.695797,15.484719,14.41477,14.8939495,18.021746,21.973335,23.926155,22.442669,17.460514,16.049232,14.690463,12.714667,10.144821,7.6898465,7.9819493,7.50277,8.464411,11.894155,17.631182,18.399181,19.524925,21.769848,24.359386,24.992823,25.458874,24.743387,25.714874,29.636925,36.17149,38.03898,36.857437,38.206364,43.542976,50.20226,56.385647,58.482876,58.564926,57.40308,54.47549,56.782772,59.1918,63.75057,70.32452,76.60308,74.03323,70.0357,66.061134,63.983593,66.09724,73.583595,71.48965,65.713234,61.630363,64.114876,73.31119,79.20575,82.95714,87.289444,96.51201,93.22339,86.40657,77.006775,66.30729,55.958977,47.599594,44.90831,41.606567,36.063183,31.310772,27.966362,26.079182,28.356926,33.391594,35.682465,33.686977,33.447388,35.918774,39.17457,38.409847,35.636517,34.85867,35.570873,36.299488,34.596104,30.493542,27.844925,25.40636,23.049849,21.746874,21.461334,21.999592,21.822361,20.434053,18.376207,16.000002,14.27036,13.200411,12.481642,11.474052,10.758565,9.682052,8.63836,7.8441033,7.3616414,6.921847,6.3212314,5.8453336,5.622154,5.648411,4.7589746,4.2863593,3.7874875,3.1671798,2.6945643,2.0808206,1.5589745,1.1191796,0.78769237,0.6268718,0.35446155,0.25271797,0.21989745,0.2297436,0.33805132,0.12471796,0.052512825,0.036102567,0.029538464,0.029538464,0.02297436,0.016410258,0.02297436,0.036102567,0.049230773,0.06235898,0.09189744,0.12143591,0.13784617,0.14769232,0.1148718,0.108307704,0.15753847,0.25928208,0.37415388,0.32164106,0.26256412,0.2100513,0.17723078,0.19692309,0.24943592,0.25271797,0.26256412,0.27897438,0.24615386,0.24287182,0.2231795,0.34789747,0.6104616,0.8533334,1.3456411,3.5216413,4.57518,3.9351797,3.2689233,3.0982566,4.640821,5.2644105,4.06318,1.8510771,1.8313848,1.5622566,1.148718,0.6826667,0.22646156,0.20348719,0.20348719,0.3052308,0.5349744,0.8566154,1.1815386,1.6672822,2.0151796,2.2416413,2.674872,3.2754874,3.0293336,2.4976413,2.15959,2.3926156,2.3368206,2.5993848,2.7602053,2.7536411,2.8947694,2.2350771,1.847795,1.7624617,1.8084104,1.6213335,1.7296412,1.204513,0.65969235,0.380718,0.3249231,0.25928208,0.2855385,0.3117949,0.30194873,0.25928208,0.23958977,0.24615386,0.25928208,0.27897438,0.3117949,0.32820517,0.3708718,0.4266667,0.47261542,0.48574364,0.48574364,0.43323082,0.37743592,0.33805132,0.318359,0.26584616,0.2100513,0.17394873,0.17066668,0.18707694,0.2100513,0.23630771,0.27241027,0.31507695,0.34133336,0.318359,0.27897438,0.23302566,0.18707694,0.13784617,0.12143591,0.15425642,0.19692309,0.2231795,0.21989745,0.28225642,0.36102566,0.44964105,0.50543594,0.446359,0.4004103,0.37743592,0.36430773,0.3511795,0.32820517,0.2231795,0.13456412,0.07876924,0.049230773,0.02297436,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016410258,0.08533334,0.016410258,0.01969231,0.08861539,0.15425642,0.101743594,0.01969231,0.0,0.0,0.0,0.0,0.0,0.0,0.1148718,0.27241027,0.21989745,0.28882053,0.12143591,0.026256412,0.08205129,0.14769232,0.108307704,0.128,0.27241027,0.36758977,0.0,0.0,0.006564103,0.04594872,0.11158975,0.17066668,0.4004103,1.1191796,2.0545642,2.9669745,3.6726158,3.95159,5.2676926,7.141744,8.812308,9.235693,10.026668,11.116308,12.22236,13.177437,13.932309,15.852309,16.000002,15.051488,13.98154,14.063591,12.386462,13.6008215,15.514257,16.567797,15.842463,15.497848,17.329231,19.43631,20.873848,21.651693,21.871592,21.93395,20.41436,16.761436,11.300103,8.490667,7.525744,7.3058467,6.8004107,5.041231,3.5282054,3.3805132,3.318154,2.6912823,1.4900514,1.0535386,0.86646163,0.5021539,0.055794876,0.14769232,0.33805132,0.574359,1.6311796,2.9472823,2.612513,2.3630772,1.1913847,0.5907693,0.77456415,0.69251287,0.827077,1.020718,0.9944616,0.7187693,0.38728207,0.5218462,0.5677949,0.53825647,0.5316923,0.73517954,0.7220513,0.5874872,0.47261542,0.4397949,0.508718,0.2986667,0.54482055,1.0568206,1.6278975,2.0217438,2.540308,2.5304618,2.3269746,2.2580514,2.6387694,2.356513,1.8051283,1.0994873,0.79425645,1.910154,2.228513,1.719795,1.467077,1.7394873,2.0151796,1.6902566,2.3860514,3.2262566,3.3772311,2.034872,2.2055387,2.2055387,2.5173335,2.7273848,1.5491283,1.3259488,1.1618463,1.0896411,1.1355898,1.3029745,1.4408206,1.0994873,0.9288206,1.3193847,2.3827693,2.3368206,2.4057438,2.4549747,2.3433847,1.9331284,1.6246156,2.3040001,3.1376412,3.3411283,2.2022567,1.9593848,2.5206156,3.1343591,3.2196925,2.3762052,2.737231,3.629949,4.6080003,5.7074876,7.4240007,7.509334,8.208411,10.640411,13.161027,11.35918,11.83836,12.018872,13.177437,14.378668,12.475078,9.593436,8.546462,9.547488,11.733335,13.177437,12.527591,11.631591,10.535385,9.199591,7.4896417,6.5772314,6.5345645,7.3714876,8.490667,8.664616,9.032206,9.399796,9.924924,10.883283,12.665437,9.475283,6.245744,4.670359,5.405539,8.067283,7.2861543,5.940513,5.861744,7.4436927,9.649232,9.301334,9.26195,9.032206,8.316719,7.030154,10.394258,10.850462,9.235693,6.7774363,5.110154,4.391385,4.896821,5.1659493,5.9995904,10.443488,10.676514,7.496206,4.886975,4.1780515,4.027077,6.193231,6.9349747,5.5007186,3.2820516,3.817026,3.56759,2.2121027,3.2328207,6.124308,6.380308,3.4822567,2.0742567,2.1234872,2.9111798,3.0227695,4.3618464,5.5565133,6.0685134,5.940513,5.8092313,4.6834874,3.0293336,2.6453335,3.6168208,4.309334,4.903385,7.1187696,9.225847,9.787078,7.6734366,4.8705645,4.4373336,5.687795,7.5388722,8.51036,8.651488,7.5487185,5.6943593,4.2601027,5.1167183,5.98318,5.4843082,4.1714873,3.5314875,6.0061545,6.7282057,6.5345645,9.3078985,13.489232,12.107488,5.366154,4.1091285,4.781949,4.7622566,2.3696413,2.1398976,2.9965131,4.522667,5.8125134,5.4613338,2.8882053,3.3805132,5.4416413,6.521436,3.0227695,1.3193847,1.723077,2.7076926,3.0391798,1.7723079,2.1792822,2.5271797,2.5435898,2.1497438,1.463795,1.7526156,2.2186668,2.294154,1.8412309,1.1684103,5.333334,3.570872,2.1267693,3.876103,8.339693,11.32636,11.306667,10.994873,10.35159,6.6034875,5.684513,7.3386674,9.5146675,10.203898,7.427283,7.8670774,10.489437,13.751796,19.6759,33.847797,33.7198,25.298054,18.343386,16.75159,18.566566,15.694771,14.690463,14.614976,15.202463,16.853334,18.875078,18.560001,16.042667,12.760616,11.428103,10.118565,9.846154,8.874667,6.8660517,4.886975,4.9854364,5.2644105,4.650667,3.3017437,2.5764105,2.5206156,2.2022567,1.9429746,1.8379488,1.7493335,1.3784616,1.5031796,1.6902566,1.7099489,1.5622566,1.6147693,1.6016412,1.4375386,1.1684103,0.95835906,1.211077,2.0578463,2.9604106,3.242667,2.0939488,2.162872,2.4582565,2.6945643,2.8389745,3.131077,4.578462,6.114462,6.5280004,5.218462,2.2219489,3.4034874,3.006359,2.487795,2.4943593,2.8717952,5.1954875,7.768616,9.281642,8.920616,6.38359,8.933744,12.33395,14.956308,15.688207,13.948719,16.964924,17.910154,18.983387,21.17908,24.297028,23.558565,22.514874,24.864822,27.559387,20.834463,20.913233,27.986053,33.040413,33.91672,35.285336,41.846157,43.47077,45.364517,48.794262,51.108105,46.263798,45.22339,38.787285,27.16554,19.977848,21.96349,23.40431,25.055182,25.554052,21.425232,20.676924,22.439386,23.785027,24.041027,24.82872,27.03754,30.995695,33.680412,33.276722,29.184002,25.823181,23.066257,19.236105,14.27036,9.701744,10.837335,11.995898,16.328207,24.18872,33.16185,33.079796,34.582977,36.74913,38.98749,41.032207,44.465233,44.97067,45.43344,46.848003,48.32821,49.765747,48.833645,47.29108,46.644516,48.12472,48.34462,52.68021,59.21149,64.13785,61.774773,61.531902,63.520824,68.5358,75.50359,81.48349,83.055595,81.31283,78.34914,77.96513,85.671394,97.739494,91.18195,76.96411,65.414566,66.241646,73.34729,82.747086,92.353645,101.014984,108.53088,106.15796,99.00308,87.34196,74.66339,67.64636,63.59303,57.93149,50.18585,41.767387,35.981133,32.512,30.181746,33.017437,40.034466,45.229954,40.579285,38.73477,40.500515,43.224617,40.76636,37.697643,37.362873,39.062977,40.82872,39.407593,36.299488,31.74072,28.399591,27.139284,27.001438,28.376617,30.53949,31.990156,31.071182,25.98072,20.263386,16.548103,14.864411,14.401642,13.5089245,12.793437,11.766154,10.729027,9.842873,9.133949,8.36595,7.643898,7.0400004,6.619898,6.419693,5.940513,5.7107697,5.3103595,4.7392826,4.4438977,3.6660516,2.8291285,2.156308,1.6771283,1.2471796,0.93866676,0.6465641,0.48574364,0.4004103,0.15097436,0.10502565,0.06235898,0.03938462,0.029538464,0.029538464,0.029538464,0.01969231,0.029538464,0.059076928,0.07876924,0.07548718,0.08205129,0.108307704,0.14769232,0.18051283,0.12471796,0.101743594,0.101743594,0.13128206,0.19692309,0.28225642,0.3117949,0.26584616,0.18379489,0.16410258,0.19364104,0.20676924,0.2100513,0.2100513,0.2231795,0.190359,0.15425642,0.23302566,0.45620516,0.761436,1.1848207,2.993231,3.8531284,3.2918978,2.7175386,3.8859491,5.290667,5.2709746,3.5314875,1.1355898,0.69251287,0.5152821,0.41025645,0.26912823,0.0951795,0.09189744,0.11158975,0.15097436,0.27897438,0.6301539,0.67610264,1.0896411,1.4539489,1.6804104,2.0217438,2.5961027,2.487795,2.3433847,2.5271797,3.1015387,2.6912823,2.5600002,2.5731285,2.612513,2.553436,2.2449234,1.8773335,1.7329233,1.7362052,1.4539489,1.5195899,1.2373334,0.8172308,0.44307697,0.27241027,0.24615386,0.28882053,0.32164106,0.3052308,0.256,0.22646156,0.26912823,0.3117949,0.3511795,0.42994875,0.42338464,0.42994875,0.42994875,0.4201026,0.4201026,0.446359,0.42338464,0.37415388,0.33805132,0.34133336,0.2986667,0.23958977,0.19692309,0.18707694,0.17066668,0.190359,0.2297436,0.29538465,0.36102566,0.36430773,0.36430773,0.3511795,0.3052308,0.24287182,0.18707694,0.12471796,0.10502565,0.12471796,0.15753847,0.17066668,0.190359,0.2855385,0.4266667,0.5349744,0.49887183,0.41025645,0.38728207,0.39056414,0.39056414,0.3708718,0.3249231,0.24287182,0.16082053,0.098461546,0.03938462,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.026256412,0.23958977,0.4660513,0.19692309,0.03938462,0.0,0.0,0.0,0.0,0.0,0.0,0.055794876,0.14769232,0.18379489,0.036102567,0.0,0.13456412,0.4135385,0.7318975,0.29210258,0.30194873,0.4660513,0.47589746,0.0,0.0,0.036102567,0.108307704,0.26912823,0.6104616,0.83035904,0.6104616,0.80738467,1.8773335,3.892513,4.7589746,5.0576415,5.540103,6.377026,7.171283,8.198565,8.342975,8.818872,10.049642,11.674257,14.982565,15.432206,14.890668,13.929027,11.841642,11.949949,15.61272,18.025026,17.769028,16.83036,15.842463,18.038155,20.394669,20.883694,18.477951,13.90277,12.547283,12.107488,11.057232,8.651488,6.9054365,5.8190775,5.7468724,6.738052,8.54318,5.2742567,4.585026,4.955898,4.8836927,2.868513,1.3784616,0.9419488,0.6071795,0.20676924,0.36758977,0.4397949,0.88943595,1.273436,1.5031796,1.8313848,0.97805136,0.8172308,1.0305642,1.1684103,0.65641034,1.1323078,0.9124103,0.49887183,0.31507695,0.7187693,0.8041026,0.8041026,0.65969235,0.44307697,0.380718,0.45620516,0.380718,0.35774362,0.38728207,0.28882053,0.26584616,0.23958977,0.23958977,0.4004103,0.9616411,1.6443079,1.6246156,1.5885129,1.7001027,1.6016412,1.5031796,1.4998976,1.401436,1.2406155,1.2504616,0.9353847,0.8172308,1.1060513,1.5753847,1.5885129,1.4276924,1.6902566,1.8937438,1.975795,2.3040001,2.7569232,2.5206156,2.2153847,2.0151796,1.6475899,1.7460514,2.2186668,2.5238976,2.3040001,1.3883078,1.401436,1.276718,1.2570257,1.394872,1.5425643,1.9922053,2.2153847,2.284308,2.176,1.785436,0.97805136,1.785436,2.425436,2.3630772,2.28759,1.9462565,2.228513,2.8258464,3.1343591,2.2416413,2.878359,4.325744,5.8092313,6.889026,7.460103,8.425026,8.530052,9.993847,12.041847,10.896411,11.286975,9.964309,9.26195,10.118565,12.084514,8.605539,7.837539,8.513641,9.563898,10.102155,10.761847,10.148104,8.89436,7.781744,7.719385,7.9524107,8.523488,9.005949,8.822155,7.24677,8.651488,10.200616,9.993847,9.344001,12.786873,13.824001,11.017847,7.709539,6.226052,7.8736415,10.266257,8.950154,6.99077,6.62318,9.245539,11.076924,10.33518,9.012513,8.116513,7.6898465,12.304411,13.328411,11.0605135,7.4043083,5.8912826,4.6933336,4.630975,5.622154,7.5881033,10.466462,11.1983595,9.140513,6.8397956,5.481026,4.8836927,5.3103595,7.0367184,6.183385,3.062154,2.1825643,1.6213335,1.782154,4.4242053,7.712821,6.2096415,3.623385,1.9035898,1.7624617,2.806154,3.5249233,3.1343591,3.751385,3.5446157,2.425436,2.0611284,0.98461545,1.6147693,3.3280003,5.543385,7.6898465,6.5050263,6.1538467,5.405539,4.279795,4.059898,5.717334,5.904411,5.3694363,5.6418467,9.048616,10.134975,7.1483083,4.4865646,4.384821,6.9120007,7.522462,7.0793853,4.827898,2.2449234,3.0523078,3.0523078,3.7842054,6.7249236,10.006975,8.408616,4.342154,2.356513,1.9035898,2.3729234,3.0654361,6.117744,6.7150774,4.923077,2.156308,1.1913847,1.5556924,3.0752823,4.535795,4.5456414,1.5556924,0.8598975,1.8215386,2.546872,2.553436,2.7602053,6.449231,7.762052,6.994052,5.1626673,4.027077,5.9569235,7.785026,7.3747697,4.647385,1.5721027,2.0841026,2.3302567,3.0096412,3.9811285,4.2896414,4.3749747,7.7456417,10.374565,10.41395,8.178872,4.273231,2.8488207,2.4746668,2.5337439,3.2032824,4.9132314,8.818872,17.509745,31.090874,47.17949,35.741543,22.94154,17.214361,18.372925,17.578669,13.952001,12.937847,14.12595,15.143386,11.628308,14.470565,16.636719,16.853334,15.018668,12.22236,10.696206,9.7214365,8.572719,7.1187696,5.8125134,5.973334,5.8847184,5.681231,5.041231,3.1737437,2.5632823,2.3105643,2.481231,2.7733335,2.5173335,1.8838975,1.7985642,1.9364104,1.9790771,1.5885129,1.8051283,2.0545642,1.9922053,1.6410258,1.3718976,1.4211283,2.5337439,3.5774362,3.5577438,1.6180514,2.6420515,6.314667,8.418462,7.7948723,6.3179493,8.283898,15.126975,17.64759,13.013334,4.7589746,2.172718,2.934154,4.069744,5.179077,8.438154,5.9470773,3.56759,2.9702566,4.4307694,6.8365135,9.278359,12.800001,16.748308,20.187899,21.894566,25.642668,24.024618,23.722668,26.532104,29.38749,32.377438,33.017437,35.574158,39.266464,38.25231,32.699078,37.930668,45.364517,51.485542,57.842876,60.56698,59.342773,60.13703,64.9518,71.83755,66.30729,65.739494,59.342773,45.492516,31.721027,25.826464,25.376822,27.526566,28.65231,24.369232,27.06708,32.482464,35.84985,35.84985,34.605953,31.445335,30.654362,32.164104,34.50749,34.835693,30.831593,27.779284,25.721437,23.62749,19.393642,21.26113,22.816822,25.764105,29.85354,32.882874,35.05559,42.371284,50.326977,57.803493,67.10483,70.452515,71.469955,69.822365,66.208824,62.37539,63.86544,67.77108,66.82585,58.742157,46.21785,50.015182,62.398365,75.7957,85.152824,87.936005,78.75611,77.1479,80.54154,85.57293,88.08698,85.001854,82.707695,82.29416,86.18339,98.1596,101.06422,94.29334,84.680214,76.00575,68.998566,68.73272,74.561646,88.605545,104.4874,107.34606,101.497444,92.81313,84.0796,76.78688,71.135185,71.34196,67.12124,58.020107,45.525337,33.05026,30.706875,32.354465,37.842052,44.911594,49.207798,43.726772,45.095387,48.078773,49.54585,48.44636,44.721233,46.355698,48.557953,49.647594,51.039185,47.13354,42.505848,40.037746,39.67344,38.390156,38.37703,39.565132,41.373543,41.045338,33.66072,24.149336,18.84554,16.873028,16.52513,15.241847,14.339283,13.682873,13.141335,12.563693,11.795693,10.889847,9.980719,9.117539,8.362667,7.752206,7.4469748,7.2336416,6.87918,6.3474874,5.799385,5.1265645,4.4012313,3.764513,3.2262566,2.6387694,2.2613335,1.6082052,1.0272821,0.65312827,0.39712822,0.24943592,0.14112821,0.06564103,0.029538464,0.029538464,0.01969231,0.016410258,0.02297436,0.04266667,0.09189744,0.07876924,0.07548718,0.108307704,0.15425642,0.16738462,0.14441027,0.118153855,0.101743594,0.08861539,0.07548718,0.16082053,0.29210258,0.3052308,0.20020515,0.15097436,0.20020515,0.23958977,0.2297436,0.18707694,0.19692309,0.23630771,0.20676924,0.2855385,0.54482055,0.94523084,1.7394873,2.8356924,3.511795,3.6463592,3.7087183,3.7809234,3.387077,2.540308,1.463795,0.6104616,0.48902568,0.32164106,0.18051283,0.0951795,0.04594872,0.032820515,0.0951795,0.15097436,0.16410258,0.15425642,0.2855385,0.5415385,0.67610264,0.75487185,1.1454359,1.4145643,1.6902566,2.228513,2.8455386,2.930872,2.6978464,2.6683078,2.6912823,2.7503593,2.9440002,2.5173335,2.1366155,1.9790771,2.0020514,1.9528207,1.8445129,1.5688206,1.0075898,0.3708718,0.19692309,0.2100513,0.21333335,0.24943592,0.32820517,0.4266667,0.32820517,0.44307697,0.5874872,0.7122052,0.86974365,0.88287187,0.81066674,0.6662565,0.50543594,0.45620516,0.446359,0.4594872,0.42338464,0.35446155,0.36758977,0.3052308,0.25271797,0.2231795,0.20676924,0.18379489,0.18379489,0.20020515,0.23958977,0.30194873,0.4135385,0.5218462,0.4660513,0.3708718,0.28225642,0.19692309,0.13784617,0.10502565,0.098461546,0.108307704,0.12143591,0.12143591,0.21333335,0.37743592,0.54482055,0.5940513,0.44964105,0.36758977,0.33476925,0.3446154,0.380718,0.40697438,0.34789747,0.26256412,0.17394873,0.07548718,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.055794876,0.09189744,0.03938462,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.029538464,0.036102567,0.006564103,0.0,0.13784617,0.46276927,0.9156924,0.7975385,0.35446155,0.17066668,0.27241027,0.108307704,0.15753847,0.07548718,0.02297436,0.09189744,0.318359,0.3117949,0.256,0.38728207,0.86974365,1.7788719,2.8816411,3.508513,3.95159,4.4110775,4.9985647,6.3376417,7.0367184,8.208411,9.888822,11.063796,11.54954,13.036308,14.700309,15.494565,14.158771,14.230975,17.926565,21.67467,23.213951,21.589334,18.58954,18.057848,18.901335,19.045746,15.451899,11.175385,10.476309,10.377847,9.32759,7.1876926,5.9995904,4.8607183,4.9394875,6.012718,6.482052,4.9099493,4.7458467,5.874872,6.665847,3.9778464,1.7690258,1.0272821,0.86646163,0.84348726,0.9517949,0.6826667,1.0765129,1.2832822,1.4473847,2.6847181,0.9911796,0.9517949,1.0929232,0.8566154,0.6071795,0.8795898,1.2438976,1.1257436,0.60061544,0.38728207,0.39384618,0.5316923,0.5677949,0.45292312,0.3314872,0.40697438,0.29538465,0.21661541,0.23630771,0.26584616,0.5546667,0.61374366,0.5218462,0.4660513,0.75487185,1.1257436,1.2603078,1.3161026,1.3620514,1.3686155,1.204513,1.3718976,1.5556924,1.6147693,1.5688206,0.636718,0.5940513,1.0010257,1.4539489,1.5753847,1.5524104,1.4834872,1.5130258,1.7460514,2.231795,2.4976413,2.3105643,2.2744617,2.356513,1.8904617,1.8248206,1.9626669,2.0512822,2.0841026,2.2908719,1.404718,1.1946667,1.2603078,1.3062565,1.1520001,1.3095386,1.4736412,1.910154,2.4188719,2.3236926,1.5163078,1.5688206,1.9790771,2.5928206,3.5938463,3.4198978,3.0162053,2.793026,3.0162053,3.8038976,5.093744,5.805949,6.5050263,7.709539,9.90195,11.247591,10.420513,10.217027,11.313231,12.274873,11.113027,8.946873,8.323282,9.275078,9.32759,8.667898,9.622975,10.512411,10.6469755,10.331899,9.527796,8.805744,7.702975,6.5969234,6.6822567,6.6822567,6.9743595,8.172308,9.714872,9.849437,11.211488,12.041847,10.873437,8.530052,8.136206,10.696206,11.096616,9.235693,6.554257,6.055385,7.568411,9.130668,8.992821,7.5388722,7.2927184,9.750975,11.296822,11.835078,11.523283,10.755282,11.900719,12.199386,10.807796,8.172308,6.0225644,5.356308,4.3552823,4.634257,6.245744,7.722667,7.515898,7.53559,7.499488,6.8955903,4.9788723,6.1308722,5.920821,4.670359,3.242667,3.0490258,2.6223593,2.2350771,2.7076926,3.7874875,4.1222568,3.6627696,2.294154,1.5524104,3.0687182,8.553026,8.700719,4.962462,2.5796926,2.5665643,1.6935385,1.6049232,3.2853336,4.8049235,5.2742567,4.8344617,4.7622566,5.182359,4.4012313,3.0030773,3.8400004,5.146257,4.4996924,4.1517954,4.644103,4.788513,4.194462,3.6069746,3.8859491,5.481026,8.438154,9.829744,7.634052,5.0904617,4.266667,6.0652313,6.4656415,5.504,4.9132314,5.172513,5.5269747,5.6320004,5.0477953,4.4438977,4.6112823,6.4590774,7.9983597,6.9743595,4.3060517,1.6311796,1.2996924,1.6968206,2.605949,2.8849232,2.4024618,2.0578463,4.6112823,5.720616,4.5423594,3.045744,5.9963083,9.780514,8.36595,5.737026,3.8334363,2.550154,3.9023592,5.6254363,5.3234878,3.0720003,1.401436,1.5622566,4.5489235,7.4043083,7.8736415,4.4110775,2.3466668,2.861949,3.9187696,4.2436924,3.308308,1.6869745,1.273436,1.9954873,3.383795,4.571898,4.8147697,10.627283,20.768822,31.72431,37.694363,26.725746,23.663591,24.598976,25.091284,20.164925,13.610668,11.385437,10.916103,10.886565,11.247591,11.690667,13.932309,15.212309,14.427898,12.114052,10.450052,10.325335,9.357129,7.7259493,8.155898,8.3364105,7.5618467,6.550975,5.4186673,3.6857438,2.7634873,2.3729234,2.2908719,2.356513,2.481231,2.2646155,2.2121027,2.2711797,2.1989746,1.5753847,1.9593848,2.2482052,2.0217438,1.5360001,1.7165129,2.1825643,2.930872,3.2032824,2.6715899,1.4342566,8.914052,24.09354,31.648823,25.961027,11.113027,8.234667,16.718771,19.777643,13.387488,6.298257,4.923077,5.3858466,5.4908724,5.408821,7.680001,7.3485136,5.3103595,4.9920006,6.5805135,7.0432825,6.2523084,8.966565,12.586668,16.009848,19.61354,23.975386,22.89231,20.522669,19.5479,21.172514,22.806976,26.692924,39.955696,57.14708,60.274876,55.794876,59.05067,65.83795,70.10462,63.973747,58.47303,62.68062,71.771904,82.45498,92.94442,81.10606,73.101135,65.250465,53.782978,34.848824,26.41395,27.776003,30.57231,31.094156,30.276926,35.521645,42.112003,45.203697,45.088825,47.202465,45.525337,42.37457,41.24554,43.057236,46.13908,45.91262,43.155697,41.73785,42.824207,44.855797,41.928207,38.485336,38.547695,41.826466,43.71036,38.84308,43.090054,53.185646,66.80288,82.55016,83.11139,79.83919,79.24513,81.273445,79.294365,84.97559,90.69621,90.32206,82.20226,69.179085,71.01375,79.99673,94.89396,110.680626,118.56083,106.19734,100.60801,100.365135,99.99426,89.98073,77.64349,69.76,65.913445,67.524925,77.84698,80.87959,78.08001,74.10216,71.6997,71.72267,67.049034,65.67713,70.94154,79.66852,82.16288,78.51324,72.98626,71.466675,74.48616,77.2037,75.36903,70.974365,62.877544,52.594875,44.28144,42.17108,45.686157,49.72308,51.085133,48.475903,47.028515,52.37826,56.451286,57.89867,62.093132,60.419285,58.919388,58.55508,58.74544,57.363697,54.47221,49.430977,48.180515,51.69231,55.955696,57.711594,63.149952,66.78647,64.42339,53.14298,34.63877,25.494976,21.448206,19.570873,18.258053,17.27672,16.938667,16.689232,16.15754,15.163078,14.437745,13.699283,12.832822,11.85477,10.912822,10.029949,9.468719,8.950154,8.402052,7.972103,7.6996927,7.02359,6.4754877,5.9963083,4.923077,4.1813335,3.4034874,2.609231,1.8576412,1.2504616,0.83035904,0.5218462,0.3052308,0.17066668,0.09189744,0.049230773,0.026256412,0.02297436,0.03938462,0.06564103,0.07548718,0.068923086,0.098461546,0.15097436,0.14441027,0.108307704,0.08205129,0.068923086,0.06564103,0.052512825,0.068923086,0.118153855,0.16738462,0.19364104,0.16410258,0.14441027,0.13128206,0.12471796,0.17066668,0.35774362,0.29538465,0.2297436,0.380718,0.764718,1.1782565,1.7165129,2.228513,2.540308,2.7109745,3.0358977,3.442872,2.858667,1.9889232,1.2406155,0.7581539,0.44964105,0.22646156,0.108307704,0.06235898,0.032820515,0.02297436,0.059076928,0.09189744,0.10502565,0.14112821,0.19692309,0.35774362,0.47261542,0.5284103,0.65641034,0.9944616,1.3751796,1.8051283,2.3302567,3.0391798,3.1409233,3.259077,3.3214362,3.190154,2.665026,2.353231,2.0020514,1.7263591,1.591795,1.6114873,2.0578463,1.7985642,1.3259488,0.90584624,0.5874872,0.36758977,0.25928208,0.24287182,0.27569234,0.3052308,0.29538465,0.32164106,0.32164106,0.318359,0.41682056,0.51856416,0.58092314,0.6629744,0.7515898,0.7515898,0.5513847,0.45620516,0.380718,0.31507695,0.318359,0.27569234,0.23630771,0.2100513,0.20020515,0.19692309,0.21333335,0.21661541,0.21989745,0.23958977,0.28882053,0.4004103,0.41025645,0.37743592,0.32164106,0.24615386,0.17723078,0.13456412,0.108307704,0.0951795,0.098461546,0.108307704,0.15753847,0.26256412,0.40369233,0.508718,0.48902568,0.49887183,0.47261542,0.41682056,0.39384618,0.38728207,0.37415388,0.36102566,0.33476925,0.24615386,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08205129,0.27241027,0.5481026,0.571077,0.2297436,0.03938462,0.13456412,0.27569234,0.256,0.15425642,0.10502565,0.21661541,0.56451285,0.51856416,0.3314872,0.2855385,0.58092314,1.3259488,2.5731285,3.0851285,3.3312824,3.5971284,3.9876926,4.6867695,5.910975,7.4797955,8.973129,9.757539,10.371283,13.961847,17.831387,19.856411,18.464823,19.22954,21.622156,24.175592,25.475285,24.17231,22.938257,20.683489,19.39036,18.563284,15.225437,10.95877,9.472001,9.156924,8.664616,6.9021544,5.671385,4.634257,4.663795,5.4613338,5.536821,4.3749747,4.4340515,5.3858466,6.048821,4.384821,2.1530259,1.211077,0.8763078,0.80738467,1.017436,1.3357949,1.1191796,0.955077,1.4441026,3.2098465,1.1881026,1.0732309,1.2406155,1.0502565,0.85005134,1.079795,1.7362052,1.7985642,1.1060513,0.3511795,0.4201026,0.47261542,0.4594872,0.4004103,0.38400003,0.37743592,0.3249231,0.35774362,0.46276927,0.47917953,0.56123084,0.48246157,0.380718,0.3708718,0.54482055,0.71548724,0.9878975,1.2209232,1.3686155,1.4867693,1.1355898,1.7362052,1.9068719,1.4145643,1.2077949,0.72861546,0.6859488,0.8992821,1.2373334,1.6278975,1.3751796,1.276718,1.2373334,1.2635899,1.4802053,1.5524104,1.6246156,1.7132308,1.7427694,1.5425643,1.394872,1.4145643,1.4145643,1.394872,1.5458462,1.2635899,0.96492314,0.81066674,0.84348726,0.9714873,1.0404103,1.1257436,1.6246156,2.4057438,2.806154,1.8018463,1.3718976,1.6246156,2.5764105,4.1583595,4.6900516,4.0533338,3.3017437,3.1967182,4.2240005,6.678975,8.129642,9.412924,11.21477,14.063591,14.670771,11.716924,9.665642,10.095591,11.703795,9.964309,7.50277,6.7872825,8.185436,9.964309,10.8537445,12.2157955,12.419283,11.132719,9.31118,8.103385,8.418462,8.887795,8.930462,8.766359,8.891078,7.7423596,7.7259493,9.485129,11.907283,14.089848,14.283488,12.324103,9.42277,8.152616,9.110975,10.371283,10.262975,8.470975,6.058667,5.937231,7.955693,9.573745,9.5835905,8.1066675,8.87795,11.053949,12.875488,13.24636,11.739899,11.559385,10.880001,9.714872,8.109949,6.1407185,5.6254363,4.568616,4.588308,5.435077,4.9821544,4.916513,5.671385,6.6133337,6.7872825,4.923077,5.211898,4.568616,3.8400004,3.3312824,2.7700515,2.9078977,2.7798977,2.3762052,2.1333334,2.934154,4.0467696,2.8389745,1.847795,2.8717952,6.9645133,5.9995904,3.4100516,2.8192823,4.096,3.3608208,2.553436,3.8367183,4.493129,3.6529233,2.281026,4.8738465,5.297231,4.1583595,3.0162053,4.3716927,5.159385,4.450462,4.4964104,5.3103595,4.6834874,5.9930263,8.772923,9.997129,9.173334,8.333129,7.827693,6.163693,4.9788723,5.211898,7.0957956,7.3452315,5.3891287,3.6594875,3.3312824,4.322462,5.2709746,4.6834874,3.8400004,3.6332312,4.59159,5.0674877,3.9942567,2.6683078,2.03159,2.681436,2.7273848,2.412308,1.9396925,1.8806155,3.1803079,5.861744,6.744616,6.0619493,4.6769233,4.096,5.100308,4.240411,3.2918978,2.7076926,1.6246156,2.1891284,2.7766156,2.4615386,1.4342566,1.0010257,1.6311796,5.395693,7.5520005,6.294975,2.7831798,2.0578463,2.793026,3.2754874,2.8816411,2.0808206,1.4998976,1.5392822,3.9023592,7.0137444,6.012718,4.096,7.515898,15.136822,23.650463,27.598772,25.583591,30.641233,34.067696,30.802053,19.403488,12.86236,11.592206,10.998155,9.911796,10.604308,10.571488,12.2157955,13.338258,13.013334,11.59877,11.21477,10.752001,9.281642,7.430565,7.397744,7.574975,6.9677954,6.36718,5.730462,4.2174363,3.3247182,3.0227695,2.737231,2.3696413,2.297436,2.0578463,1.9790771,2.028308,2.0676925,1.847795,2.5895386,2.4057438,1.7558975,1.3456411,2.1300514,3.2689233,3.2853336,2.858667,2.3926156,2.0118976,7.972103,25.009233,33.48021,26.863592,11.772718,7.017026,10.098872,11.067078,7.752206,5.7501545,7.026872,9.130668,10.184206,9.888822,9.544206,8.628513,7.181129,8.52677,11.575796,10.804514,11.730052,14.762668,17.473642,18.95713,19.849848,23.93272,23.122053,23.46667,26.466463,29.088823,29.108515,31.927797,39.253338,47.619286,48.40698,52.08944,60.452106,64.07877,59.339493,48.387287,50.783184,63.62585,80.79755,99.16719,118.60021,109.81088,96.256004,80.71549,65.21108,50.989952,44.580105,45.630363,49.759182,54.603493,59.8318,68.61457,74.4238,76.0878,75.89744,79.612724,80.99447,80.51529,79.73088,78.67406,75.861336,72.37908,70.01601,68.92308,68.82462,69.021545,67.32472,62.194878,58.975185,59.12616,60.242058,56.12308,62.621544,74.34831,86.25231,93.60739,89.17334,85.02811,86.93498,94.024216,98.78647,107.79898,110.26052,106.11857,96.265854,82.556725,81.02729,84.88042,92.00575,98.98011,101.08391,96.74175,92.48165,91.74975,91.375595,81.581955,67.387085,62.414776,60.429134,59.506878,62.020927,63.02852,60.563698,61.65334,69.06749,81.33908,77.505646,70.32452,64.55467,62.48698,63.937645,66.98995,68.31918,70.5477,73.87241,76.08452,74.18749,74.33518,73.06175,68.87385,62.257236,57.012516,57.4359,57.964314,56.155903,52.68677,54.53457,57.97416,59.68411,60.98052,67.79406,64.42339,61.95857,63.09416,65.581955,62.23098,58.043083,55.893337,58.31549,64.42339,69.90442,72.49724,73.28493,70.59364,63.002262,49.362057,34.182568,27.303387,24.103386,22.166977,21.274258,20.762259,20.394669,19.951591,19.265642,18.22195,17.575386,16.95836,16.239592,15.396104,14.496821,13.83713,13.51877,13.013334,12.133744,11.040821,10.341744,9.5835905,8.933744,8.28718,7.250052,6.419693,5.5663595,4.637539,3.6627696,2.7470772,1.9954873,1.3883078,0.92225647,0.58420515,0.35446155,0.2231795,0.13456412,0.09189744,0.08205129,0.068923086,0.08205129,0.072205134,0.09189744,0.13456412,0.13784617,0.09189744,0.06564103,0.052512825,0.049230773,0.04594872,0.03938462,0.052512825,0.098461546,0.15753847,0.17723078,0.13456412,0.108307704,0.098461546,0.14441027,0.3249231,0.40697438,0.35446155,0.41025645,0.85005134,2.0053334,2.3433847,2.228513,1.9035898,1.6672822,1.8904617,2.487795,2.8750772,2.9702566,2.6354873,1.6804104,0.764718,0.28225642,0.08533334,0.03938462,0.029538464,0.01969231,0.036102567,0.059076928,0.08205129,0.101743594,0.12143591,0.26256412,0.42338464,0.5677949,0.7089231,0.86317956,1.0633847,1.3653334,1.8281027,2.5173335,2.9997952,3.117949,3.1507695,3.1277952,2.8225644,2.425436,2.1169233,1.8182565,1.5163078,1.2603078,1.5327181,1.7296412,1.782154,1.6311796,1.2274873,0.74830776,0.45620516,0.3446154,0.36102566,0.39384618,0.28225642,0.28225642,0.2986667,0.29210258,0.26912823,0.318359,0.4004103,0.56123084,0.7253334,0.6859488,0.5677949,0.4955898,0.4135385,0.3249231,0.2855385,0.24943592,0.2297436,0.21333335,0.19364104,0.18051283,0.19692309,0.20348719,0.20020515,0.20020515,0.2231795,0.29538465,0.3511795,0.4004103,0.41682056,0.3511795,0.23958977,0.17066668,0.12471796,0.101743594,0.101743594,0.09189744,0.118153855,0.20348719,0.3314872,0.4594872,0.4955898,0.574359,0.58420515,0.5021539,0.40697438,0.4004103,0.39384618,0.39384618,0.38400003,0.33476925,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.026256412,0.098461546,0.23302566,0.21333335,0.08533334,0.009846155,0.128,0.5481026,0.6235898,0.37415388,0.3511795,0.61374366,0.72861546,0.49887183,0.26256412,0.2297436,0.53825647,1.270154,2.4746668,3.2032824,3.9253337,4.4340515,3.8531284,3.8629746,5.149539,6.6428723,7.834257,8.743385,12.389745,19.19672,24.264208,25.091284,21.586054,22.065233,22.09149,22.672413,23.952412,25.216002,26.22031,23.177849,19.945026,17.732924,15.126975,11.093334,8.687591,8.3134365,8.710565,6.9645133,5.5893335,4.709744,4.4832826,4.667077,4.6145644,4.9132314,4.7458467,4.8607183,5.169231,4.7589746,2.809436,1.5491283,0.9419488,0.9321026,1.4605129,1.4506668,0.92553854,0.7581539,1.2471796,2.1431797,1.0633847,1.7788719,2.2678976,1.8248206,1.0699488,1.7723079,2.0545642,1.8346668,1.2406155,0.62030774,0.5218462,0.40369233,0.318359,0.33805132,0.5316923,0.33476925,0.29210258,0.45620516,0.69251287,0.67282057,0.57764107,0.56123084,0.5907693,0.6301539,0.6268718,0.57764107,0.827077,1.1979488,1.4408206,1.2176411,1.1651284,1.6804104,1.6771283,1.1388719,1.1224617,1.1027694,0.97805136,0.90256417,0.97805136,1.2603078,1.1848207,1.3587693,1.3029745,0.9944616,0.86317956,1.024,1.1552821,1.2242053,1.2438976,1.2898463,1.0404103,0.93866676,0.9321026,0.90912825,0.7056411,1.3587693,1.3915899,1.2307693,1.1815386,1.4342566,1.6705642,1.6114873,1.9659488,2.6617439,2.8521028,1.9922053,1.5753847,1.6738462,2.5304618,4.568616,5.933949,5.723898,4.84759,4.2272825,4.778667,7.3714876,9.531077,11.657847,13.74195,15.38954,14.119386,10.912822,9.938052,11.913847,14.119386,11.1983595,8.086975,6.770872,7.860513,10.610872,11.254155,12.49477,12.596514,10.9915905,8.2904625,7.141744,8.303591,10.230155,11.579078,11.21477,11.772718,10.801231,10.427077,11.487181,13.545027,15.258258,15.222155,13.643488,11.457642,10.331899,9.225847,9.527796,10.223591,10.059488,7.522462,5.8847184,6.5345645,8.635077,10.436924,9.271795,8.608821,10.112,11.690667,11.96636,10.246565,10.308924,9.567181,8.4283085,7.240206,6.298257,6.560821,5.733744,5.3234878,5.2644105,3.9154875,3.8596926,4.6244106,5.7107697,6.2129235,4.8114877,4.2240005,3.4002054,3.3017437,3.56759,2.5206156,2.989949,3.2065644,2.9440002,2.4320002,2.3663592,3.5380516,2.934154,2.1398976,2.1825643,3.5216413,2.4352822,3.308308,6.7938466,10.236719,7.6734366,5.113436,6.9743595,7.3353853,4.781949,2.3827693,8.041026,7.525744,4.8049235,3.0687182,4.713026,5.3924108,4.827898,4.8836927,5.5991797,5.1922054,8.530052,13.138052,13.873232,10.154668,5.979898,5.1232824,4.57518,4.388103,4.7327185,5.8945646,5.3727183,3.9384618,3.1606157,3.4494362,4.076308,4.312616,3.761231,3.0916924,2.6978464,2.6978464,3.0752823,2.300718,1.8970258,2.3335385,3.0358977,2.7437952,2.2350771,2.3072822,3.1606157,4.394667,5.156103,4.9985647,4.588308,3.817026,1.782154,2.546872,5.9503593,7.000616,4.95918,3.3575387,4.9296412,5.904411,4.6933336,2.048,1.024,4.322462,7.2336416,7.3616414,4.827898,2.294154,3.5216413,4.650667,4.900103,3.9975388,2.172718,1.8642052,2.5862565,5.0904617,7.4469748,5.0477953,2.8422565,4.33559,9.895386,17.398155,22.226053,30.404926,41.284927,44.97067,37.48431,20.768822,13.590976,12.865642,12.941129,11.585642,10.000411,10.167795,11.346052,11.897437,11.526565,11.293539,11.651283,10.509129,9.091283,8.018052,7.328821,7.456821,6.8529234,6.4656415,6.422975,6.0192823,4.6178465,4.2994876,3.9056413,3.2196925,2.9440002,2.4681027,2.172718,1.9922053,1.9954873,2.3893335,3.2229745,2.674872,1.8149745,1.5261539,2.4582565,3.4592824,3.5840003,3.1671798,2.7798977,3.2131286,5.8978467,15.041642,19.649643,16.160822,8.448001,6.009436,6.557539,6.442667,5.543385,7.250052,8.395488,10.010257,11.030975,11.113027,10.633847,9.7673855,9.705027,11.073642,12.987078,13.08554,17.109335,19.96472,21.497438,22.357334,23.985233,28.41272,32.43323,37.24472,41.938053,43.51016,38.820107,36.00739,34.06441,34.405746,40.864822,52.562054,58.095592,55.17785,48.50872,49.775593,59.78913,69.182365,80.02954,93.70914,110.89068,109.64021,100.57519,86.74134,74.1678,71.87036,73.577034,74.11529,75.874466,79.921234,86.009445,92.31426,92.23878,89.81334,89.88226,98.11365,102.39673,104.31673,104.45129,101.92739,94.43775,88.07057,86.186676,84.55878,81.98237,80.259285,85.490875,85.41211,82.62565,79.08103,76.06811,71.473236,75.703804,83.47242,89.288216,87.463394,84.76555,85.809235,90.11529,95.0876,96.01314,103.07611,102.485344,96.99447,88.126366,76.16657,71.79816,70.05539,71.59139,74.63713,74.99488,75.54298,73.50154,72.52677,71.71283,65.581955,56.549747,53.782978,53.792824,53.750156,51.442875,53.622158,52.44718,56.42503,69.40226,90.561646,88.71057,81.05354,70.76759,62.45088,62.116108,70.272,74.87344,76.31754,75.26401,72.62852,71.37806,75.67754,80.51857,82.04144,77.55488,68.516106,65.7756,65.95939,66.720825,66.76678,67.48554,63.27139,59.250877,59.152416,65.2997,63.62257,64.86975,67.76452,69.497444,65.746056,63.28452,65.03057,69.507286,75.36575,81.404724,80.610466,72.113235,61.14134,50.18585,39.0039,30.802053,26.916105,24.999386,24.136208,24.818874,26.515694,27.401848,27.500309,26.922668,25.882257,24.067284,23.3879,22.885746,21.960207,20.391386,19.121233,18.057848,16.810667,15.254975,13.545027,12.458668,11.874462,11.109744,10.069334,9.238976,8.467693,7.6176414,6.7085133,5.720616,4.565334,3.564308,2.6847181,1.9429746,1.3423591,0.8960001,0.6170257,0.41682056,0.28882053,0.21333335,0.15425642,0.14441027,0.11158975,0.11158975,0.14112821,0.13784617,0.08861539,0.06564103,0.055794876,0.049230773,0.03938462,0.032820515,0.032820515,0.055794876,0.098461546,0.14769232,0.17066668,0.16082053,0.128,0.12143591,0.21333335,0.43323082,0.44964105,0.47261542,1.0075898,2.8356924,3.058872,3.045744,2.4681027,1.5688206,1.1618463,2.038154,3.5938463,5.0674877,5.5072823,3.7809234,1.847795,0.6859488,0.15753847,0.03938462,0.01969231,0.009846155,0.01969231,0.036102567,0.052512825,0.052512825,0.059076928,0.20348719,0.37743592,0.5415385,0.7089231,1.0305642,1.3489232,1.5655385,1.7001027,1.8773335,2.1956925,2.3401027,2.4024618,2.4155898,2.353231,2.1070771,2.0053334,1.8445129,1.5589745,1.204513,1.1552821,1.4539489,1.7723079,1.8806155,1.6607181,1.3784616,0.96492314,0.62030774,0.4660513,0.5415385,0.33476925,0.2986667,0.32164106,0.32164106,0.26256412,0.25271797,0.2855385,0.4135385,0.58420515,0.6695385,0.67610264,0.6268718,0.56123084,0.47917953,0.35446155,0.25271797,0.21333335,0.19364104,0.17723078,0.16082053,0.17394873,0.18707694,0.18707694,0.17723078,0.18707694,0.21661541,0.256,0.318359,0.3708718,0.3446154,0.26912823,0.20348719,0.15097436,0.12143591,0.108307704,0.108307704,0.10502565,0.14441027,0.23630771,0.3511795,0.42338464,0.5481026,0.60061544,0.5546667,0.4594872,0.4660513,0.446359,0.4201026,0.38728207,0.34789747,0.029538464,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.059076928,0.029538464,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.026256412,0.13456412,0.026256412,0.026256412,0.16082053,0.4201026,0.7515898,0.9419488,0.51856416,0.571077,1.0305642,0.67610264,0.20020515,0.2100513,0.39712822,0.6498462,1.0371283,2.300718,3.7284105,5.3005133,6.183385,4.7261543,4.1911798,4.7228723,5.533539,6.6461544,8.910769,16.866463,25.265232,29.039593,27.008001,21.897848,21.336617,19.498669,18.668308,20.279797,24.923899,26.850464,23.732515,19.695591,16.676104,14.441027,10.738873,7.9983597,7.8047185,8.87795,7.066257,5.618872,4.7950773,4.164923,3.6332312,3.4264617,5.9995904,5.504,4.7392826,4.778667,4.972308,3.4855387,2.0742567,1.3259488,1.3686155,1.8707694,1.0732309,0.85005134,0.88287187,0.81394875,0.25271797,0.79097444,2.540308,3.442872,2.8356924,1.4703591,2.6223593,2.3302567,1.7099489,1.2931283,1.020718,0.58420515,0.34133336,0.23630771,0.29210258,0.6268718,0.3314872,0.29210258,0.50543594,0.78769237,0.761436,0.69579494,0.8369231,1.024,1.083077,0.8566154,0.79097444,0.90256417,1.1651284,1.2635899,0.56123084,1.0043077,1.020718,0.9124103,0.92553854,1.2504616,1.3029745,1.214359,1.1946667,1.204513,0.9353847,1.1520001,1.4933335,1.4211283,0.9714873,0.75487185,1.0699488,1.142154,1.1257436,1.1093334,1.1323078,0.9156924,0.73517954,0.7122052,0.72861546,0.42338464,1.4211283,1.9561027,2.0512822,1.9528207,2.1464617,2.546872,2.4024618,2.5238976,2.937436,2.8816411,2.2219489,2.0217438,2.0184617,2.5632823,4.604718,6.442667,7.1122055,6.488616,5.398975,5.6320004,7.062975,9.202872,11.657847,13.512206,13.3251295,10.571488,9.527796,11.713642,16.12472,19.236105,14.352411,10.469745,8.39877,8.247795,9.429334,8.973129,11.119591,12.419283,11.575796,9.4457445,8.444718,9.55077,11.562668,13.010053,12.1698475,13.174155,14.214565,15.084309,15.553642,15.360002,15.379693,15.514257,15.172924,14.247386,13.088821,10.86359,9.403078,9.481847,10.259693,9.281642,7.27959,6.4032826,7.6603084,9.833026,9.478565,9.009232,9.458873,9.590155,8.914052,7.6635904,8.661334,8.710565,7.702975,6.3507695,6.2096415,7.4404106,7.1154876,6.449231,5.691077,4.1058464,3.9286156,4.3716927,5.024821,5.2709746,4.279795,3.4100516,2.487795,2.7831798,3.7185643,2.8914874,3.3280003,3.3542566,3.5544617,3.7054362,2.7437952,2.8192823,2.9440002,2.412308,1.4605129,1.2865642,1.6114873,5.159385,11.346052,15.90154,10.909539,7.253334,10.417232,11.011283,7.1548724,4.457026,11.812103,10.098872,5.5958977,2.865231,4.7589746,5.5072823,4.95918,4.598154,4.7622566,4.6145644,7.88677,11.388719,11.011283,6.7216415,2.5731285,3.5544617,4.128821,4.201026,4.0402055,4.276513,2.9833848,2.9243078,3.564308,4.20759,3.9778464,3.5216413,3.6135387,3.4002054,2.7634873,2.3335385,3.5380516,2.993231,2.3335385,2.169436,2.100513,2.038154,2.5074873,3.639795,4.781949,4.5029745,3.255795,2.15959,1.5688206,1.4441026,1.3489232,4.8738465,12.803283,14.191591,8.487385,5.5269747,9.639385,12.337232,9.993847,4.125539,1.3915899,7.515898,8.989539,7.351795,4.70318,3.7218463,6.055385,6.498462,6.1308722,5.031385,2.284308,2.1169233,3.3542566,4.391385,4.1714873,2.1956925,1.5425643,3.2722054,8.100103,15.186052,22.12431,37.986465,50.543594,51.8039,40.598976,22.596926,14.851283,13.8075905,14.201437,12.882052,8.825437,9.508103,10.643693,10.768411,10.187488,10.9686165,10.919386,9.255385,8.828718,9.593436,8.585847,8.65477,7.702975,6.8430777,6.75118,7.6701546,6.166975,5.904411,5.35959,4.3651285,4.089436,3.636513,3.2098465,2.678154,2.294154,2.6847181,3.245949,2.92759,2.4188719,2.3401027,3.2328207,3.5446157,4.1682053,4.0303593,3.43959,4.07959,5.2676926,3.8728209,3.4658465,4.9329233,6.449231,7.817847,9.235693,9.3078985,8.953437,11.437949,9.412924,8.516924,8.356103,9.140513,11.697231,13.072412,14.404924,13.929027,12.924719,15.694771,21.093744,23.82113,25.793644,28.757336,34.287594,38.288414,47.11713,53.037952,53.395695,50.61908,41.22913,33.112617,27.536413,29.751797,49.014156,62.8677,57.767387,48.557953,48.67939,70.13416,79.31734,73.6197,67.15734,66.64862,71.41744,75.549545,77.60739,75.34934,72.82544,80.3676,89.81334,91.26073,89.47857,87.33211,85.7797,84.860725,77.88637,72.123085,73.3998,86.12103,90.233444,92.205956,93.18729,91.93683,84.831184,78.290054,77.32185,76.12062,73.422775,72.51036,83.83016,91.26729,91.359184,84.88698,76.855804,70.1079,67.390366,67.9319,68.98544,65.8117,69.474464,75.66113,79.01211,76.507904,67.49539,69.71078,68.181335,65.00103,60.48821,53.22175,48.31508,43.854774,45.26277,51.53149,55.204105,55.276314,54.63303,53.0478,50.707695,48.23303,46.834877,43.073643,43.008003,45.96513,44.530876,50.497646,52.414364,56.766365,67.82687,87.643906,87.936005,84.97559,78.5559,71.89006,71.611084,81.11919,84.48985,82.34995,76.16985,68.25683,66.868515,71.6997,78.299904,83.18359,83.82688,74.35816,70.90216,73.54749,79.602875,83.59057,80.49888,69.14298,61.042877,59.91385,61.65334,62.769234,68.37498,71.620926,71.03016,70.508316,74.69949,78.129234,81.37847,85.06421,89.8396,82.54031,65.581955,49.35549,39.01375,34.432003,31.448618,29.574566,29.184002,30.388515,33.043694,38.052105,41.373543,42.39754,41.294773,39.030155,34.819286,33.040413,31.993439,30.306463,26.942362,23.945848,21.477745,19.209848,17.056822,15.159796,14.050463,13.6467705,12.826258,11.546257,10.843898,10.197334,9.373539,8.553026,7.6734366,6.4065647,5.3103595,4.269949,3.2984617,2.425436,1.7165129,1.2307693,0.8730257,0.6170257,0.4397949,0.3314872,0.26912823,0.20676924,0.18707694,0.19364104,0.15097436,0.0951795,0.08205129,0.072205134,0.052512825,0.036102567,0.04266667,0.03938462,0.032820515,0.04594872,0.098461546,0.22646156,0.23958977,0.19692309,0.15753847,0.16738462,0.35446155,0.4397949,0.7187693,1.4900514,3.0752823,3.1113849,3.5741541,3.3444104,2.2908719,1.2406155,2.1267693,4.073026,6.3277955,7.515898,5.6385646,2.9669745,1.1520001,0.256,0.049230773,0.0032820515,0.0,0.006564103,0.013128206,0.013128206,0.016410258,0.013128206,0.128,0.256,0.3708718,0.51856416,1.2274873,1.782154,1.9232821,1.6738462,1.3357949,1.1257436,1.3522053,1.5064616,1.4441026,1.3686155,1.4834872,1.7033848,1.8182565,1.7296412,1.463795,1.204513,1.1651284,1.3456411,1.6180514,1.7362052,1.913436,1.595077,1.0962052,0.6859488,0.60389745,0.446359,0.37415388,0.33476925,0.30194873,0.29210258,0.26584616,0.23630771,0.27241027,0.4201026,0.7089231,0.8172308,0.764718,0.7056411,0.65312827,0.48246157,0.31507695,0.20348719,0.15425642,0.14769232,0.14769232,0.15425642,0.16410258,0.16410258,0.16082053,0.16082053,0.16410258,0.15425642,0.17066668,0.20676924,0.23958977,0.26912823,0.23630771,0.18707694,0.14441027,0.108307704,0.13456412,0.11158975,0.101743594,0.13128206,0.19364104,0.28882053,0.4201026,0.5284103,0.58092314,0.5481026,0.571077,0.5349744,0.4660513,0.39384618,0.3249231,0.15097436,0.04266667,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.059076928,0.28882053,0.15425642,0.049230773,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13784617,0.7122052,1.2373334,0.45620516,0.23958977,0.072205134,0.41025645,0.9714873,0.761436,0.48246157,1.0535386,1.4080001,1.1848207,0.7318975,2.8455386,4.9821544,6.3573337,6.875898,7.1548724,5.691077,4.417641,3.8038976,5.2381544,11.047385,21.372719,24.195284,22.229336,19.10154,19.334566,19.114668,18.78318,18.028309,18.343386,23.056412,24.336412,21.464617,18.819284,17.322668,14.404924,10.400822,8.008205,7.6767187,8.349539,7.4469748,5.8223596,4.713026,3.6857438,2.7798977,2.487795,5.3431797,5.2348723,4.5062566,4.2141542,4.1058464,3.4198978,2.802872,2.2514873,1.6016412,0.5021539,1.2603078,1.6869745,1.2373334,0.32820517,0.3511795,1.2307693,1.6968206,2.4910772,3.3017437,2.7766156,2.9111798,3.1638978,3.0720003,2.412308,1.204513,0.7187693,0.55794877,0.41682056,0.27241027,0.380718,0.5152821,0.6859488,0.80738467,0.8467693,0.82379496,0.78769237,0.57764107,0.6432821,0.892718,0.6859488,1.332513,1.467077,1.083077,0.47589746,0.24287182,0.20676924,0.318359,0.45620516,0.54482055,0.51856416,0.5316923,1.0108719,2.048,2.9144619,2.0611284,1.3259488,0.9353847,0.76800007,0.8041026,1.083077,0.9124103,1.3456411,1.3522053,0.7778462,0.3511795,0.72861546,0.81394875,0.6301539,0.38728207,0.47261542,0.5218462,0.8008206,1.024,1.2537436,1.8773335,1.8904617,2.0118976,1.9331284,2.172718,4.089436,2.5993848,2.0184617,2.1267693,2.6518977,3.249231,4.630975,6.0258465,5.832206,4.7556925,5.8289237,5.792821,7.2664623,9.147078,10.650257,11.323078,10.541949,12.09436,14.772514,17.939693,21.530258,15.133539,11.730052,9.819899,8.234667,6.1341543,6.1472826,12.511181,16.278976,15.622565,15.852309,14.9628725,15.031796,14.752822,13.367796,10.679795,11.595488,14.122667,16.548103,17.99549,18.448412,17.824821,18.15631,18.28431,17.545847,15.763694,13.528616,11.001437,9.317744,8.87795,9.353847,9.366975,9.53436,9.711591,9.55077,8.513641,10.075898,10.587898,9.616411,7.8703594,7.1876926,8.615385,8.999385,8.395488,7.017026,5.2348723,5.7698464,6.764308,7.351795,6.5083084,3.0687182,3.8498464,3.8071797,3.4822567,3.0818465,2.4713848,1.591795,1.5556924,2.1431797,3.0490258,3.892513,4.3290257,3.131077,2.9965131,4.2830772,4.9887185,4.4898467,4.197744,3.117949,1.654154,1.6180514,3.3247182,5.76,7.6012316,7.686565,4.9887185,3.5971284,5.8781543,5.927385,3.6496413,4.7622566,10.095591,8.464411,4.893539,3.0490258,5.2348723,5.172513,4.4438977,3.748103,3.3575387,3.1113849,3.2098465,2.3827693,1.3718976,0.79097444,1.1454359,3.170462,5.435077,6.314667,5.924103,6.117744,5.3727183,5.362872,4.9821544,4.013949,3.0982566,3.367385,4.420923,4.1517954,2.481231,1.3587693,3.761231,3.761231,2.7766156,1.8543591,1.6475899,3.1015387,4.342154,4.630975,3.6758976,1.6475899,1.1126155,1.4900514,2.3991797,3.131077,2.6551797,7.4404106,12.819694,12.166565,5.917539,1.5721027,7.200821,10.06277,8.375795,3.7710772,1.2832822,4.9427695,6.170257,4.663795,2.8192823,5.737026,8.264206,7.3583593,5.179077,3.190154,2.1530259,2.7733335,2.7634873,2.5764105,2.156308,0.9616411,1.0699488,3.8531284,6.557539,10.896411,23.04,43.854774,50.88821,44.192825,29.06585,16.052513,12.87877,12.3306675,11.122872,8.362667,5.5532312,7.604513,8.914052,9.048616,8.674462,9.55077,8.674462,6.7774363,7.827693,10.587898,8.621949,8.730257,7.752206,6.1341543,4.788513,5.080616,6.6560006,7.204103,6.1505647,4.345436,4.089436,4.6145644,4.818052,4.33559,3.1737437,1.7099489,1.8674873,2.7667694,3.383795,3.892513,5.661539,6.294975,5.7501545,4.644103,3.5183592,2.8225644,5.142975,4.8804107,5.8125134,9.6984625,16.265848,16.265848,13.115078,11.536411,12.937847,15.442053,10.925949,9.796924,9.91836,11.59877,17.591797,23.207386,23.798155,22.229336,22.006155,27.267284,29.709131,35.078568,42.525543,49.926567,53.891285,52.40452,52.033646,48.50544,41.04862,32.39713,27.378874,24.356104,25.376822,34.402466,57.327595,63.30749,55.05313,47.986874,52.653954,74.735596,74.689644,58.446774,44.711388,40.546463,41.353848,40.26749,45.095387,49.611492,51.13108,50.507492,52.818054,57.94462,60.90175,56.651493,40.08698,36.76882,33.237335,33.22421,37.5598,44.176414,40.956722,41.806774,44.688416,46.3918,42.55836,35.77108,36.90339,41.27508,45.059284,45.28903,49.09949,54.55426,53.293953,45.58113,40.33313,37.90113,33.046978,32.833645,38.383595,44.878773,46.342567,42.745438,36.83118,31.766977,31.130259,34.7799,32.98462,31.474874,31.602875,30.319592,28.842669,29.94872,31.766977,32.817234,32.000004,36.11241,37.06749,36.164925,35.784206,39.384617,39.322258,35.616825,34.146465,35.974567,37.353027,43.21477,47.123695,50.261337,53.293953,56.382362,61.108517,63.744003,64.51201,65.92329,72.782776,81.69682,84.7918,80.78442,71.309135,60.944416,56.94031,57.330875,60.56698,66.78647,77.820724,76.6359,75.02113,77.010056,81.84452,83.96801,81.552414,75.93026,75.375595,77.88965,71.21067,64.47262,64.50216,67.18031,71.91303,81.60165,95.83591,94.58872,94.10626,97.115906,92.8197,81.417854,63.46175,48.751595,42.17108,43.684105,42.000412,43.11631,46.585438,50.93744,53.710773,60.67857,65.79201,66.19898,61.663185,54.53457,47.88185,42.36472,38.468925,34.97682,28.944412,24.159182,21.874874,20.207592,18.38277,16.722052,15.711181,14.614976,13.761642,13.124924,12.343796,11.85477,10.935796,10.016821,9.140513,7.9786673,6.941539,5.8945646,4.8147697,3.7316926,2.7306669,1.9987694,1.4506668,1.0469744,0.761436,0.56451285,0.44307697,0.36758977,0.34133336,0.32164106,0.19692309,0.12471796,0.108307704,0.08205129,0.049230773,0.06235898,0.098461546,0.108307704,0.08205129,0.06235898,0.12143591,0.23302566,0.26912823,0.3052308,0.3511795,0.3511795,0.25271797,0.32164106,1.3226668,2.612513,2.1366155,1.5261539,1.3718976,1.8740515,2.5009232,1.9987694,1.6804104,2.2416413,3.2623591,4.125539,4.027077,2.2350771,0.92553854,0.23630771,0.052512825,0.016410258,0.0032820515,0.0,0.0,0.0032820515,0.016410258,0.0032820515,0.0,0.055794876,0.20020515,0.45620516,0.92225647,0.88287187,0.80738467,0.85005134,0.82379496,0.6892308,0.88615394,1.079795,1.148718,1.1585642,1.3423591,1.7624617,2.166154,2.2711797,1.7690258,1.3423591,1.1520001,1.2274873,1.4572309,1.6016412,1.6640002,1.8051283,1.7460514,1.3128207,0.45620516,0.54482055,0.51856416,0.4397949,0.35446155,0.3052308,0.26912823,0.2231795,0.20348719,0.256,0.4266667,0.6826667,0.67282057,0.571077,0.4955898,0.51856416,0.46933338,0.256,0.128,0.13456412,0.12143591,0.108307704,0.108307704,0.11158975,0.12471796,0.13784617,0.15097436,0.14441027,0.13784617,0.15425642,0.2297436,0.3249231,0.29538465,0.21661541,0.14441027,0.108307704,0.108307704,0.13456412,0.15097436,0.14441027,0.108307704,0.15425642,0.24943592,0.43323082,0.6235898,0.6104616,0.67282057,0.6235898,0.5316923,0.43651286,0.3511795,0.2986667,0.12143591,0.08205129,0.052512825,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.068923086,0.3511795,0.44964105,0.190359,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.32164106,0.7778462,1.0108719,0.48246157,1.2307693,1.9003079,1.8838975,1.2209232,0.5907693,0.3117949,0.58092314,1.1520001,2.100513,3.8465643,6.0652313,8.65477,13.466257,17.847795,14.651078,9.252103,5.7632823,4.7622566,6.1013336,8.923898,13.5778475,17.536001,19.465847,19.419899,18.83241,19.140924,20.201027,19.685745,18.103796,18.819284,19.895796,18.720821,17.132309,15.53395,12.891898,9.783795,7.837539,7.1614366,7.1089234,6.2752824,4.7392826,3.7087183,2.7503593,1.9659488,1.975795,4.128821,4.634257,4.141949,3.3312824,2.9078977,3.436308,3.4921029,2.4582565,0.96492314,0.88287187,1.1126155,1.0043077,1.3029745,1.8806155,1.7165129,2.5271797,1.9823592,1.529436,1.6213335,1.6902566,1.8248206,1.8806155,1.7493335,1.4506668,1.1191796,1.020718,0.9911796,0.761436,0.41025645,0.3446154,0.47917953,0.5415385,0.60389745,0.7450257,1.0305642,0.9944616,0.8795898,0.56123084,0.23958977,0.44307697,0.8467693,0.8763078,0.67610264,0.4955898,0.6826667,0.40369233,0.5546667,0.7778462,0.86317956,0.7515898,0.88943595,1.1224617,1.6082052,2.0873847,1.8773335,1.5064616,0.9616411,0.5973334,0.5284103,0.6432821,0.764718,0.8763078,0.86974365,0.76800007,0.7417436,0.7581539,0.827077,0.73517954,0.5513847,0.6071795,0.77456415,1.0962052,1.6147693,2.0939488,2.0217438,1.9364104,2.3433847,3.2361028,3.9614363,3.2229745,2.1431797,2.4615386,3.6004105,4.630975,4.263385,3.826872,4.7327185,6.042257,7.5454364,9.770667,8.300308,6.2720003,5.9503593,7.197539,7.4896417,9.442462,11.913847,11.976206,10.587898,12.596514,9.586872,9.353847,9.527796,8.63836,6.11118,6.0619493,11.644719,14.54277,12.970668,11.680821,11.716924,12.809847,14.040616,14.158771,11.559385,10.581334,10.033232,10.459898,11.579078,12.2847185,11.749744,12.291283,12.58995,12.228924,11.684103,10.70277,10.282667,10.584617,10.9686165,10.000411,8.605539,9.002667,10.056206,10.748719,10.151385,9.426052,9.088,8.264206,7.0826674,6.6625648,7.066257,7.003898,6.6034875,5.835488,4.5029745,4.8147697,4.97559,4.4307694,3.2623591,2.2121027,3.0720003,2.9538465,2.9702566,3.1638978,2.484513,2.044718,2.4320002,2.9111798,3.2361028,3.6594875,4.0992823,2.5928206,1.8510771,3.3542566,7.3321033,7.896616,5.917539,3.446154,2.3433847,4.279795,3.9745643,4.1189747,4.5587697,5.028103,5.1232824,4.1517954,4.273231,5.0543594,6.163693,7.3714876,7.8637953,6.0619493,4.5029745,4.276513,5.024821,4.086154,4.637539,5.431795,5.152821,2.428718,1.7558975,1.6377437,1.9429746,2.5698464,3.4527183,4.315898,4.7655387,5.041231,5.481026,6.5444107,7.1187696,6.163693,4.5456414,3.114667,2.7076926,3.5905645,4.023795,3.370667,2.1530259,2.0545642,2.6420515,2.6847181,2.540308,2.4155898,2.3433847,3.817026,4.082872,3.245949,1.9692309,1.4769232,1.7690258,2.5764105,3.1540515,3.045744,2.0808206,3.2328207,4.594872,4.082872,1.9790771,0.92553854,2.7536411,3.114667,2.6683078,2.7995899,5.602462,6.9710774,4.7589746,2.7503593,2.9702566,5.7140517,5.113436,4.466872,3.5971284,3.0030773,3.8596926,4.9821544,4.9788723,5.0051284,4.391385,0.65641034,1.2438976,3.6726158,7.02359,12.757335,24.687592,36.214157,38.006157,32.676105,22.954668,11.670976,11.004719,10.57477,9.380103,7.768616,7.4207187,8.779488,8.530052,7.7325134,7.1220517,7.1122055,8.329846,9.012513,8.631796,7.788308,8.205129,9.83959,10.082462,7.824411,4.7655387,5.412103,5.3924108,5.3103595,5.7796926,6.5247183,6.3967185,4.5390773,3.948308,3.570872,2.8914874,1.9528207,2.8849232,2.9965131,2.7766156,3.0720003,5.0871797,7.821129,6.987488,4.6572313,2.793026,3.249231,5.208616,5.0838976,5.8978467,8.946873,13.774771,15.642258,16.33477,17.03713,18.438566,20.716309,14.976001,12.826258,12.455385,13.505642,17.06995,19.216412,20.647387,22.62318,26.098873,31.72431,32.758156,35.426464,39.909748,44.471798,45.472824,42.322056,38.52472,37.697643,38.409847,34.189133,34.21867,37.044518,38.324516,39.663593,48.623592,48.833645,38.2359,31.40595,33.72636,41.363697,34.901337,26.919386,23.082668,24.356104,26.998156,32.062363,34.76021,32.32821,26.883284,25.409643,31.993439,37.034668,39.46995,37.540104,28.757336,30.516516,34.244926,35.91549,34.753643,33.22421,34.54359,35.620106,34.605953,31.054771,25.944618,23.617643,24.960001,28.514463,32.019695,32.39713,34.067696,35.5118,34.6519,31.251696,26.902977,25.557335,24.392206,22.849644,22.147284,25.271797,26.200617,23.824411,19.994259,17.493334,20.033642,20.969027,17.51631,15.481437,16.922258,20.151796,26.262976,29.06585,28.66872,26.528822,25.46872,28.009027,27.96308,28.481644,30.454157,32.512,32.820515,32.07221,32.534977,34.1399,34.471386,31.766977,33.67713,34.517338,33.043694,32.43323,37.89785,40.64821,42.88985,46.116108,51.081852,55.30585,57.06175,54.770878,51.154057,53.24144,53.251286,52.302773,52.8279,55.502773,59.24103,59.99262,62.066875,65.7756,70.642876,75.4117,75.008,74.574776,74.13826,73.97744,74.6437,72.55303,70.33765,71.18442,77.90278,92.90832,111.72103,116.95591,117.021545,116.00411,113.68042,97.073235,79.744,70.72165,68.32575,60.153442,54.531284,58.098877,65.94626,74.15467,79.79652,76.58011,72.15262,67.46257,62.050465,54.035698,45.66318,38.242466,32.68595,28.58995,24.257643,21.464617,20.115694,19.252514,18.520617,18.189129,18.31713,18.028309,17.499899,16.649847,15.113848,13.797745,12.727796,11.71036,10.660104,9.616411,8.4512825,7.3714876,6.370462,5.362872,4.194462,3.1507695,2.3171284,1.6672822,1.1782565,0.8566154,0.6662565,0.53825647,0.46933338,0.4135385,0.27241027,0.17066668,0.12143591,0.108307704,0.15097436,0.32820517,0.67938465,1.020718,0.80738467,0.2100513,0.13456412,0.29210258,0.5677949,0.95835906,1.1913847,0.7417436,0.4201026,1.7558975,4.017231,5.5269747,3.6726158,3.5807183,4.4373336,4.6145644,3.6004105,1.9856411,1.5524104,1.4112822,1.6049232,1.9396925,1.9889232,1.1815386,0.56451285,0.19364104,0.04266667,0.016410258,0.0032820515,0.0,0.0,0.0032820515,0.016410258,0.013128206,0.013128206,0.029538464,0.08205129,0.20020515,0.4397949,0.8369231,1.1716924,1.1815386,0.54482055,0.41025645,0.44307697,0.5218462,0.61374366,0.7811283,1.0929232,1.463795,1.7887181,1.9429746,1.7952822,1.6804104,1.5458462,1.3751796,1.2406155,1.3095386,1.4473847,1.4441026,1.3718976,1.2340513,0.94523084,0.8369231,0.6104616,0.46276927,0.4135385,0.3052308,0.26912823,0.24615386,0.21661541,0.19692309,0.23302566,0.32164106,0.31507695,0.2986667,0.3446154,0.4955898,0.4660513,0.32820517,0.19692309,0.118153855,0.098461546,0.08533334,0.08205129,0.08205129,0.08861539,0.101743594,0.11158975,0.108307704,0.0951795,0.0951795,0.118153855,0.13784617,0.16082053,0.16082053,0.13456412,0.108307704,0.108307704,0.13456412,0.15097436,0.14112821,0.0951795,0.1148718,0.15097436,0.21989745,0.32164106,0.4266667,0.5874872,0.6268718,0.60389745,0.5481026,0.47261542,0.16082053,0.06235898,0.04594872,0.029538464,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.029538464,0.14769232,0.2100513,0.09189744,0.0,0.013128206,0.06564103,0.049230773,0.01969231,0.0,0.01969231,0.101743594,0.04266667,0.009846155,0.0,0.0,0.0,0.0,0.16738462,0.33805132,0.446359,0.52512825,1.7920002,1.9659488,1.6377437,1.1585642,0.6301539,0.6071795,1.4309745,3.370667,5.937231,7.9097443,7.8703594,10.745437,16.088617,19.951591,14.867694,10.482873,6.62318,5.1364107,5.910975,6.882462,9.435898,14.621539,18.435284,19.577436,19.449438,18.642054,18.763489,17.795284,16.150976,16.689232,17.801847,16.804104,14.880821,12.724514,10.551796,8.411898,6.810257,5.901129,5.467898,4.9296412,4.023795,3.259077,2.5107694,1.9298463,1.9200002,3.114667,3.5610259,3.639795,3.3444104,2.281026,3.1376412,3.3608208,2.4024618,0.9189744,0.764718,1.6246156,1.8281027,2.1989746,2.9636924,3.7448208,2.4516926,1.8445129,1.657436,1.6147693,1.4112822,1.5885129,1.7591796,2.0512822,2.2121027,1.6213335,1.2996924,1.4605129,1.332513,0.827077,0.51856416,0.5513847,0.43651286,0.36430773,0.4594872,0.79097444,0.76800007,0.7122052,0.67938465,0.69251287,0.74830776,0.81066674,0.7515898,0.55794877,0.40697438,0.65641034,0.76800007,0.8172308,0.8205129,0.88943595,1.2307693,1.4441026,1.4408206,1.5753847,1.7329233,1.3193847,1.1388719,0.8566154,0.75487185,0.86317956,0.96492314,0.99774367,1.0929232,1.2012309,1.2406155,1.0962052,0.8992821,0.92553854,0.82379496,0.6170257,0.69579494,1.1027694,1.4900514,1.9528207,2.3269746,2.1792822,2.3335385,2.5173335,2.7634873,3.131077,3.7120004,2.6683078,3.1343591,4.2174363,5.1364107,5.221744,4.95918,5.477744,6.088206,6.7216415,7.9458466,7.3747697,6.0947695,5.3070774,5.182359,4.8640003,5.684513,7.3058467,7.7456417,7.1187696,7.634052,6.6002054,8.149334,9.53436,9.238976,6.9809237,6.744616,9.741129,10.912822,9.586872,9.481847,10.161232,10.761847,11.428103,11.9860525,11.936821,10.220308,8.976411,8.474257,8.89436,10.328616,9.291488,9.028924,9.596719,10.518975,10.7848215,9.219283,8.960001,9.895386,11.264001,11.654565,11.001437,10.896411,10.916103,10.709334,10.010257,8.467693,7.1614366,6.3474874,6.042257,6.009436,6.0980515,5.737026,4.95918,3.9384618,3.0096412,3.8728209,4.854154,4.5587697,3.190154,2.546872,3.1573336,3.3476925,4.8640003,6.9152827,6.1768208,4.785231,4.9821544,5.07077,4.716308,4.9362054,5.691077,4.0402055,2.934154,3.7021542,6.0258465,6.3212314,4.9920006,4.141949,4.6572313,6.2162056,4.7524104,4.2830772,4.890257,5.9569235,6.163693,4.70318,4.962462,5.802667,6.4722056,6.5969234,5.4908724,5.7665644,6.701949,7.312411,6.3573337,4.266667,4.3585644,4.699898,4.0992823,2.0939488,3.0884104,3.7415388,4.010667,4.4964104,6.4557953,5.7764106,4.414359,3.9647183,4.84759,6.340924,5.9930263,4.781949,3.5347695,2.9111798,3.4133337,3.5741541,3.4002054,3.131077,2.9768207,3.1343591,3.0260515,2.9407182,2.917744,2.8750772,2.6190772,2.8225644,2.5632823,2.0939488,1.7920002,2.156308,2.5107694,2.4648206,2.3630772,2.5074873,3.1638978,3.006359,3.6562054,4.345436,4.781949,5.1200004,4.2502565,2.556718,1.6344616,3.0490258,8.329846,8.077128,4.70318,2.3762052,2.537026,3.9023592,3.623385,4.1714873,4.598154,4.6145644,4.598154,4.4734364,3.889231,3.626667,3.2065644,0.8992821,0.9485129,3.7251284,7.9163084,12.721231,17.867489,25.170053,26.643694,22.849644,15.839181,9.156924,12.471796,12.547283,12.3076935,12.438975,11.369026,9.849437,7.8834877,6.75118,6.449231,5.677949,6.889026,8.792616,8.211693,5.989744,6.994052,7.90318,7.141744,5.156103,4.2174363,8.457847,8.533334,6.0750775,4.4045134,4.7655387,6.314667,4.519385,4.6867695,5.0051284,4.7261543,4.1846156,6.3606157,6.3474874,5.2348723,4.2535386,4.7622566,6.1308722,5.225026,4.2962055,4.821334,7.4863596,9.176616,11.08677,13.131488,15.307488,17.667284,18.730669,18.471386,18.028309,18.241642,19.636515,16.90913,15.465027,14.775796,14.87754,16.351181,18.182566,22.38031,26.758566,31.002258,36.673645,38.242466,36.877132,35.380516,34.435284,32.59077,30.644516,30.900515,34.69785,38.754463,35.160618,32.600616,33.82154,33.66072,31.497849,31.261541,28.422565,21.024822,16.072206,15.82277,17.785437,14.12595,11.510155,11.195078,12.983796,15.205745,18.819284,20.841026,20.397951,18.793028,19.51836,24.982977,28.36349,30.595284,30.690464,25.760822,25.51467,29.689438,33.217644,32.899284,27.43795,28.009027,30.933336,30.792208,26.361439,20.598156,18.694565,18.369642,20.25354,22.934977,22.967796,26.725746,30.165335,31.379694,29.472822,24.579285,20.86072,17.641027,15.419078,15.333745,19.154053,21.812515,18.87836,14.65436,12.219078,13.423591,13.971693,12.176412,11.034257,12.777026,18.86195,23.906464,26.423798,27.733335,27.615181,24.346258,23.302567,23.427284,25.127386,28.182976,31.744003,31.041643,30.864412,31.320618,32.01641,32.068924,27.910566,26.952208,26.197336,25.127386,25.682053,28.583387,30.286772,31.071182,31.573336,32.784412,33.667286,36.16821,38.52472,41.06503,46.208004,47.218876,47.38954,47.218876,47.13354,47.481438,47.104004,48.196926,50.43857,52.64739,52.785236,50.304005,51.25908,54.400005,59.024414,64.95508,66.68472,64.58421,63.63898,67.93519,80.65642,93.88637,104.0837,112.0197,117.53683,119.57498,108.83611,98.46811,95.22216,96.07877,88.24452,81.82483,86.52473,91.11303,89.73457,81.92329,75.2476,68.28636,62.720005,58.21375,52.42749,44.862362,37.993027,33.375183,30.595284,27.250874,24.237951,22.44595,21.668104,21.651693,22.107899,22.87918,23.184412,23.243488,22.856207,21.382566,19.035898,16.17395,13.899488,12.484924,11.362462,10.295795,9.189744,8.090257,6.997334,5.861744,4.709744,3.6496413,2.7241027,1.972513,1.4441026,1.1257436,0.8795898,0.69251287,0.5415385,0.380718,0.24287182,0.14769232,0.10502565,0.15425642,0.36102566,0.58092314,0.8369231,0.69579494,0.27897438,0.256,0.46276927,0.6662565,0.9714873,1.2964103,1.3784616,2.737231,5.0609236,6.377026,6.619898,7.637334,8.172308,7.026872,5.221744,3.6529233,3.1015387,2.789744,2.1989746,1.8871796,1.9495386,2.0217438,1.4966155,0.8467693,0.33805132,0.07876924,0.02297436,0.0032820515,0.0,0.0,0.0,0.006564103,0.006564103,0.006564103,0.009846155,0.026256412,0.08205129,0.21333335,1.3653334,2.359795,2.428718,1.1946667,0.85005134,0.6859488,0.5152821,0.34789747,0.40369233,0.5973334,0.85005134,1.1224617,1.3587693,1.4900514,1.6443079,1.6443079,1.5064616,1.3226668,1.2537436,1.273436,1.1454359,1.0108719,0.892718,0.7122052,0.53825647,0.38400003,0.28882053,0.24615386,0.20348719,0.190359,0.18379489,0.17066668,0.15425642,0.14769232,0.16738462,0.16410258,0.17723078,0.23302566,0.3511795,0.34133336,0.28225642,0.2231795,0.17066668,0.101743594,0.07548718,0.06564103,0.06235898,0.059076928,0.06564103,0.07548718,0.07548718,0.07548718,0.07548718,0.072205134,0.072205134,0.08861539,0.09189744,0.08205129,0.07876924,0.072205134,0.108307704,0.13784617,0.13456412,0.09189744,0.10502565,0.12471796,0.15753847,0.20348719,0.28225642,0.43323082,0.56123084,0.6629744,0.7089231,0.65969235,0.026256412,0.006564103,0.006564103,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.06564103,0.049230773,0.01969231,0.0,0.01969231,0.101743594,0.04266667,0.052512825,0.07876924,0.07876924,0.0,0.0,0.02297436,0.02297436,0.06564103,0.32820517,1.8116925,2.1825643,2.2547693,2.3630772,2.353231,1.8838975,2.4385643,4.6867695,7.8080006,9.472001,7.1647186,10.66995,16.164104,18.609232,11.772718,10.157949,7.9885135,6.5247183,6.0750775,6.0028725,7.857231,11.881026,15.750566,18.067694,18.379488,17.46708,16.971489,15.832617,14.585437,15.360002,15.868719,14.408206,12.071385,9.737847,8.064001,6.8529234,5.7632823,5.0215387,4.667077,4.532513,4.096,3.4231799,2.7175386,2.166154,1.9265642,2.284308,2.4910772,2.989949,3.3247182,2.103795,2.5665643,2.868513,2.3466668,1.2406155,0.69251287,1.6246156,1.7920002,1.8576412,2.3368206,3.5872824,2.0611284,1.6902566,1.6869745,1.6147693,1.3915899,1.4441026,1.6147693,1.972513,2.3171284,2.1891284,2.4648206,2.4943593,1.9462565,1.079795,0.7318975,0.58420515,0.45620516,0.36758977,0.41025645,0.73517954,0.69907695,0.67610264,0.86317956,1.1257436,1.017436,0.90256417,0.80738467,0.67610264,0.571077,0.6432821,0.85005134,0.86974365,0.8336411,0.9682052,1.6082052,2.156308,1.8707694,1.6147693,1.6049232,1.4145643,1.5392822,1.4834872,1.3784616,1.2964103,1.2635899,0.98461545,1.0371283,1.2537436,1.3883078,1.1191796,0.81066674,0.84348726,0.8992821,0.86646163,0.82379496,1.079795,1.3784616,1.9429746,2.6157951,2.8324106,3.6562054,3.117949,2.540308,2.8882053,4.7655387,3.0391798,2.9735386,3.8432825,5.0182567,5.9470773,6.619898,6.8332314,6.1472826,5.1626673,5.5302567,5.9602056,6.042257,5.618872,4.824616,4.1025643,3.9778464,4.4274874,4.95918,5.2578464,5.159385,4.634257,6.564103,8.162462,8.274052,7.39118,7.64718,9.074872,9.396514,8.809027,9.987283,10.824206,9.970873,8.89436,8.710565,10.220308,10.266257,10.253129,9.189744,7.9852314,9.475283,8.585847,8.083693,8.651488,10.108719,11.418258,10.072617,8.65477,8.454565,9.741129,11.746463,11.707078,11.034257,10.269539,9.494975,8.342975,7.578257,5.8486156,4.8640003,5.074052,5.684513,5.330052,4.9362054,4.325744,3.754667,3.9318976,4.5587697,5.5762057,5.737026,5.0149746,4.598154,4.824616,5.152821,6.8332314,8.841846,7.8670774,6.11118,6.229334,6.626462,6.482052,5.756718,5.9634876,5.9963083,6.5247183,7.020308,5.7731285,4.562052,5.0838976,6.4656415,7.565129,6.9743595,4.644103,4.4340515,5.277539,5.9667697,5.169231,4.1747694,5.290667,6.1046157,5.8945646,5.61559,4.8738465,6.124308,7.5388722,7.90318,6.6133337,4.1124105,3.820308,3.7349746,3.2131286,2.9472823,7.5552826,9.137232,7.640616,5.4941545,7.6012316,6.616616,4.322462,3.3017437,4.138667,5.4383593,4.854154,3.4888208,2.5698464,2.6617439,3.6463592,3.121231,2.6026669,2.5993848,3.0818465,3.4625645,3.5183592,3.2196925,2.8849232,2.6584618,2.5074873,2.15959,1.7690258,1.7493335,2.1989746,2.9013336,2.737231,2.0250258,2.0250258,3.3411283,5.8912826,5.861744,5.3398976,5.290667,5.7435904,5.8125134,4.3060517,2.5304618,1.6377437,2.6683078,6.554257,5.8781543,3.570872,2.038154,1.9331284,2.162872,4.315898,6.9054365,7.315693,5.586052,4.414359,3.2722054,2.7602053,2.8521028,2.9472823,1.8773335,1.5885129,5.5597954,9.977437,12.20595,10.774975,14.624822,17.106052,15.737437,11.67754,9.728001,13.5778475,12.763899,11.648001,11.835078,12.179693,10.738873,8.480822,7.4929237,7.4207187,5.4514875,6.3179493,8.457847,7.9261546,5.477744,6.560821,6.5312824,5.431795,4.886975,7.1515903,15.117129,14.309745,10.640411,6.9087186,5.1232824,6.498462,5.0871797,5.477744,5.7829747,5.5663595,5.8453336,8.086975,9.321027,8.835282,7.240206,6.4689236,5.5105643,5.1331286,5.7764106,7.525744,10.112,11.713642,14.92677,17.184822,18.067694,19.27877,19.551182,18.297438,18.028309,19.606976,22.239182,21.96349,20.447182,18.346668,16.538258,16.114874,19.042463,23.870361,28.032001,31.40595,36.34544,37.58277,32.564514,27.707079,25.892105,26.473028,24.293745,28.015593,32.515285,33.207798,26.04308,23.683285,22.86277,21.320208,18.425438,15.195899,12.49477,9.570462,7.430565,6.5870776,7.056411,6.370462,6.0192823,6.1505647,6.7544622,7.64718,9.032206,10.384411,11.976206,13.853539,15.839181,19.695591,22.278566,23.929438,24.415182,22.915283,19.794052,22.117744,26.256413,28.586668,25.504822,25.649233,27.858053,27.812105,24.448002,19.977848,17.769028,15.05477,14.641232,16.338053,16.945232,20.407797,23.210669,24.185438,22.767591,18.98995,15.363283,12.199386,11.529847,14.503386,21.372719,24.49395,20.801643,15.970463,12.852514,11.480617,12.2387705,11.464206,11.076924,13.308719,20.686771,24.71713,29.049438,32.564514,33.35549,28.734362,25.189745,22.849644,22.629745,24.625233,28.09436,30.578875,33.122463,34.048004,32.92554,30.578875,27.270567,24.976412,23.758772,23.88677,25.823181,26.450054,27.300104,26.998156,25.554052,24.359386,25.85272,28.281439,31.130259,34.034874,36.785233,36.545643,37.72062,38.741337,39.03672,39.023594,37.855183,37.264412,37.438362,37.576206,35.895798,32.656414,33.28985,37.333336,43.700516,50.691284,54.239185,52.059902,49.02072,49.39816,56.864826,65.414566,76.045135,87.3157,97.25375,103.34196,97.887184,94.23426,94.89724,98.38934,99.23611,102.974365,108.74422,106.93581,96.07221,82.82257,78.10954,73.36698,67.40678,60.94113,56.546467,50.284313,44.66872,40.799183,38.265438,35.144207,31.734156,29.4039,28.517746,28.79672,29.321848,29.919182,30.211285,29.974977,29.078976,27.474054,24.87795,20.847591,17.253744,14.841437,13.210258,12.176412,11.122872,10.033232,8.933744,7.8834877,6.7938466,5.5597954,4.391385,3.4166157,2.674872,2.1136413,1.5688206,1.0994873,0.7417436,0.5021539,0.3314872,0.19692309,0.12143591,0.128,0.256,0.3117949,0.40369233,0.37743592,0.30194873,0.47589746,0.69907695,0.79425645,1.2504616,2.3204105,4.027077,6.9087186,8.740103,8.467693,7.752206,10.95877,11.605334,8.257642,4.667077,3.0260515,3.948308,3.6135387,3.0227695,2.8356924,3.1442053,3.4855387,2.0873847,1.0568206,0.42338464,0.13456412,0.036102567,0.006564103,0.0032820515,0.006564103,0.0032820515,0.0,0.0,0.0032820515,0.006564103,0.02297436,0.08205129,0.44307697,1.5819489,2.5009232,2.5304618,1.3128207,1.083077,1.020718,0.761436,0.34133336,0.19692309,0.318359,0.45292312,0.60061544,0.7581539,0.9156924,1.1913847,1.332513,1.3620514,1.3128207,1.1979488,1.1355898,1.0043077,0.88615394,0.77128214,0.5349744,0.3314872,0.24287182,0.18379489,0.13128206,0.12471796,0.13456412,0.15097436,0.16082053,0.15097436,0.128,0.1148718,0.101743594,0.1148718,0.15753847,0.21661541,0.2297436,0.23630771,0.23958977,0.22646156,0.14441027,0.072205134,0.052512825,0.04594872,0.03938462,0.03938462,0.04594872,0.052512825,0.059076928,0.06235898,0.055794876,0.055794876,0.055794876,0.052512825,0.049230773,0.055794876,0.04266667,0.06564103,0.08861539,0.09189744,0.072205134,0.07548718,0.098461546,0.13128206,0.16082053,0.18379489,0.27241027,0.40697438,0.56451285,0.6892308,0.69579494,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08205129,0.15753847,0.15753847,0.0,0.0,0.006564103,0.006564103,0.0,0.0,1.6869745,3.1245131,3.9023592,4.1714873,4.644103,3.4560003,3.2295387,5.0149746,7.817847,8.605539,4.8738465,8.185436,13.351386,15.07118,7.9261546,8.264206,8.237949,7.3353853,6.0750775,6.009436,7.5552826,8.845129,11.539693,14.930053,15.963899,16.423386,16.114874,14.86113,13.426873,13.51877,13.177437,11.480617,9.278359,7.282872,6.048821,5.664821,5.2348723,4.9526157,4.903385,5.0609236,4.716308,3.9089234,3.0523078,2.3860514,1.9561027,1.6836925,1.6607181,2.2711797,2.9997952,2.409026,2.0709746,2.300718,2.1792822,1.522872,0.892718,1.0371283,0.73517954,0.5546667,0.82379496,1.6213335,1.6804104,1.5163078,1.3817437,1.4112822,1.6410258,1.2964103,1.2832822,1.3423591,1.5524104,2.300718,3.5314875,3.2984617,2.297436,1.2832822,1.0633847,0.69251287,0.6465641,0.65641034,0.67282057,0.88615394,0.764718,0.7417436,0.86974365,1.0436924,0.9878975,1.0633847,1.0666667,1.0404103,0.9911796,0.8960001,0.77456415,0.7417436,0.8008206,1.0305642,1.595077,2.546872,2.0906668,1.5491283,1.522872,1.913436,2.2514873,2.5238976,2.281026,1.6213335,1.1815386,0.7450257,0.7056411,0.892718,1.0601027,0.88615394,0.574359,0.65969235,0.9616411,1.1913847,0.92553854,0.8041026,0.88287187,1.5524104,2.6322052,3.387077,5.549949,4.57518,3.5774362,3.9844105,5.5105643,3.6332312,2.7536411,3.0654361,4.2929235,5.677949,7.1548724,7.1515903,5.802667,4.2962055,4.8738465,5.3070774,5.668103,5.986462,6.2129235,6.23918,6.51159,5.976616,5.142975,4.4767184,4.4012313,3.5905645,5.0116925,6.117744,6.413129,7.466667,8.477539,9.173334,9.373539,9.649232,11.339488,11.88759,9.954462,7.39118,5.940513,7.2270775,10.029949,12.179693,11.32636,8.598975,8.608821,7.9950776,8.034462,8.595693,9.741129,11.749744,11.762873,9.357129,7.6077952,7.955693,10.20718,9.734565,8.953437,8.379078,7.837539,6.4623594,6.629744,5.3792825,4.598154,5.034667,6.294975,5.3858466,4.9394875,5.0904617,6.0717955,8.218257,7.1483083,6.616616,6.636308,6.941539,6.994052,7.066257,7.0826674,7.315693,7.394462,6.314667,5.159385,5.3825645,6.4557953,7.131898,5.425231,4.529231,6.7282057,9.563898,10.564924,7.213949,4.818052,6.7117953,8.835282,8.930462,6.521436,4.1222568,4.33559,4.9952826,4.7294364,2.986667,3.2065644,4.8311796,5.8978467,5.83877,5.4449234,5.602462,5.8847184,5.7829747,5.277539,4.8344617,3.0916924,3.1507695,3.4494362,3.6004105,4.397949,11.444513,13.082257,9.6984625,5.0576415,6.2884107,6.4722056,4.640821,3.43959,3.7054362,4.4964104,4.778667,3.4560003,2.5764105,2.8882053,3.8498464,2.9013336,2.0644104,1.7723079,2.1169233,2.8717952,3.4231799,3.0949745,2.5173335,2.1497438,2.2777438,2.4385643,2.2449234,2.225231,2.5698464,3.1409233,2.4320002,1.8215386,2.6715899,5.152821,8.251078,8.172308,5.930667,4.010667,3.1638978,2.412308,1.8281027,1.5360001,1.6410258,2.0020514,2.231795,1.9495386,1.9331284,2.0217438,1.9922053,1.5327181,5.7403083,10.036513,9.764103,5.7140517,4.138667,3.3247182,3.4888208,4.2469745,4.6276927,3.1015387,3.259077,8.576,12.609642,12.337232,8.155898,8.132924,10.765129,11.946668,11.178667,11.552821,12.12718,10.174359,7.4404106,6.2063594,9.301334,10.515693,9.82318,9.383386,9.127385,6.764308,7.830975,8.707283,7.8408213,6.121026,6.8594875,6.73477,6.163693,6.8496413,10.617436,19.429745,17.716515,14.401642,10.279386,6.921847,6.672411,5.8256416,5.421949,4.857436,4.417641,5.277539,6.498462,9.035488,10.013539,9.094564,8.484103,6.7610264,7.4141545,8.946873,10.223591,10.436924,10.919386,13.51877,15.261539,15.698052,16.899282,17.513027,18.018463,20.535797,24.937027,28.845951,28.468515,26.512413,23.207386,19.666052,17.8839,21.622156,24.546463,26.0759,26.896412,28.944412,29.321848,23.673437,20.109129,21.819078,27.083488,22.659285,25.219284,25.80677,20.59159,10.870154,12.649027,11.227899,8.868103,6.8233852,5.35959,4.7294364,4.630975,4.781949,5.0510774,5.4613338,5.3005133,5.431795,5.3694363,5.028103,4.709744,5.3825645,5.7074876,6.567385,8.116513,9.800206,13.088821,15.671796,16.275694,15.776822,17.23077,13.965129,14.55918,17.506462,21.001848,22.918566,24.01149,22.994053,21.126566,19.14749,17.286566,15.589745,11.772718,9.865847,10.840616,12.612924,12.829539,12.012309,11.063796,10.240001,9.156924,8.726975,8.507077,10.230155,15.451899,25.544207,26.95549,23.70954,19.373951,15.694771,12.593232,13.774771,13.397334,13.948719,17.066668,23.529028,28.310976,34.353233,37.74359,37.123283,33.690258,29.289028,23.460104,19.685745,19.032618,20.158361,28.737642,35.144207,37.120003,34.514053,29.252926,26.5879,24.802464,23.93272,24.1559,25.813335,26.187489,27.264002,27.336206,26.207182,25.19631,29.630362,31.77354,30.880823,28.209232,27.008001,24.352823,24.612104,26.673233,29.154465,30.375387,29.952002,29.013336,28.196104,28.09436,29.266054,28.278156,28.658875,30.306463,33.060104,36.716312,39.96554,36.952618,32.40698,30.191591,33.30954,41.40636,49.14216,57.2718,65.404724,72.00821,67.45929,66.3598,68.21744,73.86913,85.500725,103.279594,110.175186,105.79693,95.56678,90.706055,90.584625,87.5356,79.75385,70.331085,67.28206,64.80411,61.81416,58.210464,54.226055,50.39262,46.10626,42.824207,40.966568,39.998363,38.46236,38.127594,37.953644,37.02154,35.157337,32.938667,30.70031,26.564924,21.930668,17.8839,15.222155,14.027489,13.138052,12.2387705,11.241027,10.276103,9.409642,8.070564,6.7117953,5.5729237,4.6539493,3.7152824,2.7470772,1.8609232,1.1585642,0.7187693,0.4660513,0.2855385,0.17066668,0.12471796,0.14112821,0.15097436,0.18379489,0.23630771,0.34789747,0.6104616,0.7778462,0.85005134,1.6180514,3.5577438,6.810257,10.033232,10.394258,9.737847,9.872411,12.57354,12.662155,8.080411,3.8071797,2.5337439,4.647385,5.093744,5.4449234,5.805949,6.045539,5.8092313,2.7175386,1.1060513,0.4135385,0.18051283,0.04594872,0.013128206,0.009846155,0.013128206,0.013128206,0.0,0.0,0.006564103,0.013128206,0.052512825,0.20676924,1.3883078,1.723077,1.657436,1.3653334,0.7515898,0.98133343,1.3095386,1.2012309,0.65641034,0.23302566,0.30851284,0.3446154,0.33805132,0.31507695,0.3314872,0.5513847,0.7450257,0.90584624,0.99774367,0.9747693,0.9353847,0.9189744,0.94523084,0.9485129,0.76800007,0.5513847,0.39384618,0.27569234,0.18707694,0.128,0.14112821,0.16410258,0.17394873,0.16082053,0.13456412,0.1148718,0.08533334,0.08205129,0.108307704,0.14769232,0.19364104,0.21989745,0.24287182,0.24615386,0.18707694,0.07548718,0.03938462,0.029538464,0.029538464,0.026256412,0.026256412,0.036102567,0.04266667,0.04266667,0.04266667,0.04266667,0.04594872,0.04594872,0.04594872,0.04594872,0.032820515,0.029538464,0.029538464,0.032820515,0.04266667,0.032820515,0.055794876,0.09189744,0.12143591,0.12471796,0.15753847,0.24287182,0.380718,0.5218462,0.57764107,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.026256412,0.026256412,0.0,0.0,2.3302567,4.0402055,4.338872,3.692308,3.8137438,3.436308,4.2469745,7.5552826,11.07036,8.910769,3.9680004,3.373949,5.037949,6.413129,4.4701543,4.007385,3.121231,2.7864618,3.495385,5.2644105,7.0465646,8.15918,9.462154,11.72677,15.671796,17.283283,16.275694,13.522053,10.614155,9.856001,10.102155,9.238976,7.637334,5.9503593,5.097026,5.3760004,5.4580517,5.4153852,5.3398976,5.3398976,4.9854364,4.073026,3.1474874,2.5304618,2.3335385,1.4178462,1.0699488,1.6377437,2.7634873,3.370667,2.3236926,1.7591796,1.3915899,1.1716924,1.2832822,0.892718,0.702359,0.90256417,1.3259488,1.4506668,0.86317956,0.892718,1.4572309,2.2514873,2.7175386,1.7165129,1.6114873,1.8248206,1.8871796,1.4342566,1.5819489,1.7263591,1.9462565,2.103795,1.847795,1.2471796,1.0535386,1.0469744,0.9944616,0.64000005,0.33476925,0.24943592,0.35446155,0.56123084,0.7318975,1.4998976,1.8674873,1.7099489,1.3259488,1.4342566,1.2635899,0.73517954,0.43651286,0.571077,0.9616411,1.7066668,1.5458462,1.3423591,1.3653334,1.2668719,1.0601027,2.4910772,2.9669745,1.913436,0.7778462,0.9353847,1.0305642,0.94523084,0.77456415,0.82379496,0.6892308,0.8041026,1.0043077,1.083077,0.7778462,0.8992821,0.86646163,0.8172308,1.079795,2.166154,6.7314878,7.177847,5.8847184,4.706462,4.97559,6.3277955,5.0838976,3.1803079,2.1398976,3.0687182,4.6769233,4.588308,4.0434875,4.07959,5.5072823,4.9821544,4.768821,6.2096415,9.304616,12.711386,12.941129,11.188514,8.457847,5.9995904,5.280821,4.7917953,5.868308,6.485334,6.73477,8.835282,9.199591,6.820103,5.5893335,6.7872825,9.094564,9.193027,8.648206,6.8496413,5.0051284,6.163693,8.362667,12.06154,13.725539,12.186257,8.621949,6.0816417,6.308103,7.765334,9.222565,9.734565,10.28595,9.442462,8.854975,9.061745,9.475283,7.939283,7.899898,7.79159,7.171283,6.744616,4.9854364,5.159385,6.1374364,7.3091288,8.5891285,7.906462,6.7117953,7.1680007,10.023385,14.601848,10.57477,7.7357955,6.5837955,6.6395903,6.4689236,7.1154876,6.3901544,5.504,4.9952826,4.716308,3.9220517,3.82359,4.31918,4.8771286,4.5456414,3.7776413,4.2272825,5.674667,7.141744,6.8955903,6.675693,7.2631803,6.8529234,5.533539,5.2644105,5.1298466,5.32677,5.904411,6.088206,4.2568207,4.1846156,5.3727183,7.1089234,7.788308,4.9427695,4.955898,4.017231,2.9407182,2.15959,1.7099489,1.7329233,2.3893335,3.4625645,4.420923,4.4110775,6.9743595,5.6451287,3.8465643,3.259077,3.8465643,5.5532312,5.7534366,4.9329233,4.128821,4.896821,5.044513,4.788513,4.8049235,5.402257,6.498462,4.4373336,2.612513,1.4572309,1.2603078,2.1530259,2.7634873,3.0326157,2.9801028,2.7044106,2.412308,2.8258464,3.0752823,2.9538465,2.6026669,2.5173335,2.1530259,2.1333334,3.3476925,5.3234878,6.226052,3.5774362,2.6486156,2.3794873,2.2153847,2.1070771,2.0217438,2.4385643,3.2131286,3.5872824,2.1825643,1.8510771,3.3542566,4.414359,3.9844105,2.228513,4.4734364,7.8539495,8.832001,7.056411,5.3694363,6.5312824,6.6100516,6.5050263,5.933949,3.4166157,4.7491283,10.052924,13.860104,13.942155,11.306667,8.891078,10.052924,11.670976,11.808822,9.734565,7.427283,8.15918,8.03118,6.5903597,6.8365135,7.384616,9.38995,9.878975,9.012513,10.085744,11.85477,8.598975,6.738052,7.3616414,6.226052,6.921847,5.2742567,3.9318976,4.709744,8.592411,10.518975,7.000616,3.6069746,2.740513,3.6332312,5.366154,4.2863593,2.9997952,2.409026,1.723077,2.7011285,3.239385,3.5610259,4.1156926,5.5532312,7.200821,8.766359,11.293539,13.6467705,12.511181,8.326565,8.651488,12.100924,15.872002,15.763694,17.42113,23.256617,29.006771,31.77354,30.030771,27.85477,28.393028,27.959797,25.793644,24.047592,26.63713,28.389746,26.791388,21.960207,16.662975,19.140924,19.429745,20.25354,22.078362,23.11877,17.59836,14.336001,10.873437,7.453539,6.987488,8.697436,4.857436,1.5031796,0.9156924,1.6475899,2.0644104,1.5524104,1.2603078,1.6508719,2.5173335,4.263385,5.917539,6.5870776,6.196513,5.477744,4.7458467,4.397949,5.0018463,6.7117953,9.26195,11.155693,12.022155,11.588924,10.614155,10.896411,11.224616,10.548513,10.791386,11.933539,11.992617,11.884309,9.393231,7.0859494,5.970052,5.4941545,4.8836927,4.125539,4.132103,5.1167183,6.6067696,6.0816417,6.6100516,7.282872,7.6077952,7.522462,8.730257,8.034462,8.621949,13.203693,24.018053,23.30913,22.94154,20.578463,16.452925,13.351386,16.121437,19.498669,23.384617,27.02113,28.960823,30.9399,30.116104,28.809849,28.3799,29.220104,23.630772,20.33559,17.161848,14.260514,14.116103,23.525745,28.386463,29.80431,28.767181,26.154669,23.712822,22.52472,21.730463,21.270975,21.881437,23.860516,26.706053,27.480618,26.551796,27.588924,31.458464,37.185642,35.262363,26.899694,24.018053,19.19672,15.593027,14.605129,16.032822,18.084105,18.950565,19.065437,19.10154,19.830154,22.12431,24.359386,26.016823,26.896412,26.535387,24.218258,26.010258,22.816822,19.446156,18.737232,21.530258,28.954258,35.93518,42.423798,46.982567,46.802055,42.85703,38.915283,39.525745,46.828312,60.547287,74.24657,81.28657,87.6078,94.637955,99.28862,102.04555,91.897446,80.73518,75.77929,79.57334,89.3637,93.42032,91.84493,86.43939,80.70236,72.402054,65.84123,60.274876,54.321236,45.95857,44.373337,43.966362,44.04513,43.4478,40.543182,37.953644,33.378464,27.556105,21.704206,17.51631,16.039387,15.376411,14.693745,13.755078,12.924719,12.458668,11.116308,9.603283,8.2904625,7.2172313,5.802667,4.5128207,3.2328207,2.038154,1.2209232,0.7318975,0.4266667,0.24943592,0.16410258,0.15097436,0.16410258,0.23958977,0.39384618,0.49887183,0.3052308,0.318359,0.38400003,0.8172308,1.9626669,4.197744,6.6002054,6.73477,9.019077,13.013334,13.426873,12.609642,7.2894363,3.3575387,3.4264617,6.820103,11.152411,14.168616,14.76595,12.681848,8.484103,4.0041027,1.5458462,0.47917953,0.18051283,0.04594872,0.02297436,0.006564103,0.006564103,0.013128206,0.0,0.0,0.0,0.0,0.098461546,0.48902568,3.3575387,3.1507695,1.8248206,0.7515898,0.702359,1.214359,1.8642052,1.9987694,1.4408206,0.48902568,0.23302566,0.14112821,0.13456412,0.16082053,0.19692309,0.2100513,0.25928208,0.30194873,0.3511795,0.47261542,0.48574364,0.63343596,0.8598975,1.1093334,1.3423591,1.1848207,0.84348726,0.54482055,0.36102566,0.21333335,0.17723078,0.12143591,0.098461546,0.108307704,0.12143591,0.17066668,0.13784617,0.0951795,0.08533334,0.12143591,0.20676924,0.20020515,0.190359,0.18707694,0.13784617,0.07548718,0.04266667,0.029538464,0.026256412,0.016410258,0.016410258,0.02297436,0.029538464,0.029538464,0.029538464,0.029538464,0.03938462,0.04594872,0.04594872,0.04594872,0.032820515,0.029538464,0.029538464,0.029538464,0.029538464,0.029538464,0.049230773,0.06235898,0.06564103,0.07548718,0.13784617,0.25271797,0.40697438,0.5284103,0.5021539,0.098461546,0.01969231,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.032820515,0.068923086,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.006564103,0.37743592,1.8904617,6.626462,6.744616,4.394667,2.4976413,4.7655387,6.232616,4.9952826,4.9296412,6.498462,6.738052,5.3398976,4.384821,3.511795,2.5140514,1.332513,1.1815386,1.086359,1.5064616,2.793026,5.179077,7.722667,8.5202055,9.32759,11.047385,13.728822,14.647796,13.833847,12.107488,10.292514,9.222565,8.802463,7.9491286,6.892308,5.9569235,5.5597954,5.536821,5.717334,5.8945646,5.9667697,5.927385,5.796103,5.152821,3.698872,2.103795,2.0184617,2.4681027,1.591795,1.2471796,2.0020514,3.1409233,3.0391798,4.132103,5.1265645,5.1954875,3.9680004,1.7394873,1.1881026,0.97805136,0.67938465,0.7417436,0.7811283,0.8763078,0.96492314,1.0043077,0.9714873,1.1913847,1.719795,1.6968206,1.0699488,0.6301539,1.467077,2.5632823,3.0129232,2.6322052,1.9561027,1.2209232,1.1093334,1.1126155,0.9616411,0.6301539,0.5677949,0.6235898,0.6892308,0.7384616,0.84348726,1.3292309,1.8871796,2.103795,1.9265642,1.654154,1.6016412,1.2471796,1.1355898,1.332513,1.4506668,1.3161026,1.1815386,1.1618463,1.1520001,0.8402052,0.6695385,1.4244103,1.7788719,1.4080001,0.98461545,0.8795898,0.9517949,0.90584624,0.7384616,0.7384616,0.7220513,0.827077,1.017436,1.148718,0.9616411,1.0633847,0.9156924,0.7844103,0.9189744,1.5556924,3.8564105,4.562052,4.3716927,4.128821,4.8147697,7.312411,7.650462,6.557539,5.0116925,4.240411,3.8596926,3.5840003,4.2863593,5.677949,6.3277955,6.7577443,6.8430777,7.3649235,8.592411,10.269539,9.416205,7.7292314,5.5138464,3.9745643,5.2053337,6.1440005,7.6143594,7.351795,5.504,4.6244106,5.976616,5.225026,5.0051284,6.0750775,7.3485136,5.796103,4.7228723,4.017231,3.8367183,4.6276927,6.921847,10.738873,14.27036,15.9573345,14.49354,10.8307705,9.091283,8.923898,9.189744,7.965539,7.39118,7.397744,8.218257,9.642668,11.0145645,9.173334,8.283898,8.116513,8.277334,8.2215395,7.1876926,7.0137444,7.174565,7.53559,8.3593855,7.4010262,5.5302567,5.333334,7.5454364,11.0375395,7.975385,5.8190775,5.297231,5.9602056,6.189949,6.2785645,5.7796926,4.9394875,4.3618464,5.0215387,5.5072823,5.9995904,7.748924,10.210463,11.053949,6.2227697,5.4941545,6.124308,6.770872,7.496206,5.8880005,6.114462,6.432821,6.419693,6.961231,5.7731285,4.210872,5.0477953,7.2664623,6.052103,3.4198978,3.6036925,4.7228723,5.3431797,4.493129,5.4613338,5.1856413,5.72718,6.8562055,6.055385,4.5554876,3.8432825,3.757949,3.9351797,3.7874875,3.56759,2.6354873,1.8838975,1.8707694,2.806154,4.6145644,5.723898,5.536821,4.4340515,3.7874875,4.568616,5.2315903,5.2611284,5.074052,6.0356927,4.33559,2.9669745,2.2088206,2.044718,2.162872,2.228513,1.9364104,1.9167181,2.231795,2.3860514,2.5074873,2.540308,2.422154,2.28759,2.4582565,2.5796926,3.4658465,3.9187696,3.9056413,4.565334,4.640821,4.4898467,4.4110775,4.3552823,3.9253337,4.06318,4.1189747,3.9056413,3.2623591,2.0709746,2.3269746,2.8192823,3.045744,2.6715899,1.5195899,1.9593848,2.5600002,2.6617439,2.2646155,2.0250258,2.8455386,3.8137438,5.730462,7.5618467,6.432821,4.923077,8.937026,11.881026,11.431385,9.537642,8.067283,7.1876926,7.7718983,9.373539,10.246565,8.027898,7.8834877,7.515898,6.5805135,6.688821,6.5345645,5.720616,6.5837955,8.27077,6.7183595,5.5171285,6.0980515,7.2631803,7.6898465,5.920821,6.2063594,7.837539,7.7456417,6.058667,6.11118,7.788308,6.997334,7.5191803,10.312206,13.505642,11.237744,13.272616,15.058052,14.519796,12.087796,10.066052,6.889026,5.106872,5.8518977,8.825437,10.765129,11.877745,11.392001,9.77395,8.717129,10.955488,14.060308,15.924514,15.858873,14.565744,13.052719,18.25477,23.867079,26.899694,27.67426,27.385439,30.831593,32.308514,29.216824,22.071796,20.233849,20.795078,22.610052,24.385643,24.681028,20.900105,17.78872,17.23077,18.825848,19.882668,16.006565,14.263796,11.753027,8.641642,8.149334,6.75118,3.748103,1.654154,1.1552821,1.086359,1.0535386,0.8763078,1.2668719,2.228513,3.05559,2.993231,2.9735386,2.9013336,2.8455386,3.0260515,2.2613335,2.3991797,3.2656412,4.3585644,4.8311796,7.571693,9.947898,10.548513,9.970873,10.807796,11.539693,10.604308,10.368001,11.076924,10.834052,9.6,7.50277,6.042257,5.7534366,6.2129235,6.432821,6.770872,8.891078,11.808822,11.890873,11.053949,9.997129,8.579283,6.9743595,5.677949,7.463385,7.0498466,6.8463597,9.07159,15.766975,20.164925,22.793848,21.622156,17.841232,15.852309,14.483693,15.212309,15.921232,16.006565,16.36431,16.672821,16.344616,16.15754,16.190361,15.829334,15.366566,14.372104,13.781334,14.057027,15.199181,16.292105,17.857643,19.035898,20.903387,26.482874,29.042873,28.297848,25.094566,21.313643,19.90236,19.908924,20.26995,19.80718,19.157335,20.801643,23.479797,26.148104,26.742155,24.937027,22.17354,17.174976,12.58995,10.771693,11.825232,13.6008215,15.064616,16.46277,17.27672,17.591797,18.110361,19.22954,20.588308,21.760002,22.032412,20.407797,20.424206,19.347694,18.336823,17.864206,17.723078,19.695591,22.583797,25.03877,26.476309,27.073643,26.38113,26.377848,27.818668,31.806362,39.794876,45.357952,52.78195,61.68944,71.135185,79.625854,83.370674,79.85888,74.555084,72.3397,77.52534,91.211494,101.07734,108.64575,112.8796,110.168625,98.254776,90.1317,83.400215,75.57909,64.12144,55.778465,51.741543,50.103798,48.29867,43.119595,42.29908,39.138466,34.3598,29.30872,25.951181,25.32431,24.01149,22.262156,19.682463,15.232001,14.14236,12.832822,11.552821,10.420513,9.412924,8.155898,6.685539,5.1954875,3.817026,2.6486156,1.719795,1.0568206,0.636718,0.40697438,0.2855385,0.16082053,0.17394873,0.26912823,0.33805132,0.21989745,0.21333335,0.3249231,0.8467693,2.3926156,5.917539,10.8996935,11.401847,11.080206,10.834052,8.789334,6.944821,4.59159,3.3411283,4.086154,6.99077,12.593232,17.67713,19.006361,15.547078,8.448001,3.7316926,1.4145643,0.46933338,0.16082053,0.04594872,0.02297436,0.006564103,0.009846155,0.02297436,0.0,0.0,0.0,0.0,0.06235898,0.318359,1.3587693,1.5163078,1.4867693,1.6869745,2.2646155,1.9954873,1.7394873,1.9922053,2.540308,2.477949,2.6420515,2.3926156,2.0184617,1.6278975,1.1257436,0.6301539,0.3314872,0.21989745,0.24287182,0.3249231,0.4660513,0.64000005,0.761436,0.8402052,0.96492314,1.148718,1.1979488,1.1716924,1.024,0.60389745,0.36102566,0.24287182,0.16738462,0.11158975,0.08533334,0.0951795,0.0951795,0.08205129,0.06235898,0.06235898,0.07876924,0.09189744,0.0951795,0.09189744,0.101743594,0.08861539,0.059076928,0.03938462,0.032820515,0.03938462,0.049230773,0.052512825,0.04594872,0.029538464,0.029538464,0.029538464,0.032820515,0.032820515,0.036102567,0.04594872,0.032820515,0.029538464,0.029538464,0.029538464,0.01969231,0.029538464,0.04266667,0.049230773,0.055794876,0.07548718,0.108307704,0.15753847,0.21661541,0.25928208,0.23630771,0.049230773,0.06235898,0.026256412,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016410258,0.032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.16410258,0.92225647,2.9702566,8.67118,7.752206,4.1485133,1.522872,3.2853336,4.59159,3.7973337,3.373949,4.44718,6.7905645,4.6966157,4.650667,4.141949,2.678154,1.785436,1.3981539,0.9944616,1.3751796,2.8882053,5.4416413,7.5618467,9.032206,10.666668,12.317539,12.905026,12.859077,12.137027,10.794667,9.206155,8.067283,8.562873,8.4053335,7.830975,7.1614366,6.7840004,6.370462,6.304821,6.482052,6.672411,6.51159,6.226052,5.910975,4.391385,2.2514873,1.8084104,2.3171284,1.8773335,1.5524104,2.0512822,3.7218463,5.7042055,6.3540516,5.474462,3.8038976,3.0194874,2.281026,1.6640002,1.0568206,0.5874872,0.60061544,0.56123084,0.60389745,1.1651284,2.0020514,2.2186668,2.0611284,2.0217438,1.6246156,0.9517949,0.6301539,1.1454359,1.782154,2.231795,2.2744617,1.7723079,1.4276924,1.2996924,1.332513,1.3817437,1.2209232,1.6311796,1.6935385,1.7362052,1.6475899,0.8598975,1.020718,1.4408206,1.7165129,1.7362052,1.6902566,1.782154,1.6246156,1.5031796,1.4408206,1.204513,1.1881026,1.1913847,1.3193847,1.4375386,1.1913847,0.8402052,1.276718,1.4375386,1.2570257,1.6869745,2.1398976,1.9790771,1.5163078,1.0075898,0.6432821,1.1979488,1.4145643,1.5622566,1.595077,1.1815386,1.0502565,1.0994873,1.1158975,1.1355898,1.404718,2.5435898,3.5314875,4.2207184,4.5423594,4.5029745,5.835488,7.171283,7.1909747,6.009436,5.172513,5.280821,5.5565133,6.048821,6.6461544,7.0531287,6.918565,6.557539,5.8945646,5.35959,5.8880005,5.6352825,5.07077,4.06318,3.43959,4.9854364,6.229334,7.6143594,6.997334,4.70318,3.5347695,6.245744,6.8955903,6.5280004,6.1013336,6.5017443,5.654975,4.9985647,4.4964104,4.352,5.0116925,6.0619493,8.100103,11.52,15.199181,16.49231,14.299898,11.0605135,8.910769,7.9294367,6.157129,5.5236926,5.87159,6.705231,7.9491286,9.970873,9.399796,8.851693,8.769642,8.815591,7.8408213,7.79159,7.39118,7.020308,6.774154,6.47877,6.5017443,6.0061545,5.9930263,6.9349747,8.766359,7.571693,6.4032826,5.979898,6.2720003,6.4754877,5.8912826,4.965744,4.2305646,4.027077,4.493129,6.3310776,6.872616,7.026872,7.466667,8.615385,6.892308,5.8453336,5.910975,6.8299494,7.6635904,5.7534366,5.651693,5.651693,5.366154,5.737026,4.5029745,3.3280003,4.312616,6.7314878,7.003898,4.516103,4.0303593,4.0303593,3.9844105,4.332308,7.276308,7.4797955,6.885744,6.180103,4.8082056,4.023795,4.0402055,4.06318,3.879385,3.8432825,3.0818465,3.05559,2.865231,2.5238976,2.934154,4.141949,5.7107697,5.796103,4.384821,3.3280003,4.332308,4.896821,4.5390773,3.7907696,4.197744,3.4166157,2.9407182,2.6256413,2.359795,2.0742567,2.044718,1.8182565,1.8018463,1.9495386,1.7591796,1.719795,1.8740515,1.9856411,2.041436,2.2678976,2.9210258,3.8367183,4.1156926,4.073026,5.211898,5.1922054,5.3825645,5.3727183,5.0018463,4.342154,4.5456414,4.309334,3.761231,3.131077,2.7602053,2.297436,2.281026,2.412308,2.4484105,2.1956925,2.3729234,2.0053334,1.5458462,1.3161026,1.5097437,3.3411283,7.8145647,11.943385,13.075693,8.917334,5.2315903,6.6002054,7.397744,6.373744,6.678975,7.7456417,6.8660517,7.181129,10.243283,16.01641,13.620514,11.047385,9.074872,7.5421543,5.3431797,5.139693,4.352,4.903385,6.665847,7.456821,5.612308,5.6352825,6.5083084,7.1187696,6.265436,6.2785645,7.499488,7.315693,5.5762057,4.578462,4.95918,4.2502565,4.95918,7.5552826,10.456616,9.616411,12.491488,15.396104,15.990155,13.259488,9.82318,7.3550773,6.8397956,7.906462,8.838565,11.621744,13.50236,11.667693,8.093539,9.55077,9.091283,12.232206,14.628103,15.100719,15.632411,11.999181,15.16636,19.321438,21.523693,21.720617,21.382566,24.641644,26.98831,24.979694,16.249437,17.457232,18.313848,18.86195,18.763489,17.302977,14.191591,14.027489,16.177233,18.225233,15.960617,13.344822,13.249642,13.321847,12.629334,11.661129,10.453334,6.048821,2.409026,1.1651284,1.6147693,1.4736412,1.6147693,1.6804104,1.7165129,2.1825643,2.1891284,2.4451284,2.3466668,1.8806155,1.6311796,1.5885129,1.9396925,2.2613335,2.2678976,1.8018463,3.5183592,4.926359,5.622154,6.1341543,7.9327188,9.202872,9.32759,9.813334,10.81436,11.113027,9.728001,9.032206,8.470975,7.890052,7.5388722,8.096821,8.684308,11.71036,15.937642,16.472616,14.693745,12.363488,10.276103,9.032206,9.035488,9.616411,8.533334,7.9950776,8.592411,9.291488,13.141335,16.131283,16.443079,14.290052,11.884309,8.996103,8.28718,8.054154,7.64718,7.50277,7.574975,7.824411,8.51036,9.373539,9.642668,10.768411,11.201642,11.119591,10.778257,10.528821,10.44677,14.900514,23.555285,33.857643,41.00267,37.077335,29.696003,22.738052,18.372925,17.066668,16.49559,16.469334,16.160822,15.829334,16.833643,17.42113,18.326975,19.094976,18.70113,15.53395,10.909539,8.293744,7.722667,8.73354,10.338462,11.539693,13.164309,14.483693,15.232001,15.61272,16.390566,17.588514,18.62236,19.006361,18.376207,17.480206,16.705643,16.580925,16.955078,17.007591,16.827078,17.165129,17.716515,18.33354,19.009642,19.380514,20.660515,22.419695,24.477541,26.90954,29.367798,33.536003,38.623184,44.47508,51.61026,56.98626,60.04185,63.72431,70.26872,81.19467,91.98934,104.36596,114.93745,121.33088,122.1875,115.222984,110.20801,105.78052,98.97026,85.21519,63.36657,52.42421,47.090874,44.90503,46.208004,49.532722,53.454773,57.99713,61.026466,58.243286,45.14134,34.43857,27.329643,22.695387,17.06995,14.982565,13.610668,12.547283,11.592206,10.752001,9.757539,8.480822,7.1122055,5.7698464,4.4898467,3.4822567,2.5961027,1.8871796,1.3522053,0.9353847,0.60061544,0.48246157,0.48574364,0.5218462,0.48246157,0.39056414,0.45620516,1.142154,3.1638978,7.4929237,12.422565,13.131488,11.61518,9.271795,6.889026,6.685539,7.2205133,7.7981544,7.890052,7.145026,9.842873,12.504617,13.078976,10.834052,6.377026,2.477949,0.88943595,0.34133336,0.108307704,0.036102567,0.013128206,0.0032820515,0.0032820515,0.009846155,0.0,0.0,0.0,0.0,0.04266667,0.21989745,0.5349744,0.67610264,1.079795,1.7690258,2.3696413,1.6443079,1.0666667,1.1881026,1.9331284,2.6289232,3.754667,4.4340515,4.5423594,4.2436924,4.0041027,4.164923,3.1737437,1.7788719,0.6170257,0.19692309,0.28225642,0.42338464,0.574359,0.69907695,0.761436,1.0666667,1.4473847,1.6771283,1.6246156,1.270154,0.97805136,0.90584624,0.8533334,0.69251287,0.3708718,0.19364104,0.1148718,0.07876924,0.059076928,0.04594872,0.04594872,0.049230773,0.04594872,0.04594872,0.055794876,0.06235898,0.068923086,0.07548718,0.07876924,0.08205129,0.21989745,0.24615386,0.19692309,0.118153855,0.0951795,0.059076928,0.03938462,0.029538464,0.032820515,0.036102567,0.032820515,0.036102567,0.03938462,0.03938462,0.04266667,0.049230773,0.04594872,0.04266667,0.03938462,0.059076928,0.08205129,0.08861539,0.098461546,0.1148718,0.10502565,0.0,0.052512825,0.026256412,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.049230773,0.22646156,0.827077,2.3335385,8.470975,7.4797955,4.194462,2.3729234,4.673641,5.435077,4.4077954,3.9876926,4.8804107,6.0816417,5.182359,4.5423594,3.8301542,3.058872,2.553436,1.9561027,1.1979488,1.4112822,3.0752823,6.038975,7.4010262,9.426052,11.697231,13.2562065,12.593232,11.595488,10.420513,9.107693,7.9852314,7.650462,8.608821,8.835282,8.720411,8.539898,8.480822,7.962257,7.506052,7.2631803,7.194257,7.0498466,6.9743595,6.75118,5.5729237,3.6857438,2.3958976,2.169436,1.9429746,1.8445129,2.1136413,3.1113849,5.297231,5.546667,4.023795,2.028308,1.9790771,2.3893335,1.8773335,1.2340513,0.8730257,0.827077,0.5152821,0.6235898,1.4244103,2.409026,2.2908719,1.6968206,1.3456411,1.0371283,0.73517954,0.5546667,0.7778462,0.90912825,1.2832822,1.7624617,1.7362052,1.7099489,1.8904617,2.03159,1.9659488,1.5983591,2.3204105,2.4155898,2.297436,1.9954873,1.142154,1.0502565,1.2012309,1.3522053,1.394872,1.3554872,1.6475899,1.7329233,1.8379488,1.9003079,1.5655385,1.6180514,1.5360001,1.6082052,1.6508719,1.0010257,0.8992821,1.3128207,1.3423591,1.1257436,1.8281027,2.300718,2.03159,1.4867693,0.9878975,0.7220513,1.5753847,1.8149745,1.8642052,1.8346668,1.5425643,1.3423591,1.4375386,1.5753847,1.7329233,2.1300514,2.6157951,3.564308,4.8607183,5.87159,5.428513,5.1200004,7.0432825,8.349539,7.830975,5.924103,6.0225644,6.091488,5.9602056,5.8486156,6.370462,5.930667,5.5236926,5.146257,5.4416413,7.6931286,4.9427695,4.9952826,5.7796926,6.363898,6.9382567,6.770872,6.8529234,6.193231,4.8705645,4.0336413,6.928411,7.6570263,7.128616,6.189949,5.6287184,5.5236926,5.5565133,4.824616,3.757949,4.096,4.640821,5.034667,6.892308,10.151385,13.08554,13.574565,10.594462,7.5552826,5.658257,3.895795,3.751385,4.378257,5.3136415,6.5050263,8.297027,8.421744,8.576,8.507077,7.9228725,6.47877,6.997334,7.3649235,7.702975,7.6176414,6.2030773,5.72718,5.865026,6.121026,6.554257,7.752206,8.109949,7.6931286,7.2336416,6.99077,6.764308,5.4383593,4.8738465,5.3760004,6.432821,6.7117953,7.39118,6.7150774,5.4843082,4.634257,5.2512827,6.5706673,6.2490263,6.160411,6.8365135,7.466667,5.9503593,5.284103,4.7228723,4.2929235,4.8147697,4.017231,3.387077,3.7120004,5.0051284,6.491898,6.121026,5.225026,4.1091285,3.626667,5.175795,9.193027,8.4972315,6.189949,4.1058464,2.8356924,3.3444104,4.138667,4.263385,3.8400004,4.066462,3.9318976,4.2305646,4.2207184,3.7809234,3.4100516,5.142975,6.488616,6.363898,5.1167183,4.516103,4.634257,4.1747694,3.3247182,2.550154,2.5993848,2.7208207,2.9078977,2.8488207,2.550154,2.3368206,2.7437952,2.6486156,2.3204105,1.8806155,1.3128207,1.1815386,1.4998976,1.8018463,1.9396925,2.0906668,2.7634873,3.3247182,3.8334363,4.342154,4.900103,4.164923,4.4800005,4.8836927,4.7556925,3.8432825,4.1911798,3.754667,3.2196925,2.9210258,2.8488207,2.3926156,2.2186668,2.3138463,2.6223593,3.0194874,3.0884104,2.5600002,1.8313848,1.4342566,2.028308,4.4996924,10.614155,15.028514,14.605129,8.418462,4.640821,4.7950773,4.71959,3.9942567,5.927385,7.394462,7.145026,8.241231,12.891898,22.465643,21.868309,16.764719,11.690667,8.093539,4.342154,3.9614363,4.352,5.093744,6.0947695,7.5913854,6.426257,5.651693,5.973334,6.7249236,5.8945646,5.9667697,5.920821,5.277539,4.2568207,3.7842054,3.95159,4.059898,4.312616,5.211898,7.5487185,9.645949,11.844924,13.279181,13.236514,11.16554,9.074872,9.793642,11.565949,12.652308,11.32636,13.778052,13.797745,11.437949,9.032206,11.204924,10.256411,10.971898,12.524308,14.194873,15.376411,12.750771,14.592001,16.534975,16.725334,15.816206,15.061335,17.050259,18.491077,17.158566,11.884309,14.677335,14.129231,12.422565,10.610872,8.63836,7.8473854,13.262771,18.628925,19.659489,14.03077,12.314258,12.084514,12.816411,13.184001,11.080206,9.4457445,5.3169236,2.1464617,1.1946667,1.5425643,1.5195899,1.9396925,1.8642052,1.2603078,0.98133343,1.270154,1.9987694,2.231795,1.7263591,0.9616411,1.079795,1.2964103,1.2931283,0.9682052,0.45292312,1.0338463,1.3883078,1.7624617,2.540308,4.269949,5.654975,7.000616,8.3593855,9.504821,9.921641,9.173334,9.708308,9.642668,8.503796,7.207385,8.342975,9.193027,11.602052,15.281232,17.811693,17.240616,15.094155,13.059283,12.324103,13.587693,11.050668,8.04759,6.76759,7.017026,6.226052,8.28718,10.174359,10.509129,9.028924,6.6100516,4.414359,3.8104618,3.9384618,4.1222568,3.892513,4.020513,4.529231,5.2742567,6.0717955,6.7150774,8.297027,9.298052,9.140513,8.083693,7.197539,8.864821,15.24513,25.787079,36.309338,39.02031,32.712208,24.159182,17.769028,14.900514,13.856822,12.993642,13.308719,13.797745,14.024206,14.099693,13.692719,14.020925,14.129231,12.947693,9.284924,6.0816417,5.6320004,6.3376417,7.466667,9.16677,9.803488,10.873437,12.032001,13.036308,13.768207,14.263796,14.907078,15.524104,16.091898,16.764719,16.932104,16.984617,17.59836,18.891489,20.417643,19.531488,17.45395,15.842463,15.330462,15.51754,16.31836,17.575386,18.898052,19.984411,20.608002,22.885746,25.291489,27.90072,30.838156,34.254772,39.67344,44.639183,51.36739,60.849236,72.84842,81.273445,94.58872,105.885544,111.793236,112.51857,110.92678,110.7758,108.57683,100.703186,83.39365,58.15467,45.151184,39.59795,40.064003,48.469337,58.09231,69.08062,79.1598,83.41334,74.30565,49.99221,34.386055,25.993849,21.943796,17.985641,15.963899,14.749539,13.8075905,12.898462,12.074668,11.218052,10.131693,8.937026,7.7357955,6.5936418,5.7632823,5.0871797,4.4701543,3.7743592,2.8127182,1.8674873,1.3850257,1.1848207,1.0929232,0.92225647,0.7122052,0.8566154,1.6836925,3.5610259,6.8693337,9.537642,9.865847,8.704,7.1680007,6.6560006,9.035488,11.805539,13.39077,12.727796,9.281642,8.1066675,8.060719,7.5421543,6.038975,4.125539,1.4736412,0.5152821,0.21661541,0.059076928,0.02297436,0.0032820515,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0032820515,0.03938462,0.17723078,0.29538465,0.40369233,0.97805136,1.8313848,2.097231,1.0502565,0.55794877,0.7253334,1.5031796,2.674872,4.4701543,5.5893335,6.413129,7.7718983,10.935796,9.563898,6.4590774,3.3476925,1.2504616,0.4594872,0.3052308,0.26256412,0.33476925,0.4660513,0.5152821,0.83035904,1.6377437,2.3368206,2.6026669,2.3991797,1.9790771,1.7099489,1.4933335,1.2176411,0.75487185,0.43651286,0.2100513,0.09189744,0.059076928,0.052512825,0.04266667,0.032820515,0.029538464,0.026256412,0.036102567,0.059076928,0.09189744,0.1148718,0.128,0.14441027,0.29538465,0.31507695,0.256,0.20676924,0.30851284,0.27569234,0.17394873,0.118153855,0.118153855,0.07876924,0.068923086,0.07548718,0.14441027,0.24287182,0.24943592,0.21661541,0.14769232,0.098461546,0.08205129,0.07548718,0.08533334,0.07876924,0.068923086,0.068923086,0.072205134,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016410258,0.032820515,0.0,0.0,0.16738462,0.21333335,0.26256412,0.8763078,6.2227697,5.835488,4.342154,4.634257,7.8703594,7.719385,5.687795,4.8640003,5.2512827,3.757949,5.6418467,3.5577438,1.9593848,2.1366155,2.2055387,1.6804104,0.97805136,1.1782565,2.92759,6.432821,7.3321033,9.104411,11.063796,12.304411,11.697231,10.322052,8.684308,7.6012316,7.4141545,7.9852314,8.4283085,8.904206,9.619693,10.400822,10.66995,10.059488,9.212719,8.316719,7.5979495,7.322257,7.719385,7.4436927,6.741334,5.536821,3.4231799,2.297436,1.782154,1.7887181,2.0086155,1.9167181,2.3860514,2.6026669,2.2547693,1.6869745,1.8937438,1.913436,1.522872,1.1618463,0.99774367,0.92553854,0.52512825,0.7417436,1.1979488,1.3653334,0.574359,0.15425642,0.13456412,0.27241027,0.36102566,0.23302566,0.46276927,0.508718,0.761436,1.2603078,1.6869745,1.8707694,2.556718,2.7569232,2.2678976,1.6410258,2.172718,2.3040001,2.0611284,1.6738462,1.5983591,1.3883078,1.2209232,1.1946667,1.2406155,1.1060513,1.5524104,1.7624617,2.1103592,2.5074873,2.4024618,2.1070771,1.910154,1.9823592,1.8806155,0.56123084,0.92553854,1.1848207,1.1093334,0.93866676,1.404718,1.2307693,1.0043077,0.8008206,0.81066674,1.3292309,1.6968206,1.6902566,1.6607181,1.8149745,2.2186668,2.3794873,2.1792822,2.0841026,2.4024618,3.3017437,3.4034874,3.8990772,5.35959,7.131898,7.3386674,6.482052,8.418462,10.817642,11.191795,6.8955903,5.8847184,4.9854364,4.3290257,4.1583595,4.8311796,5.0838976,5.2742567,6.701949,9.810052,14.17518,6.806975,6.373744,8.930462,11.247591,10.7848215,7.75877,5.720616,4.9952826,5.159385,5.0215387,6.6100516,6.5772314,6.5411286,6.564103,5.142975,4.706462,5.0871797,4.06318,2.0118976,1.9462565,3.1638978,2.917744,2.7864618,3.826872,6.6034875,9.334154,8.205129,5.720616,3.4100516,1.8248206,2.2580514,3.1277952,4.647385,6.4557953,7.6307697,7.8539495,8.434873,7.9885135,6.491898,5.2578464,5.671385,7.581539,9.645949,10.43036,8.421744,5.835488,5.146257,5.32677,5.930667,7.1089234,8.155898,8.073847,7.637334,7.243488,6.9087186,5.4843082,5.7468724,8.018052,10.95877,11.54954,9.055181,6.436103,5.0018463,4.7622566,4.4438977,5.733744,6.2030773,6.0652313,5.796103,6.12759,5.7665644,4.906667,4.086154,3.9680004,5.333334,5.35959,5.1167183,4.204308,3.446154,4.8771286,7.243488,6.3376417,4.4767184,3.7415388,5.989744,9.03877,6.994052,4.315898,2.9965131,2.5731285,3.501949,4.4274874,4.2896414,3.5282054,4.059898,4.7360005,4.8049235,4.824616,4.7917953,4.1517954,7.194257,7.7259493,6.8496413,5.7796926,5.8453336,5.0215387,3.5872824,2.4582565,1.9692309,1.8904617,2.4320002,2.7306669,2.7503593,2.6518977,2.7995899,3.8859491,3.8071797,3.0227695,2.03159,1.394872,1.1881026,1.529436,1.847795,1.9528207,2.041436,2.3794873,2.6354873,3.3050258,3.9318976,3.1113849,2.2908719,2.737231,3.6693337,4.1517954,3.0752823,3.4822567,3.131077,2.7995899,2.6584618,2.2711797,2.8258464,2.4910772,2.3040001,2.6256413,3.1540515,3.006359,2.6978464,2.100513,1.719795,2.674872,4.3618464,8.536616,10.962052,9.688616,5.044513,3.3312824,4.066462,4.532513,4.5029745,6.2523084,6.3606157,7.207385,9.796924,15.875283,27.930258,29.797747,22.367182,13.768207,7.8441033,4.1682053,3.7218463,5.4580517,7.1614366,7.512616,6.11118,5.907693,6.048821,6.701949,6.994052,5.0215387,4.9460516,4.2305646,3.43959,2.9997952,3.1770258,4.604718,7.3682055,8.050873,6.961231,8.116513,11.188514,12.1238985,11.536411,10.14154,8.736821,9.284924,12.678565,15.707899,16.57436,14.903796,15.579899,12.041847,10.095591,11.286975,12.87877,15.140103,12.422565,11.625027,13.732103,13.820719,13.3940525,14.601848,14.8020525,13.640206,13.042872,12.064821,12.416001,11.687386,9.964309,9.819899,11.024411,8.996103,6.5969234,5.3366156,5.353026,6.6100516,16.918976,23.857233,22.3639,14.742975,12.803283,10.686359,10.06277,10.138257,7.6603084,3.6463592,1.657436,1.2865642,1.5885129,1.0765129,0.98133343,1.5327181,1.6738462,1.214359,0.8008206,0.5546667,1.204513,1.7460514,1.6607181,0.9124103,0.6235898,0.5481026,0.54482055,0.508718,0.36430773,0.5546667,0.85005134,0.9747693,1.0371283,1.5360001,2.4057438,4.125539,5.832206,7.0432825,7.64718,8.024616,9.019077,9.084719,8.0377445,7.0400004,8.792616,9.754257,10.6469755,12.770463,18.01518,20.539078,19.840002,18.008617,16.705643,17.155283,10.709334,5.504,3.3772311,4.197744,5.8453336,7.0957956,7.650462,7.056411,5.4974365,3.8104618,3.114667,3.5183592,4.2601027,4.716308,4.4012313,4.788513,5.395693,5.681231,5.602462,5.6320004,7.450257,8.448001,8.231385,7.3452315,7.276308,10.187488,14.5952835,19.062155,21.32677,18.294155,16.633438,13.929027,12.232206,11.766154,10.935796,9.754257,10.266257,11.398565,12.232206,12.005745,11.943385,12.2157955,11.559385,9.334154,5.5072823,4.2568207,5.044513,6.3376417,7.643898,9.511385,9.741129,10.338462,11.149129,12.071385,13.046155,13.233232,12.980514,12.947693,13.66318,15.527386,17.969233,19.492104,20.79836,22.488617,25.048616,24.237951,20.22072,16.02954,13.410462,12.813129,13.794462,14.50995,14.982565,15.671796,17.483488,20.23713,23.190975,26.377848,29.105232,29.974977,33.920002,37.25785,41.488415,47.36657,54.908722,63.737442,76.22237,86.04226,89.79693,87.0236,87.08267,89.915085,87.97211,77.46298,58.34503,43.231182,34.642056,34.628925,42.548515,55.062977,66.75365,76.045135,80.436516,76.45539,59.638157,35.823593,24.421745,20.243694,19.226257,18.395899,17.552412,16.853334,16.082052,15.182771,14.276924,13.364513,12.2157955,11.001437,9.842873,8.815591,8.408616,8.828718,9.133949,8.644924,6.954667,4.857436,3.4297438,2.609231,2.1366155,1.5556924,1.3489232,1.7066668,2.6354873,3.8531284,4.781949,4.6211286,4.3749747,4.3651285,4.9460516,6.4754877,9.8592825,13.282462,15.002257,14.290052,11.444513,8.54318,7.3780518,6.0947695,4.2272825,2.7175386,1.1651284,0.44964105,0.15097436,0.026256412,0.016410258,0.006564103,0.0,0.0,0.0,0.006564103,0.02297436,0.029538464,0.026256412,0.04594872,0.15097436,0.23630771,0.40369233,1.0699488,1.8838975,1.7132308,0.6629744,0.47589746,0.8566154,1.719795,3.1967182,5.3891287,6.816821,9.26195,13.88636,21.22831,14.657642,8.14277,3.6430771,1.5983591,0.9288206,0.5677949,0.28225642,0.15753847,0.18379489,0.23958977,0.51856416,1.7296412,3.1048207,4.1189747,4.4767184,4.1747694,3.5971284,2.7733335,1.8806155,1.2307693,0.9189744,0.5021539,0.19692309,0.07548718,0.06235898,0.03938462,0.032820515,0.026256412,0.02297436,0.04266667,0.07876924,0.1148718,0.13784617,0.15753847,0.19364104,0.23302566,0.2231795,0.20348719,0.25928208,0.512,0.508718,0.3446154,0.24615386,0.24287182,0.15753847,0.17723078,0.19364104,0.31507695,0.48246157,0.48246157,0.4201026,0.2986667,0.21989745,0.20348719,0.17066668,0.13784617,0.12143591,0.101743594,0.08205129,0.09189744,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08533334,0.17066668,0.0,0.0,0.36758977,0.4397949,0.4004103,1.2668719,2.3171284,2.231795,3.6036925,5.8912826,5.4186673,2.4155898,1.6180514,1.0929232,0.49887183,1.083077,0.5940513,0.33476925,0.40369233,0.7417436,1.1454359,0.9124103,0.56123084,0.8041026,2.284308,5.5532312,6.675693,7.1581545,7.824411,8.621949,8.621949,8.2904625,7.706257,7.8506675,8.425026,7.827693,7.79159,9.714872,12.422565,14.378668,13.673027,12.097642,10.935796,9.701744,8.283898,6.941539,7.125334,7.125334,6.5706673,5.32677,3.508513,2.03159,1.3718976,1.4506668,2.15959,3.3575387,3.1113849,2.1924105,1.5327181,1.3784616,1.2832822,0.65969235,0.23958977,0.06564103,0.08205129,0.108307704,0.068923086,0.02297436,0.0,0.0,0.0,0.19692309,0.45620516,0.58420515,0.48902568,0.18379489,0.20676924,0.15753847,0.18379489,0.39384618,0.86974365,1.6869745,2.3762052,2.2678976,1.6771283,1.9232821,1.4572309,1.4441026,1.6082052,1.7460514,1.7099489,1.4769232,0.92553854,0.8041026,1.2996924,2.044718,2.3860514,2.225231,1.9561027,1.8642052,2.1202054,1.3751796,1.7591796,2.556718,2.9046156,1.7690258,1.7329233,0.955077,0.571077,0.90256417,1.463795,1.086359,0.73517954,0.69907695,1.3193847,2.989949,1.7952822,1.1093334,1.1848207,2.034872,3.4625645,4.562052,3.7842054,2.740513,2.5074873,3.629949,3.7415388,3.5216413,4.4077954,6.449231,8.316719,9.304616,10.200616,12.918155,14.844719,8.848411,7.397744,6.2194877,5.139693,4.4406157,4.8672824,6.4656415,7.250052,10.371283,14.565744,14.17518,6.8266673,5.182359,8.379078,13.115078,13.640206,7.453539,4.027077,2.7536411,3.3378465,5.8289237,5.5597954,5.979898,7.273026,8.339693,6.7905645,5.044513,4.9099493,3.7809234,1.8116925,1.9232821,3.8038976,3.623385,2.5895386,2.0020514,3.2361028,5.8486156,6.564103,5.3005133,3.0096412,1.6771283,2.3269746,3.045744,4.900103,7.5585647,9.291488,11.136001,11.395283,9.783795,7.1614366,5.540103,5.356308,8.277334,11.664412,13.354668,11.657847,7.8014364,6.232616,5.858462,5.7403083,5.080616,6.0685134,6.1078978,5.7829747,5.8486156,7.200821,7.702975,7.141744,9.442462,13.892924,15.153232,11.073642,7.584821,6.0225644,5.943795,5.1265645,4.5423594,3.7448208,2.8914874,2.2088206,2.0151796,4.1124105,4.886975,4.397949,4.0041027,6.3474874,7.9327188,9.245539,7.6964107,4.266667,3.508513,7.243488,7.0990777,5.110154,3.367385,4.013949,3.6824617,2.8980515,2.8521028,3.5971284,4.013949,3.2918978,4.338872,4.1189747,2.7536411,3.508513,4.315898,4.7458467,5.0018463,5.287385,5.8125134,8.425026,8.008205,5.8157954,3.5380516,3.2820516,4.2929235,3.7973337,2.9538465,2.3072822,1.7690258,1.8806155,1.7329233,1.9035898,2.409026,2.7011285,4.07959,4.076308,3.3214362,2.409026,1.9068719,1.6147693,1.7788719,1.9200002,1.9561027,2.2121027,2.737231,3.0982566,3.121231,2.7602053,2.0742567,2.1103592,2.8914874,3.5807183,3.6496413,2.868513,2.6486156,3.0424619,3.121231,2.6847181,2.2580514,3.370667,2.356513,1.6836925,2.0053334,2.1530259,2.5435898,2.9965131,3.1671798,3.1376412,3.4166157,2.540308,2.2547693,1.8116925,1.2603078,1.4802053,2.678154,3.7809234,3.8859491,3.0687182,2.3958976,3.8596926,7.3386674,11.208206,17.847795,33.631184,33.78872,23.381334,13.121642,7.39118,4.240411,5.0838976,8.096821,10.860309,10.909539,5.720616,5.674667,8.195283,9.288206,7.8047185,5.4482055,3.751385,2.9965131,2.789744,2.6157951,1.847795,4.6900516,10.765129,12.744206,9.42277,5.737026,4.821334,4.9952826,6.5903597,8.041026,5.904411,6.245744,7.788308,9.284924,10.266257,11.047385,9.691898,6.626462,7.1089234,11.805539,16.784412,17.591797,13.059283,11.634872,14.309745,14.601848,11.588924,10.742155,11.54954,13.459693,15.898257,14.470565,12.228924,9.810052,7.7456417,6.439385,8.4053335,11.237744,11.142565,8.257642,6.6822567,11.113027,22.721643,28.868925,25.412926,16.708925,11.88759,8.100103,7.496206,9.40636,10.345026,3.2656412,1.723077,2.2908719,2.7995899,2.3335385,1.273436,1.6016412,1.4441026,1.1454359,3.2820516,1.2668719,1.522872,1.9626669,1.8149745,1.6311796,1.657436,1.5721027,1.0896411,0.44964105,0.4135385,0.88943595,1.913436,2.3335385,1.8773335,1.1454359,1.0108719,1.4080001,2.6387694,4.841026,7.965539,9.563898,10.200616,10.555078,11.264001,12.924719,14.217847,13.974976,14.011078,16.475899,23.850668,28.025438,28.49149,26.584618,23.318975,19.364103,10.633847,5.156103,3.5577438,4.57518,5.0510774,6.514872,6.7905645,7.1089234,7.315693,5.874872,5.0674877,5.7829747,6.229334,5.8289237,5.218462,7.062975,8.320001,8.789334,8.464411,7.5388722,8.759795,9.7673855,9.170052,7.6176414,7.8112826,8.851693,8.605539,7.653744,6.3901544,5.037949,5.330052,6.042257,7.1056414,8.274052,9.140513,8.113232,8.306872,9.065026,9.990565,10.955488,11.040821,10.587898,9.042052,6.4000006,3.190154,2.8849232,4.46359,6.294975,7.778462,9.353847,9.7214365,11.329642,12.973949,14.181745,15.241847,15.632411,14.788924,13.817437,13.830565,15.931078,19.203283,20.73272,21.556515,22.472206,24.047592,24.635078,21.238155,16.128002,11.690667,10.420513,10.545232,10.427077,10.538668,11.073642,11.979488,13.443283,15.796514,18.244925,20.857437,24.566156,27.936823,32.915695,38.95467,45.092106,49.988926,59.168823,66.93744,69.37273,66.37949,61.692722,59.506878,59.090057,55.19098,46.431183,35.311592,33.772312,31.199183,41.636105,63.10729,77.62052,74.6437,61.650055,46.32944,33.555695,25.363695,20.06318,17.959387,17.985641,18.95713,19.590565,19.715284,19.846565,19.643078,19.049026,18.281027,17.240616,15.675078,14.020925,12.47836,11.001437,11.355898,14.391796,16.918976,17.14872,14.693745,10.9456415,7.463385,5.097026,3.7907696,2.5928206,2.7766156,3.2984617,4.3290257,5.2709746,4.7458467,4.086154,4.279795,4.585026,4.585026,4.1813335,3.6693337,4.896821,5.7435904,6.0750775,7.722667,8.257642,7.1122055,5.543385,4.0500517,2.3663592,1.1946667,0.46933338,0.12143591,0.026256412,0.016410258,0.016410258,0.006564103,0.0,0.006564103,0.029538464,0.06564103,0.12143591,0.108307704,0.052512825,0.07548718,0.12471796,0.3117949,0.7384616,1.1027694,0.6859488,0.4660513,0.6498462,0.9419488,1.6344616,3.6004105,6.8004107,10.748719,17.657436,26.17108,31.369848,16.344616,6.4623594,1.7329233,0.7811283,0.8533334,0.7581539,0.45620516,0.23302566,0.16738462,0.16738462,0.38728207,1.6049232,3.626667,6.052103,8.283898,9.225847,8.838565,6.695385,3.6824617,1.9987694,1.8642052,1.2373334,0.56451285,0.13456412,0.06235898,0.049230773,0.036102567,0.029538464,0.029538464,0.029538464,0.06564103,0.0951795,0.118153855,0.14441027,0.16738462,0.18051283,0.18379489,0.20676924,0.256,0.3052308,0.23302566,0.23958977,0.23958977,0.20676924,0.18379489,0.36758977,0.4397949,0.38400003,0.27569234,0.27569234,0.3117949,0.32820517,0.36102566,0.39056414,0.36758977,0.256,0.18379489,0.128,0.09189744,0.09189744,0.0,0.0,0.0,0.0,0.0,0.0,0.118153855,0.059076928,0.0,0.0,0.0,0.059076928,0.029538464,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016410258,0.032820515,0.0,0.0,0.22646156,0.26584616,0.128,0.25271797,1.214359,1.3554872,1.7887181,2.9735386,4.7327185,6.1538467,3.8137438,1.2406155,0.11158975,0.2297436,0.12143591,0.06564103,0.17723078,0.85005134,2.7569232,3.062154,1.782154,1.332513,2.4648206,4.2601027,4.827898,5.139693,5.943795,7.000616,7.1089234,6.7577443,7.830975,8.956718,9.248821,8.280616,8.937026,10.643693,12.796719,14.162052,12.87877,11.956513,12.117334,12.005745,11.136001,9.872411,9.048616,7.8539495,6.5312824,5.4449234,5.07077,2.3269746,1.1848207,0.8008206,0.7581539,1.0732309,1.339077,1.6935385,2.733949,3.826872,3.1245131,3.3608208,1.6410258,0.3708718,0.23302566,0.18051283,0.18379489,0.27897438,0.4004103,0.44307697,0.26912823,0.2986667,0.39712822,0.571077,0.7811283,0.96492314,0.73517954,0.65969235,0.5316923,0.4397949,0.761436,1.9200002,2.1891284,2.2547693,2.422154,2.605949,2.5632823,2.3072822,2.409026,2.806154,2.8192823,2.9111798,2.4155898,2.3040001,2.6584618,2.678154,2.2777438,2.034872,2.3236926,2.8160002,2.487795,3.56759,2.7503593,1.8116925,1.5786668,1.9298463,2.3105643,1.9396925,1.5983591,1.8346668,2.9407182,2.2219489,1.529436,1.5622566,2.2219489,2.6256413,2.2383592,1.522872,1.204513,1.5195899,2.1956925,5.481026,4.8607183,3.4592824,3.4133337,5.865026,5.7009234,4.923077,4.969026,5.8223596,6.0225644,5.2315903,6.426257,8.536616,9.42277,5.87159,4.8672824,4.850872,5.097026,5.149539,4.8049235,3.8071797,3.6562054,4.6769233,6.1472826,6.314667,6.485334,7.890052,9.160206,9.012513,6.2555904,4.1682053,3.170462,2.6486156,2.7437952,4.315898,4.604718,5.080616,6.180103,7.24677,6.5444107,4.841026,4.854154,4.57518,4.096,5.622154,5.8814363,6.048821,5.87159,5.717334,6.5805135,7.1122055,7.0826674,5.979898,4.164923,2.861949,4.1747694,5.169231,6.550975,7.77518,7.059693,7.5552826,8.1066675,8.726975,9.176616,8.969847,6.294975,6.8004107,8.113232,8.730257,8.021334,7.0925136,7.5585647,7.5520005,6.488616,5.0674877,5.7632823,5.933949,6.0061545,6.3376417,7.213949,6.1997952,6.1341543,8.146052,11.306667,12.612924,10.440206,8.297027,6.7085133,5.5893335,4.2371287,4.276513,3.7152824,2.6847181,1.6804104,1.5622566,2.793026,3.9417439,4.8672824,5.3366156,5.0051284,7.1483083,9.170052,7.9524107,4.3651285,3.2656412,6.452513,8.067283,7.4010262,5.428513,4.8049235,3.9581542,4.161641,6.409847,8.923898,7.1515903,4.1846156,4.9920006,5.4449234,4.2896414,3.1442053,3.3542566,3.3936412,3.4330258,3.6004105,3.9581542,5.280821,5.1856413,4.5456414,4.092718,4.4045134,3.8334363,2.9407182,2.484513,2.5600002,2.5862565,2.0053334,1.3981539,1.1290257,1.3981539,2.2482052,3.259077,3.95159,4.1222568,3.5905645,2.2121027,1.6475899,1.785436,2.048,2.2580514,2.6518977,3.1474874,3.367385,3.242667,2.934154,2.8553848,2.8455386,3.2000003,3.7152824,4.1682053,4.332308,3.2065644,3.0490258,3.1376412,3.0752823,2.7831798,3.0162053,2.733949,2.5600002,2.4746668,1.8084104,1.9462565,1.8838975,2.0676925,2.5961027,3.1967182,2.6026669,2.5140514,2.284308,2.5173335,5.080616,3.4855387,2.5862565,2.2678976,2.6945643,4.348718,6.741334,8.283898,10.758565,14.739694,19.603693,16.853334,13.2562065,10.489437,8.41518,5.07077,6.091488,8.39877,8.684308,6.5739493,4.647385,6.2588725,6.186667,5.907693,5.7468724,4.886975,3.82359,5.395693,6.2194877,4.896821,2.028308,5.2545643,13.403898,14.608412,7.9425645,3.4067695,5.4383593,8.992821,11.090053,10.134975,5.917539,8.641642,11.34277,13.213539,13.13477,9.668923,11.680821,16.905848,18.162872,14.972719,13.538463,13.63036,15.02195,17.11918,18.763489,18.215385,16.305231,13.925745,12.356924,11.946668,12.104206,10.47959,9.104411,7.837539,6.8463597,6.5870776,7.75877,9.590155,10.889847,11.83836,13.994668,19.236105,23.972105,23.88349,19.715284,17.270155,12.3995905,8.864821,6.5444107,5.346462,5.182359,2.858667,2.4910772,3.2886157,4.1911798,3.8859491,5.4580517,5.789539,3.9942567,1.7657437,3.367385,2.3368206,1.9331284,1.7624617,1.6213335,1.4867693,1.3062565,0.9189744,0.5513847,0.3511795,0.4135385,0.8795898,1.214359,1.4966155,1.8904617,2.6322052,2.7536411,2.546872,2.6289232,3.7940516,7.0367184,11.858052,14.496821,14.552616,13.147899,12.924719,12.928001,11.431385,10.374565,11.218052,14.9398985,18.947283,19.02277,18.487797,19.219694,21.622156,17.365335,11.503591,7.4010262,5.7534366,4.598154,5.225026,6.0291286,6.3310776,5.832206,4.6178465,4.571898,5.2742567,5.1954875,4.781949,6.426257,8.749949,8.441437,7.4010262,6.8594875,7.3682055,8.342975,7.9950776,7.3386674,6.8955903,6.701949,6.9677954,6.4722056,5.9602056,5.6352825,5.169231,6.488616,7.026872,7.4830775,8.021334,8.274052,8.303591,8.598975,9.189744,9.750975,9.613129,9.941334,9.101129,7.8080006,6.2785645,4.240411,4.450462,5.481026,6.961231,8.569437,10.036513,10.617436,11.162257,11.021129,10.617436,11.434668,12.097642,12.42913,12.438975,12.448821,13.072412,13.748514,14.460719,16.600616,19.580719,20.86072,19.787489,16.466053,12.363488,9.104411,8.467693,8.356103,8.480822,8.684308,9.081436,10.072617,10.8537445,12.33395,14.431181,17.09949,20.33231,23.03672,25.924925,29.784618,35.026054,41.688618,47.058056,51.905643,52.8279,49.608208,45.22339,48.380722,50.835697,51.01949,49.726364,50.126774,52.017235,62.6478,78.72657,95.38955,106.233444,97.89375,73.232414,50.021748,34.789745,22.820105,20.676924,20.775387,22.340925,24.362669,25.622976,27.014566,26.87672,25.550772,23.702976,22.321232,21.379284,19.859694,18.497643,17.6279,17.165129,19.784206,26.17108,32.482464,35.876106,34.517338,29.440002,20.867283,13.000206,8.008205,6.012718,4.7589746,4.716308,5.605744,6.636308,6.5017443,5.297231,4.926359,5.2578464,5.5696416,4.571898,3.318154,3.1048207,3.045744,3.1638978,4.414359,4.089436,3.6726158,3.69559,3.6102567,1.7788719,0.6465641,0.19692309,0.059076928,0.016410258,0.016410258,0.016410258,0.013128206,0.016410258,0.036102567,0.07876924,0.15425642,0.21333335,0.21333335,0.15097436,0.03938462,0.059076928,0.09189744,0.18707694,0.3249231,0.41682056,1.6738462,3.7185643,5.3924108,6.4656415,7.6307697,10.368001,15.067899,22.550976,29.9159,30.506668,13.778052,4.857436,1.2012309,0.45292312,0.4397949,0.3708718,0.256,0.29210258,0.5415385,0.9124103,2.3335385,4.1813335,6.6002054,9.826463,14.168616,12.678565,9.058462,5.366154,2.7142565,1.3029745,1.2077949,0.9911796,0.65641034,0.2986667,0.108307704,0.068923086,0.049230773,0.049230773,0.055794876,0.055794876,0.06235898,0.08861539,0.1148718,0.13128206,0.15425642,0.14769232,0.13128206,0.118153855,0.12143591,0.17066668,0.16738462,0.16410258,0.16738462,0.17394873,0.15753847,0.2231795,0.27569234,0.30851284,0.33805132,0.39712822,0.37415388,0.33476925,0.3446154,0.4397949,0.6104616,0.6268718,0.5349744,0.36758977,0.190359,0.10502565,0.14769232,0.029538464,0.0,0.0,0.068923086,0.34789747,0.3117949,0.12143591,0.068923086,0.23958977,0.5021539,0.43651286,0.41682056,0.39384618,0.29210258,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.068923086,0.34789747,0.068923086,0.30851284,1.2504616,2.0578463,0.8598975,0.6071795,1.0272821,1.4408206,2.169436,4.5522056,5.037949,2.6880002,0.6301539,0.013128206,0.006564103,0.0,0.0,0.4135385,1.8838975,5.2644105,5.221744,3.1540515,2.2383592,2.917744,2.9111798,2.92759,3.245949,4.0369234,4.972308,5.208616,5.464616,7.256616,8.973129,9.714872,9.288206,10.843898,11.185231,11.588924,11.98277,10.948924,10.57477,10.656821,10.279386,9.278359,8.251078,8.077128,7.0957956,5.622154,4.33559,4.273231,2.034872,1.0535386,0.60061544,0.33476925,0.29210258,0.5513847,1.0272821,1.785436,2.5042052,2.4681027,2.6420515,1.7558975,1.142154,1.0732309,0.7581539,0.46276927,0.38400003,0.45620516,0.5284103,0.380718,0.3708718,0.5677949,0.72861546,0.761436,0.7384616,0.9156924,1.0633847,1.0765129,0.90912825,0.60389745,1.2274873,1.401436,1.6147693,2.0053334,2.3729234,2.0775387,2.0742567,2.3040001,2.809436,3.7185643,3.6627696,3.5905645,3.6069746,3.6693337,3.5610259,2.9965131,2.989949,3.2000003,3.314872,3.0358977,3.18359,2.3893335,1.6475899,1.5064616,2.0512822,2.7733335,2.9768207,2.9013336,2.7470772,2.6880002,2.3729234,2.3893335,2.6026669,2.7437952,2.4057438,2.4713848,2.15959,1.9429746,2.048,2.4615386,4.069744,4.1189747,3.8400004,4.2568207,6.2030773,5.0116925,4.2929235,4.571898,5.4416413,5.5565133,5.5171285,6.9842057,7.466667,6.363898,4.9427695,4.8804107,5.3136415,6.042257,6.695385,6.75118,7.6209235,7.958975,7.4830775,7.0826674,8.815591,11.109744,11.080206,9.826463,7.650462,4.07959,3.2000003,2.4188719,2.1234872,2.6518977,4.3027697,3.4625645,3.5183592,4.5128207,5.6976414,5.5236926,4.325744,4.352,4.1747694,3.895795,5.146257,7.634052,7.3485136,6.8233852,7.3025646,8.723693,8.914052,8.713847,7.9852314,7.000616,6.445949,7.4765134,8.100103,8.139488,7.5881033,6.6100516,6.87918,6.6428723,6.8594875,7.788308,8.976411,8.717129,9.114257,9.481847,9.216001,7.778462,7.3550773,8.28718,8.224821,7.0334363,6.7774363,8.710565,8.257642,7.0826674,6.314667,6.5312824,5.8945646,5.2676926,6.012718,7.778462,8.52677,7.7390776,7.5881033,7.1876926,6.121026,4.4340515,4.388103,3.9417439,3.0752823,2.1924105,2.1070771,4.059898,5.156103,5.4449234,4.9394875,3.6168208,4.962462,6.009436,5.421949,3.7907696,3.6529233,5.861744,7.1680007,6.8496413,5.4843082,4.9329233,3.7415388,5.0642056,7.7948723,9.580308,6.806975,3.764513,4.073026,5.1922054,5.2709746,3.1442053,3.629949,3.2918978,3.1015387,3.3214362,3.5216413,3.761231,3.7907696,4.017231,4.342154,4.161641,2.8980515,2.0184617,1.8313848,2.2022567,2.5632823,2.2744617,1.8707694,1.6049232,1.585231,1.7624617,2.2383592,2.806154,3.370667,3.4855387,2.3269746,1.5163078,1.463795,1.7329233,2.0808206,2.4516926,2.9538465,3.1638978,3.308308,3.4330258,3.4264617,2.9407182,2.8192823,3.1934361,3.9876926,4.9099493,3.892513,3.3378465,3.0358977,2.806154,2.4746668,2.4943593,2.4385643,2.409026,2.3269746,1.9068719,1.7099489,1.2077949,1.1093334,1.6344616,2.540308,2.3302567,2.3072822,2.9407182,4.1156926,5.149539,4.1124105,4.138667,4.775385,5.5729237,6.1013336,6.7249236,6.5870776,6.987488,8.339693,10.184206,10.410667,12.511181,13.216822,11.241027,7.276308,6.163693,6.921847,6.747898,5.540103,5.917539,6.961231,6.7938466,6.3245134,6.114462,6.36718,4.135385,6.2129235,9.701744,11.382154,7.6964107,7.4732313,9.225847,7.821129,3.5478978,2.1530259,6.0619493,7.955693,7.571693,5.7435904,4.391385,8.868103,11.661129,12.744206,11.516719,6.7971287,18.625643,39.246773,44.061543,31.271387,21.897848,17.447386,18.474669,18.86195,16.370872,12.655591,11.467488,10.397539,9.567181,8.973129,8.500513,7.896616,7.250052,6.6625648,6.3606157,6.705231,5.2512827,5.5138464,7.5388722,11.158976,15.996719,21.691078,22.442669,19.081848,14.171899,12.028719,7.650462,5.280821,3.9187696,3.1540515,3.1770258,2.481231,2.166154,2.7011285,3.8629746,4.7294364,5.9667697,7.026872,5.7435904,3.1507695,3.4789746,1.9364104,1.2898463,1.148718,1.2242053,1.3292309,1.083077,0.6465641,0.39712822,0.37743592,0.29210258,0.6235898,0.9517949,1.2931283,1.6672822,2.0808206,2.2646155,2.7864618,3.3509746,4.1025643,5.61559,9.110975,12.002462,13.062565,12.583385,12.347078,11.67754,10.374565,9.242257,9.147078,11.027693,12.665437,12.150155,11.776001,13.082257,16.866463,16.820515,14.191591,10.988309,8.260923,6.1078978,4.926359,4.6112823,4.673641,4.5456414,3.6069746,3.6594875,4.1124105,4.414359,4.8672824,6.6002054,8.178872,7.9294367,7.2270775,6.626462,5.858462,6.3868723,6.2555904,6.1407185,6.186667,6.012718,5.799385,5.674667,5.681231,5.7107697,5.4974365,6.009436,6.166975,6.4722056,6.889026,6.8496413,6.7905645,7.026872,7.0793853,6.8594875,6.685539,6.564103,5.835488,5.1331286,4.6933336,4.3552823,4.7983594,5.425231,6.160411,6.892308,7.453539,7.890052,8.218257,8.356103,8.546462,9.337437,9.908514,10.371283,10.587898,10.581334,10.528821,10.515693,11.434668,13.505642,15.691488,15.698052,12.970668,10.624001,8.539898,7.003898,6.688821,6.547693,7.003898,7.322257,7.450257,8.024616,8.464411,9.475283,10.952206,12.937847,15.619284,18.576412,21.746874,24.864822,27.910566,31.126976,32.725334,34.527184,34.999798,33.906876,32.292107,36.26995,40.03118,45.298874,52.194466,59.234467,72.4677,85.7436,95.19262,97.19467,88.37908,75.01457,58.88985,47.317337,39.79159,27.989336,26.305643,26.643694,27.608618,29.000208,31.809643,38.95795,43.17867,43.88431,42.003696,39.972107,38.95467,36.58503,35.14749,34.517338,32.164104,31.747284,35.879387,41.49826,46.027493,47.35672,43.136,35.93518,27.0999,18.30072,11.526565,8.802463,7.762052,7.7292314,8.03118,8.021334,7.1647186,5.874872,5.1232824,4.818052,3.8071797,2.9111798,2.737231,2.8914874,3.2032824,3.7415388,3.190154,2.9801028,2.993231,2.6486156,0.892718,0.318359,0.101743594,0.032820515,0.013128206,0.032820515,0.07876924,0.08205129,0.07876924,0.10502565,0.21989745,0.36430773,0.4266667,0.39384618,0.27897438,0.10502565,0.049230773,0.026256412,0.026256412,0.06235898,0.18707694,1.142154,3.2754874,5.6287184,7.6734366,9.29477,11.670976,16.489027,22.232616,25.682053,21.920822,9.5606165,3.245949,0.7811283,0.29210258,0.23630771,0.18707694,0.15425642,0.38728207,1.142154,2.681436,4.9526157,7.5454364,10.089026,12.360206,14.28677,11.254155,7.0925136,3.7054362,1.7788719,0.7811283,0.7089231,0.65641034,0.5218462,0.318359,0.15753847,0.118153855,0.098461546,0.0951795,0.101743594,0.1148718,0.12471796,0.12471796,0.118153855,0.10502565,0.1148718,0.10502565,0.09189744,0.07548718,0.06564103,0.09189744,0.10502565,0.1148718,0.13128206,0.14769232,0.14441027,0.15753847,0.18051283,0.20676924,0.23958977,0.2986667,0.32164106,0.318359,0.33476925,0.39056414,0.47917953,0.5349744,0.5316923,0.50543594,0.446359,0.2986667,0.14769232,0.029538464,0.12143591,0.21333335,0.37415388,0.94523084,0.41025645,0.18707694,0.14769232,0.3117949,0.86317956,0.47917953,0.4004103,0.39384618,0.29210258,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.029538464,0.10502565,0.30194873,0.7515898,0.21333335,0.3446154,1.6771283,3.0260515,1.4900514,0.9616411,1.5491283,2.0873847,2.6256413,4.4242053,2.8127182,1.083077,0.12143591,0.006564103,0.0,0.0,0.006564103,0.6235898,2.5140514,6.3934364,5.4449234,3.764513,2.8488207,2.7470772,2.0250258,1.8248206,2.1202054,2.7175386,3.3378465,3.6102567,4.1222568,5.7468724,7.4404106,8.608821,9.088,11.575796,12.035283,11.595488,10.94236,10.308924,9.7903595,8.923898,7.6996927,6.51159,6.163693,6.665847,5.940513,4.522667,3.1671798,2.8488207,1.6738462,1.0404103,0.65969235,0.37743592,0.15753847,0.24615386,0.56123084,1.024,1.5524104,2.041436,2.0184617,1.9561027,1.8248206,1.5819489,1.1585642,0.67938465,0.5677949,0.6498462,0.7122052,0.5284103,0.5677949,0.88287187,1.0043077,0.7811283,0.39056414,0.97805136,1.4145643,1.6311796,1.4834872,0.7811283,0.7778462,0.94523084,1.1881026,1.4802053,1.8740515,1.6935385,2.2646155,3.117949,3.9844105,4.8049235,4.466872,4.4110775,4.4110775,4.414359,4.5390773,3.9384618,3.4592824,3.0490258,2.7963078,2.937436,2.546872,1.9495386,1.5622566,1.5261539,1.7033848,2.1924105,3.1934361,3.9942567,3.9187696,2.3401027,2.231795,2.5238976,2.7142565,2.5731285,2.1300514,2.5632823,2.6420515,2.5140514,2.425436,2.7175386,2.9636924,3.95159,4.969026,5.8092313,6.770872,5.0477953,4.699898,5.0543594,5.5926156,5.98318,6.698667,7.9524107,7.571693,5.9536414,6.0717955,5.8781543,5.8486156,6.62318,7.8736415,8.283898,9.7214365,10.683078,10.643693,10.387693,12.002462,12.655591,10.738873,8.14277,5.6352825,2.8521028,2.540308,2.028308,1.8740515,2.3236926,3.3214362,2.4352822,3.4888208,5.208616,6.4032826,5.9569235,5.2020516,4.5095387,3.8334363,3.498667,4.2174363,7.2172313,7.0400004,6.8627696,7.9195905,9.504821,9.93477,9.6754875,9.29477,8.92718,8.293744,7.821129,7.8047185,7.53559,7.5487185,9.626257,12.081232,10.768411,8.539898,7.2927184,7.9917955,9.314463,9.787078,9.878975,9.504821,8.054154,8.513641,9.219283,8.700719,7.4797955,8.083693,10.545232,9.094564,7.026872,6.235898,7.200821,6.6560006,5.356308,5.100308,5.9995904,6.4623594,5.9470773,7.145026,7.762052,6.941539,5.2348723,4.5095387,5.0674877,5.179077,4.516103,4.164923,6.1078978,6.3474874,5.4941545,4.082872,2.6026669,3.2853336,3.892513,4.0041027,3.764513,3.8728209,4.9099493,5.366154,5.330052,4.9526157,4.450462,3.4691284,4.841026,6.619898,7.062975,4.6112823,2.9965131,3.2787695,4.532513,5.182359,3.0162053,4.027077,3.8596926,3.892513,4.4701543,4.900103,4.457026,3.8629746,3.7710772,3.9680004,3.370667,2.2908719,1.529436,1.4441026,1.8871796,2.2022567,2.15959,2.100513,2.100513,2.0545642,1.6640002,1.6836925,1.9626669,2.4615386,2.7634873,2.0873847,1.394872,1.2635899,1.4539489,1.7329233,1.8937438,2.4024618,2.733949,2.9833848,3.170462,3.2262566,2.553436,2.1825643,2.422154,3.2820516,4.4898467,4.2338467,3.69559,3.1409233,2.7306669,2.546872,2.2547693,2.2088206,2.1366155,1.9790771,1.8707694,1.7526156,1.4309745,1.4408206,2.1234872,3.6069746,3.9384618,3.314872,3.5577438,4.663795,4.781949,4.7917953,5.1626673,5.474462,5.7042055,6.235898,4.8147697,4.713026,5.179077,6.2687182,8.835282,10.082462,12.340514,12.662155,10.427077,7.3550773,5.3202057,5.32677,5.7403083,6.163693,7.460103,8.320001,8.392206,7.9163084,7.1844106,6.5378466,3.9318976,4.630975,7.6701546,10.295795,7.965539,8.648206,6.1407185,2.92759,1.273436,3.2032824,5.986462,6.695385,6.5903597,6.7971287,8.310155,11.421539,13.958565,13.820719,10.322052,4.201026,23.305847,48.50544,54.79713,40.004925,24.786053,18.22195,19.790771,18.999796,13.351386,8.346257,7.1220517,6.314667,5.8157954,5.5138464,5.287385,6.1505647,6.514872,6.3540516,6.0028725,6.157129,4.125539,3.8006158,6.2818465,11.963078,20.539078,25.32431,22.42954,16.131283,10.387693,8.841846,5.8092313,3.7448208,2.6518977,2.2646155,2.0545642,1.7690258,1.5360001,1.6771283,2.4024618,3.8465643,4.9952826,5.8223596,4.923077,2.917744,2.4615386,1.1355898,0.69579494,0.62030774,0.6465641,0.77456415,0.6268718,0.42338464,0.37743592,0.45292312,0.36102566,0.45292312,0.7417436,1.1191796,1.3915899,1.2931283,1.5688206,2.484513,3.3345644,3.8006158,3.9384618,5.1331286,7.4863596,9.097847,9.521232,9.760821,9.199591,8.900924,8.687591,8.704,9.432616,8.805744,7.5421543,6.518154,6.9152827,10.233437,14.503386,16.239592,14.8480015,11.119591,7.240206,5.077334,4.4767184,4.8377438,5.2447186,4.460308,3.5347695,3.1803079,3.2918978,3.8137438,4.7261543,5.6451287,6.1407185,6.2884107,5.858462,4.315898,4.6080003,4.9920006,5.362872,5.720616,6.163693,5.687795,5.5597954,5.72718,5.98318,5.973334,5.8223596,5.664821,5.914257,6.3245134,5.9930263,5.5105643,5.0609236,4.5423594,4.1222568,4.2207184,3.8531284,3.501949,3.4592824,3.6857438,3.82359,4.391385,4.8640003,5.172513,5.32677,5.4186673,5.609026,5.7698464,6.124308,6.672411,7.207385,7.5585647,7.8736415,7.958975,7.748924,7.312411,7.125334,7.752206,8.818872,9.6,9.015796,6.8266673,5.805949,5.2545643,4.8738465,4.7491283,4.7327185,5.211898,5.5302567,5.5597954,5.677949,6.160411,6.961231,8.356103,10.440206,13.115078,15.9573345,19.193438,21.874874,23.492926,23.985233,24.362669,24.365952,23.939283,23.414156,23.5159,28.52431,34.021748,42.0759,52.453747,62.61498,79.65539,90.8439,91.854774,81.66072,62.53621,51.7678,46.63139,45.70585,44.757336,36.755695,36.43077,39.079388,43.06708,47.901543,54.222775,60.081234,62.92021,63.730877,63.793236,64.70564,64.18052,61.679596,60.731083,61.525337,60.908314,55.88349,54.38031,55.118774,56.277336,55.506054,50.56985,45.298874,38.839798,31.044926,22.439386,16.403694,13.039591,11.946668,12.199386,12.373334,10.896411,8.050873,5.668103,4.3027697,3.239385,2.4648206,2.4910772,3.0096412,3.5807183,3.6496413,3.5511796,3.446154,2.9013336,1.8248206,0.48902568,0.22646156,0.15425642,0.20020515,0.24943592,0.14441027,0.26584616,0.3446154,0.32164106,0.27241027,0.4135385,0.6235898,0.72861546,0.6826667,0.49887183,0.26912823,0.101743594,0.029538464,0.006564103,0.016410258,0.052512825,0.36430773,1.5130258,3.1606157,4.923077,6.36718,7.9130263,11.204924,14.329437,15.064616,10.893129,4.781949,1.6475899,0.42338464,0.17723078,0.118153855,0.098461546,0.101743594,0.35774362,1.4703591,4.414359,7.1122055,10.19077,13.423591,15.556924,14.303181,9.724719,5.477744,2.6453335,1.3259488,0.6301539,0.4397949,0.38400003,0.34789747,0.28225642,0.19692309,0.18707694,0.20020515,0.20348719,0.190359,0.16410258,0.15097436,0.14112821,0.12471796,0.101743594,0.09189744,0.07876924,0.07876924,0.072205134,0.059076928,0.06235898,0.072205134,0.10502565,0.13128206,0.13784617,0.13784617,0.15097436,0.15753847,0.15097436,0.14769232,0.18379489,0.2297436,0.25271797,0.27241027,0.29538465,0.31507695,0.34133336,0.36102566,0.4004103,0.4266667,0.34789747,0.43651286,0.42994875,0.636718,0.8763078,1.1913847,1.847795,0.6268718,0.34133336,0.21333335,0.14441027,0.7187693,0.14441027,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.059076928,0.23630771,0.5349744,0.9321026,0.42338464,0.2986667,1.0765129,2.0808206,1.463795,1.6771283,2.15959,2.6190772,2.9965131,3.4724104,1.2471796,0.28225642,0.006564103,0.0,0.0,0.072205134,0.19692309,0.8566154,2.412308,5.110154,3.754667,3.2295387,2.674872,1.9528207,1.6377437,1.529436,1.7132308,2.0184617,2.3401027,2.6322052,3.0293336,4.2962055,5.6451287,6.76759,7.834257,10.581334,12.186257,12.150155,11.024411,10.387693,10.400822,8.408616,6.1538467,4.8705645,5.277539,5.687795,4.9493337,3.7218463,2.550154,1.8806155,1.4769232,1.1290257,0.83035904,0.5546667,0.23958977,0.26912823,0.57764107,1.214359,1.9823592,2.409026,2.4385643,2.484513,2.4746668,2.281026,1.7099489,0.93866676,0.9485129,1.2012309,1.2504616,0.7318975,0.79097444,1.1191796,1.1881026,0.8336411,0.26584616,0.8992821,1.4572309,1.7887181,1.7657437,1.2668719,1.1126155,1.2373334,1.3817437,1.522872,1.8740515,1.9922053,3.2689233,5.0543594,6.3245134,5.6976414,5.395693,5.149539,4.97559,5.0084105,5.4941545,4.84759,3.5840003,2.4188719,1.8576412,2.1989746,2.3138463,1.8313848,1.4933335,1.4605129,1.3029745,1.4309745,3.1770258,4.772103,4.906667,2.733949,2.3269746,2.156308,2.0512822,1.9167181,1.7362052,2.353231,2.678154,2.674872,2.5304618,2.665026,3.5905645,4.965744,6.4032826,7.4732313,7.716103,6.560821,6.669129,6.73477,6.4722056,6.62318,7.069539,7.384616,7.0990777,6.675693,7.509334,6.5936418,5.7764106,6.301539,7.722667,7.9097443,7.6012316,8.914052,10.496001,11.392001,11.063796,9.242257,6.9710774,4.7589746,2.8914874,1.4244103,1.7755898,2.038154,2.166154,2.0545642,1.5261539,1.9200002,4.525949,7.00718,8.04759,7.3682055,6.9120007,5.142975,3.757949,3.4822567,4.073026,5.031385,5.9963083,7.1483083,8.362667,9.235693,9.370257,9.216001,9.442462,9.662359,8.448001,6.183385,5.093744,5.395693,8.008205,14.532925,21.264412,19.862976,14.805334,9.803488,7.7981544,8.01477,8.0377445,8.165744,8.385642,8.375795,10.587898,10.607591,9.061745,7.4108725,7.9261546,9.176616,7.204103,5.4974365,5.8223596,8.208411,7.433847,5.976616,5.477744,6.114462,6.5837955,5.8781543,7.2927184,8.129642,7.4436927,6.058667,5.402257,6.9710774,8.057437,7.7292314,6.8496413,7.145026,6.173539,5.0084105,3.9909747,2.7109745,3.1113849,4.1058464,4.71959,4.5587697,3.8301542,4.027077,3.8498464,3.9253337,4.1156926,3.508513,3.4034874,4.017231,4.342154,3.8859491,2.6715899,2.809436,3.367385,4.076308,4.2469745,2.7602053,4.069744,4.571898,5.0215387,5.691077,6.377026,5.737026,4.3716927,3.4658465,3.170462,2.6190772,2.1267693,1.5327181,1.4473847,1.8084104,1.8707694,1.6475899,1.7624617,2.048,2.2416413,1.9922053,1.9659488,2.1497438,2.2383592,2.0808206,1.6705642,1.394872,1.3751796,1.4867693,1.5589745,1.3784616,1.7394873,2.156308,2.297436,2.2416413,2.4746668,2.041436,1.8084104,1.9364104,2.5009232,3.511795,4.023795,3.7448208,3.18359,2.7634873,2.8225644,2.3926156,2.359795,2.1989746,1.8937438,1.9396925,2.0118976,2.0873847,2.4451284,3.3903592,5.2512827,5.9470773,4.5522056,3.442872,3.5249233,4.240411,4.4996924,4.1156926,3.1671798,2.802872,5.2315903,3.8629746,4.8082056,6.488616,8.4053335,11.155693,10.440206,9.645949,8.707283,7.571693,6.2194877,4.71959,4.857436,5.7074876,6.997334,9.074872,9.353847,9.045334,8.6580515,7.8670774,5.5269747,3.8432825,2.8356924,2.681436,2.9538465,2.6190772,6.928411,5.5105643,2.8192823,1.9593848,4.667077,5.074052,8.293744,13.164309,17.792002,19.554462,19.232822,19.472412,17.729643,12.71795,4.4077954,19.954874,34.87508,39.085953,30.762669,16.347898,12.425847,15.839181,15.619284,10.187488,7.3485136,6.3376417,4.1780515,2.7634873,2.674872,3.190154,5.2742567,6.9645133,7.578257,7.282872,7.076103,6.514872,6.2096415,8.904206,16.167385,28.389746,30.802053,24.425028,15.264822,8.418462,8.057437,7.000616,4.8607183,3.4133337,2.9833848,2.4582565,2.034872,1.4998976,0.9353847,0.761436,1.723077,3.3509746,3.1540515,2.1530259,1.148718,0.7187693,0.5284103,0.47261542,0.33805132,0.14112821,0.08861539,0.07548718,0.18051283,0.37743592,0.571077,0.60061544,0.446359,0.45620516,0.7122052,1.0404103,0.9944616,1.3981539,1.975795,2.422154,2.556718,2.297436,2.2580514,3.8071797,5.0182567,5.395693,5.8781543,5.9569235,6.692103,7.650462,8.39877,8.467693,6.7249236,4.772103,3.0720003,2.6486156,5.077334,11.808822,16.15754,16.144411,12.225642,7.282872,5.1987696,5.398975,6.47877,7.4207187,7.5881033,5.5565133,3.7743592,2.6617439,2.3105643,2.4681027,2.9013336,3.6824617,4.2141542,4.194462,3.620103,3.9614363,4.532513,5.024821,5.5729237,6.73477,6.2720003,5.72718,5.6385646,6.009436,6.311385,6.2129235,6.045539,6.23918,6.564103,6.121026,5.3858466,4.1452312,3.308308,3.0949745,3.062154,2.7667694,2.8389745,3.1606157,3.3903592,2.9407182,3.5314875,3.9975388,4.273231,4.4242053,4.673641,4.6802053,4.650667,4.70318,4.824616,4.8705645,4.9099493,5.0510774,4.9329233,4.4734364,3.8564105,3.5971284,3.436308,3.3805132,3.3280003,3.0982566,2.930872,2.9243078,2.9144619,2.858667,2.8225644,2.9111798,3.1540515,3.3641028,3.442872,3.373949,4.2896414,5.3037953,7.250052,10.138257,13.161027,15.442053,17.831387,19.662771,20.54236,20.378258,21.927387,21.848618,20.201027,18.034874,17.401438,23.70954,31.149952,39.5159,48.653133,58.459904,69.645134,77.34811,74.0398,60.5079,45.853542,44.100925,45.167595,47.166363,47.957336,45.1479,47.22872,54.898876,67.8039,82.82585,94.06032,92.37334,88.428314,85.61231,85.819084,89.46216,91.34934,91.4117,91.25088,91.864624,93.650055,84.78524,77.952,73.419495,69.93067,64.66626,57.028927,50.835697,46.15221,42.39426,38.327797,29.282463,22.82995,19.74154,19.416616,19.86954,17.460514,12.84595,8.470975,5.586052,4.2371287,2.6551797,2.5206156,3.1343591,3.7415388,3.5249233,3.8104618,3.6890259,2.7470772,1.3423591,0.6170257,0.33476925,0.3117949,0.4955898,0.65312827,0.380718,0.67282057,1.024,1.1027694,0.9124103,0.7844103,0.892718,1.0108719,0.9714873,0.75487185,0.47917953,0.21989745,0.068923086,0.009846155,0.013128206,0.013128206,0.02297436,0.068923086,0.27569234,0.6432821,1.0633847,1.5261539,2.3893335,3.255795,3.4855387,2.1989746,0.9682052,0.39384618,0.16738462,0.07548718,0.036102567,0.03938462,0.06235898,0.19364104,1.3029745,5.031385,7.259898,10.230155,14.381949,17.660719,15.540514,9.878975,5.35959,2.793026,1.8412309,1.020718,0.46933338,0.256,0.21333335,0.21661541,0.18707694,0.2231795,0.28882053,0.31507695,0.27569234,0.18379489,0.13784617,0.12471796,0.118153855,0.10502565,0.09189744,0.09189744,0.0951795,0.0951795,0.101743594,0.14441027,0.11158975,0.14441027,0.16410258,0.14769232,0.14769232,0.17394873,0.17066668,0.14769232,0.128,0.14441027,0.16082053,0.16738462,0.18379489,0.21333335,0.25271797,0.2231795,0.18051283,0.15753847,0.16738462,0.21333335,2.1825643,2.1464617,1.972513,2.2383592,2.8980515,3.2656412,1.5425643,0.7384616,0.29210258,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.12471796,0.35774362,0.6268718,0.67282057,0.37415388,0.2231795,0.45292312,1.0371283,1.0732309,1.0371283,1.2832822,1.4342566,0.39712822,0.10502565,0.013128206,0.0,0.0,0.0,0.36758977,0.90584624,1.6869745,2.2514873,1.6180514,2.1169233,1.7132308,1.4145643,1.4572309,1.2964103,1.2373334,1.2832822,1.401436,1.657436,2.2416413,3.0490258,5.1364107,6.6067696,7.066257,7.6143594,8.713847,8.914052,9.110975,9.107693,7.6307697,12.133744,9.724719,6.245744,4.6178465,4.8377438,4.44718,4.138667,3.4921029,2.540308,1.7690258,1.4145643,1.2274873,1.0075898,0.72861546,0.5349744,0.827077,1.2931283,1.5622566,1.6508719,1.9692309,2.2744617,2.4582565,3.761231,5.225026,3.7218463,1.6836925,1.5130258,2.044718,2.172718,0.8533334,0.65969235,0.892718,0.9189744,0.571077,0.16738462,0.4135385,0.6301539,0.92225647,1.2898463,1.6311796,2.1333334,2.156308,2.1464617,2.4352822,3.2656412,2.4352822,4.332308,6.7150774,7.5881033,5.2348723,5.8814363,6.3901544,6.1341543,5.5893335,6.3474874,5.799385,5.284103,3.9778464,2.2482052,1.6640002,1.4441026,1.5425643,1.8445129,2.1333334,2.1202054,3.1573336,4.9920006,5.5171285,4.565334,3.9056413,3.0391798,2.5107694,2.0118976,1.5163078,1.2964103,1.4441026,2.0939488,2.8324106,3.31159,3.249231,6.180103,5.9963083,6.1440005,7.2631803,7.200821,7.6898465,8.178872,8.421744,8.149334,7.0498466,6.695385,5.3169236,4.6933336,5.1922054,5.7534366,6.058667,5.5302567,5.3169236,5.4941545,5.0674877,4.457026,6.308103,7.857231,7.755488,6.058667,5.156103,4.013949,3.190154,2.6453335,1.7558975,2.097231,2.2744617,2.8160002,3.1737437,1.7099489,2.4155898,3.4822567,4.4274874,5.280821,6.560821,6.62318,4.778667,3.1245131,2.6945643,3.4625645,3.757949,6.439385,8.576,9.074872,8.697436,6.928411,7.6110773,9.521232,11.23118,11.109744,8.923898,5.602462,5.1626673,9.124104,16.508718,27.654566,28.901747,23.397745,15.241847,9.504821,8.004924,7.7292314,7.9819493,8.743385,10.696206,13.686155,12.137027,8.67118,5.874872,6.301539,4.788513,4.07959,3.8071797,4.069744,5.4613338,6.232616,5.481026,5.211898,5.72718,5.6320004,6.166975,6.997334,7.3649235,7.02359,6.242462,8.963283,8.756514,8.713847,9.202872,7.8736415,5.408821,4.132103,4.637539,5.8486156,5.0051284,4.516103,5.100308,5.674667,5.4908724,4.135385,4.634257,4.020513,2.934154,2.1070771,2.349949,3.629949,4.4012313,4.266667,3.6102567,3.5872824,4.086154,4.1485133,3.8859491,3.4198978,2.8849232,3.9089234,4.962462,5.0116925,4.2535386,4.1189747,3.7415388,3.2361028,2.8750772,2.6551797,2.28759,1.8248206,1.6278975,1.6278975,1.723077,1.785436,1.2603078,1.2471796,1.522872,1.9331284,2.3958976,3.1409233,3.4724104,3.0227695,2.0709746,1.5721027,1.5589745,1.6935385,1.913436,1.9659488,1.404718,1.1979488,1.3554872,1.6475899,1.9364104,2.1825643,1.9626669,2.281026,2.4057438,2.3663592,2.9768207,3.3411283,2.930872,2.3138463,1.8576412,1.723077,2.6518977,2.7733335,2.6026669,2.5993848,3.1737437,2.4549747,1.7887181,1.6968206,2.2383592,3.006359,3.1638978,2.3893335,1.4244103,0.8205129,0.9321026,0.9682052,1.1782565,1.3981539,2.3138463,5.4613338,8.585847,8.700719,7.9130263,6.8955903,4.8672824,5.0018463,7.059693,9.780514,11.30995,9.186462,6.672411,6.3277955,6.0685134,6.806975,12.419283,7.5618467,6.51159,7.128616,7.6996927,6.941539,5.904411,5.9930263,5.4186673,3.7907696,2.1070771,1.2898463,2.156308,2.6978464,2.2613335,1.5425643,3.7251284,14.076719,26.784822,35.813747,34.911182,33.690258,25.465437,21.097027,20.105848,10.679795,4.2371287,3.9253337,4.397949,3.436308,1.9692309,3.8367183,4.010667,2.7733335,1.6377437,3.3575387,5.1889234,2.8455386,1.0929232,1.7001027,3.4330258,5.8978467,8.87795,11.588924,13.5089245,14.388514,13.436719,11.457642,13.771488,21.83549,33.24718,32.613747,25.094566,15.261539,6.8004107,2.5042052,3.2722054,3.4264617,4.4898467,6.488616,7.965539,6.2785645,3.0490258,0.7975385,0.25928208,0.380718,0.45620516,0.46276927,0.446359,0.38728207,0.2297436,0.21661541,0.15753847,0.15753847,0.2100513,0.19692309,0.07548718,0.118153855,0.41682056,0.77128214,0.6859488,0.45620516,0.2231795,0.16738462,0.3708718,0.82379496,1.1782565,1.5589745,1.7788719,1.6640002,1.0535386,1.332513,1.9167181,2.556718,3.117949,3.570872,4.1682053,4.9854364,5.933949,6.8332314,7.430565,5.5007186,3.3280003,2.0808206,2.1234872,2.989949,6.0192823,7.9195905,8.67118,8.342975,7.1122055,4.850872,4.9920006,6.196513,8.274052,12.1928215,11.201642,7.5881033,4.7917953,4.007385,4.164923,3.1507695,2.3762052,2.2055387,2.8258464,4.240411,4.630975,5.106872,5.405539,5.674667,6.4557953,6.47877,6.0258465,5.612308,5.5532312,5.979898,5.835488,6.1374364,6.449231,6.6461544,6.928411,6.3179493,5.723898,5.0215387,4.0992823,2.8521028,2.2547693,2.5829747,2.5632823,2.0512822,2.0151796,2.3794873,2.674872,2.7470772,2.6945643,2.8521028,2.8422565,3.242667,3.698872,3.9318976,3.7218463,3.186872,2.858667,2.5665643,2.2580514,2.0151796,2.3696413,2.428718,2.3072822,2.1333334,2.0611284,1.8149745,1.7001027,1.723077,1.7723079,1.6016412,1.4572309,1.7132308,1.8412309,1.7755898,1.9232821,3.6562054,5.792821,8.300308,11.0375395,13.748514,16.164104,17.99549,18.228514,16.850052,14.8480015,17.129026,18.267899,16.856617,13.410462,10.345026,13.617231,20.742565,29.879797,38.452515,43.152412,50.051285,53.71734,51.61026,44.035286,34.133335,38.114464,43.897438,48.180515,49.726364,49.345646,51.557747,64.19365,90.71262,122.246574,137.61642,135.27304,130.19241,121.49827,111.70134,106.67324,114.85211,122.49929,121.93806,113.581955,105.941345,94.97929,88.257645,85.40555,84.88042,83.9516,74.528824,63.678364,53.441647,48.278976,55.05313,49.375183,41.10113,32.836926,27.451078,28.06154,27.585644,22.09149,15.189335,9.803488,8.178872,4.821334,4.4406157,5.0215387,5.1856413,4.197744,3.2328207,2.5042052,1.719795,0.9353847,0.58092314,0.5316923,0.508718,0.6432821,0.8336411,0.74830776,1.4178462,2.428718,3.0030773,2.737231,1.6016412,1.1749744,1.0765129,1.0272821,0.88287187,0.6268718,0.40697438,0.16738462,0.026256412,0.0,0.0,0.0,0.009846155,0.016410258,0.02297436,0.06235898,0.18379489,0.2231795,0.2297436,0.20676924,0.12143591,0.072205134,0.13456412,0.13456412,0.049230773,0.0,0.013128206,0.016410258,0.02297436,0.7122052,3.4330258,3.4330258,5.402257,9.156924,13.24636,14.953027,10.535385,6.4623594,4.4110775,3.8662567,2.1202054,0.86317956,0.29210258,0.10502565,0.07548718,0.07548718,0.11158975,0.2231795,0.28225642,0.256,0.18379489,0.14769232,0.09189744,0.06235898,0.06564103,0.09189744,0.14112821,0.13456412,0.13456412,0.21661541,0.47261542,0.26584616,0.23958977,0.23630771,0.19692309,0.18379489,0.17066668,0.15753847,0.14769232,0.14441027,0.16738462,0.15425642,0.17066668,0.19692309,0.21661541,0.2297436,0.18051283,0.14112821,0.14112821,0.16410258,0.15097436,3.6594875,1.0732309,0.39384618,0.44964105,0.58092314,0.65312827,0.30851284,0.14769232,0.059076928,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03938462,0.15097436,0.27897438,0.28225642,0.21661541,0.17394873,0.13784617,0.13456412,0.23302566,0.34789747,0.41025645,0.42338464,0.34789747,0.09189744,0.02297436,0.0032820515,0.0,0.013128206,0.06235898,2.2908719,3.0424619,2.3302567,1.1290257,1.3718976,1.7460514,1.3226668,0.9911796,0.97805136,0.86974365,0.9747693,1.3718976,1.5425643,1.4867693,1.7296412,3.308308,6.114462,8.224821,9.015796,9.163487,8.700719,7.5520005,6.6822567,6.9152827,8.937026,10.197334,8.41518,6.5870776,5.7829747,5.142975,4.4307694,3.761231,3.1113849,2.4943593,1.9889232,1.7624617,1.4966155,1.2373334,1.079795,1.1552821,1.204513,1.0994873,1.1290257,1.591795,2.7995899,4.7327185,3.7743592,2.9768207,3.3411283,3.820308,2.2121027,1.4441026,1.5327181,1.972513,1.7591796,1.8149745,1.1618463,0.6498462,0.6432821,1.020718,1.0043077,0.9124103,1.0108719,1.2471796,1.2668719,1.0436924,0.8369231,0.9124103,1.3817437,2.1924105,2.993231,5.1364107,6.5312824,6.452513,5.549949,6.560821,6.5805135,6.232616,6.042257,6.4590774,5.7042055,5.028103,4.4274874,3.9253337,3.6036925,2.3696413,2.1924105,2.1891284,2.0939488,2.2678976,2.934154,4.9099493,5.5072823,4.3618464,3.4297438,2.681436,2.1234872,2.228513,2.7044106,2.5042052,2.0939488,2.8553848,4.2272825,5.1232824,3.9089234,6.301539,6.672411,6.1505647,5.6385646,5.8223596,6.4590774,6.5870776,6.8594875,7.2237954,6.9152827,6.7774363,7.4929237,6.9087186,5.5597954,6.669129,6.114462,4.8082056,4.4373336,5.720616,8.39877,6.265436,5.3202057,5.8190775,6.629744,5.21518,5.474462,4.8344617,3.6102567,2.3105643,1.6443079,1.5261539,1.6475899,2.7470772,3.882667,2.4155898,2.3138463,2.6945643,3.318154,4.450462,6.8660517,6.633026,4.571898,3.2164104,3.3345644,3.9286156,3.7710772,4.4964104,5.356308,6.226052,7.5881033,7.565129,9.235693,11.490462,13.138052,12.87877,10.732308,9.93477,12.1468725,16.981335,22.002874,22.57067,18.907898,14.25395,10.499283,8.139488,8.503796,8.956718,9.110975,8.956718,8.891078,10.230155,9.26195,7.076103,4.886975,4.056616,4.6605134,5.7074876,7.312411,8.411898,6.7577443,5.024821,4.850872,5.3234878,5.8190775,5.98318,7.4010262,6.948103,6.426257,7.1647186,10.023385,10.06277,7.7259493,7.506052,9.363693,8.726975,6.009436,6.38359,8.4512825,10.003693,8.021334,5.7435904,5.7403083,5.7731285,5.3136415,5.549949,6.012718,5.5630774,4.33559,3.2065644,3.8038976,4.673641,4.7983594,4.565334,4.3684106,4.598154,4.161641,4.1124105,4.6802053,5.4580517,5.398975,4.197744,3.6332312,3.7251284,4.342154,5.1954875,4.31918,3.6857438,3.3805132,3.2164104,2.7536411,2.1431797,1.8281027,1.7329233,1.6672822,1.2964103,1.1520001,1.0732309,1.0601027,1.1684103,1.5031796,2.169436,2.5731285,2.5796926,2.2744617,1.9495386,1.6640002,1.4211283,1.2242053,1.0994873,1.1355898,1.3193847,1.6344616,2.2547693,3.0030773,3.367385,2.930872,2.487795,2.2744617,2.2777438,2.2416413,1.9462565,1.9003079,2.3433847,3.114667,3.6660516,3.1967182,2.8160002,2.4188719,2.1234872,2.2580514,1.4408206,1.0010257,0.8730257,0.9747693,1.1881026,1.1618463,1.394872,2.0250258,3.6463592,7.3025646,6.0291286,5.028103,4.6080003,6.0685134,11.687386,15.593027,12.166565,6.994052,4.6605134,8.736821,10.601027,13.587693,15.353437,15.648822,16.324924,13.059283,9.780514,6.770872,4.8607183,5.4383593,4.4865646,5.349744,6.157129,6.045539,5.159385,4.092718,3.515077,2.8980515,2.2613335,2.1792822,1.6836925,3.9056413,9.042052,13.3940525,9.353847,6.557539,12.970668,22.15713,28.488207,27.136002,19.8039,14.145642,10.482873,7.860513,4.0533338,2.2744617,2.5665643,3.0260515,2.865231,2.3958976,2.172718,1.5622566,0.88943595,0.5218462,0.86646163,1.1454359,0.6826667,0.9714873,1.975795,2.1267693,5.8125134,7.003898,10.692924,16.367592,17.979078,13.636924,11.280411,14.221129,20.230566,21.56636,17.913437,13.193847,8.27077,4.0467696,1.4276924,1.2898463,2.793026,3.6102567,3.1277952,2.4484105,2.481231,3.6036925,2.7503593,0.3117949,0.16082053,0.23630771,0.24287182,0.21661541,0.16082053,0.068923086,0.059076928,0.036102567,0.032820515,0.04266667,0.03938462,0.08205129,0.190359,0.23630771,0.20020515,0.17394873,0.27569234,0.19692309,0.108307704,0.118153855,0.2855385,0.4266667,0.6071795,0.75487185,0.86646163,1.017436,1.083077,1.4736412,1.8215386,2.3794873,4.023795,4.6605134,3.8990772,3.2065644,3.1770258,3.511795,3.2623591,3.1409233,3.1507695,3.2853336,3.5282054,3.751385,5.3103595,6.3376417,6.626462,7.6603084,6.445949,5.3694363,5.0084105,5.681231,7.430565,8.474257,9.179898,8.070564,5.83877,5.3727183,4.4373336,4.0500517,4.141949,4.516103,4.841026,5.1331286,4.6572313,4.4701543,4.8771286,5.4547696,4.919795,4.821334,4.844308,5.0904617,6.055385,6.229334,6.5312824,6.741334,6.701949,6.3179493,4.955898,3.383795,2.3926156,2.0151796,1.5097437,1.6147693,2.0020514,1.7920002,1.148718,1.270154,1.6640002,2.097231,2.3762052,2.3991797,2.156308,1.9298463,1.8084104,1.6902566,1.5491283,1.4276924,1.595077,1.7591796,1.8281027,1.8116925,1.8313848,2.5173335,2.6912823,2.674872,2.6617439,2.7076926,2.7963078,2.7766156,2.6584618,2.4418464,2.1136413,1.9889232,1.9265642,1.8248206,1.8937438,2.6551797,6.0980515,9.655796,13.00677,15.862155,17.99549,18.888206,17.417847,14.201437,10.262975,7.02359,7.899898,9.147078,9.744411,9.189744,7.512616,8.674462,12.2847185,19.465847,28.360207,34.14318,38.334362,38.498463,35.140926,30.592003,28.983797,33.939693,39.79159,45.42359,50.093952,53.43508,57.472004,69.986465,92.3077,119.38134,139.7793,149.85847,157.33499,155.59879,145.15529,133.66154,114.37949,111.19591,107.48062,96.03939,79.11057,74.85703,72.88123,73.66893,76.38975,78.90052,76.9477,72.64821,63.888416,54.304825,53.297234,61.11508,62.5559,56.155903,45.380928,38.6199,37.888004,35.108105,27.91713,17.742771,9.7903595,8.677744,8.162462,8.3134365,8.192,5.85518,3.6726158,2.2678976,1.6738462,1.8970258,2.9111798,2.9013336,2.4648206,2.0775387,1.8445129,1.5031796,1.5983591,2.6551797,3.9286156,4.338872,2.481231,1.3784616,0.9616411,0.7975385,0.6629744,0.5021539,0.3511795,0.19692309,0.07548718,0.009846155,0.0,0.0,0.0032820515,0.0032820515,0.0032820515,0.013128206,0.04594872,0.101743594,0.12471796,0.10502565,0.049230773,0.049230773,0.16738462,0.15753847,0.02297436,0.013128206,0.0032820515,0.0032820515,0.0032820515,0.16410258,0.7975385,1.0108719,2.044718,3.508513,4.841026,5.3103595,3.9876926,2.917744,2.8521028,3.2098465,2.0611284,0.71548724,0.20348719,0.072205134,0.049230773,0.03938462,0.055794876,0.08861539,0.10502565,0.10502565,0.108307704,0.101743594,0.08533334,0.068923086,0.06564103,0.07876924,0.13784617,0.18707694,0.26256412,0.3446154,0.33805132,0.25928208,0.23630771,0.21989745,0.2100513,0.256,0.36102566,0.36430773,0.30194873,0.23630771,0.23958977,0.2100513,0.20348719,0.23958977,0.27897438,0.25271797,0.16410258,0.12471796,0.128,0.16082053,0.190359,1.6114873,0.32164106,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02297436,0.068923086,0.10502565,0.07876924,0.049230773,0.07548718,0.20020515,0.45292312,0.8533334,0.50543594,0.29210258,0.13784617,0.029538464,0.006564103,0.0,0.0,0.0032820515,0.06235898,0.27897438,1.723077,2.6683078,2.6486156,1.8510771,1.1290257,1.0765129,0.88287187,0.81394875,0.8566154,0.73517954,1.020718,1.975795,3.0720003,3.7152824,3.2131286,4.20759,5.4416413,6.0160003,6.045539,6.6592827,7.3419495,6.5050263,5.402257,5.0904617,6.422975,6.7150774,6.38359,6.2030773,6.2916927,6.088206,5.0674877,4.0008206,3.2032824,2.8389745,2.934154,2.3433847,1.6804104,1.211077,1.0305642,1.083077,1.9265642,2.3368206,1.9987694,1.7329233,3.4921029,3.9745643,3.1113849,2.359795,2.4681027,3.4527183,2.9833848,2.2416413,1.8707694,2.0644104,2.5796926,2.2186668,1.3456411,1.0404103,1.3751796,1.4276924,1.2537436,1.401436,1.6836925,1.8838975,1.7427694,1.339077,1.1454359,1.3095386,1.6508719,1.657436,3.4231799,4.7392826,5.3891287,5.7796926,6.948103,8.024616,7.8047185,7.6570263,7.7456417,6.997334,5.737026,4.97559,4.7327185,5.031385,5.901129,4.896821,3.9614363,3.0916924,2.487795,2.5238976,3.259077,3.876103,4.2240005,4.3684106,4.57518,3.8400004,2.9078977,2.612513,3.0358977,3.5216413,3.2065644,4.3585644,6.117744,7.2172313,5.976616,6.7216415,6.918565,6.6002054,6.265436,6.8693337,6.948103,6.1472826,5.5565133,5.691077,6.488616,7.8736415,9.353847,9.412924,8.605539,9.544206,9.4916935,7.702975,6.0225644,5.674667,7.253334,5.435077,3.8695388,4.0434875,5.225026,4.4832826,4.709744,4.1780515,3.2623591,2.4188719,2.176,1.9429746,2.028308,3.190154,4.315898,2.4188719,2.5337439,3.058872,3.5314875,4.2141542,6.091488,6.994052,5.4580517,4.2371287,4.201026,4.3552823,3.9023592,4.3618464,5.284103,6.4590774,7.893334,9.107693,11.346052,12.737642,12.550565,11.188514,10.9915905,11.995898,14.55918,17.371899,17.444103,14.953027,12.038565,9.4457445,7.748924,7.3747697,8.549745,8.303591,7.686565,7.6931286,9.235693,10.676514,9.816616,8.297027,7.000616,6.058667,5.874872,7.0990777,9.481847,11.004719,7.8769236,5.5630774,5.720616,6.3212314,7.0400004,9.248821,10.482873,8.395488,7.2205133,9.344001,15.320617,11.835078,7.4436927,5.927385,7.427283,8.418462,6.0685134,5.7074876,6.5870776,7.5881033,7.207385,6.413129,6.377026,6.1308722,5.5105643,5.1626673,5.211898,4.916513,4.2896414,3.6168208,3.442872,3.6693337,4.023795,4.1517954,4.1091285,4.3585644,4.713026,5.579488,5.933949,5.533539,4.919795,3.892513,3.0949745,3.058872,3.6430771,4.023795,3.3542566,3.2689233,3.4855387,3.5741541,2.9702566,2.2416413,1.8674873,1.6935385,1.5622566,1.2832822,1.3226668,0.99774367,0.77128214,0.86317956,1.2635899,1.7362052,1.8018463,1.7329233,1.654154,1.5491283,1.5327181,1.7755898,1.9495386,2.038154,2.3302567,2.281026,2.4451284,2.6584618,2.930872,3.4231799,3.1277952,2.665026,2.2022567,1.8445129,1.657436,1.9856411,2.1267693,2.4943593,3.0227695,3.1803079,2.5961027,2.4451284,2.4484105,2.487795,2.6157951,2.1333334,1.723077,1.4736412,1.4802053,1.8313848,4.312616,6.2063594,7.174565,7.680001,8.969847,6.806975,5.3760004,5.159385,7.0367184,12.301129,15.379693,12.370052,7.9261546,5.930667,9.511385,10.512411,11.881026,13.545027,15.753847,19.072002,18.504206,16.810667,12.435693,6.7905645,4.2601027,5.10359,7.1581545,8.480822,8.041026,5.7042055,5.5597954,5.5696416,5.7074876,6.262154,7.8539495,7.00718,8.251078,14.795488,22.514874,19.968002,10.19077,9.7673855,12.849232,14.956308,12.970668,7.5881033,4.900103,3.387077,2.28759,1.6278975,1.7427694,2.3827693,2.9538465,3.0030773,2.228513,1.4605129,0.8172308,0.67938465,0.80738467,0.3446154,0.16082053,0.12471796,0.7417436,1.6968206,1.8543591,8.54318,9.442462,10.134975,12.07795,12.603078,8.530052,7.3091288,9.110975,11.644719,10.161232,7.1515903,4.8377438,3.4888208,2.9210258,2.4976413,2.7963078,2.865231,2.3269746,1.394872,0.8402052,1.0896411,1.9593848,1.7558975,0.58092314,0.318359,0.16410258,0.0951795,0.06235898,0.04266667,0.013128206,0.006564103,0.0032820515,0.0,0.01969231,0.101743594,0.39056414,0.32164106,0.14769232,0.026256412,0.036102567,0.21989745,0.18707694,0.128,0.12471796,0.18051283,0.20020515,0.23630771,0.32820517,0.4660513,0.60389745,0.8008206,1.1585642,1.5556924,2.1267693,3.2853336,3.6824617,3.7316926,3.6791797,3.508513,2.934154,3.2229745,3.820308,4.352,4.6211286,4.604718,4.972308,6.242462,6.747898,6.3901544,6.6625648,6.091488,5.5105643,5.149539,5.074052,5.1987696,6.4032826,7.6012316,7.282872,5.832206,5.5105643,5.041231,5.277539,5.76,6.340924,7.1876926,6.5772314,6.2162056,5.9963083,5.858462,5.799385,5.037949,4.8836927,4.916513,5.1265645,5.917539,6.2752824,5.7403083,5.106872,4.598154,3.8564105,2.7175386,1.7624617,1.2898463,1.3456411,1.7165129,1.7329233,1.7788719,1.5064616,1.0535386,1.0732309,1.1848207,1.2931283,1.3653334,1.3554872,1.1979488,1.083077,1.0371283,0.9616411,0.86646163,0.86317956,0.97805136,1.1191796,1.2603078,1.4605129,1.8773335,2.6157951,3.0358977,3.370667,3.6069746,3.4822567,3.314872,3.3214362,3.2065644,2.9669745,2.8553848,2.7109745,2.7306669,2.7011285,2.681436,3.0030773,5.208616,8.1066675,12.035283,16.15754,18.464823,16.758156,13.124924,8.848411,5.169231,3.2722054,3.8859491,4.886975,5.7435904,6.0717955,5.6352825,6.232616,8.78277,13.968411,20.578463,25.527798,28.691694,28.967386,27.51672,26.230156,27.703796,32.134567,35.728413,38.994053,42.738876,48.08862,55.230362,68.64739,87.41088,108.07468,124.67529,136.84842,147.09827,147.37724,136.13293,118.31139,99.33457,89.52452,81.47037,70.38031,54.065235,54.69211,62.336006,78.011086,96.48575,106.30893,102.334366,94.69375,83.03262,70.482056,63.678364,67.40021,66.907906,58.771698,45.71898,36.627697,34.192413,30.972721,25.947899,19.971283,15.766975,14.060308,12.20595,10.971898,10.026668,7.936001,4.670359,2.7109745,1.8871796,2.0545642,3.0654361,4.8377438,3.7382567,2.4648206,2.0578463,1.9035898,1.8346668,2.484513,3.239385,3.3805132,2.0873847,1.2800001,0.9321026,0.764718,0.62030774,0.46276927,0.35774362,0.23302566,0.10502565,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.029538464,0.04266667,0.055794876,0.10502565,0.6662565,0.5284103,0.20676924,0.006564103,0.006564103,0.0,0.006564103,0.009846155,0.02297436,0.08205129,0.24943592,0.67610264,1.1191796,1.4178462,1.4802053,1.2012309,1.0272821,1.1782565,1.3981539,0.955077,0.34133336,0.128,0.068923086,0.03938462,0.013128206,0.02297436,0.029538464,0.03938462,0.055794876,0.06564103,0.06564103,0.072205134,0.07876924,0.07876924,0.07548718,0.19692309,0.3314872,0.4201026,0.4266667,0.3708718,0.38728207,0.42994875,0.44307697,0.42338464,0.44964105,0.48902568,0.4594872,0.40697438,0.380718,0.43323082,0.33805132,0.29210258,0.26584616,0.23958977,0.20348719,0.15097436,0.17394873,0.21661541,0.23302566,0.190359,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.006564103,0.0,0.0,0.026256412,0.052512825,0.25271797,0.7056411,1.404718,0.761436,0.2986667,0.059076928,0.0,0.0,0.01969231,0.15097436,0.43323082,0.7450257,0.81394875,1.3850257,2.156308,2.4582565,2.0184617,0.96492314,0.69251287,0.7844103,1.2504616,1.6311796,1.0108719,1.0469744,2.3433847,3.7842054,4.31918,2.9636924,3.2525132,3.3509746,3.0687182,2.8521028,3.7776413,5.156103,5.2020516,4.7950773,4.562052,4.8738465,4.6769233,5.0018463,5.4482055,5.756718,5.8125134,5.097026,4.2305646,3.4888208,3.0949745,3.2262566,2.4549747,1.654154,1.1323078,0.9517949,0.9321026,1.8445129,2.3827693,2.03159,1.5163078,2.8127182,2.92759,2.9505644,2.5928206,2.2350771,2.9505644,3.121231,2.6584618,2.176,2.0512822,2.4385643,2.0709746,1.9068719,1.8937438,1.8707694,1.5688206,1.4244103,1.5327181,1.7033848,1.8248206,1.8576412,1.6935385,1.8051283,1.9232821,1.9200002,1.8084104,3.4297438,3.7776413,3.8990772,4.6933336,6.9120007,7.653744,7.466667,7.936001,8.937026,8.644924,7.653744,7.062975,6.9677954,7.213949,7.3714876,6.0750775,4.6080003,3.4560003,2.7963078,2.5107694,3.3345644,3.43959,3.7907696,4.601436,5.3366156,4.9887185,4.315898,3.6430771,3.442872,4.338872,4.900103,6.2030773,7.1548724,7.1187696,5.924103,5.533539,5.477744,5.5302567,5.8092313,6.7971287,7.8014364,7.2270775,6.921847,7.499488,8.342975,8.805744,8.953437,8.707283,8.572719,9.622975,10.811078,9.5606165,7.53559,5.986462,5.733744,3.9548721,2.8488207,3.0654361,4.013949,3.879385,3.6824617,3.1048207,2.5337439,2.1825643,2.0841026,1.9889232,2.041436,3.0523078,4.1156926,2.6322052,3.1015387,3.2262566,3.1540515,3.4166157,4.9329233,6.8594875,5.8125134,4.6244106,4.33559,4.1911798,3.9089234,5.100308,6.3540516,7.0859494,7.529026,9.517949,11.641437,12.258463,11.152411,9.521232,10.794667,13.305437,15.379693,15.563488,12.635899,10.893129,9.885539,8.743385,7.496206,7.1023593,8.129642,7.3780518,6.7872825,7.4010262,9.373539,10.834052,9.672206,8.247795,7.4863596,6.882462,6.0947695,6.9152827,8.605539,9.501539,7.0104623,5.658257,6.058667,6.5280004,7.433847,11.191795,11.900719,8.960001,7.3386674,9.590155,15.839181,11.782565,7.243488,5.1659493,6.298257,9.176616,8.753231,8.004924,7.1056414,6.314667,5.9634876,7.02359,7.634052,7.273026,6.124308,5.0543594,4.824616,4.345436,3.9023592,3.5282054,3.0096412,3.383795,4.6966157,6.0783596,6.6494365,5.536821,5.4908724,7.427283,8.018052,6.3606157,3.9909747,3.6463592,3.1409233,2.9078977,2.9243078,2.7175386,2.6518977,3.1048207,3.498667,3.4297438,2.665026,1.9626669,1.6246156,1.4933335,1.4178462,1.2668719,1.2504616,0.92553854,0.7975385,1.0272821,1.3981539,1.5622566,1.3423591,1.1684103,1.1749744,1.2012309,1.3751796,2.044718,2.793026,3.3017437,3.3575387,2.7076926,2.487795,2.3893335,2.4746668,3.1671798,3.1048207,2.8750772,2.4155898,1.9167181,1.8281027,2.6322052,2.9111798,3.121231,3.3411283,3.2525132,2.8750772,2.793026,2.8553848,2.9243078,2.865231,2.8258464,2.8127182,2.865231,3.0293336,3.3509746,5.8880005,7.722667,8.342975,7.8047185,6.7117953,4.824616,3.7284105,3.6857438,5.106872,8.55959,11.247591,10.315488,9.005949,8.677744,8.79918,7.571693,8.132924,10.640411,14.450873,18.120207,18.36308,17.539284,13.436719,7.6734366,5.6943593,6.675693,7.6931286,7.90318,7.0432825,5.421949,5.832206,7.460103,9.012513,9.8592825,10.059488,8.851693,9.488411,14.03077,19.643078,18.609232,9.133949,5.930667,5.802667,5.8847184,3.626667,2.1103592,2.1497438,2.5961027,3.121231,4.2338467,3.882667,3.2722054,2.8521028,2.540308,1.719795,1.1290257,0.6071795,0.54482055,0.71548724,0.25271797,0.118153855,0.07548718,0.380718,0.9485129,1.3554872,7.643898,9.009232,7.975385,6.518154,6.0717955,3.7448208,3.3312824,3.7973337,4.0500517,2.92759,1.5491283,0.9485129,1.1913847,1.9692309,2.5895386,4.388103,3.892513,2.4910772,1.1782565,0.5513847,0.5415385,0.508718,0.52512825,0.5284103,0.32820517,0.11158975,0.02297436,0.0,0.0,0.0,0.0,0.0,0.0,0.02297436,0.108307704,0.36758977,0.24615386,0.108307704,0.10502565,0.15097436,0.18051283,0.12471796,0.098461546,0.16082053,0.3314872,0.34133336,0.28225642,0.24615386,0.25271797,0.23302566,0.52512825,0.8402052,1.1815386,1.6377437,2.3794873,2.8356924,4.06318,4.699898,4.4012313,3.826872,3.9056413,4.4406157,4.972308,5.353026,5.7698464,6.5312824,7.515898,7.6242056,6.6461544,5.2644105,5.32677,5.618872,5.7665644,5.668103,5.4908724,6.0160003,6.62318,6.7610264,6.701949,7.5388722,6.157129,6.0160003,6.616616,7.5881033,8.694155,7.50277,7.1548724,6.918565,6.49518,6.0291286,4.709744,4.3552823,4.5029745,4.772103,4.8607183,4.522667,3.4789746,2.605949,2.103795,1.5195899,1.0305642,0.83035904,0.80738467,0.96492314,1.4276924,1.2996924,1.1749744,0.97805136,0.75487185,0.67610264,0.6104616,0.5284103,0.46933338,0.43651286,0.4135385,0.4201026,0.48246157,0.5218462,0.5284103,0.55794877,0.574359,0.65312827,0.78769237,1.0404103,1.5360001,2.1464617,2.8914874,3.7809234,4.453744,4.1583595,4.2141542,4.2535386,4.141949,3.9745643,4.082872,3.9581542,3.9909747,3.9811285,3.895795,3.8498464,4.5587697,5.901129,8.470975,11.634872,13.515489,11.172104,7.7259493,4.6867695,2.878359,2.4484105,2.8750772,3.3411283,3.7940516,4.2338467,4.7228723,6.426257,10.043077,14.519796,18.786463,21.766565,23.906464,24.42831,24.320002,24.65149,26.551796,29.663181,31.153233,32.36431,34.87508,40.493954,48.610466,60.622772,76.95098,95.49129,111.612724,128.24945,137.26524,135.07283,121.85929,101.56309,85.179085,70.02914,57.475285,47.9639,41.00267,47.481438,62.588722,87.59467,116.371704,135.41089,126.56247,115.77109,103.51263,90.81437,79.24185,73.32431,66.63221,54.41313,39.007183,29.817438,25.793644,22.468925,20.128822,18.95713,19.058874,18.17272,16.741745,15.143386,13.436719,11.355898,7.830975,5.182359,3.5216413,2.7864618,2.7273848,4.6178465,3.4166157,2.1333334,1.847795,1.7099489,1.7394873,2.0151796,2.1300514,1.9593848,1.6246156,1.3784616,1.1618463,0.9321026,0.71548724,0.6301539,0.8402052,0.508718,0.17066668,0.04266667,0.006564103,0.006564103,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.026256412,0.09189744,0.6662565,0.4660513,0.14441027,0.0,0.0,0.0,0.006564103,0.009846155,0.013128206,0.026256412,0.101743594,0.21989745,0.318359,0.36430773,0.3708718,0.30194873,0.24287182,0.21333335,0.19692309,0.15097436,0.08205129,0.128,0.128,0.052512825,0.013128206,0.013128206,0.016410258,0.01969231,0.029538464,0.032820515,0.03938462,0.055794876,0.068923086,0.07876924,0.07548718,0.2100513,0.4004103,0.54482055,0.5907693,0.5513847,0.6629744,0.8467693,0.90912825,0.827077,0.74830776,0.761436,0.73517954,0.6826667,0.6432821,0.6892308,0.52512825,0.42338464,0.3314872,0.23958977,0.16738462,0.13784617,0.17066668,0.21333335,0.2231795,0.16410258,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0,0.0,0.0,0.0032820515,0.013128206,0.13784617,0.14769232,0.24943592,0.56123084,1.142154,0.6498462,0.21989745,0.013128206,0.013128206,0.032820515,0.1148718,0.48902568,1.2832822,2.0545642,1.8051283,2.034872,2.176,1.8182565,1.1224617,0.82379496,0.67610264,0.9419488,1.8116925,2.5337439,1.4080001,0.90256417,1.9396925,2.7602053,2.484513,1.1257436,1.1585642,1.1749744,1.2307693,1.5163078,2.356513,3.2754874,4.135385,4.824616,5.395693,6.052103,5.930667,5.3070774,4.8016415,4.585026,4.381539,4.31918,4.1124105,3.6463592,3.0391798,2.6518977,2.041436,1.4802053,1.1323078,1.014154,0.9682052,1.1027694,1.211077,1.1979488,1.1618463,1.3915899,2.7700515,3.7284105,3.446154,2.4615386,2.6880002,2.8553848,2.5140514,2.1136413,1.8609232,1.6902566,1.7558975,2.5665643,2.740513,2.1070771,1.6804104,1.7165129,1.5360001,1.3554872,1.3554872,1.7033848,1.785436,2.2022567,2.103795,1.6869745,2.1956925,2.9669745,2.802872,2.674872,3.308308,5.182359,5.5072823,5.6418467,6.8004107,8.822155,10.194052,10.069334,9.961026,9.91836,9.363693,7.0990777,5.024821,3.69559,3.0916924,2.8225644,2.1333334,2.9636924,3.6004105,4.096,4.5095387,4.890257,5.7468724,5.7632823,4.8311796,3.8334363,4.6276927,6.2588725,7.141744,6.6592827,5.159385,3.9778464,3.5052311,3.3903592,3.4756925,3.892513,5.080616,7.7390776,8.267488,9.288206,10.932513,10.843898,8.39877,6.675693,5.651693,5.5762057,6.9645133,8.832001,8.553026,7.450257,6.294975,5.284103,3.058872,2.7602053,3.1967182,3.6332312,3.761231,3.1245131,2.5173335,2.1267693,1.9429746,1.7723079,1.8281027,1.6836925,2.297436,3.2820516,2.8947694,3.6036925,3.0326157,2.297436,2.353231,3.9909747,6.117744,5.536821,4.640821,4.309334,3.9318976,3.7054362,5.3891287,6.8463597,7.1647186,6.6494365,8.582564,9.941334,10.473026,10.203898,9.429334,10.538668,13.699283,15.514257,14.582155,11.503591,11.001437,10.912822,10.28595,8.986258,7.6996927,7.837539,7.2631803,7.3091288,8.044309,8.267488,8.845129,7.8014364,6.685539,6.0849237,5.6287184,5.398975,5.8486156,6.1440005,6.009436,5.733744,6.3573337,6.485334,6.186667,6.5837955,9.829744,10.499283,8.293744,6.5837955,7.3386674,11.132719,10.44677,8.533334,7.2237954,7.7981544,10.981745,13.082257,13.249642,11.37559,8.441437,6.5247183,8.188719,9.268514,8.848411,7.240206,6.0225644,5.297231,4.322462,3.570872,3.255795,3.3345644,4.4110775,6.6527185,9.284924,10.532104,7.6209235,6.038975,8.490667,9.816616,7.9458466,3.9023592,3.6693337,3.3608208,2.9538465,2.537026,2.3138463,2.802872,3.3903592,3.4724104,2.9078977,2.0217438,1.5130258,1.2800001,1.2242053,1.211077,1.0666667,0.9714873,0.90256417,1.020718,1.2865642,1.4834872,1.3620514,1.1224617,1.0732309,1.2570257,1.4572309,1.5753847,2.1825643,3.1343591,3.892513,3.501949,2.409026,1.8609232,1.7723079,2.1431797,3.0424619,3.1442053,3.1540515,2.9243078,2.5895386,2.5895386,3.1376412,3.511795,3.8728209,4.20759,4.342154,4.1189747,3.7776413,3.4231799,3.05559,2.556718,2.7175386,3.170462,3.7021542,4.1124105,4.2338467,4.315898,4.493129,4.4964104,4.056616,2.9046156,2.2449234,2.0118976,2.0086155,2.425436,3.8334363,6.6560006,7.634052,9.494975,11.237744,8.119796,4.6539493,5.85518,9.26195,12.78359,14.693745,13.892924,12.747488,10.469745,8.260923,9.321027,9.659078,7.53559,5.8781543,5.8453336,6.820103,6.6067696,8.792616,10.338462,9.777231,7.210667,7.056411,8.385642,8.861539,7.906462,6.7117953,3.945026,2.8225644,3.1803079,3.698872,1.8904617,2.6945643,4.5489235,6.0619493,7.017026,8.372514,6.2720003,3.7382567,2.0250258,1.394872,1.1191796,0.86317956,0.39712822,0.08861539,0.02297436,0.02297436,0.026256412,0.03938462,0.08205129,0.19364104,0.44964105,2.8389745,4.4077954,4.194462,2.7864618,2.3072822,1.4834872,1.1454359,0.9616411,0.7515898,0.48246157,0.20020515,0.43651286,0.6695385,0.8008206,1.1618463,3.9844105,4.3716927,3.2065644,1.4933335,0.34133336,0.17394873,0.12143591,0.15425642,0.19364104,0.118153855,0.04266667,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.02297436,0.009846155,0.072205134,0.20020515,0.27241027,0.101743594,0.02297436,0.016410258,0.12471796,0.45620516,0.5973334,0.5677949,0.43323082,0.27569234,0.2100513,0.37743592,0.53825647,0.6629744,0.9321026,1.723077,2.5665643,4.0369234,4.7392826,4.6145644,4.9394875,4.6900516,4.7458467,4.775385,4.916513,5.7764106,6.3967185,7.1154876,7.3353853,6.5936418,4.5554876,4.9887185,5.76,6.3245134,6.6560006,7.259898,7.4141545,7.6734366,7.955693,8.592411,10.325335,7.683283,6.482052,6.8562055,8.096821,8.635077,6.8955903,6.183385,5.9569235,5.7764106,5.290667,3.56759,3.0391798,3.3411283,3.7185643,3.0227695,1.7558975,0.8795898,0.5284103,0.512,0.3446154,0.38400003,0.46276927,0.4955898,0.46276927,0.38400003,0.31507695,0.28882053,0.23958977,0.15753847,0.08861539,0.055794876,0.04594872,0.03938462,0.029538464,0.029538464,0.04266667,0.059076928,0.07876924,0.08861539,0.08205129,0.16410258,0.26584616,0.38400003,0.5349744,0.764718,1.1552821,2.0118976,3.2328207,4.2896414,4.2305646,4.965744,5.179077,5.1167183,5.0543594,5.290667,5.2315903,5.0838976,4.97559,4.962462,5.034667,5.1364107,5.142975,5.1987696,5.4514875,6.0685134,5.142975,3.6036925,2.7831798,2.8914874,2.9801028,3.1113849,3.1409233,3.2623591,3.6594875,4.4865646,7.4075904,12.314258,17.142155,20.52595,21.812515,22.656002,22.367182,21.891283,21.976618,23.161438,24.799181,25.72472,27.30995,30.57231,36.194466,42.925953,51.124516,65.398155,85.52698,106.45334,128.50873,135.95898,130.97684,116.94278,98.44514,80.47262,60.209236,43.201645,34.79303,40.09026,53.38257,72.21498,96.96493,124.521034,148.30606,137.07487,127.451904,118.53458,108.511185,94.654366,81.70667,69.61231,53.441647,35.639797,26.020105,21.40554,18.94072,18.15631,18.527182,19.442873,20.437334,21.051079,20.824617,19.531488,17.207796,13.8765135,10.384411,7.4043083,5.156103,3.3969233,3.3608208,2.4582565,1.7493335,1.4933335,1.1388719,1.273436,1.3489232,1.214359,1.0633847,1.4441026,1.5753847,1.3915899,1.083077,0.8566154,0.9517949,1.4441026,0.86974365,0.3052308,0.13128206,0.036102567,0.02297436,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03938462,0.01969231,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.032820515,0.055794876,0.07548718,0.0951795,0.10502565,0.08205129,0.06235898,0.049230773,0.036102567,0.026256412,0.032820515,0.16082053,0.18051283,0.08533334,0.09189744,0.052512825,0.02297436,0.006564103,0.0032820515,0.013128206,0.026256412,0.03938462,0.049230773,0.06564103,0.08861539,0.17723078,0.36430773,0.5973334,0.8008206,0.88287187,1.1257436,1.3620514,1.3883078,1.2209232,1.0929232,1.1913847,1.2373334,1.2012309,1.1126155,1.0666667,0.81394875,0.6170257,0.4660513,0.33805132,0.20676924,0.16738462,0.12471796,0.11158975,0.118153855,0.118153855,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.0032820515,0.0,0.0,0.013128206,0.06235898,0.49887183,0.46276927,0.24943592,0.07876924,0.09189744,0.01969231,0.009846155,0.02297436,0.059076928,0.16738462,0.37415388,0.92225647,2.1070771,3.3805132,3.3575387,2.4418464,1.6902566,1.024,0.54482055,0.51856416,0.6170257,0.78769237,1.1355898,1.4572309,1.2373334,0.6268718,0.4266667,0.36758977,0.60061544,1.723077,1.8346668,1.3226668,1.0896411,1.4998976,2.3794873,3.4560003,4.8672824,5.904411,6.7971287,8.713847,11.178667,7.9950776,4.8836927,3.9680004,3.7842054,3.6135387,3.6069746,3.3017437,2.674872,2.1530259,1.6869745,1.4244103,1.2832822,1.1979488,1.1126155,1.1520001,1.3883078,1.595077,1.6836925,1.7099489,2.930872,3.8301542,3.8038976,3.1540515,3.0654361,3.5183592,2.6880002,1.9200002,1.7526156,1.9232821,1.8116925,2.3072822,2.8455386,2.9144619,2.0611284,2.281026,2.425436,2.4451284,2.4352822,2.6551797,2.28759,2.3794873,1.9593848,1.270154,1.7690258,2.2449234,2.3105643,2.353231,2.7273848,3.754667,4.352,5.0674877,6.193231,7.5552826,8.546462,8.461129,9.078155,9.061745,7.5979495,4.4242053,2.937436,2.5829747,2.740513,2.681436,1.5721027,2.546872,2.809436,2.806154,2.937436,3.570872,6.892308,6.6395903,4.71959,3.0752823,3.7218463,5.346462,5.0838976,4.6145644,4.4898467,4.135385,4.073026,3.9680004,3.4789746,3.114667,4.2272825,5.5565133,5.789539,6.9120007,8.585847,8.132924,5.4843082,5.225026,5.4580517,5.609026,6.439385,6.452513,5.684513,5.2578464,5.2447186,4.6834874,3.2328207,3.7120004,4.516103,4.8738465,4.8377438,3.6890259,3.1474874,3.0490258,3.190154,3.31159,3.1507695,2.3171284,1.9692309,2.1891284,1.9692309,3.1638978,3.4921029,3.1113849,2.7700515,3.7842054,5.3825645,6.0849237,6.377026,6.23918,5.1265645,3.370667,3.5249233,5.3431797,7.515898,7.6767187,7.906462,8.1755905,9.206155,10.541949,10.528821,9.91836,11.332924,13.810873,15.192616,12.114052,10.381129,10.459898,10.571488,10.19077,10.056206,8.89436,8.487385,7.962257,7.069539,6.180103,5.1659493,6.2851286,7.2270775,6.994052,5.920821,6.2851286,6.6428723,6.7282057,7.076103,9.019077,11.933539,10.256411,7.456821,5.618872,5.4482055,7.4732313,8.100103,6.9710774,5.4449234,6.5936418,11.414975,14.7790785,14.900514,12.655591,11.58236,13.925745,15.471591,14.057027,10.771693,9.977437,10.627283,10.164514,9.590155,8.999385,7.584821,4.9362054,3.5413337,3.0030773,3.2131286,4.348718,5.1922054,6.948103,8.608821,9.025641,6.9120007,5.691077,7.5454364,8.707283,7.565129,4.6834874,3.757949,3.1507695,2.678154,2.4352822,2.7766156,3.1803079,3.4002054,3.1967182,2.556718,1.6771283,1.4834872,1.3062565,1.0994873,0.8960001,0.82379496,1.0666667,1.1388719,1.0404103,0.8960001,0.94523084,0.82379496,0.81066674,1.1290257,1.785436,2.5796926,2.6880002,2.8160002,3.0654361,3.2722054,2.989949,2.4057438,2.048,1.9331284,2.1989746,3.1277952,3.239385,3.5314875,3.5183592,3.190154,3.006359,2.809436,3.1474874,3.6758976,4.1485133,4.378257,4.4898467,4.1058464,3.5314875,2.8980515,2.166154,1.8871796,1.7329233,1.9167181,2.425436,3.0358977,3.2065644,2.7569232,2.1136413,1.6246156,1.5261539,1.8313848,2.556718,3.131077,3.3936412,3.6004105,5.211898,6.5772314,9.593436,12.3076935,8.92718,4.6769233,5.868308,8.375795,10.020103,10.545232,12.251899,13.889642,14.552616,14.976001,17.499899,17.719797,12.081232,11.513436,16.695797,18.051283,15.753847,13.459693,9.573745,5.4186673,5.2348723,9.737847,12.209231,9.45559,3.5741541,1.9396925,1.2406155,1.7263591,2.3729234,2.5764105,2.1366155,2.930872,4.9788723,6.882462,7.5520005,6.2096415,2.793026,0.86646163,0.38400003,0.7187693,0.65641034,0.5940513,0.29538465,0.08205129,0.04594872,0.04594872,0.02297436,0.1148718,0.24943592,0.28882053,0.04594872,0.032820515,0.23302566,0.6826667,1.1979488,1.3423591,0.49887183,0.53825647,0.5973334,0.38400003,0.15097436,0.055794876,0.18707694,0.20348719,0.11158975,0.25928208,0.8467693,1.0469744,0.8402052,0.4397949,0.3052308,0.24287182,0.14769232,0.14112821,0.18051283,0.04594872,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.0032820515,0.0,0.006564103,0.04266667,0.15097436,0.60389745,0.90912825,0.9878975,0.88287187,0.74830776,0.5513847,0.4397949,0.512,0.77128214,1.1126155,2.1530259,2.3729234,3.4002054,5.110154,5.661539,5.8190775,5.1364107,4.020513,2.9702566,2.5796926,3.629949,4.210872,4.900103,5.605744,5.5696416,5.1922054,5.8912826,6.6067696,7.1876926,8.408616,9.764103,9.80677,9.442462,9.078155,8.651488,8.247795,7.1515903,7.194257,8.231385,8.132924,4.1780515,3.3444104,3.6332312,3.7907696,3.3280003,3.0096412,2.409026,2.2055387,2.2186668,1.3883078,0.99774367,0.49887183,0.41682056,0.6498462,0.44307697,0.3446154,0.4397949,0.3708718,0.14112821,0.09189744,0.09189744,0.08205129,0.07548718,0.07548718,0.07548718,0.06564103,0.052512825,0.03938462,0.029538464,0.029538464,0.04266667,0.04594872,0.03938462,0.032820515,0.04594872,0.059076928,0.068923086,0.07548718,0.08205129,0.108307704,0.25271797,0.49230772,0.98133343,1.7887181,2.8980515,3.692308,4.3684106,4.673641,4.7655387,5.218462,5.2053337,4.919795,4.7917953,4.97559,5.3398976,5.353026,5.2742567,4.890257,4.2371287,3.6004105,3.2853336,2.9111798,2.7766156,2.868513,2.868513,3.2853336,3.6627696,3.9351797,4.1189747,4.3027697,5.3398976,8.283898,12.731078,17.19795,19.088411,19.505232,18.464823,17.335796,16.738462,16.554668,17.129026,19.350975,23.899899,30.726566,39.062977,45.042873,50.13662,60.7639,78.805336,101.60903,114.50093,121.63283,121.41293,113.34893,98.05457,86.86934,62.516518,40.500515,31.520823,41.458874,59.67098,82.37621,106.04965,126.71017,139.96965,132.89027,126.91693,121.85601,116.01724,106.21703,93.09211,79.16637,62.838158,45.830566,33.171696,29.154465,26.266258,24.576002,23.850668,23.545437,22.505028,23.538874,25.833027,27.743181,26.77826,22.675694,18.372925,14.020925,9.892103,6.363898,5.0084105,3.7185643,2.356513,1.1881026,0.86974365,0.7122052,0.5973334,0.50543594,0.56451285,1.0535386,1.1749744,0.9321026,0.77128214,0.892718,1.2209232,1.0371283,0.77128214,0.5152821,0.3052308,0.12143591,0.06235898,0.026256412,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.016410258,0.026256412,0.04266667,0.029538464,0.01969231,0.02297436,0.02297436,0.016410258,0.016410258,0.03938462,0.06564103,0.06564103,0.10502565,0.33476925,0.190359,0.06235898,0.0,0.0,0.0,0.02297436,0.029538464,0.036102567,0.06564103,0.13784617,0.18707694,0.33476925,0.5481026,0.8566154,1.3587693,1.847795,1.7132308,1.401436,1.2274873,1.3718976,1.5688206,1.7624617,1.8970258,1.910154,1.7394873,1.2996924,0.92553854,0.67282057,0.52512825,0.36758977,0.3052308,0.18051283,0.08205129,0.04594872,0.04594872,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.068923086,0.08533334,0.052512825,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.049230773,0.02297436,0.0,0.01969231,0.101743594,0.098461546,0.03938462,0.059076928,0.13784617,0.108307704,0.48246157,0.93866676,0.81394875,0.24287182,0.17723078,0.18051283,0.14112821,0.37743592,0.9156924,1.4867693,0.9714873,1.1684103,1.8412309,2.300718,1.4276924,1.2438976,1.2274873,0.97805136,0.56123084,0.50543594,1.142154,1.4112822,1.2832822,1.024,1.1749744,0.56451285,0.23302566,0.118153855,0.23302566,0.6629744,0.7515898,0.88615394,1.3784616,2.172718,2.8553848,2.681436,4.969026,6.7774363,7.9983597,11.349334,8.41518,6.0291286,4.716308,4.1911798,3.3444104,2.802872,2.8127182,2.6683078,2.166154,1.6016412,1.6082052,1.4178462,1.3062565,1.273436,1.0535386,1.0010257,1.3193847,2.0545642,2.6847181,2.1234872,1.8510771,1.9823592,2.044718,1.9528207,1.9922053,2.9440002,2.609231,2.2186668,2.1398976,1.910154,1.9659488,3.3805132,3.9975388,3.114667,1.4998976,1.719795,2.0053334,2.2121027,2.422154,2.9243078,3.045744,2.2186668,1.4506668,1.1979488,1.3686155,1.6082052,1.7526156,1.8445129,2.3368206,4.096,4.8705645,5.7042055,6.813539,7.860513,7.972103,6.8693337,5.8092313,4.84759,3.9122055,2.789744,2.5107694,2.8127182,3.7349746,4.522667,3.5971284,3.0424619,2.5042052,2.409026,2.737231,3.0227695,5.3760004,7.1548724,7.5487185,6.8693337,6.5312824,6.1997952,6.5772314,7.8080006,8.976411,8.113232,6.1013336,5.76,5.83877,6.0028725,6.8496413,5.3398976,4.640821,5.7731285,7.8112826,7.8769236,5.218462,5.093744,5.5138464,5.733744,6.2818465,5.668103,4.6145644,4.0336413,4.2962055,5.208616,3.318154,3.7743592,5.3136415,6.294975,4.716308,4.1058464,3.3280003,3.2065644,4.125539,6.0324106,5.2676926,3.4100516,2.0906668,1.8445129,2.103795,2.176,2.294154,2.1989746,2.15959,2.9669745,3.9417439,4.962462,5.405539,5.464616,6.1407185,5.3891287,4.916513,5.5236926,6.695385,6.6002054,5.904411,5.874872,7.2336416,9.55077,11.247591,10.161232,11.526565,12.78359,12.583385,10.7848215,9.284924,9.475283,9.573745,9.636104,11.533129,11.408411,9.025641,6.7216415,5.421949,4.630975,5.1200004,6.170257,6.7249236,6.5083084,6.0291286,8.086975,8.507077,8.004924,8.021334,10.7158985,11.661129,10.167795,8.418462,6.7577443,3.7251284,6.9349747,10.016821,9.898667,7.506052,7.762052,17.99549,21.819078,19.012924,12.242052,7.076103,9.537642,12.675283,14.017642,13.131488,11.61518,8.969847,8.04759,7.8145647,7.6964107,7.5585647,5.5171285,5.218462,5.4941545,5.917539,6.7905645,6.265436,6.186667,6.2752824,6.1374364,5.2644105,5.536821,6.7840004,7.026872,5.8289237,4.3060517,4.345436,4.2272825,3.8038976,3.2065644,2.8750772,2.868513,2.793026,2.5928206,2.228513,1.6902566,1.4375386,1.0633847,0.92225647,1.0896411,1.3489232,1.5425643,1.3226668,1.0272821,0.84348726,0.82379496,1.2471796,1.8871796,2.4484105,2.8488207,3.2000003,3.0490258,3.0129232,2.7700515,2.2613335,1.6968206,1.2668719,1.2340513,1.4211283,1.8773335,2.8849232,3.4231799,3.2951798,3.1770258,2.989949,1.9200002,1.6475899,1.9035898,2.4155898,2.9538465,3.3411283,3.3542566,2.7766156,2.428718,2.5304618,2.7175386,2.484513,2.1103592,2.0775387,2.3762052,2.5009232,2.7175386,2.989949,2.9013336,2.4451284,2.0151796,3.6069746,4.0041027,4.315898,4.4406157,3.0752823,4.197744,5.3103595,6.7577443,8.231385,8.756514,9.340718,10.466462,9.862565,8.546462,10.801231,12.235488,12.908309,13.751796,15.133539,16.879591,15.038361,10.217027,7.0432825,6.304821,4.965744,4.1846156,4.522667,7.2960005,12.928001,20.969027,11.1064625,7.768616,6.9021544,6.482052,6.514872,9.101129,12.836103,12.317539,7.3321033,2.8816411,2.9997952,3.0851285,2.8947694,2.4713848,2.1464617,1.4211283,1.7526156,2.353231,2.4320002,1.1815386,0.38728207,0.08861539,0.016410258,0.009846155,0.009846155,0.013128206,0.08533334,0.16738462,0.18379489,0.04594872,0.013128206,0.04594872,0.14112821,0.25271797,0.28225642,0.13128206,0.13784617,0.16410258,0.16082053,0.16410258,0.055794876,0.055794876,0.059076928,0.049230773,0.08861539,0.26584616,0.47261542,0.508718,0.40369233,0.4135385,0.33476925,0.28225642,0.19364104,0.07876924,0.032820515,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0,0.0,0.0,0.009846155,0.029538464,0.2297436,0.55794877,0.8763078,1.1618463,1.5163078,1.3620514,1.3292309,1.2832822,1.0929232,0.67610264,1.4080001,2.5074873,3.698872,5.106872,7.24677,7.1515903,5.989744,4.9887185,4.8016415,5.4974365,4.388103,4.9362054,5.717334,5.874872,5.106872,6.2129235,6.948103,7.4240007,7.680001,7.6996927,6.5444107,6.052103,6.1407185,6.4722056,6.4557953,6.3934364,6.7117953,6.5936418,6.3376417,7.3649235,5.8289237,4.8771286,3.757949,2.3762052,1.2865642,1.214359,1.0043077,0.955077,0.96492314,0.5349744,0.47589746,0.571077,1.1126155,1.6902566,1.1979488,0.45620516,0.20020515,0.128,0.0951795,0.1148718,0.12471796,0.118153855,0.108307704,0.098461546,0.08861539,0.07548718,0.055794876,0.03938462,0.029538464,0.029538464,0.032820515,0.032820515,0.032820515,0.036102567,0.059076928,0.068923086,0.068923086,0.068923086,0.07876924,0.08205129,0.11158975,0.38728207,0.8008206,1.3653334,2.2022567,3.4658465,3.9122055,3.9154875,3.7087183,3.387077,3.170462,2.993231,2.9768207,3.2000003,3.692308,3.9187696,3.95159,3.7776413,3.436308,3.0260515,2.6617439,2.6945643,2.9735386,3.259077,3.2098465,3.3805132,3.9122055,4.414359,4.9394875,5.9634876,6.76759,8.067283,9.734565,11.536411,13.144616,14.496821,14.181745,12.773745,11.227899,10.880001,11.785847,13.220103,16.183796,21.418669,29.394054,34.008617,38.445953,44.389748,54.04226,70.11446,77.8798,77.16103,73.56062,71.791595,75.65457,78.39836,66.4517,50.763493,40.4119,42.594463,51.022774,64.65642,83.203285,104.1756,122.893135,121.5639,114.98011,107.83836,103.4076,103.50606,103.624214,94.87426,77.794464,57.869133,45.512207,40.60882,37.10031,35.488823,34.95713,33.381744,32.64657,32.94195,33.614773,34.46154,35.715286,33.94626,29.545029,23.988514,18.6519,14.821745,11.592206,8.720411,6.3507695,4.3618464,2.3466668,1.6508719,0.96492314,0.48574364,0.2986667,0.35774362,0.4004103,0.37743592,0.5973334,1.1158975,1.7591796,1.4375386,0.9911796,0.65312827,0.43651286,0.14769232,0.07548718,0.03938462,0.02297436,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.013128206,0.009846155,0.01969231,0.036102567,0.032820515,0.02297436,0.016410258,0.016410258,0.029538464,0.052512825,0.055794876,0.098461546,0.3117949,0.08533334,0.013128206,0.0,0.0,0.0,0.013128206,0.01969231,0.029538464,0.06564103,0.15097436,0.24615386,0.5481026,1.024,1.723077,2.7602053,2.2547693,1.6147693,1.5655385,2.1431797,2.678154,2.3171284,2.7634873,3.1803079,3.05559,2.1924105,1.467077,1.3161026,1.1585642,0.81394875,0.48902568,0.30851284,0.17066668,0.08861539,0.055794876,0.04594872,0.47589746,0.0951795,0.0,0.0,0.016410258,0.08205129,0.20676924,0.22646156,0.13128206,0.0,0.0,0.04266667,0.052512825,0.029538464,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03938462,0.01969231,0.0,0.009846155,0.049230773,0.049230773,0.16082053,0.3117949,0.45620516,0.5874872,0.6432821,1.2537436,1.5524104,1.2898463,0.8402052,0.71548724,0.5316923,0.5218462,0.702359,0.88287187,0.6826667,0.7089231,0.9353847,1.1224617,0.827077,0.92225647,1.0601027,1.017436,0.98461545,1.5753847,1.1782565,0.92225647,0.7253334,0.69907695,1.142154,0.45620516,0.14769232,0.0951795,0.21333335,0.42338464,0.53825647,1.1388719,1.782154,2.2678976,2.6551797,3.1474874,4.128821,4.7622566,5.5204105,8.192,6.0291286,4.893539,4.309334,4.2601027,5.2020516,4.706462,3.9187696,3.0391798,2.2383592,1.6213335,1.529436,1.273436,1.1355898,1.1782565,1.2307693,1.1257436,1.1946667,1.5589745,1.9298463,1.5885129,1.3784616,1.4933335,1.6640002,1.8346668,2.172718,2.740513,2.484513,2.15959,2.0053334,1.7427694,2.0512822,2.5304618,2.6518977,2.281026,1.6705642,2.034872,2.3171284,2.6420515,3.0949745,3.7152824,3.255795,2.1398976,1.3653334,1.2931283,1.6410258,1.5983591,1.591795,1.6049232,2.1891284,4.4373336,4.8804107,4.9821544,5.5302567,6.560821,7.351795,6.554257,5.2578464,4.384821,4.0533338,3.5872824,3.8104618,5.3070774,7.463385,8.992821,7.9327188,7.00718,6.2162056,5.349744,4.9887185,6.518154,7.5979495,7.640616,7.499488,7.3485136,6.7216415,7.0432825,7.8769236,8.864821,9.498257,9.117539,7.75877,7.0367184,6.6560006,6.6822567,7.5454364,6.163693,5.7009234,6.229334,7.2205133,7.5454364,6.482052,5.618872,5.4875903,6.114462,7.000616,5.858462,4.601436,3.7349746,3.7316926,5.0215387,3.5380516,4.020513,4.972308,5.1922054,3.767795,4.010667,3.6660516,3.308308,3.7185643,5.861744,5.1889234,3.6332312,2.665026,2.5173335,2.1924105,2.3794873,2.6453335,2.6912823,2.6683078,3.1540515,3.3509746,4.1813335,4.824616,4.9887185,4.9099493,5.9995904,5.8453336,5.717334,5.9963083,6.157129,5.156103,4.634257,5.159385,6.6494365,8.372514,8.848411,11.083488,12.609642,12.3536415,10.663385,9.590155,8.887795,8.283898,8.100103,9.238976,9.783795,8.500513,6.889026,5.8945646,5.907693,6.6494365,6.9710774,7.2927184,8.214975,10.505847,12.068104,11.211488,9.508103,8.809027,11.221334,10.407386,9.212719,7.785026,5.979898,3.3608208,4.7983594,7.059693,7.030154,5.2053337,5.6943593,12.86236,15.947489,14.641232,10.745437,8.1755905,10.584617,12.232206,12.87877,12.274873,10.138257,8.4512825,7.9425645,7.7259493,7.5552826,7.817847,9.412924,10.627283,10.423796,8.726975,6.419693,6.961231,6.7807183,6.298257,5.7468724,5.1626673,5.208616,5.8847184,5.914257,5.097026,4.3290257,3.7120004,3.1409233,2.6584618,2.3171284,2.176,2.0086155,1.8576412,1.7394873,1.595077,1.2832822,1.020718,0.82379496,0.9288206,1.3522053,1.8838975,1.8313848,1.585231,1.332513,1.1257436,0.8763078,2.0742567,3.511795,4.31918,4.201026,3.4198978,2.9243078,3.0260515,2.989949,2.5993848,2.169436,2.4910772,2.8488207,2.930872,2.7634873,2.7044106,2.917744,3.2328207,4.066462,4.7327185,3.4231799,1.6968206,1.332513,1.6935385,2.2514873,2.605949,2.7109745,2.4385643,2.1924105,2.1431797,2.2219489,2.0086155,1.6968206,1.6049232,1.7362052,1.7788719,2.0545642,2.412308,2.6453335,2.7634873,2.9965131,3.764513,3.7284105,4.6211286,6.0192823,5.353026,4.46359,4.9296412,6.0160003,6.9710774,7.000616,6.3343596,6.173539,5.5269747,5.287385,8.228104,9.186462,9.005949,9.540924,10.971898,11.798975,8.848411,6.8627696,5.970052,6.0619493,6.7938466,8.674462,9.787078,9.754257,10.584617,16.672821,12.438975,6.885744,3.9023592,4.338872,5.98318,7.3025646,9.412924,8.477539,4.529231,1.4834872,1.5819489,1.3423591,0.9419488,0.5940513,0.571077,1.8904617,3.7874875,4.6572313,3.6332312,0.5874872,0.15425642,0.029538464,0.06235898,0.13784617,0.18379489,0.108307704,0.06564103,0.059076928,0.06235898,0.01969231,0.0032820515,0.0,0.009846155,0.02297436,0.02297436,0.055794876,0.072205134,0.10502565,0.15753847,0.19692309,0.24615386,0.27241027,0.24615386,0.17723078,0.108307704,0.072205134,0.17394873,0.256,0.28225642,0.3314872,0.23958977,0.18051283,0.12471796,0.059076928,0.013128206,0.006564103,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.052512825,0.23630771,0.47917953,0.7581539,1.0962052,1.5261539,1.6968206,1.5688206,1.3095386,1.2800001,1.7165129,2.8816411,3.748103,4.3651285,5.8518977,6.452513,6.0619493,5.4186673,5.218462,6.114462,5.0477953,5.034667,5.353026,5.648411,5.933949,6.0192823,6.669129,7.1515903,7.312411,7.5585647,6.567385,6.2687182,7.6964107,10.171078,11.296822,12.596514,12.419283,10.640411,8.169026,6.941539,5.421949,4.647385,3.7874875,2.6945643,1.9035898,1.4539489,1.1585642,0.9878975,0.9156924,0.9156924,0.8533334,0.6662565,0.69251287,0.83035904,0.5546667,0.2100513,0.07548718,0.052512825,0.072205134,0.0951795,0.12143591,0.1148718,0.0951795,0.07876924,0.08205129,0.06235898,0.049230773,0.03938462,0.029538464,0.029538464,0.029538464,0.029538464,0.032820515,0.04266667,0.052512825,0.055794876,0.059076928,0.06235898,0.06564103,0.06564103,0.07548718,0.20020515,0.4004103,0.7056411,1.2340513,2.0939488,2.6945643,2.934154,2.8258464,2.4910772,2.9472823,3.3509746,3.498667,3.4297438,3.436308,3.3936412,3.0884104,2.737231,2.4976413,2.4713848,2.1956925,2.228513,2.7011285,3.3805132,3.6627696,4.161641,4.1550775,4.0303593,4.2141542,5.159385,6.2555904,7.5913854,8.848411,9.970873,11.162257,11.995898,10.272821,7.975385,6.436103,6.3376417,7.4141545,9.179898,11.844924,15.881847,22.016,24.06072,25.59672,28.160002,33.716515,44.68185,55.118774,58.23016,59.346054,61.43672,65.11919,63.56021,59.4478,52.98216,45.620518,40.083694,42.765133,49.765747,62.66421,80.19693,98.28104,95.90811,88.14278,80.620316,77.003494,78.962875,85.40555,86.88903,81.72308,73.62955,71.76862,70.54442,70.797134,68.91324,64.36103,59.700516,54.925133,51.715286,47.84575,42.96862,38.61662,36.24698,32.60718,28.314259,24.185438,21.241438,17.657436,14.155488,11.024411,8.310155,5.802667,4.1058464,2.5829747,1.3751796,0.6268718,0.4660513,0.37415388,0.3249231,0.46933338,0.84348726,1.3522053,1.0994873,0.7515898,0.48246157,0.32164106,0.14441027,0.14441027,0.14112821,0.1148718,0.068923086,0.026256412,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.0,0.12471796,0.15425642,0.098461546,0.016410258,0.006564103,0.118153855,0.18707694,0.16082053,0.068923086,0.02297436,0.02297436,0.02297436,0.036102567,0.0951795,0.24943592,0.055794876,0.0032820515,0.0,0.0,0.0,0.013128206,0.016410258,0.04266667,0.1148718,0.24287182,0.39712822,1.0338463,1.4506668,1.6213335,2.169436,2.2186668,2.0775387,2.1169233,2.353231,2.4484105,3.0227695,5.398975,7.4896417,7.273026,2.7700515,1.5819489,1.1881026,1.017436,0.764718,0.4004103,0.26584616,0.16082053,0.098461546,0.068923086,0.06564103,0.47589746,0.0951795,0.0,0.0,0.016410258,0.08205129,1.8609232,2.8521028,1.9889232,0.118153855,0.0,0.006564103,0.009846155,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.04266667,0.032820515,0.013128206,0.0,0.006564103,0.036102567,0.19364104,0.73517954,1.3718976,1.7788719,1.5885129,0.92553854,1.1716924,1.5425643,1.6114873,1.3226668,1.0469744,0.761436,0.5907693,0.5677949,0.61374366,0.7417436,0.6629744,0.57764107,0.5973334,0.74830776,0.8730257,1.0502565,1.1257436,1.1848207,1.5491283,0.81394875,0.41682056,0.32164106,0.5513847,1.1913847,0.7515898,0.30851284,0.14112821,0.25928208,0.4004103,0.56451285,1.0338463,1.4933335,1.8018463,1.972513,2.7175386,2.8553848,3.170462,4.164923,6.048821,5.0116925,4.417641,3.8662567,4.0303593,6.636308,6.0160003,4.781949,3.5741541,2.6518977,1.913436,1.5360001,1.2668719,1.1979488,1.3095386,1.4867693,1.2865642,1.1716924,1.1454359,1.1749744,1.214359,1.3292309,1.4441026,1.5753847,1.7952822,2.2350771,2.3926156,2.2777438,2.2350771,2.2678976,2.0545642,2.03159,1.723077,1.6311796,1.8576412,2.1103592,2.3138463,2.3368206,2.4681027,2.7667694,3.062154,2.484513,1.9823592,1.7526156,1.7624617,1.7394873,1.782154,1.6804104,1.8576412,2.7208207,4.663795,4.493129,4.089436,4.2568207,5.10359,6.038975,5.98318,5.21518,4.962462,5.297231,5.146257,6.5083084,8.201847,10.180923,11.720206,11.392001,11.073642,10.633847,9.668923,9.301334,12.199386,11.759591,11.858052,11.398565,9.987283,7.9163084,7.2205133,7.1909747,7.39118,7.7423596,8.52677,8.805744,8.536616,8.254359,8.329846,8.976411,7.9950776,7.460103,6.820103,6.2194877,6.498462,6.7610264,6.0061545,5.681231,6.245744,7.1483083,6.0717955,5.1364107,4.141949,3.498667,4.197744,3.4625645,3.442872,3.6036925,3.6102567,3.3247182,3.9023592,3.7054362,3.1081028,2.8849232,4.2338467,3.8728209,3.308308,3.045744,3.1113849,3.0523078,3.4724104,3.3805132,2.92759,2.6157951,3.2853336,3.7218463,4.204308,4.397949,4.4110775,4.8114877,6.058667,6.0258465,5.481026,5.146257,5.730462,5.156103,5.097026,5.146257,5.1200004,5.0642056,6.564103,11.782565,15.90154,16.233027,12.225642,9.734565,7.709539,6.7905645,7.177847,8.628513,8.4053335,7.2664623,6.363898,6.4722056,7.9786673,7.893334,7.9163084,8.612103,10.394258,13.522053,13.571283,12.160001,10.443488,9.45559,10.085744,8.480822,6.744616,5.2545643,4.4012313,4.5817437,4.9394875,4.9427695,4.1550775,3.373949,4.630975,8.103385,10.098872,10.466462,10.043077,10.633847,13.289026,13.377642,12.265027,10.686359,8.740103,8.260923,8.083693,7.906462,7.6931286,7.653744,10.052924,11.687386,11.0605135,8.474257,6.012718,7.8736415,8.241231,7.3321033,5.858462,5.028103,4.640821,4.95918,5.024821,4.571898,4.0500517,2.8422565,1.9823592,1.6738462,1.7887181,1.8707694,1.5425643,1.4244103,1.3850257,1.2996924,1.0568206,0.8336411,0.7844103,1.0371283,1.5622566,2.176,2.2908719,1.9561027,1.6147693,1.3456411,0.8566154,2.3138463,4.092718,5.156103,4.9920006,3.5807183,2.7700515,2.7963078,2.930872,2.9833848,3.2853336,4.027077,4.240411,4.007385,3.4494362,2.7208207,2.609231,3.0424619,4.2141542,5.3727183,4.821334,2.487795,1.6836925,1.6475899,1.8806155,2.15959,2.3138463,2.3893335,2.2219489,1.9232821,1.847795,1.8018463,1.5983591,1.4769232,1.5360001,1.7066668,1.8543591,2.281026,2.740513,3.1606157,3.6135387,3.6036925,4.663795,8.418462,13.029744,13.213539,7.8080006,5.9634876,5.8847184,6.0258465,5.097026,3.190154,2.4057438,2.5862565,3.7382567,6.0619493,6.0061545,5.799385,6.550975,7.7981544,7.4699492,5.4449234,6.7183595,8.434873,9.330873,9.718155,11.053949,11.021129,8.644924,6.0356927,8.408616,8.884514,4.71959,2.1956925,3.1573336,5.037949,5.85518,7.1023593,6.3474874,3.5511796,1.086359,0.9682052,0.5973334,0.28225642,0.256,0.6629744,2.7044106,5.169231,5.540103,3.3247182,0.068923086,0.026256412,0.14112821,0.45292312,0.80738467,0.8598975,0.52512825,0.2100513,0.032820515,0.0,0.0,0.013128206,0.009846155,0.013128206,0.029538464,0.055794876,0.21989745,0.15425642,0.15097436,0.24287182,0.21333335,0.24943592,0.27241027,0.26584616,0.21661541,0.10502565,0.055794876,0.098461546,0.16082053,0.20020515,0.18051283,0.13456412,0.0951795,0.06564103,0.04594872,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.052512825,0.17723078,0.3708718,0.6268718,1.2438976,1.4998976,1.5458462,1.5261539,1.585231,1.8871796,3.1015387,3.7054362,3.4724104,3.4888208,4.263385,4.8804107,4.841026,4.601436,5.5729237,5.481026,5.0871797,4.84759,5.031385,5.737026,5.6943593,5.8190775,6.0652313,6.49518,7.2861543,6.5805135,6.564103,8.530052,11.835078,13.90277,16.449642,16.311796,13.90277,11.011283,10.794667,7.4863596,5.7042055,4.821334,4.276513,3.5872824,2.605949,1.9593848,1.7558975,1.8412309,1.782154,1.8412309,1.529436,0.88943595,0.2100513,0.006564103,0.01969231,0.032820515,0.04594872,0.06564103,0.08205129,0.108307704,0.098461546,0.07876924,0.068923086,0.07548718,0.052512825,0.04594872,0.04266667,0.036102567,0.029538464,0.029538464,0.032820515,0.03938462,0.04594872,0.04594872,0.04594872,0.052512825,0.055794876,0.06235898,0.06235898,0.068923086,0.08533334,0.13128206,0.24287182,0.48902568,0.82379496,1.2964103,1.591795,1.6114873,1.4703591,2.1333334,2.7569232,2.989949,2.8455386,2.7044106,2.612513,2.3138463,2.041436,1.9528207,2.1234872,1.9561027,1.8445129,2.100513,2.6486156,3.0326157,3.764513,3.6135387,3.239385,3.18359,3.8662567,4.95918,6.088206,6.944821,7.50277,8.027898,8.254359,6.196513,4.266667,3.5446157,3.767795,4.4832826,6.11118,8.349539,11.10318,14.454155,15.136822,15.028514,15.944206,19.26236,25.918362,36.470158,43.798977,50.143185,56.717133,63.734158,57.458878,53.39898,50.113644,45.380928,36.18462,34.724106,38.908722,46.93334,57.327595,68.978874,64.83365,57.327595,51.616825,50.264618,53.26113,64.48247,77.35139,86.505035,92.48165,101.71406,106.06934,110.69704,109.72883,102.4197,93.14462,82.707695,72.92062,62.690468,52.25026,43.17539,38.7118,34.658463,30.962873,27.72349,25.183182,21.914259,18.921026,15.908104,12.868924,10.105436,7.7390776,5.533539,3.7120004,2.3302567,1.2800001,0.90256417,0.6301539,0.51856416,0.58420515,0.8041026,0.69251287,0.5940513,0.7515898,1.2242053,1.8773335,1.5097437,0.84348726,0.32820517,0.12143591,0.07548718,0.036102567,0.036102567,0.029538464,0.013128206,0.013128206,0.013128206,0.009846155,0.013128206,0.02297436,0.01969231,0.03938462,0.20348719,0.36430773,0.41025645,0.2855385,0.27897438,0.24287182,0.17066668,0.10502565,0.128,0.18051283,0.25271797,0.21661541,0.09189744,0.036102567,0.01969231,0.006564103,0.013128206,0.055794876,0.13456412,0.04266667,0.009846155,0.006564103,0.01969231,0.02297436,0.06564103,0.26256412,0.48574364,0.88943595,1.9167181,1.522872,2.2777438,2.9801028,3.3214362,3.895795,3.5413337,2.7142565,2.353231,2.5961027,2.802872,4.519385,8.205129,11.149129,10.624001,3.876103,1.6508719,0.8566154,0.6498462,0.5152821,0.26584616,0.19364104,0.14112821,0.098461546,0.068923086,0.06564103,0.0,0.19364104,0.190359,0.0951795,0.009846155,0.0,3.442872,5.362872,3.757949,0.23302566,0.0,0.0,0.0,0.0,0.006564103,0.02297436,0.009846155,0.0032820515,0.0,0.0,0.0,0.0032820515,0.04266667,0.03938462,0.016410258,0.08533334,0.052512825,0.04594872,0.026256412,0.013128206,0.072205134,0.45292312,1.5622566,2.8160002,3.4724104,2.6322052,1.3784616,1.020718,1.0010257,1.211077,1.9823592,1.5753847,0.9419488,0.6071795,0.7089231,0.9944616,1.1618463,1.1552821,1.1290257,1.1093334,1.017436,0.9288206,1.0043077,1.0568206,0.93866676,0.5349744,0.36758977,0.380718,0.48246157,0.86317956,1.9659488,1.5622566,0.6859488,0.3708718,0.7220513,0.9321026,0.6268718,0.4660513,0.64000005,1.014154,1.1355898,1.2964103,1.7591796,2.9210258,4.6244106,6.1768208,5.0149746,4.2371287,3.4789746,3.5544617,6.445949,5.5236926,4.644103,3.9154875,3.239385,2.300718,1.6672822,1.4802053,1.5688206,1.7526156,1.8248206,1.5261539,1.3653334,1.1913847,1.0568206,1.2242053,1.3686155,1.3751796,1.4342566,1.6311796,1.9495386,1.9167181,1.9823592,2.2678976,2.5796926,2.3991797,1.9232821,1.6672822,1.7394873,2.044718,2.28759,2.1300514,1.8970258,1.7558975,1.657436,1.3554872,1.339077,1.7755898,2.3105643,2.4615386,1.595077,1.9659488,2.0808206,2.5993848,3.6463592,4.821334,4.2469745,4.0533338,4.4242053,5.0510774,5.106872,5.5302567,5.3924108,5.5138464,5.973334,6.1046157,8.651488,9.557334,10.400822,11.756309,13.197129,13.702565,14.060308,13.948719,14.391796,17.749334,16.692514,18.566566,18.58954,15.425642,11.195078,7.4765134,5.874872,5.717334,6.498462,7.8670774,9.222565,9.728001,10.000411,10.35159,10.79795,9.95118,8.907488,7.1844106,5.4383593,5.467898,6.0225644,6.124308,6.0225644,5.986462,6.298257,5.789539,5.4875903,4.709744,3.6036925,3.1507695,3.0916924,2.349949,2.1333334,2.733949,3.5183592,3.6463592,3.1638978,2.5961027,2.3302567,2.6157951,2.553436,2.8521028,3.1376412,3.4888208,4.420923,4.5554876,3.6496413,2.4320002,1.847795,3.045744,4.3290257,4.673641,4.1813335,3.9023592,5.8125134,6.2030773,5.7764106,5.0018463,4.578462,5.464616,5.4153852,6.2720003,6.698667,5.9930263,4.1025643,5.100308,12.921437,19.465847,20.14195,13.88636,9.29477,6.245744,5.930667,8.237949,11.766154,9.622975,7.131898,6.445949,8.027898,10.643693,8.55959,8.39877,9.6,11.336206,12.517745,11.316514,10.706052,10.272821,9.517949,7.8506675,6.4065647,4.2601027,3.170462,3.9975388,6.705231,7.450257,5.4482055,3.9614363,4.604718,7.322257,9.258667,9.7903595,9.747693,10.029949,11.61518,15.041642,15.205745,13.000206,10.010257,8.507077,7.8506675,7.958975,8.267488,8.303591,7.6964107,7.6734366,8.477539,8.070564,6.6822567,6.810257,8.421744,8.861539,7.604513,5.35959,4.073026,3.7382567,4.017231,4.273231,4.1878977,3.7316926,2.6256413,1.719795,1.5589745,1.9298463,1.8806155,1.4276924,1.3915899,1.4276924,1.3423591,1.086359,1.020718,1.0371283,1.2832822,1.7624617,2.3138463,2.7831798,2.281026,1.7165129,1.3489232,0.8172308,1.8018463,3.2722054,4.5587697,5.024821,4.069744,3.0030773,2.546872,2.5238976,2.937436,3.948308,4.3552823,4.020513,3.564308,3.186872,2.6387694,2.4976413,2.5731285,3.2065644,4.1780515,4.709744,3.131077,2.3401027,1.9396925,1.8051283,2.0644104,2.1956925,2.3466668,2.2088206,1.9068719,1.9987694,2.1464617,2.0611284,1.9856411,2.0676925,2.3368206,2.1989746,2.5140514,2.9965131,3.3903592,3.495385,3.2000003,6.0816417,13.39077,21.376001,21.27754,11.969642,7.318975,5.4416413,4.772103,4.076308,2.8258464,2.3368206,2.9144619,4.2535386,5.428513,4.519385,4.9099493,6.1374364,7.0400004,5.7435904,6.166975,10.522257,13.433437,12.553847,8.5891285,6.3245134,4.5587697,3.3575387,2.9013336,3.4888208,2.1103592,1.0765129,1.8609232,4.1222568,5.691077,7.5946674,9.580308,9.278359,6.449231,2.9669745,2.5140514,1.4736412,0.571077,0.3708718,1.273436,3.2951798,5.4908724,4.9394875,1.9429746,0.016410258,0.013128206,0.3249231,0.9747693,1.657436,1.723077,1.0568206,0.42338464,0.06564103,0.0,0.0,0.036102567,0.036102567,0.02297436,0.032820515,0.08533334,0.39056414,0.25271797,0.190359,0.28225642,0.17066668,0.052512825,0.016410258,0.055794876,0.108307704,0.04594872,0.12471796,0.19692309,0.23958977,0.2231795,0.08205129,0.08861539,0.08205129,0.055794876,0.01969231,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.07876924,0.23302566,0.4660513,0.7515898,0.97805136,1.3161026,1.6016412,1.3423591,1.5327181,2.740513,3.2131286,2.546872,1.6738462,1.8674873,2.8291285,3.383795,3.511795,4.342154,5.0215387,4.9526157,4.6900516,4.535795,4.529231,5.3005133,4.775385,4.706462,5.5597954,6.5050263,5.658257,6.308103,8.008205,10.272821,12.576821,15.392821,16.331488,14.972719,13.371078,16.091898,12.041847,8.694155,6.8299494,6.091488,4.9854364,3.8301542,2.986667,2.8356924,3.0523078,2.6289232,3.0129232,2.9472823,1.9331284,0.46933338,0.052512825,0.026256412,0.032820515,0.049230773,0.068923086,0.0951795,0.10502565,0.09189744,0.07876924,0.07548718,0.072205134,0.052512825,0.04594872,0.04594872,0.04266667,0.032820515,0.032820515,0.03938462,0.04594872,0.049230773,0.049230773,0.04594872,0.04594872,0.052512825,0.06235898,0.06235898,0.06235898,0.07548718,0.08861539,0.11158975,0.16410258,0.2297436,0.28225642,0.33805132,0.37743592,0.36102566,0.5546667,0.8763078,1.0568206,1.0929232,1.2176411,1.3620514,1.4998976,1.6213335,1.723077,1.8084104,1.7066668,1.5589745,1.463795,1.4867693,1.6508719,2.3335385,2.4320002,2.3236926,2.3762052,2.92759,3.56759,3.9844105,4.066462,3.8564105,3.5577438,3.570872,2.7634873,2.359795,2.7273848,3.3772311,3.7185643,4.630975,5.9569235,7.3058467,8.034462,8.690872,8.854975,9.619693,11.575796,14.828309,20.315899,26.532104,33.634464,43.559387,60.051697,58.801235,51.86298,45.522057,40.382362,31.38626,27.02113,30.959593,35.380516,37.730465,40.720413,37.16267,32.462772,30.529644,32.89272,38.68226,53.645134,73.724724,91.82195,105.921646,119.131905,126.59529,131.74155,130.9637,123.51016,111.465034,98.82913,84.64082,70.64616,58.51898,49.88062,44.501335,39.824413,35.59057,31.776823,28.583387,25.622976,23.552002,21.287386,18.379488,14.998976,12.42913,9.869129,7.6176414,5.5007186,2.878359,1.9823592,1.2931283,0.86317956,0.67282057,0.636718,0.65969235,0.8763078,1.7920002,3.370667,5.0609236,4.056616,2.428718,1.0272821,0.2855385,0.2297436,0.15753847,0.12471796,0.08205129,0.032820515,0.032820515,0.055794876,0.055794876,0.07548718,0.12471796,0.16410258,0.34133336,0.7253334,1.0436924,1.1290257,0.90912825,0.5907693,0.39712822,0.3117949,0.318359,0.39056414,0.2100513,0.18379489,0.14441027,0.06235898,0.04266667,0.01969231,0.0032820515,0.0,0.009846155,0.03938462,0.03938462,0.016410258,0.01969231,0.06235898,0.108307704,0.20676924,0.7220513,1.3554872,2.353231,4.4996924,3.889231,4.70318,6.0258465,7.325539,8.487385,6.0849237,3.4756925,2.4681027,3.18359,4.066462,5.9995904,9.301334,11.34277,10.154668,4.4307694,1.5097437,0.5349744,0.32164106,0.2297436,0.16738462,0.12143591,0.10502565,0.09189744,0.072205134,0.052512825,0.0,0.97805136,0.94523084,0.48246157,0.049230773,0.0,0.65969235,0.5481026,0.21989745,0.0,0.0,0.0,0.0,0.006564103,0.032820515,0.108307704,0.04594872,0.013128206,0.0,0.0,0.0,0.013128206,0.20676924,0.20020515,0.0,0.0,0.072205134,0.17394873,0.13784617,0.0,0.0,0.32820517,1.9035898,3.1967182,3.4494362,2.6551797,2.1530259,1.7001027,1.3095386,1.7033848,4.3027697,3.6791797,1.7394873,0.48246157,0.38400003,0.39712822,0.7384616,1.3259488,2.1136413,2.6518977,2.0906668,1.3587693,0.67282057,0.32820517,0.43651286,0.8992821,0.4135385,0.702359,1.1716924,2.1103592,4.699898,2.6847181,1.0929232,1.1716924,2.5665643,3.31159,0.955077,0.28225642,0.27897438,0.40369233,0.6104616,0.83035904,1.5721027,2.537026,3.4921029,4.273231,4.3716927,3.826872,3.117949,3.0884104,4.9427695,4.1517954,4.0992823,4.197744,3.8990772,2.7175386,1.9462565,1.782154,1.9889232,2.300718,2.412308,2.1924105,1.8445129,1.4342566,1.0765129,0.9321026,1.017436,1.3029745,1.6443079,1.9626669,2.2416413,1.8904617,1.6082052,1.4244103,1.3259488,1.2504616,1.8018463,1.8084104,1.7788719,1.8116925,1.6180514,1.5556924,1.6771283,1.8904617,1.9298463,1.3423591,1.4539489,1.7099489,2.3696413,2.8914874,1.9364104,2.169436,3.0424619,3.6036925,3.9318976,5.1265645,5.139693,5.72718,6.9776416,8.086975,7.3550773,7.463385,7.4469748,6.6395903,5.467898,5.431795,6.6527185,7.3780518,8.881231,11.562668,14.969437,15.199181,16.41354,17.322668,18.103796,20.384823,21.848618,21.546669,20.900105,19.495386,15.074463,9.974154,8.43159,8.914052,9.685334,8.818872,9.199591,8.809027,8.3134365,8.369231,9.613129,10.322052,9.554052,8.067283,6.738052,6.5903597,6.7249236,6.49518,6.0619493,5.5532312,5.0674877,4.919795,4.699898,4.5423594,4.1124105,2.6256413,2.8816411,2.3762052,2.3236926,2.9078977,3.31159,2.481231,1.9068719,2.0217438,2.553436,2.5173335,2.737231,2.793026,3.4034874,4.44718,4.95918,4.1156926,2.9078977,1.9265642,1.7394873,2.8980515,3.6069746,4.4077954,4.5423594,4.1911798,4.4701543,6.8496413,6.009436,5.106872,5.405539,6.2720003,5.477744,5.5269747,6.6560006,8.057437,7.8736415,7.4469748,11.329642,14.280207,14.165335,11.992617,8.953437,6.088206,7.2960005,12.438975,17.332514,13.745232,11.372309,11.825232,14.293334,15.563488,9.924924,7.975385,8.41518,9.330873,8.208411,7.427283,8.165744,8.717129,8.093539,6.042257,4.9329233,5.395693,6.51159,7.584821,8.132924,8.631796,6.422975,6.0324106,9.229129,15.015386,15.320617,13.098668,10.289231,8.635077,9.6754875,14.39836,16.66954,15.117129,11.047385,8.421744,6.944821,8.333129,10.043077,10.663385,9.91836,9.3078985,9.255385,9.517949,9.557334,8.54318,6.8365135,5.7140517,4.9427695,4.0500517,2.3040001,2.3893335,2.9702566,3.8432825,4.598154,4.6244106,3.8301542,2.166154,1.3062565,1.3554872,0.8533334,0.6465641,0.7220513,0.9321026,1.0732309,0.9156924,1.270154,1.5589745,1.8215386,2.1530259,2.7175386,2.6683078,2.2055387,1.6443079,1.2209232,1.0994873,1.1848207,1.9462565,3.3214362,4.778667,5.3398976,3.9975388,2.793026,2.4188719,2.802872,3.0818465,2.484513,2.041436,1.8707694,1.8707694,1.723077,1.7001027,1.8116925,2.1924105,2.7076926,2.9768207,2.3171284,1.8116925,1.7690258,2.1234872,2.4418464,2.6617439,2.4681027,2.1464617,1.9856411,2.3040001,2.2678976,2.477949,2.7175386,2.8750772,2.9604106,2.605949,1.7132308,1.6278975,2.3958976,2.7634873,1.394872,3.5905645,10.548513,17.956104,15.990155,10.620719,6.265436,4.33559,4.4800005,4.578462,3.5413337,2.878359,3.0424619,4.023795,5.356308,5.4547696,5.9634876,6.3901544,6.2555904,5.097026,7.4174366,15.07118,18.802874,15.238565,6.928411,2.6912823,1.3029745,0.98461545,0.764718,0.47261542,0.31507695,0.38400003,1.3357949,3.5807183,7.27959,8.205129,8.546462,8.480822,7.9228725,6.5312824,6.616616,4.3749747,1.8379488,0.41682056,0.9321026,4.020513,5.723898,4.4865646,1.3587693,0.016410258,0.0032820515,0.35774362,0.9747693,1.6016412,1.847795,1.0535386,0.34133336,0.0,0.0,0.0,0.036102567,0.06564103,0.059076928,0.036102567,0.06235898,0.17066668,0.2986667,0.28225642,0.12143591,0.0,0.0,0.0,0.006564103,0.032820515,0.108307704,0.31507695,0.42994875,0.45620516,0.37415388,0.16738462,0.04594872,0.02297436,0.01969231,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.03938462,0.101743594,0.19692309,0.35774362,0.6629744,0.9321026,1.1355898,1.404718,1.086359,1.3456411,1.4178462,1.2373334,1.4178462,1.3095386,1.1552821,1.7591796,2.681436,2.2416413,2.4615386,3.7349746,4.7983594,5.0674877,4.637539,3.8564105,3.515077,3.9056413,4.7491283,5.1889234,5.1889234,8.146052,10.469745,11.441232,13.200411,14.723283,16.331488,16.459488,14.992412,13.259488,14.588719,11.85477,8.6580515,6.5378466,4.97559,4.571898,4.332308,3.9318976,3.4100516,3.190154,3.8006158,3.767795,2.553436,0.77128214,0.19692309,0.06564103,0.029538464,0.04266667,0.068923086,0.108307704,0.108307704,0.098461546,0.08533334,0.072205134,0.06235898,0.06235898,0.052512825,0.04594872,0.04594872,0.04594872,0.04594872,0.04594872,0.052512825,0.06235898,0.06235898,0.049230773,0.04594872,0.052512825,0.06235898,0.06235898,0.072205134,0.0951795,0.11158975,0.128,0.15097436,0.17723078,0.19364104,0.2231795,0.26256412,0.27569234,0.27569234,0.27569234,0.2855385,0.30194873,0.28882053,0.37415388,0.761436,1.0502565,1.0896411,0.9911796,0.9189744,1.0929232,1.2570257,1.3226668,1.3587693,1.9922053,1.6672822,1.404718,1.6082052,2.0611284,2.3269746,2.917744,3.4494362,3.4855387,2.5337439,2.300718,2.1431797,2.349949,3.1573336,4.7458467,6.1013336,7.0990777,7.709539,7.9491286,7.890052,7.6931286,7.8736415,9.058462,11.044104,12.803283,13.180719,12.826258,13.830565,19.403488,33.890465,49.857643,50.067696,42.96862,33.765747,24.415182,20.079592,22.459078,24.25436,23.217232,22.14072,21.641848,22.485334,25.380104,30.818464,39.108925,52.401234,68.79836,85.1036,97.54913,101.822365,103.82442,100.44391,93.75508,85.97662,79.471596,75.5758,69.96021,62.526363,55.217236,52.017235,50.80944,49.250465,45.54503,40.142773,35.734978,32.610462,30.217848,28.20267,25.655796,21.103592,18.271181,15.622565,12.806565,9.531077,5.540103,3.7940516,2.422154,1.6114873,1.2832822,1.1126155,1.2242053,1.7624617,3.498667,5.937231,7.3550773,6.2916927,4.97559,2.917744,0.8402052,0.65641034,0.54482055,0.28882053,0.101743594,0.04594872,0.04594872,0.15425642,0.19364104,0.24615386,0.38400003,0.64000005,1.3357949,1.585231,1.6147693,1.6049232,1.6771283,1.3981539,1.0535386,0.8041026,0.69579494,0.67282057,0.256,0.098461546,0.049230773,0.029538464,0.029538464,0.006564103,0.0,0.006564103,0.03938462,0.13784617,0.08861539,0.029538464,0.02297436,0.108307704,0.3052308,0.45292312,1.0666667,2.2383592,3.764513,5.156103,7.13518,8.664616,10.262975,11.844924,12.711386,7.778462,4.640821,3.5544617,4.017231,4.7622566,5.0051284,6.38359,6.114462,3.895795,1.8937438,0.8172308,0.33805132,0.17394873,0.13128206,0.108307704,0.068923086,0.068923086,0.101743594,0.12471796,0.07548718,1.2832822,1.7099489,1.1552821,0.43323082,0.118153855,0.53825647,1.8904617,1.8937438,1.0043077,0.190359,0.9517949,1.8609232,1.2603078,0.4266667,0.006564103,0.02297436,0.4594872,0.42338464,0.19692309,0.0,0.0,0.0032820515,0.47261542,0.56451285,0.18707694,0.0,1.4408206,2.8356924,2.1136413,0.0,0.0,0.12471796,0.86317956,1.6344616,2.1792822,2.556718,4.1452312,2.7273848,1.4572309,1.3883078,1.4605129,1.4802053,1.1815386,0.71548724,0.28882053,0.16410258,0.7122052,0.79425645,1.0075898,1.404718,1.5163078,0.67610264,0.31507695,0.20348719,0.27897438,0.65641034,0.73517954,2.8488207,3.4855387,2.166154,1.4539489,0.86317956,0.7778462,1.6475899,2.6486156,1.6640002,0.6071795,0.34133336,0.37743592,0.46276927,0.574359,0.508718,0.9911796,1.6607181,2.3269746,2.9407182,3.0293336,2.6453335,2.2547693,2.1956925,2.674872,2.6715899,2.8816411,3.0523078,2.9833848,2.5206156,2.044718,1.8445129,1.9331284,2.2350771,2.5698464,2.0184617,1.719795,1.6410258,1.6082052,1.2832822,1.1158975,1.1848207,1.3226668,1.4703591,1.6804104,1.6902566,1.5786668,1.4605129,1.4966155,1.910154,2.3433847,2.5796926,2.674872,2.6354873,2.412308,2.477949,2.6453335,3.1573336,3.56759,2.7470772,2.3860514,1.8018463,1.9232821,2.605949,2.609231,2.6256413,3.1737437,3.9056413,4.916513,6.738052,6.75118,6.8332314,7.3583593,7.6635904,6.0717955,6.262154,6.4590774,6.1472826,5.5958977,5.87159,6.2916927,6.2916927,6.8004107,8.205129,10.331899,11.0605135,11.641437,12.4685135,13.472821,14.122667,15.218873,14.230975,13.590976,14.093129,14.867694,12.773745,9.537642,7.3386674,6.5739493,5.8518977,6.5444107,7.0826674,7.0465646,7.026872,8.612103,7.8539495,7.5585647,7.2992826,6.944821,6.6395903,6.3442054,6.189949,6.2523084,6.554257,7.0432825,5.5696416,5.0609236,4.923077,4.522667,3.2098465,3.623385,2.9669745,2.2646155,1.9561027,1.9200002,1.3128207,1.4834872,1.723077,1.7526156,1.723077,3.5741541,3.5249233,3.9351797,5.172513,5.618872,4.4340515,3.0949745,2.0217438,1.7526156,2.9735386,5.221744,6.665847,6.1440005,4.6080003,5.093744,5.481026,4.8377438,4.240411,4.2535386,4.916513,4.71959,5.290667,6.2096415,7.1909747,8.080411,8.103385,9.800206,10.052924,8.723693,8.648206,8.03118,5.904411,6.432821,10.358154,14.979283,13.029744,11.611898,12.251899,13.988104,13.354668,10.742155,8.904206,7.3452315,6.3868723,7.1581545,8.1066675,7.9458466,7.4404106,6.925129,6.298257,8.516924,11.651283,13.22995,12.081232,8.36595,5.330052,4.397949,5.2020516,7.834257,12.829539,11.953232,9.888822,8.146052,7.939283,10.197334,12.86236,12.097642,9.757539,7.9261546,8.937026,9.16677,9.547488,10.801231,12.389745,12.49477,11.85477,10.916103,9.737847,8.454565,7.276308,5.9470773,6.1440005,7.003898,7.2960005,5.405539,4.844308,4.7589746,5.044513,5.221744,4.414359,4.0336413,3.0358977,2.0644104,1.4080001,1.024,0.98461545,1.5195899,1.585231,1.1323078,1.1093334,1.7788719,2.034872,2.038154,1.9954873,2.166154,2.156308,1.7723079,1.4736412,1.4145643,1.4408206,2.930872,4.0533338,4.637539,4.919795,5.5597954,4.1189747,2.9111798,2.5731285,2.8422565,2.556718,1.8806155,1.6246156,1.5458462,1.5031796,1.4441026,1.1946667,1.3095386,1.5163078,1.6016412,1.401436,1.5327181,2.0118976,2.2613335,2.2646155,2.5632823,2.5009232,2.3466668,2.228513,2.3105643,2.806154,2.6420515,2.6880002,3.4724104,4.309334,3.3017437,2.353231,1.8084104,2.1891284,3.2853336,4.128821,2.665026,2.1103592,3.5544617,5.677949,4.7491283,4.1911798,3.9056413,4.1780515,4.84759,5.284103,4.2568207,3.5380516,3.245949,3.5413337,4.647385,5.4186673,4.919795,4.1780515,3.8038976,3.9614363,9.347282,17.375181,19.331284,13.6697445,5.9995904,2.162872,0.9714873,0.6695385,0.4135385,0.26584616,0.52512825,1.4112822,2.809436,4.516103,6.2523084,7.240206,7.7292314,7.6668725,7.131898,6.3343596,6.380308,4.4242053,2.2088206,1.0108719,1.6508719,3.5183592,4.1878977,3.0358977,0.88943595,0.016410258,0.013128206,0.10502565,0.508718,1.0896411,1.3817437,0.65641034,0.20348719,0.04266667,0.06235898,0.013128206,0.049230773,0.13456412,0.17723078,0.13456412,0.013128206,0.06235898,0.14769232,0.15753847,0.08205129,0.0,0.0,0.0,0.009846155,0.029538464,0.04594872,0.108307704,0.28882053,0.51856416,0.6465641,0.44964105,0.15097436,0.032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.049230773,0.13784617,0.3052308,0.69251287,0.8205129,0.6826667,0.7581539,0.7220513,1.1552821,1.3620514,1.2865642,1.529436,1.5360001,1.2635899,1.4572309,2.028308,2.048,1.719795,1.9035898,2.540308,3.5314875,4.7228723,4.0303593,3.748103,4.0992823,4.955898,5.835488,7.7292314,11.503591,13.344822,13.472821,16.128002,15.31077,17.161848,17.302977,15.638975,16.347898,15.540514,13.8075905,11.684103,9.350565,6.6461544,4.7491283,4.460308,3.8531284,2.7700515,2.8225644,3.7054362,3.9187696,3.3247182,2.1464617,0.9682052,0.3249231,0.08533334,0.032820515,0.03938462,0.059076928,0.07876924,0.0951795,0.101743594,0.0951795,0.072205134,0.072205134,0.06564103,0.052512825,0.04594872,0.04594872,0.036102567,0.032820515,0.036102567,0.036102567,0.036102567,0.032820515,0.03938462,0.04594872,0.052512825,0.06235898,0.06235898,0.08205129,0.10502565,0.12471796,0.14112821,0.16410258,0.18707694,0.2231795,0.26584616,0.2855385,0.2855385,0.3314872,0.37743592,0.39712822,0.37415388,0.35446155,0.5152821,0.69907695,0.761436,0.57764107,0.5513847,0.702359,0.827077,0.90912825,1.1027694,1.5983591,1.211077,1.0896411,1.4080001,1.3522053,1.3456411,1.5589745,1.9003079,2.2482052,2.4484105,2.7241027,2.9833848,3.3280003,3.95159,5.149539,8.093539,9.865847,10.650257,10.791386,10.768411,10.57477,10.886565,11.45436,12.015591,12.288001,11.418258,9.580308,8.753231,11.638155,21.648413,31.90154,32.521847,26.151386,17.270155,12.196103,12.773745,15.711181,18.898052,21.014977,21.543386,22.633028,24.192001,26.148104,29.689438,37.264412,48.26585,58.29252,65.52944,68.5719,66.44842,61.105236,59.828518,60.550568,62.595287,66.67487,71.71611,72.85498,70.669136,66.93744,64.64001,67.76452,67.92206,65.424416,60.356926,52.58175,45.538464,40.021336,35.83016,32.561234,29.610668,26.535387,24.402054,22.75118,20.276514,14.841437,10.70277,7.936001,5.7403083,3.95159,3.0293336,2.7503593,2.4976413,2.6223593,3.0916924,3.4724104,3.308308,2.793026,1.9528207,1.083077,0.75487185,0.61374366,0.47589746,0.39384618,0.4397949,0.69251287,1.5261539,1.214359,0.9321026,1.276718,2.2777438,2.4155898,2.2153847,1.8937438,1.5130258,0.9714873,0.5907693,0.4201026,0.36102566,0.34133336,0.318359,0.41025645,1.3883078,1.4900514,0.56123084,0.055794876,0.009846155,0.006564103,0.01969231,0.06564103,0.2100513,0.25928208,0.13128206,0.04266667,0.09189744,0.256,0.5284103,0.80738467,1.7624617,3.754667,6.8660517,9.235693,11.306667,12.868924,13.735386,13.771488,10.043077,6.9120007,5.3858466,4.70318,2.3302567,3.2984617,7.640616,10.955488,10.709334,6.226052,2.6322052,0.86317956,0.21661541,0.10502565,0.068923086,0.052512825,0.04266667,0.06564103,0.12471796,0.2231795,1.0699488,0.9911796,0.8598975,1.1454359,1.9823592,3.170462,2.6322052,2.1103592,1.2274873,0.5284103,1.4736412,1.7887181,1.3784616,0.6301539,0.0,0.0,0.23958977,0.41025645,0.6268718,0.7089231,0.18379489,0.6662565,2.1136413,2.6978464,1.8838975,0.42994875,0.98133343,3.3542566,3.8859491,2.103795,0.7056411,0.24943592,0.28225642,0.6268718,1.1585642,1.8018463,2.412308,1.972513,2.4057438,3.186872,1.3522053,2.2153847,1.4375386,1.3784616,1.9331284,0.49887183,1.9626669,2.048,1.913436,1.7493335,0.76800007,0.35774362,0.20020515,0.46276927,1.2898463,2.802872,1.1257436,1.5524104,2.0906668,1.8116925,0.85005134,0.4594872,0.636718,1.2373334,1.6246156,0.69251287,0.44964105,0.3708718,0.37743592,0.42994875,0.49887183,0.33805132,0.5481026,0.99774367,1.5360001,1.9856411,1.9200002,1.7001027,1.5556924,1.5425643,1.5392822,1.6147693,1.8642052,2.166154,2.4385643,2.6190772,2.4582565,2.0873847,1.7887181,1.6771283,1.7033848,1.4998976,1.5130258,1.5425643,1.4309745,1.079795,0.94523084,0.94523084,0.9682052,0.9747693,1.0108719,1.2898463,1.4933335,1.5655385,1.6836925,2.2580514,2.6256413,2.7011285,2.6420515,2.4976413,2.2055387,2.1136413,2.1924105,3.1507695,4.1911798,2.9965131,3.8400004,3.4658465,2.9702566,2.8947694,3.2361028,4.3027697,4.7524104,4.916513,5.6254363,8.165744,7.030154,6.49518,6.547693,6.669129,5.8453336,5.077334,5.2480006,5.2480006,4.900103,4.9460516,4.7360005,4.3651285,4.5128207,5.481026,7.2205133,8.779488,9.747693,10.47959,10.781539,9.911796,10.282667,10.689642,11.365745,12.2387705,12.921437,12.383181,10.436924,8.057437,6.0980515,5.2676926,6.1013336,6.875898,6.806975,6.554257,8.241231,8.789334,9.4457445,9.393231,8.759795,8.602257,7.788308,6.488616,6.294975,7.194257,7.574975,6.0160003,5.7140517,5.5565133,4.8836927,3.4756925,3.0490258,2.5862565,2.0775387,1.6147693,1.3883078,1.4605129,1.9429746,2.0709746,1.9396925,2.487795,4.2830772,3.8990772,3.5216413,3.7940516,3.8334363,3.370667,2.5140514,1.6771283,1.5163078,2.917744,7.496206,8.89436,7.955693,5.917539,4.4340515,5.4974365,6.370462,6.229334,5.4153852,5.4482055,5.287385,5.4153852,5.9536414,6.8955903,8.067283,8.027898,8.792616,7.890052,5.8978467,6.4656415,6.550975,5.874872,6.2720003,7.765334,8.585847,7.4141545,7.269744,8.507077,10.095591,9.6065645,9.626257,8.973129,7.076103,5.4580517,7.7292314,9.4457445,8.697436,7.056411,5.989744,6.8562055,11.34277,14.913642,15.084309,11.588924,6.373744,4.6145644,4.4406157,4.955898,6.363898,9.96759,10.8307705,10.427077,9.334154,8.421744,8.848411,9.317744,8.759795,8.937026,10.673231,13.833847,14.601848,11.460924,9.373539,9.655796,9.980719,9.829744,10.157949,10.023385,9.133949,7.8473854,6.554257,6.3934364,6.7807183,6.9710774,6.0619493,5.3858466,5.218462,4.9099493,4.1189747,2.8356924,2.7011285,2.4418464,2.0611284,1.6705642,1.4703591,1.4342566,1.6738462,1.7263591,1.5163078,1.3522053,1.6935385,2.048,2.6289232,3.2886157,3.4855387,2.8980515,2.294154,2.0184617,2.156308,2.5337439,3.314872,3.5511796,3.7316926,3.9975388,4.1583595,3.0030773,1.910154,1.4802053,1.6147693,1.5031796,1.2242053,1.2209232,1.2504616,1.1979488,1.079795,0.9353847,0.83035904,0.8960001,1.1323078,1.401436,1.7526156,1.7788719,1.719795,1.8149745,2.2908719,2.4057438,2.484513,2.5009232,2.484513,2.5074873,1.9265642,1.6869745,2.7733335,4.4701543,4.3684106,3.2886157,3.0030773,3.1934361,3.6758976,4.397949,3.3411283,2.0644104,1.7493335,2.2055387,1.8642052,2.0873847,2.6715899,3.4002054,4.279795,5.536821,5.4482055,4.240411,3.5183592,4.2207184,6.629744,7.8802056,7.893334,7.6996927,7.9261546,8.802463,11.779283,14.8020525,13.617231,8.247795,3.0030773,1.2077949,0.571077,0.4201026,0.48902568,0.9288206,1.529436,1.9954873,2.934154,4.4800005,6.2818465,6.432821,7.3419495,7.24677,6.1505647,5.8486156,6.4032826,5.4843082,4.1124105,3.446154,4.7589746,5.034667,3.9286156,2.1398976,0.508718,0.016410258,0.006564103,0.016410258,0.21333335,0.5940513,0.96492314,0.32164106,0.07876924,0.026256412,0.03938462,0.04266667,0.04266667,0.068923086,0.08205129,0.06235898,0.0,0.12471796,0.108307704,0.06235898,0.029538464,0.009846155,0.0032820515,0.0,0.0032820515,0.013128206,0.013128206,0.02297436,0.101743594,0.27569234,0.4201026,0.26256412,0.08861539,0.02297436,0.016410258,0.026256412,0.026256412,0.101743594,0.14112821,0.108307704,0.029538464,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.01969231,0.06564103,0.18707694,0.4397949,0.56451285,0.69251287,1.3456411,1.4572309,1.3883078,1.2406155,1.1585642,1.3554872,1.4572309,1.1946667,1.4178462,2.0676925,2.172718,1.6049232,1.6640002,2.041436,2.6584618,3.6660516,3.9023592,3.892513,4.201026,5.2381544,7.259898,6.698667,9.577026,11.057232,10.801231,12.970668,13.801026,16.311796,15.993437,12.980514,12.058257,12.281437,11.930258,10.755282,8.756514,6.166975,3.9844105,2.986667,2.1103592,1.339077,1.6869745,2.5731285,2.300718,1.7033848,1.1815386,0.702359,0.256,0.06564103,0.013128206,0.013128206,0.01969231,0.04266667,0.06564103,0.07876924,0.07548718,0.06564103,0.06564103,0.068923086,0.06564103,0.052512825,0.04594872,0.032820515,0.029538464,0.029538464,0.029538464,0.02297436,0.02297436,0.026256412,0.029538464,0.03938462,0.04266667,0.04266667,0.049230773,0.06235898,0.08205129,0.101743594,0.118153855,0.14441027,0.18379489,0.21989745,0.24287182,0.25928208,0.32164106,0.40369233,0.46933338,0.48902568,0.49230772,0.49887183,0.54482055,0.58420515,0.49887183,0.4660513,0.512,0.56451285,0.6268718,0.77128214,1.0469744,0.88287187,0.8172308,0.92553854,0.8467693,0.86646163,1.014154,1.2800001,1.6640002,2.1956925,3.0391798,3.8137438,4.604718,5.346462,5.8157954,7.8637953,9.67877,10.886565,11.457642,11.71036,11.88759,11.930258,11.661129,10.965334,9.7903595,9.03877,8.277334,8.986258,12.540719,20.197744,21.910976,18.011898,11.877745,6.672411,5.3398976,8.457847,12.973949,17.929848,22.600206,26.50913,29.682875,30.391798,32.725334,38.85949,49.069954,49.16185,46.208004,43.602055,42.0759,39.686565,35.96472,35.91549,39.122055,45.876514,57.16021,70.00288,79.40267,84.46688,85.61888,84.61129,85.9077,87.3157,88.930466,88.3758,80.79755,71.25334,61.47611,53.42195,47.379696,41.96431,37.779694,34.835693,32.62031,30.12267,25.816618,20.466873,16.57436,13.243078,10.010257,6.8693337,5.691077,4.240411,3.117949,2.5173335,2.1989746,1.9889232,1.6410258,1.2373334,0.8730257,0.6695385,0.6695385,0.6498462,0.92553854,1.4998976,2.0709746,2.3236926,1.7132308,1.3554872,1.5622566,1.8609232,1.5327181,1.1651284,0.892718,0.69579494,0.41682056,0.21989745,0.15425642,0.14441027,0.19364104,0.36758977,0.98133343,1.4933335,1.3292309,0.5907693,0.052512825,0.016410258,0.052512825,0.21333335,0.58420515,1.2635899,1.1093334,0.571077,0.30851284,0.446359,0.5907693,0.8533334,1.2176411,1.9396925,3.7940516,8.080411,10.699488,12.432411,12.698257,12.3306675,13.581129,10.509129,6.941539,4.4767184,3.5478978,3.436308,9.271795,14.378668,17.634462,16.630156,7.6668725,3.436308,1.1881026,0.28882053,0.11158975,0.052512825,0.03938462,0.026256412,0.036102567,0.07876924,0.16738462,0.9189744,0.764718,0.7417436,1.3522053,2.4516926,3.2689233,2.0250258,1.6377437,1.3981539,1.1815386,1.4441026,1.4572309,1.5360001,0.9616411,0.01969231,0.0,0.013128206,0.27569234,1.1027694,1.847795,0.9156924,1.0436924,2.7437952,3.442872,2.3827693,0.6498462,1.2603078,3.131077,3.9384618,3.2000003,2.2547693,0.63343596,0.12143591,0.42994875,1.086359,1.4342566,2.048,1.8248206,2.2022567,2.7241027,1.0535386,1.8445129,1.0404103,1.3128207,2.674872,2.4910772,3.511795,3.6102567,3.0490258,1.9528207,0.3117949,0.25928208,0.21661541,0.57764107,1.5360001,3.0818465,0.90256417,0.26256412,0.6892308,1.2964103,0.79097444,0.42338464,0.48574364,0.69251287,0.761436,0.42994875,0.8041026,0.67282057,0.50543594,0.4955898,0.56123084,0.4266667,0.446359,0.67282057,1.0010257,1.1881026,1.0469744,1.014154,1.0502565,1.083077,1.014154,0.99774367,1.1979488,1.5753847,2.038154,2.422154,2.550154,2.3433847,1.8510771,1.2865642,1.0371283,1.1585642,1.2931283,1.2603078,1.0436924,0.77456415,0.75487185,0.75487185,0.7417436,0.7220513,0.77128214,1.2832822,1.6738462,1.9298463,2.1070771,2.349949,2.5698464,2.5665643,2.4549747,2.2711797,1.9790771,1.7263591,1.6246156,2.2678976,3.0523078,2.1792822,3.564308,4.194462,4.33559,4.3552823,4.6933336,6.0750775,6.7216415,7.125334,7.9097443,9.833026,7.9195905,6.8430777,6.741334,7.1122055,6.820103,5.9963083,6.0947695,6.12759,5.756718,5.293949,4.5095387,4.096,4.201026,4.8344617,5.8518977,7.9425645,9.649232,10.246565,9.800206,9.160206,9.275078,10.082462,10.840616,11.158976,10.985026,11.011283,10.443488,8.907488,6.806975,5.32677,5.920821,6.8496413,6.8496413,6.3540516,7.4863596,8.539898,9.563898,9.655796,8.900924,8.36595,7.712821,6.554257,6.6034875,7.5585647,7.1220517,5.8190775,5.717334,5.5532312,4.6834874,3.1113849,2.3401027,2.4516926,2.5042052,2.2678976,2.231795,2.2711797,2.802872,2.8127182,2.422154,2.9013336,4.013949,3.9844105,3.4330258,2.9111798,2.8882053,3.1343591,2.4615386,1.9298463,2.28759,3.9614363,9.353847,10.348309,8.835282,6.51159,4.854154,5.927385,7.702975,7.650462,6.0258465,5.8880005,5.61559,5.425231,5.920821,7.072821,8.208411,7.571693,7.529026,6.6428723,5.4416413,6.4295387,6.121026,6.0750775,6.232616,6.2063594,5.3070774,6.0258465,7.9195905,9.593436,10.006975,8.490667,8.900924,8.897642,8.01477,7.2664623,9.127385,9.895386,8.425026,6.5805135,5.677949,6.498462,10.765129,14.427898,14.355694,10.499283,5.8945646,5.648411,5.366154,5.5958977,6.8988724,9.83959,10.965334,10.226872,8.897642,7.785026,7.194257,7.059693,7.680001,9.248821,11.552821,13.961847,14.946463,11.690667,9.573745,9.905231,9.911796,10.397539,11.093334,11.109744,10.246565,8.992821,7.7456417,6.961231,6.698667,6.619898,5.9569235,5.152821,4.598154,3.9023592,3.0326157,2.3171284,2.2350771,2.0939488,1.9954873,1.9429746,1.8379488,1.7427694,1.7558975,1.7788719,1.6607181,1.1979488,1.276718,1.6344616,2.4188719,3.442872,4.1878977,2.9965131,2.3401027,2.231795,2.487795,2.7175386,2.8422565,3.117949,3.4691284,3.5610259,2.809436,1.7165129,1.2077949,1.204513,1.3915899,1.2274873,1.1158975,1.332513,1.4276924,1.2242053,0.82379496,0.8402052,0.7417436,0.7450257,1.0305642,1.7427694,1.8445129,1.7755898,2.0250258,2.477949,2.4024618,2.5796926,2.6945643,2.5140514,2.1267693,1.9659488,1.5327181,1.1093334,2.044718,4.06318,5.2709746,4.0336413,3.6758976,3.5282054,3.3411283,3.2853336,2.6190772,1.8937438,1.6049232,1.6640002,1.394872,1.4998976,2.6912823,3.895795,4.8114877,5.901129,6.196513,4.923077,3.6726158,3.8564105,6.7183595,8.756514,9.734565,10.033232,10.075898,10.33518,10.082462,9.101129,6.7577443,3.56759,1.1848207,0.6826667,0.39712822,0.4135385,0.76800007,1.4211283,2.0086155,2.0151796,2.4451284,3.5872824,4.9985647,4.844308,5.8518977,5.83877,4.7917953,4.890257,5.7764106,5.8190775,5.786257,6.2720003,7.6668725,6.1538467,3.7940516,1.6410258,0.318359,0.016410258,0.0032820515,0.0,0.06235898,0.22646156,0.52512825,0.128,0.04594872,0.072205134,0.08861539,0.049230773,0.049230773,0.029538464,0.009846155,0.0,0.0,0.1148718,0.068923086,0.009846155,0.0032820515,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.06564103,0.14441027,0.07876924,0.23958977,0.380718,0.5874872,0.7975385,0.8041026,0.47589746,0.27569234,0.13456412,0.029538464,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.02297436,0.0951795,0.20676924,0.36430773,0.69251287,1.4572309,1.9429746,1.7952822,1.5425643,1.4769232,1.654154,1.3718976,1.1257436,1.3489232,1.9298463,2.1858463,1.7394873,1.595077,1.7558975,2.2678976,3.2196925,3.4560003,3.7382567,3.895795,4.457026,6.619898,6.052103,8.0377445,9.298052,9.32759,10.371283,12.704822,15.602873,15.872002,12.895181,8.6580515,8.470975,8.710565,8.392206,7.1483083,5.208616,3.114667,1.6410258,0.7384616,0.38728207,0.6268718,1.2373334,0.8008206,0.56123084,0.7975385,0.83035904,0.2231795,0.029538464,0.0,0.0,0.0,0.01969231,0.03938462,0.052512825,0.055794876,0.06235898,0.06235898,0.06235898,0.06235898,0.059076928,0.052512825,0.03938462,0.032820515,0.029538464,0.029538464,0.02297436,0.016410258,0.016410258,0.01969231,0.026256412,0.029538464,0.026256412,0.029538464,0.032820515,0.03938462,0.059076928,0.06564103,0.08861539,0.118153855,0.14441027,0.16410258,0.18379489,0.24287182,0.3117949,0.36758977,0.40369233,0.44307697,0.45292312,0.5677949,0.7384616,0.7187693,0.69907695,0.8041026,0.76800007,0.6170257,0.6629744,0.77128214,0.8172308,0.8402052,0.8467693,0.8402052,0.8598975,0.96492314,1.1454359,1.4244103,1.8806155,2.8291285,3.817026,4.9427695,6.045539,6.695385,7.512616,8.477539,9.245539,9.734565,10.121847,10.33518,10.837335,11.23118,11.008,9.540924,8.421744,8.04759,9.472001,12.855796,17.480206,14.01436,8.310155,3.8006158,1.9922053,2.477949,5.5532312,9.944616,14.76595,19.958155,26.285952,33.152004,38.052105,46.047184,57.22585,66.733955,52.548927,36.230568,26.262976,24.523489,26.289232,27.72349,29.456413,33.22421,40.10667,50.52062,63.737442,76.80329,87.282875,94.20473,98.10052,99.97457,100.94278,102.25232,103.0236,100.2437,96.80739,88.86154,78.35898,67.508514,58.755287,52.772106,47.51426,43.53313,40.49067,37.16267,31.61272,27.411694,23.936003,20.38154,15.766975,12.409437,8.644924,5.8945646,4.4340515,3.3772311,2.166154,1.3883078,0.9189744,0.6662565,0.58420515,0.6235898,0.6170257,0.88615394,1.4178462,1.8707694,1.7033848,1.2176411,0.97805136,1.014154,0.84348726,0.508718,0.24943592,0.12471796,0.11158975,0.11158975,0.07548718,0.059076928,0.055794876,0.118153855,0.32820517,0.88287187,0.88287187,0.6465641,0.3708718,0.12471796,0.18707694,0.27241027,0.62030774,1.3128207,2.2646155,1.9331284,1.1881026,0.8467693,1.0371283,1.1651284,1.4966155,2.281026,2.861949,4.007385,7.9228725,10.059488,10.745437,9.882257,9.065026,11.608616,9.974154,6.3376417,3.370667,2.5206156,4.017231,10.916103,14.119386,14.966155,12.872206,5.333334,2.5042052,0.9288206,0.256,0.10502565,0.04594872,0.029538464,0.01969231,0.016410258,0.029538464,0.068923086,1.086359,1.1848207,0.827077,0.83035904,1.1224617,0.74830776,0.571077,0.88287187,1.394872,1.6738462,1.1520001,1.5130258,1.8248206,1.2012309,0.049230773,0.04594872,0.026256412,0.16082053,1.1913847,2.4352822,1.8182565,1.1881026,2.1202054,2.4976413,1.7099489,0.63343596,2.2613335,2.674872,2.537026,2.5042052,3.245949,0.86317956,0.16738462,0.6268718,1.4080001,1.3850257,3.0260515,2.100513,0.7844103,0.118153855,0.0,0.0,0.04594872,0.48902568,1.7099489,4.125539,3.7218463,3.7710772,3.0523078,1.591795,0.64000005,0.45620516,0.574359,0.8172308,1.0338463,1.0962052,0.26256412,0.24943592,0.5940513,0.82379496,0.4660513,0.3314872,0.3314872,0.4135385,0.53825647,0.6892308,1.5327181,1.2504616,0.8402052,0.7253334,0.76800007,0.69251287,0.6170257,0.6235898,0.65969235,0.5481026,0.46933338,0.5907693,0.7187693,0.77128214,0.761436,0.7417436,0.8730257,1.2012309,1.6049232,1.8215386,2.15959,2.3269746,1.9232821,1.1815386,0.9714873,1.1257436,1.1027694,0.95835906,0.75487185,0.571077,0.6498462,0.69251287,0.74830776,0.8992821,1.2832822,1.8543591,2.162872,2.4155898,2.553436,2.2449234,2.2777438,2.422154,2.4418464,2.294154,2.1267693,2.1300514,1.8379488,1.5195899,1.3095386,1.2012309,2.2186668,3.761231,5.1659493,6.0816417,6.47877,6.813539,7.7325134,9.051898,10.282667,10.640411,8.933744,7.64718,7.716103,8.674462,8.65477,8.740103,8.690872,8.457847,7.939283,6.9809237,5.8190775,5.5926156,5.8880005,6.232616,6.1078978,8.15918,10.072617,10.417232,9.701744,10.377847,10.43036,10.157949,9.747693,9.409642,9.383386,9.330873,9.104411,8.425026,7.177847,5.412103,5.402257,6.498462,6.8266673,6.232616,6.2785645,6.4590774,7.381334,7.8670774,7.3747697,5.9930263,6.0750775,6.235898,6.8266673,7.328821,6.3277955,5.4908724,5.172513,4.7950773,3.9876926,2.605949,2.3171284,2.934154,3.4002054,3.4822567,3.761231,3.1277952,3.7218463,3.761231,2.993231,2.6880002,3.1277952,3.889231,3.8990772,3.2918978,3.4133337,3.9187696,3.255795,3.006359,3.9286156,5.9470773,10.276103,10.896411,8.786052,6.0980515,6.1538467,6.12759,7.394462,7.059693,5.284103,5.284103,4.9952826,5.0871797,5.924103,7.2205133,8.054154,6.770872,5.8978467,5.5958977,6.0783596,7.5913854,7.0957956,6.422975,5.8223596,5.5762057,5.986462,9.278359,12.78359,14.27036,12.960821,9.508103,8.746667,8.789334,9.176616,9.596719,9.878975,8.726975,7.069539,6.2194877,6.1997952,5.7665644,8.018052,11.428103,12.097642,9.5606165,6.7905645,6.8233852,5.858462,6.0356927,8.011488,10.932513,10.354873,7.77518,6.180103,6.4065647,7.125334,8.283898,10.029949,11.053949,11.221334,11.605334,13.095386,12.698257,12.914873,13.938873,13.682873,14.720001,14.634667,13.384206,11.47077,9.961026,9.314463,8.786052,8.717129,8.612103,7.1548724,5.9503593,4.6966157,3.698872,3.2164104,3.4592824,3.2689233,2.6912823,2.3335385,2.3368206,2.356513,2.225231,2.2646155,2.0873847,1.5819489,0.8992821,1.0568206,1.3489232,1.6836925,2.1891284,3.2131286,2.3860514,1.9200002,2.034872,2.428718,2.2711797,2.4746668,3.7218463,4.417641,3.8596926,2.2449234,1.2832822,1.7788719,2.409026,2.4910772,1.9790771,1.5819489,1.7690258,1.7558975,1.3029745,0.7056411,0.88615394,0.98461545,0.9714873,1.0896411,1.8740515,1.8379488,2.3072822,3.1671798,3.7743592,2.9735386,2.8389745,2.6847181,2.1792822,1.6902566,2.28759,3.0424619,2.665026,2.8356924,4.096,5.8190775,5.0904617,4.650667,4.06318,3.1638978,2.044718,1.4080001,1.4998976,1.5458462,1.2635899,0.8566154,1.4408206,3.4888208,5.113436,5.72718,6.0225644,6.432821,5.986462,4.667077,3.6332312,5.221744,7.0334363,8.208411,8.3593855,7.653744,6.813539,5.172513,3.511795,2.2383592,1.4998976,1.1815386,0.74830776,0.5907693,0.761436,1.1388719,1.4244103,1.6705642,1.7296412,2.038154,2.550154,2.7470772,2.9013336,3.6529233,3.8071797,3.3903592,3.636513,4.4373336,5.0182567,6.2523084,7.9294367,8.763078,6.055385,3.6758976,1.7493335,0.4660513,0.06235898,0.013128206,0.006564103,0.013128206,0.04266667,0.14441027,0.072205134,0.10502565,0.19364104,0.22646156,0.03938462,0.06564103,0.052512825,0.02297436,0.0,0.0032820515,0.009846155,0.0032820515,0.006564103,0.016410258,0.026256412,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.009846155,0.032820515,0.08533334,0.5218462,0.9682052,1.4178462,1.7165129,1.5688206,0.7515898,0.27241027,0.052512825,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.059076928,0.055794876,0.026256412,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.06235898,0.11158975,0.256,0.49887183,0.761436,1.654154,2.0611284,2.166154,2.1792822,2.3466668,1.3883078,1.3062565,1.467077,1.6475899,2.0151796,1.9035898,1.4506668,1.4703591,2.2646155,3.6069746,2.9965131,3.2656412,3.2164104,3.0949745,4.5817437,7.0793853,8.513641,9.67877,10.633847,10.71918,12.2847185,14.720001,16.439796,15.638975,10.312206,7.8145647,6.7971287,6.413129,5.8486156,4.309334,2.2350771,0.9485129,0.36758977,0.2231795,0.06564103,0.27569234,0.16738462,0.5284103,1.2537436,1.332513,0.30194873,0.01969231,0.0,0.0,0.0,0.009846155,0.02297436,0.032820515,0.04594872,0.059076928,0.055794876,0.049230773,0.052512825,0.06235898,0.06235898,0.049230773,0.03938462,0.032820515,0.029538464,0.032820515,0.02297436,0.01969231,0.01969231,0.01969231,0.029538464,0.01969231,0.02297436,0.02297436,0.016410258,0.026256412,0.029538464,0.03938462,0.055794876,0.07548718,0.09189744,0.10502565,0.13784617,0.16082053,0.16410258,0.17723078,0.21661541,0.3052308,0.58420515,0.9189744,0.90256417,1.1027694,1.3292309,1.2209232,0.8730257,0.827077,0.8960001,1.014154,1.1323078,1.2176411,1.2406155,1.1979488,1.1716924,1.2012309,1.3226668,1.5786668,2.1924105,3.045744,4.194462,5.684513,7.525744,8.769642,8.845129,8.342975,7.788308,7.6603084,7.578257,8.759795,10.456616,11.69395,11.257437,9.728001,8.746667,8.960001,10.066052,10.817642,6.9054365,3.495385,1.654154,1.463795,2.0250258,3.515077,5.98318,9.084719,13.35795,20.233849,29.909336,41.012516,55.440414,69.4318,73.567184,48.94195,27.024412,15.944206,16.873028,24.018053,31.461746,36.804924,41.590157,46.29662,50.33026,56.42503,65.19139,74.85375,84.67693,94.959595,101.56637,102.84309,102.009445,101.98975,105.41293,113.71652,113.7756,105.00596,91.083496,79.92452,71.24677,63.021954,56.76308,52.394672,48.275696,42.57149,38.311386,35.252514,32.341335,27.720207,21.799387,15.448617,10.817642,8.231385,6.166975,3.5610259,1.9889232,1.1191796,0.7122052,0.6268718,0.5513847,0.45292312,0.3708718,0.3314872,0.3314872,0.29538465,0.21989745,0.15097436,0.12143591,0.12471796,0.108307704,0.072205134,0.03938462,0.02297436,0.02297436,0.029538464,0.02297436,0.02297436,0.052512825,0.11158975,0.16082053,0.15097436,0.128,0.16082053,0.3446154,0.5415385,0.764718,1.3554872,2.2744617,3.1245131,3.0162053,2.3762052,1.9495386,1.9495386,2.0545642,2.4582565,3.6857438,4.1189747,4.1452312,6.173539,7.9491286,8.241231,7.1089234,6.2129235,8.815591,8.730257,5.651693,3.2131286,2.6551797,2.806154,5.733744,5.9602056,4.4800005,2.4516926,1.2012309,0.6235898,0.28225642,0.12471796,0.072205134,0.04266667,0.01969231,0.016410258,0.009846155,0.0032820515,0.016410258,0.5481026,0.5973334,0.46276927,0.41025645,0.39384618,0.07548718,0.12471796,0.2297436,0.49230772,0.892718,1.2964103,1.5885129,1.2340513,0.5677949,0.04594872,0.2297436,0.13128206,0.04266667,0.22646156,0.80738467,1.7690258,2.1858463,2.1234872,2.4352822,2.6486156,0.97805136,1.3915899,1.6147693,1.723077,1.5622566,0.7318975,0.18379489,0.036102567,0.13456412,0.3249231,0.45620516,0.16410258,0.036102567,0.0,0.0,0.0,0.0,0.009846155,0.026256412,0.098461546,0.3052308,0.28225642,0.5874872,1.0075898,1.5195899,2.28759,1.214359,1.8051283,2.2711797,1.7427694,0.28882053,0.27897438,0.5940513,0.7220513,0.5513847,0.380718,0.380718,0.380718,0.44964105,0.65312827,1.0666667,2.0578463,1.8182565,1.3259488,1.0502565,0.97805136,0.83035904,0.7122052,0.62030774,0.512,0.3052308,0.29210258,0.41025645,0.52512825,0.5874872,0.6268718,0.67282057,0.7220513,0.8402052,1.017436,1.1749744,1.5885129,1.6311796,1.3259488,0.95835906,1.0666667,1.1651284,0.9878975,0.8172308,0.69251287,0.4135385,0.55794877,0.7220513,1.0469744,1.6475899,2.6256413,2.7963078,2.7175386,2.5731285,2.3794873,2.0151796,2.0250258,2.3401027,2.4615386,2.359795,2.4582565,3.6890259,3.3017437,2.5435898,2.044718,1.8018463,3.3641028,4.240411,4.9099493,5.684513,6.698667,5.3924108,6.12759,7.250052,7.896616,7.9819493,7.1515903,6.311385,6.8299494,8.690872,10.499283,10.679795,10.112,9.386667,8.631796,7.506052,6.518154,6.6002054,7.4174366,8.155898,7.522462,9.048616,9.540924,9.380103,9.061745,9.170052,8.011488,7.282872,6.9349747,6.882462,7.003898,6.491898,6.2063594,5.865026,5.605744,5.9963083,5.3136415,6.166975,6.764308,6.413129,5.5072823,5.83877,7.466667,8.283898,7.5191803,5.737026,6.1538467,6.0652313,5.85518,5.792821,6.012718,6.5017443,5.211898,3.9548721,3.436308,3.2656412,3.4231799,3.5446157,3.761231,4.017231,4.089436,3.4658465,4.4734364,4.7983594,3.9351797,3.190154,3.190154,3.7743592,4.086154,3.8531284,3.4034874,3.879385,4.2174363,4.338872,4.9099493,7.3386674,10.282667,11.044104,8.937026,5.717334,5.5696416,5.7632823,5.4482055,4.972308,4.4406157,3.7087183,3.5872824,4.414359,5.5696416,6.416411,6.3310776,5.3431797,4.44718,4.453744,5.504,7.0793853,8.54318,6.685539,4.667077,4.1189747,5.156103,8.868103,10.712616,11.053949,10.023385,7.506052,7.213949,8.149334,8.15918,7.3025646,7.827693,6.0225644,6.5312824,7.397744,7.5881033,6.987488,8.234667,9.114257,8.136206,5.8880005,5.0215387,5.7764106,4.493129,3.8038976,4.7556925,6.806975,5.976616,4.532513,4.8114877,7.3452315,10.84718,14.096412,17.14872,18.497643,18.720821,20.49313,23.151592,21.812515,18.58954,15.91795,16.54154,17.956104,18.500925,16.886156,13.512206,10.499283,11.756309,13.279181,14.322873,14.162052,12.100924,10.220308,8.871386,7.181129,5.425231,5.034667,4.670359,3.892513,3.3050258,3.259077,3.8465643,3.7842054,3.639795,2.92759,1.8642052,1.3883078,1.8281027,2.2482052,2.169436,1.5786668,0.9321026,2.8488207,2.4648206,2.28759,2.989949,3.4166157,3.6004105,4.6178465,4.84759,3.8334363,2.2580514,2.6715899,4.1517954,4.3684106,3.245949,2.930872,2.0742567,1.6410258,1.142154,0.6071795,0.5940513,1.1093334,1.0699488,0.9747693,1.1782565,1.9232821,2.9111798,3.3247182,3.249231,3.058872,3.387077,2.6190772,2.041436,1.785436,2.4582565,5.156103,8.195283,8.132924,6.8266673,5.85518,6.514872,8.884514,9.209436,7.640616,5.1331286,3.4494362,2.3138463,2.2219489,1.9396925,1.3095386,1.2373334,2.737231,3.9745643,4.0533338,3.56759,4.59159,6.9382567,8.300308,8.618668,8.12636,7.3682055,4.7589746,4.013949,3.9876926,4.0434875,4.0434875,3.495385,2.7798977,1.9331284,1.1946667,1.020718,0.86317956,1.1618463,1.5031796,1.6082052,1.3259488,1.2406155,1.7887181,2.3729234,2.6617439,2.5632823,2.4155898,3.0752823,3.2656412,2.806154,2.6256413,3.1606157,3.9909747,5.297231,6.73477,7.430565,5.5269747,4.5095387,3.0391798,1.148718,0.24287182,0.06235898,0.032820515,0.03938462,0.032820515,0.04594872,0.08205129,0.16410258,0.2855385,0.3314872,0.07548718,0.052512825,0.026256412,0.009846155,0.0032820515,0.016410258,0.0032820515,0.0,0.029538464,0.08861539,0.13784617,0.052512825,0.013128206,0.0,0.0,0.0,0.0,0.0,0.01969231,0.072205134,0.18379489,0.4135385,1.1323078,1.3686155,0.8730257,0.09189744,0.01969231,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.04594872,0.30194873,0.28225642,0.13784617,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.049230773,0.068923086,0.108307704,0.190359,0.33476925,0.88615394,1.8281027,2.425436,2.5173335,2.5173335,1.4441026,2.0644104,2.484513,2.172718,1.9528207,2.038154,2.1234872,2.2777438,2.6551797,3.508513,3.1442053,2.6683078,2.550154,3.2754874,5.32677,8.402052,8.602257,9.708308,11.979488,12.160001,10.561642,11.224616,13.367796,15.829334,17.073233,14.060308,8.992821,5.930667,5.0904617,2.868513,0.69579494,0.20676924,0.23302566,0.17394873,0.016410258,0.0032820515,0.0,0.0,0.15097436,0.74830776,0.28225642,0.06564103,0.0,0.0,0.0,0.0,0.009846155,0.02297436,0.032820515,0.04594872,0.032820515,0.03938462,0.052512825,0.06235898,0.06235898,0.049230773,0.055794876,0.049230773,0.032820515,0.04594872,0.04594872,0.036102567,0.029538464,0.029538464,0.029538464,0.01969231,0.016410258,0.016410258,0.016410258,0.016410258,0.026256412,0.03938462,0.052512825,0.06564103,0.09189744,0.10502565,0.1148718,0.128,0.14112821,0.15097436,0.15097436,0.190359,0.23958977,0.3052308,0.4266667,1.3292309,1.2996924,1.2012309,1.2668719,1.083077,1.2307693,1.3292309,1.3915899,1.4506668,1.5721027,1.6443079,1.4703591,1.2996924,1.2603078,1.3587693,1.7493335,2.4057438,3.3017437,4.841026,7.8441033,12.983796,14.020925,12.57354,10.161232,8.208411,8.2445135,8.182155,8.36595,8.999385,10.148104,10.893129,10.948924,10.016821,8.375795,6.9120007,3.8498464,1.9462565,1.2635899,1.5392822,2.1956925,2.8553848,4.1189747,6.806975,11.35918,17.85436,23.35836,29.96185,38.60021,45.856823,43.979492,21.930668,12.199386,10.561642,14.592001,23.650463,38.019283,49.903595,57.941338,62.194878,64.1477,61.76821,57.649235,55.32226,58.033234,68.72616,79.15324,87.5717,95.24842,101.848625,105.439186,117.95037,125.13478,124.698265,116.94934,104.766365,91.897446,81.916725,73.731285,66.42544,59.247593,51.679184,45.942158,42.213745,39.489643,35.584003,29.321848,22.472206,16.705643,12.47836,9.048616,5.7764106,3.4756925,1.9364104,1.0666667,0.86974365,0.69907695,0.508718,0.3708718,0.29538465,0.25928208,0.2231795,0.16738462,0.12471796,0.101743594,0.07548718,0.03938462,0.02297436,0.009846155,0.0,0.0,0.02297436,0.02297436,0.009846155,0.0032820515,0.016410258,0.016410258,0.016410258,0.04594872,0.2231795,0.74830776,0.955077,1.585231,2.6223593,3.820308,4.699898,5.6287184,5.100308,4.1583595,3.5183592,3.5544617,3.6660516,4.8377438,4.824616,3.5872824,3.2820516,7.125334,10.184206,9.6295395,6.889026,7.643898,6.5837955,4.394667,3.754667,4.0402055,1.3423591,0.7450257,0.5874872,0.43323082,0.190359,0.09189744,0.07876924,0.049230773,0.029538464,0.029538464,0.029538464,0.01969231,0.016410258,0.009846155,0.0032820515,0.016410258,0.512,0.6104616,0.4660513,0.2986667,0.18707694,0.07548718,0.036102567,0.04594872,0.098461546,0.18051283,0.25928208,3.255795,2.5862565,1.0929232,0.7253334,2.546872,3.9844105,1.7952822,0.10502565,0.4004103,1.5491283,2.5993848,3.1803079,3.3936412,3.0326157,1.5753847,2.917744,2.1267693,1.4375386,1.6804104,2.294154,3.0818465,2.7503593,1.5360001,0.2100513,0.09189744,0.13128206,0.128,0.072205134,0.09189744,0.46276927,0.6104616,0.78769237,0.6170257,0.51856416,1.719795,0.38728207,0.32820517,0.892718,1.4966155,1.6311796,1.3554872,1.4145643,1.3292309,0.86974365,0.08205129,0.07876924,0.2100513,0.30851284,0.30851284,0.23630771,0.36102566,0.4004103,0.46933338,0.63343596,0.92225647,1.3062565,1.2964103,1.1520001,1.020718,0.9288206,0.7811283,0.6695385,0.56451285,0.43323082,0.256,0.19692309,0.20348719,0.24287182,0.31507695,0.47917953,0.6662565,0.6892308,0.6695385,0.72861546,1.0043077,1.595077,2.0808206,1.8642052,1.276718,1.591795,1.4080001,1.3587693,1.2209232,0.9616411,0.72861546,0.90584624,1.0994873,1.3062565,1.6246156,2.2580514,2.3401027,2.425436,2.6322052,2.7109745,2.0512822,2.1300514,2.8422565,2.989949,3.0227695,5.044513,6.432821,6.042257,5.07077,4.3552823,4.3651285,5.9470773,6.439385,6.547693,6.705231,7.066257,4.8607183,4.0533338,4.6244106,5.7665644,5.8814363,7.453539,7.030154,6.764308,7.430565,8.448001,9.088,9.304616,9.324308,9.199591,8.789334,7.6635904,7.02359,7.3714876,8.369231,8.828718,9.8363085,10.029949,10.036513,10.112,10.121847,8.592411,9.18318,9.275078,8.316719,7.834257,8.152616,6.9021544,5.2315903,4.059898,4.066462,3.882667,5.0215387,6.73477,8.024616,7.6570263,6.744616,7.640616,8.605539,8.802463,8.300308,9.068309,8.474257,8.500513,8.986258,7.6242056,8.306872,7.27959,5.7042055,4.4701543,4.1813335,4.338872,3.9122055,3.570872,3.4789746,3.308308,3.3411283,4.4373336,4.7622566,4.1452312,4.092718,4.4340515,4.1156926,3.5446157,3.1113849,3.2065644,4.1025643,4.562052,4.263385,3.7152824,4.2502565,5.2020516,5.3398976,5.2414365,5.330052,5.8880005,5.156103,4.1583595,3.895795,4.381539,4.634257,3.751385,4.3027697,5.179077,5.691077,5.5762057,4.9493337,4.7491283,4.673641,5.0182567,6.701949,7.8539495,6.5772314,4.923077,4.1091285,4.522667,5.930667,6.9842057,7.466667,7.6898465,8.4972315,9.012513,8.326565,6.488616,4.525949,4.44718,4.1714873,4.4373336,5.152821,5.9470773,6.157129,6.8365135,6.636308,6.0849237,5.8781543,6.889026,7.194257,5.9963083,4.460308,3.6594875,4.5587697,3.748103,4.135385,7.128616,12.383181,17.769028,20.752413,24.050873,26.660105,29.134771,33.588516,32.97149,27.375591,21.536821,18.153027,17.906874,22.35077,23.332104,21.812515,18.970259,16.196924,13.033027,10.666668,8.4972315,6.6625648,6.0324106,6.048821,5.481026,4.8738465,4.7556925,5.6451287,4.594872,3.889231,4.1091285,4.7950773,4.4438977,3.4560003,3.826872,3.7218463,2.986667,3.1343591,3.1540515,2.6354873,1.9003079,1.2274873,0.8467693,2.4976413,2.556718,2.3204105,2.4484105,2.9538465,4.466872,5.8880005,5.937231,4.788513,4.0533338,3.5774362,3.5446157,3.1540515,2.4451284,2.284308,1.5163078,1.3095386,0.9714873,0.574359,0.9616411,1.7165129,1.4572309,1.467077,1.9954873,2.2514873,2.2449234,2.6945643,2.7766156,2.3302567,1.8510771,3.6791797,3.05559,2.9210258,4.6900516,8.257642,8.093539,7.384616,7.4830775,7.955693,6.564103,9.498257,11.805539,11.848206,9.275078,5.0215387,2.15959,1.3718976,1.7296412,2.5600002,3.446154,5.113436,4.5587697,4.263385,5.5532312,8.621949,10.65354,10.722463,8.999385,6.521436,5.1987696,5.504,5.2644105,5.169231,5.142975,4.312616,2.6584618,1.9331284,1.6114873,1.4145643,1.3029745,1.1848207,1.7788719,2.162872,1.8904617,0.98461545,0.88943595,1.339077,1.9298463,2.3762052,2.5009232,2.2088206,2.0053334,1.6968206,1.404718,1.5622566,2.412308,3.2164104,3.879385,4.4045134,4.903385,5.3234878,4.890257,3.442872,1.5130258,0.318359,0.20348719,0.118153855,0.08533334,0.07876924,0.02297436,0.03938462,0.049230773,0.068923086,0.07548718,0.016410258,0.009846155,0.006564103,0.0032820515,0.0032820515,0.016410258,0.013128206,0.128,0.21333335,0.18379489,0.026256412,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.036102567,0.08205129,0.22646156,0.27569234,0.17394873,0.01969231,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.059076928,0.055794876,0.026256412,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03938462,0.036102567,0.032820515,0.059076928,0.128,0.45292312,1.3981539,2.3433847,2.7700515,2.2744617,2.0086155,2.4648206,2.6289232,2.2055387,1.6246156,1.972513,2.7011285,2.8980515,2.3958976,1.7755898,2.356513,2.4385643,2.681436,3.3805132,4.4832826,8.681026,9.38995,9.462154,9.724719,8.999385,8.710565,8.27077,10.8537445,14.464001,11.959796,6.738052,4.5489235,3.2656412,1.913436,0.65969235,0.15753847,0.04266667,0.04594872,0.036102567,0.0032820515,0.0,0.0,0.0,0.029538464,0.15097436,0.055794876,0.013128206,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.01969231,0.02297436,0.029538464,0.032820515,0.04594872,0.06235898,0.06235898,0.059076928,0.059076928,0.059076928,0.055794876,0.059076928,0.049230773,0.04266667,0.049230773,0.052512825,0.04266667,0.03938462,0.04594872,0.04594872,0.04266667,0.052512825,0.04594872,0.059076928,0.07548718,0.0951795,0.128,0.13128206,0.14112821,0.14769232,0.15097436,0.15097436,0.16082053,0.18707694,0.21989745,0.26256412,0.3052308,0.52512825,0.5513847,0.58420515,0.6892308,0.7778462,0.9747693,1.1224617,1.2668719,1.4112822,1.522872,1.595077,1.5983591,1.5622566,1.5130258,1.4441026,1.5031796,1.8182565,2.4516926,3.5314875,5.2545643,8.910769,11.74318,12.2617445,10.532104,8.198565,7.64718,7.5618467,7.9195905,8.710565,9.915077,10.210463,10.308924,10.095591,9.219283,7.1187696,4.601436,2.537026,1.522872,1.6902566,2.7109745,3.7710772,4.210872,4.962462,7.0892315,11.785847,16.003283,17.670565,18.743795,19.029335,16.180513,10.94236,8.480822,9.025641,12.901745,20.512821,29.571285,42.23672,53.0478,60.051697,64.80739,65.1717,63.54708,58.19734,50.98667,47.363285,48.62031,51.780926,57.678772,66.33354,76.97395,91.29355,104.68432,115.885956,121.49498,115.97129,107.15898,96.06565,87.3518,80.909134,71.84739,66.15303,56.18216,48.928825,45.54831,41.37026,35.75139,29.233232,23.161438,18.15631,14.102976,10.781539,7.962257,5.5663595,3.6726158,2.5304618,1.9692309,1.6082052,1.3522053,1.1224617,0.86974365,0.636718,0.47589746,0.35446155,0.256,0.17394873,0.098461546,0.03938462,0.009846155,0.0,0.0,0.013128206,0.02297436,0.016410258,0.0,0.0032820515,0.0032820515,0.0032820515,0.049230773,0.23302566,0.69907695,0.86646163,1.5589745,2.8553848,5.10359,8.923898,9.403078,8.579283,7.9163084,7.8047185,7.5454364,5.4383593,5.4514875,6.5805135,7.8473854,8.283898,9.163487,12.2847185,16.65313,17.706669,7.3025646,5.7534366,3.9680004,3.245949,3.6069746,3.8071797,1.1881026,0.36430773,0.18051283,0.072205134,0.04266667,0.029538464,0.02297436,0.013128206,0.009846155,0.01969231,0.006564103,0.0032820515,0.006564103,0.009846155,0.0032820515,1.4998976,0.79097444,0.4004103,0.20676924,0.10502565,0.029538464,0.33476925,0.636718,0.62030774,0.4201026,0.64000005,2.3663592,2.4451284,1.4539489,0.6465641,1.9659488,2.5764105,1.1191796,0.072205134,0.45620516,1.8445129,1.719795,1.6344616,1.5360001,1.3128207,0.77128214,1.7526156,1.3193847,0.8795898,0.9616411,1.2209232,1.9331284,2.8914874,2.5435898,1.2307693,1.1716924,2.1956925,2.2482052,1.6475899,1.148718,1.9331284,1.8116925,1.7591796,2.4385643,3.1967182,2.0939488,0.56451285,0.36102566,0.9189744,1.5392822,1.3817437,1.0469744,0.7975385,0.6498462,0.48574364,0.029538464,0.02297436,0.072205134,0.118153855,0.13784617,0.12471796,0.24615386,0.38728207,0.508718,0.60061544,0.67282057,0.81066674,0.8566154,0.8369231,0.79425645,0.8041026,0.7384616,0.6071795,0.46933338,0.3511795,0.22646156,0.13128206,0.09189744,0.09189744,0.13784617,0.25928208,0.4201026,0.92553854,1.5753847,1.9922053,1.591795,1.7066668,1.8642052,2.612513,3.3805132,2.4648206,1.6246156,1.4080001,1.3193847,1.1782565,1.1552821,1.3751796,1.5983591,1.7558975,1.9495386,2.4320002,2.9111798,2.7733335,2.6256413,2.5731285,2.2055387,2.2153847,2.3401027,2.2514873,2.4615386,4.3290257,5.3169236,5.146257,4.6276927,4.2436924,4.161641,5.654975,5.796103,5.5269747,5.47118,5.937231,3.6627696,3.2131286,3.8596926,5.0018463,6.1341543,6.3212314,6.058667,6.11118,6.6592827,7.2927184,7.8080006,8.576,9.199591,9.504821,9.531077,9.088,9.061745,9.232411,9.435898,9.577026,10.761847,10.998155,10.765129,10.469745,10.433641,9.212719,9.642668,9.396514,8.041026,7.0334363,8.254359,8.192,6.9087186,5.080616,3.9975388,3.7448208,4.0434875,5.5302567,7.7948723,9.366975,8.4512825,8.169026,8.546462,9.078155,8.713847,9.964309,10.066052,10.466462,11.234463,11.063796,10.443488,9.291488,8.214975,7.2237954,5.72718,4.5554876,4.4307694,4.6966157,4.906667,4.844308,4.31918,4.6966157,4.630975,4.0533338,4.1550775,4.2601027,4.1714873,3.9712822,3.7973337,3.8531284,3.6627696,3.4560003,2.9702566,2.5206156,3.0227695,3.9712822,4.5128207,5.2053337,6.0061545,6.2687182,3.8596926,2.7864618,2.8225644,3.5610259,4.381539,4.2305646,5.0543594,5.664821,5.8486156,6.3474874,5.9634876,5.5007186,5.2709746,5.737026,7.512616,6.311385,5.024821,5.077334,6.5706673,8.2904625,8.756514,7.8145647,6.875898,6.7774363,7.79159,7.0465646,5.756718,4.460308,3.4789746,2.934154,3.3050258,4.5029745,5.865026,6.672411,6.1440005,6.62318,7.069539,7.6570263,9.199591,13.157744,14.378668,10.794667,6.3868723,4.020513,5.4449234,5.5105643,5.333334,8.277334,13.991385,18.438566,19.423182,21.30708,22.705233,23.266464,23.683285,24.503798,20.778667,16.827078,15.82277,19.797335,24.937027,25.403078,23.22708,20.79836,20.864002,16.439796,10.8307705,6.705231,5.2348723,6.1013336,6.997334,6.9809237,6.928411,7.076103,7.02359,5.7665644,6.363898,7.020308,6.616616,4.713026,3.3444104,3.757949,3.6758976,2.9407182,3.5249233,3.387077,2.5993848,1.8412309,1.3718976,1.024,2.0775387,2.5895386,2.7503593,2.9078977,3.570872,4.5062566,5.917539,6.340924,5.7829747,5.717334,4.1878977,2.6880002,1.7394873,1.4834872,1.7001027,2.0742567,2.0250258,1.4178462,0.71548724,0.9714873,1.7952822,1.4900514,1.4539489,1.8543591,1.6311796,1.4539489,1.6508719,1.9298463,2.1989746,2.553436,3.5314875,3.0818465,3.826872,6.0324106,7.5946674,6.698667,6.747898,6.8430777,6.416411,5.2315903,7.75877,8.2904625,7.282872,5.3136415,3.0916924,1.3686155,4.7556925,9.078155,10.9686165,7.890052,6.0291286,4.5062566,4.969026,7.4436927,10.325335,8.562873,8.438154,7.397744,5.3103595,4.460308,5.3891287,5.3234878,4.5817437,3.5216413,2.5107694,1.7624617,1.8281027,1.7887181,1.5031796,1.6114873,1.3029745,1.5163078,1.6049232,1.3357949,0.88287187,0.7778462,0.9124103,1.3193847,1.8379488,2.1300514,1.5819489,1.1257436,0.86646163,0.86317956,1.1585642,1.7296412,2.4484105,2.9965131,3.3805132,3.9417439,5.172513,5.2512827,4.342154,2.8553848,1.4539489,0.8730257,0.5481026,0.38400003,0.35446155,0.49887183,0.23302566,0.2231795,0.17066668,0.026256412,0.0,0.0,0.0,0.0,0.0,0.006564103,0.013128206,0.20020515,0.27897438,0.17066668,0.0,0.0,0.0,0.006564103,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.052512825,0.06564103,0.03938462,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.009846155,0.006564103,0.013128206,0.049230773,0.16410258,0.636718,1.332513,1.9200002,1.8838975,1.7493335,2.2383592,2.4582565,2.2350771,2.1267693,2.8717952,3.442872,3.5938463,3.2689233,2.6256413,3.0982566,3.5413337,4.1550775,4.5128207,3.5872824,6.7610264,7.683283,7.322257,6.8496413,7.634052,5.98318,5.32677,6.5280004,8.129642,6.3507695,4.2174363,2.7109745,1.5097437,0.5546667,0.068923086,0.013128206,0.0,0.0,0.0,0.0,0.0,0.006564103,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.006564103,0.01969231,0.032820515,0.04594872,0.052512825,0.06235898,0.06235898,0.06564103,0.068923086,0.068923086,0.068923086,0.059076928,0.055794876,0.055794876,0.059076928,0.055794876,0.055794876,0.068923086,0.07548718,0.07548718,0.07876924,0.07548718,0.08533334,0.108307704,0.13784617,0.18379489,0.190359,0.19692309,0.19692309,0.20020515,0.20676924,0.190359,0.19364104,0.21333335,0.24615386,0.28225642,0.30194873,0.318359,0.36102566,0.4397949,0.54482055,0.702359,0.86317956,1.0338463,1.2077949,1.3554872,1.4736412,1.5885129,1.6836925,1.7296412,1.6836925,1.6738462,1.8116925,2.1103592,2.6223593,3.4264617,5.3037953,7.181129,8.172308,8.103385,7.525744,6.918565,6.62318,7.1614366,8.474257,9.921641,9.458873,9.547488,9.67877,9.101129,6.806975,4.519385,2.8127182,1.8838975,1.8346668,2.6354873,3.4527183,3.6069746,3.5446157,3.9844105,5.910975,7.643898,8.1755905,8.178872,7.640616,5.861744,5.930667,6.8693337,8.339693,10.210463,12.570257,17.302977,26.368002,35.186874,42.12513,48.512005,53.96349,57.95775,58.223595,54.419697,48.118156,41.127388,40.178875,43.585644,50.166157,59.234467,71.36165,82.65847,92.196106,99.99098,107.01129,108.96739,104.618675,98.38606,91.68411,82.93416,76.977234,68.978874,61.282467,54.803696,49.030567,43.43467,36.516106,29.705849,24.182156,20.857437,17.686975,14.404924,11.346052,8.740103,6.7150774,5.2676926,4.2469745,3.495385,2.868513,2.2482052,1.719795,1.3128207,0.9878975,0.69907695,0.41682056,0.25271797,0.14769232,0.07548718,0.02297436,0.0,0.01969231,0.029538464,0.02297436,0.009846155,0.009846155,0.04594872,0.07548718,0.08205129,0.11158975,0.28225642,0.37743592,0.8205129,1.9593848,4.240411,8.231385,9.96759,9.481847,9.42277,10.509129,11.556104,9.714872,10.039796,11.565949,13.088821,13.161027,11.67754,11.959796,17.522873,22.147284,9.882257,4.525949,2.2744617,3.1507695,5.7534366,7.253334,3.3444104,1.910154,1.0962052,0.27569234,0.06564103,0.01969231,0.006564103,0.0032820515,0.0,0.006564103,0.0,0.0,0.0032820515,0.0032820515,0.0,1.4145643,0.702359,0.508718,0.41025645,0.22646156,0.01969231,0.41682056,0.8172308,0.7581539,0.4201026,0.64000005,1.4834872,1.9396925,1.394872,0.508718,1.2340513,2.1300514,0.9419488,0.04266667,0.446359,1.7952822,2.0151796,1.5425643,0.761436,0.12143591,0.11158975,0.46933338,0.45292312,0.35446155,0.2855385,0.18379489,1.0994873,2.0742567,2.3302567,2.0644104,2.428718,2.9833848,3.131077,2.605949,1.9265642,2.4057438,2.294154,2.3040001,2.878359,3.2262566,1.3193847,0.4397949,0.30194873,0.6235898,0.9944616,0.8763078,0.5481026,0.318359,0.25271797,0.256,0.06564103,0.068923086,0.08533334,0.09189744,0.08861539,0.108307704,0.190359,0.3511795,0.47261542,0.5021539,0.4660513,0.47261542,1.7099489,1.7427694,0.58092314,0.67282057,0.63343596,0.49230772,0.35446155,0.25271797,0.15753847,0.07876924,0.03938462,0.029538464,0.055794876,0.118153855,0.20676924,0.8172308,1.8642052,2.8258464,2.7470772,2.1825643,1.972513,2.8389745,3.8334363,2.3630772,1.6869745,1.5163078,1.4703591,1.4211283,1.5097437,1.7657437,2.03159,2.225231,2.484513,3.1638978,3.383795,2.9243078,2.5600002,2.4976413,2.3663592,2.2219489,1.9659488,1.7690258,1.8773335,2.6190772,3.1245131,3.2295387,3.2754874,3.3575387,3.3280003,4.4077954,4.2436924,3.7349746,3.495385,3.8400004,2.809436,3.0194874,3.7710772,4.716308,5.858462,4.919795,4.6112823,4.9427695,5.61559,6.0291286,6.1341543,7.017026,7.8670774,8.457847,9.140513,10.069334,10.512411,10.374565,10.010257,10.197334,11.953232,12.599796,12.5374365,12.20595,12.100924,11.162257,10.725744,10.033232,8.674462,6.5837955,7.748924,8.034462,7.397744,6.235898,5.3825645,5.5171285,5.297231,6.0258465,8.0377445,10.7158985,10.601027,10.541949,10.666668,10.673231,9.82318,9.344001,9.435898,10.345026,11.690667,12.445539,11.569232,10.65354,9.921641,9.081436,7.322257,5.5762057,5.2348723,5.2578464,5.2512827,5.47118,5.0182567,4.8049235,4.585026,4.352,4.348718,3.9351797,4.0467696,4.381539,4.667077,4.6539493,3.5807183,2.8455386,2.4155898,2.3991797,3.0227695,3.754667,4.493129,5.481026,6.1407185,5.0674877,3.1803079,2.4713848,2.7831798,3.6758976,4.4077954,4.089436,4.824616,5.5236926,5.901129,6.4689236,6.4590774,5.668103,5.549949,6.5411286,8.080411,5.3234878,3.9680004,5.024821,8.01477,10.939077,9.685334,7.387898,6.091488,6.370462,7.3091288,5.435077,4.1517954,4.06318,4.6276927,4.1517954,4.2436924,5.8157954,7.1548724,7.4896417,7.0104623,6.7938466,6.9809237,7.4830775,8.809027,12.041847,13.259488,9.7673855,5.7107697,3.8596926,5.609026,6.363898,5.3760004,6.5969234,10.47959,13.978257,14.614976,15.750566,16.282257,15.563488,13.397334,15.281232,14.473847,13.643488,15.563488,23.115488,25.862566,24.109951,20.611284,18.176,19.656206,15.553642,11.273847,8.2215395,7.3485136,9.15036,9.409642,8.635077,7.936001,7.6668725,7.4174366,7.194257,8.205129,8.352821,7.0367184,5.1331286,4.132103,4.5817437,4.5456414,3.8038976,3.8596926,3.820308,2.8521028,2.3729234,2.4582565,1.8379488,2.793026,3.8137438,4.2994876,4.240411,4.2371287,4.673641,6.0356927,6.4065647,5.5958977,5.152821,3.8498464,2.3269746,1.5491283,1.5655385,1.5097437,2.2416413,2.3138463,1.7723079,1.142154,1.4473847,2.5238976,2.03159,1.4080001,1.1782565,0.9353847,1.5064616,1.910154,2.4057438,3.0785644,3.8596926,3.2787695,2.6322052,3.190154,4.562052,4.667077,4.4898467,5.277539,5.6418467,5.3005133,5.0642056,5.943795,5.481026,4.644103,3.817026,2.8160002,2.041436,7.1581545,13.715693,17.017437,12.100924,6.422975,4.0500517,4.906667,7.322257,8.03118,5.146257,6.1997952,7.27959,6.5772314,4.4012313,5.533539,4.906667,3.4297438,2.034872,1.6804104,2.2350771,2.861949,2.7306669,1.9856411,1.7460514,1.2570257,1.2340513,1.1388719,0.8598975,0.7056411,0.6301539,0.65969235,1.0043077,1.5753847,1.9954873,1.1158975,0.5907693,0.42994875,0.5546667,0.81066674,1.1224617,1.5721027,2.034872,2.6157951,3.6496413,4.4767184,4.716308,4.3290257,3.4592824,2.4352822,1.4769232,0.94523084,0.67938465,0.56451285,0.50543594,0.22646156,0.21661541,0.16410258,0.02297436,0.0,0.0,0.0,0.0,0.0,0.0,0.032820515,0.31507695,0.40697438,0.21333335,0.0,0.0,0.0,0.009846155,0.01969231,0.0,0.0,0.0,0.0,0.0,0.006564103,0.06564103,0.08861539,0.055794876,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.01969231,0.029538464,0.13456412,0.42994875,0.86974365,1.2406155,1.5195899,1.9200002,2.172718,2.356513,2.9078977,3.4231799,3.5577438,3.7120004,3.764513,3.0752823,3.7940516,5.1659493,5.723898,5.2480006,4.788513,5.668103,6.0685134,5.8125134,5.4875903,6.436103,4.6211286,4.06318,3.9220517,3.698872,3.239385,3.1507695,2.044718,0.94523084,0.30851284,0.026256412,0.006564103,0.0,0.0,0.0,0.0,0.0,0.006564103,0.006564103,0.006564103,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.02297436,0.036102567,0.04266667,0.055794876,0.059076928,0.06564103,0.068923086,0.072205134,0.07548718,0.068923086,0.06235898,0.059076928,0.055794876,0.06235898,0.06564103,0.08205129,0.0951795,0.098461546,0.10502565,0.10502565,0.108307704,0.13128206,0.17066668,0.21333335,0.2297436,0.24615386,0.256,0.25928208,0.26256412,0.23630771,0.2231795,0.22646156,0.25271797,0.29538465,0.33476925,0.380718,0.41025645,0.4266667,0.45620516,0.5481026,0.6892308,0.85005134,1.0108719,1.142154,1.2209232,1.3161026,1.4309745,1.5392822,1.591795,1.6705642,1.785436,1.910154,2.1202054,2.5895386,3.6660516,4.604718,5.421949,6.1308722,6.7249236,7.128616,6.6822567,6.514872,7.026872,7.9195905,7.90318,8.953437,10.049642,10.187488,8.385642,6.0652313,4.5522056,3.4888208,2.7602053,2.477949,3.058872,3.6463592,3.6824617,3.18359,2.7306669,2.8324106,3.2098465,3.6562054,3.826872,3.2328207,3.4067695,4.4307694,5.431795,5.8781543,5.546667,7.9294367,12.71795,17.506462,21.950361,27.785849,34.727386,40.89108,45.42031,47.310772,45.41703,38.583797,37.270977,39.076107,42.499287,46.923492,53.983185,61.328415,67.534775,74.249855,86.19324,97.51303,104.34627,105.104416,100.8837,95.465034,87.52575,80.20021,72.766365,65.50975,59.72021,54.39672,47.799797,40.42503,33.329235,28.114054,24.923899,21.786259,18.770052,15.904821,13.174155,10.843898,8.966565,7.4207187,6.088206,4.84759,3.7710772,2.9046156,2.2022567,1.6114873,1.0601027,0.6695385,0.41025645,0.23630771,0.118153855,0.049230773,0.029538464,0.029538464,0.032820515,0.03938462,0.06564103,0.17723078,0.25271797,0.2231795,0.12143591,0.052512825,0.072205134,0.2297436,0.86317956,2.2514873,4.637539,6.744616,7.312411,8.6580515,11.720206,16.055796,15.199181,14.424617,14.204719,14.516514,14.834873,12.35036,10.06277,12.422565,15.921232,9.088,3.114667,1.0043077,2.4549747,5.549949,6.747898,3.7021542,2.3827693,1.3817437,0.36758977,0.072205134,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.65312827,0.6268718,0.8467693,0.8402052,0.508718,0.17066668,0.2231795,0.43323082,0.3446154,0.009846155,0.006564103,1.3554872,1.4998976,0.9944616,0.58420515,1.2242053,3.2000003,1.4867693,0.009846155,0.21989745,1.0994873,2.8455386,2.678154,1.4506668,0.22646156,0.25928208,0.21661541,0.2297436,0.34133336,0.4955898,0.508718,1.7033848,1.3292309,1.2274873,1.9265642,2.6551797,1.7723079,2.1858463,2.5829747,2.4549747,2.0873847,2.0873847,2.1136413,1.5491283,0.574359,0.14769232,0.10502565,0.190359,0.20348719,0.14112821,0.20348719,0.23630771,0.23958977,0.18379489,0.1148718,0.15097436,0.17394873,0.17723078,0.17066668,0.16082053,0.16410258,0.20676924,0.2855385,0.3314872,0.3314872,0.32164106,0.3052308,2.9604106,3.0227695,0.47589746,0.54482055,0.49230772,0.37743592,0.256,0.15097436,0.068923086,0.03938462,0.02297436,0.029538464,0.059076928,0.12143591,0.13456412,0.4201026,1.3259488,2.678154,3.7940516,2.6683078,2.3762052,2.4681027,2.4385643,1.7329233,1.8740515,1.8970258,1.8116925,1.6968206,1.6771283,2.1398976,2.5304618,2.8914874,3.3969233,4.3585644,3.2951798,2.5928206,2.477949,2.7273848,2.674872,2.4681027,2.428718,2.425436,2.3335385,2.038154,2.0184617,2.1136413,2.4713848,2.9801028,3.2754874,3.764513,3.370667,2.7634873,2.3105643,2.0709746,2.605949,3.006359,3.5807183,4.197744,4.2863593,3.692308,3.2918978,3.4297438,3.9647183,4.279795,4.128821,4.8738465,5.677949,6.4590774,7.88677,9.757539,9.964309,9.435898,9.097847,9.852718,11.943385,13.092104,13.653335,13.843694,13.74195,13.216822,12.091078,11.221334,10.226872,7.4830775,7.6668725,6.931693,6.422975,6.5280004,6.87918,7.830975,7.9195905,8.073847,8.963283,10.988309,11.776001,13.075693,13.561437,12.977232,12.137027,9.143796,7.9786673,8.694155,10.266257,10.604308,10.630565,10.387693,9.793642,8.969847,8.2445135,7.030154,5.9930263,5.0018463,4.3585644,4.8049235,5.0543594,4.7983594,4.9788723,5.4514875,4.9854364,3.8596926,3.5774362,3.945026,4.588308,4.919795,3.879385,3.0916924,2.8127182,3.0030773,3.318154,3.2754874,3.7284105,4.6966157,5.169231,3.0982566,3.2196925,3.0654361,3.4494362,4.2863593,4.59159,3.2295387,3.2886157,4.0336413,4.788513,4.919795,5.723898,5.402257,5.5663595,6.547693,7.4108725,5.3136415,4.2469745,4.9329233,7.0367184,9.176616,6.3343596,4.46359,4.562052,6.245744,7.755488,5.7140517,4.6966157,5.346462,6.774154,6.5870776,5.664821,6.3442054,6.665847,6.3474874,6.7872825,6.038975,5.1298466,4.6802053,4.772103,4.962462,5.2742567,4.388103,3.4133337,3.1934361,4.3060517,5.1626673,4.1222568,3.5610259,4.906667,8.65477,10.440206,11.894155,12.737642,12.563693,10.834052,11.303386,11.690667,12.918155,16.308514,23.561848,23.072823,19.377232,15.258258,12.757335,13.184001,10.781539,10.9226675,10.663385,9.872411,11.237744,10.266257,8.5202055,7.059693,6.5936418,7.4863596,8.605539,8.598975,7.6274877,6.294975,5.661539,5.4547696,6.180103,6.370462,5.546667,4.210872,4.1846156,3.3903592,3.5577438,4.3027697,3.1113849,4.20759,5.284103,5.668103,5.221744,4.345436,4.9362054,6.160411,6.058667,4.44718,2.9046156,2.7602053,2.4943593,2.4418464,2.3630772,1.4441026,1.5622566,1.7690258,1.7296412,1.6147693,2.1103592,3.3805132,3.114667,2.0644104,1.0568206,0.97805136,2.3105643,3.2164104,3.820308,4.1189747,3.9909747,2.7536411,1.8313848,1.4408206,1.6311796,2.2711797,3.2623591,4.1878977,5.175795,6.038975,6.2884107,5.211898,5.5762057,6.6133337,7.026872,4.97559,3.564308,6.4295387,11.703795,15.563488,12.209231,5.658257,3.1507695,3.9253337,5.664821,4.493129,3.764513,5.976616,8.274052,8.3364105,4.3749747,5.353026,3.9548721,2.3269746,1.7460514,2.605949,3.876103,4.4734364,4.06318,2.878359,1.7296412,1.1323078,1.0896411,0.98133343,0.6465641,0.39384618,0.39384618,0.65312827,1.1224617,1.6738462,2.100513,1.0535386,0.41682056,0.17723078,0.22646156,0.35446155,0.61374366,0.73517954,0.9911796,1.6738462,3.0523078,3.0851285,3.2131286,3.1245131,2.789744,2.4681027,1.5885129,0.99774367,0.69579494,0.49230772,0.02297436,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.029538464,0.06564103,0.0951795,0.40697438,0.49887183,0.26256412,0.0,0.0,0.0,0.0032820515,0.009846155,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.032820515,0.052512825,0.036102567,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.026256412,0.055794876,0.17066668,0.49887183,1.3292309,1.5458462,1.8248206,2.481231,3.4560003,3.05559,2.917744,3.1803079,3.3542566,2.3236926,3.446154,5.648411,6.0652313,5.2611284,7.213949,5.87159,5.218462,5.228308,5.464616,5.0543594,4.4767184,3.9122055,3.255795,2.6715899,2.609231,2.041436,1.5753847,1.017436,0.40369233,0.009846155,0.006564103,0.0032820515,0.0,0.0,0.006564103,0.009846155,0.009846155,0.013128206,0.01969231,0.016410258,0.006564103,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.01969231,0.026256412,0.036102567,0.049230773,0.052512825,0.052512825,0.055794876,0.06564103,0.068923086,0.06235898,0.052512825,0.049230773,0.059076928,0.068923086,0.08205129,0.09189744,0.10502565,0.1148718,0.1148718,0.11158975,0.13128206,0.16410258,0.19692309,0.2297436,0.27241027,0.30194873,0.30851284,0.2986667,0.29538465,0.27897438,0.26912823,0.27897438,0.30194873,0.39712822,0.512,0.55794877,0.5349744,0.5284103,0.5284103,0.6268718,0.764718,0.88943595,0.9616411,0.95835906,0.955077,0.9878975,1.0699488,1.1815386,1.3456411,1.5130258,1.657436,1.8871796,2.4484105,3.5216413,4.4767184,5.172513,5.5696416,5.723898,7.194257,6.7577443,5.612308,4.6900516,4.670359,5.9634876,8.2904625,10.476309,11.621744,11.109744,9.373539,8.044309,6.889026,5.5565133,3.5807183,4.266667,6.170257,7.145026,6.340924,4.194462,3.498667,3.249231,3.1573336,2.986667,2.5764105,1.7952822,1.339077,1.2176411,1.401436,1.8116925,3.43959,5.4416413,6.810257,8.201847,11.9171295,16.180513,19.859694,23.61436,27.454361,30.733131,30.815182,32.52513,34.783184,36.801643,38.052105,40.44472,45.390774,50.77662,56.3758,63.86544,78.36883,94.40821,104.42175,107.46421,109.22996,100.90668,92.28801,84.496414,77.827286,71.71611,67.14421,62.546055,55.972107,47.405952,38.757748,33.942978,30.198156,27.168823,24.405334,21.349745,18.409027,15.734155,13.302155,11.08677,9.03877,7.200821,5.6287184,4.33559,3.2820516,2.3696413,1.5885129,1.0075898,0.6071795,0.3511795,0.18379489,0.08205129,0.049230773,0.049230773,0.07876924,0.15425642,0.36430773,0.4660513,0.4397949,0.3117949,0.14441027,0.09189744,0.068923086,0.14441027,0.38400003,0.84348726,2.4418464,4.5522056,7.702975,12.419283,19.24595,19.140924,15.753847,12.337232,10.866873,12.032001,10.28595,7.4141545,5.1298466,4.210872,4.5029745,2.038154,0.93866676,1.4145643,2.6354873,2.7142565,1.847795,1.2307693,0.6892308,0.22646156,0.03938462,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,2.1070771,1.5819489,1.3128207,1.0666667,0.8041026,0.67282057,0.24287182,0.36758977,0.33476925,0.055794876,0.029538464,0.92225647,0.84348726,0.6465641,0.7122052,0.9321026,0.6498462,0.27897438,0.04594872,0.0,0.0,0.4397949,0.5218462,0.4660513,0.5284103,0.9911796,0.7220513,0.77456415,1.4966155,2.4024618,2.1825643,1.6082052,1.1093334,0.7417436,0.58092314,0.702359,0.4955898,1.4769232,2.9735386,4.027077,3.4166157,2.540308,1.2012309,0.29210258,0.072205134,0.18379489,0.12143591,0.48246157,0.51856416,0.20348719,0.2297436,0.58420515,0.71548724,0.5349744,0.22646156,0.27569234,0.2855385,0.28225642,0.29210258,0.2986667,0.21333335,0.17723078,0.15097436,0.13784617,0.13784617,0.13784617,0.45620516,1.6246156,1.5983591,0.45620516,0.39712822,0.43323082,0.37743592,0.24943592,0.108307704,0.04594872,0.032820515,0.029538464,0.055794876,0.12143591,0.24287182,0.15753847,0.45620516,1.2438976,2.4024618,3.5872824,2.2055387,1.9987694,2.0906668,2.2350771,2.806154,2.8816411,2.6157951,2.2678976,1.9462565,1.6180514,2.8488207,3.5511796,4.279795,5.139693,5.799385,2.8324106,2.0250258,2.4484105,3.2262566,3.5544617,3.639795,4.020513,4.4898467,4.772103,4.516103,3.5413337,2.8488207,3.0720003,4.0303593,4.716308,4.923077,4.4438977,3.9253337,3.4888208,2.7306669,2.6715899,2.8192823,2.930872,2.8947694,2.7634873,2.3729234,2.0709746,1.8346668,1.8018463,2.28759,2.6190772,3.5347695,4.4800005,5.431795,6.8955903,7.177847,6.810257,6.294975,6.058667,6.422975,7.6931286,8.825437,9.728001,10.33518,10.604308,11.641437,10.985026,10.30236,10.108719,9.764103,9.130668,7.9195905,6.9054365,6.3901544,6.196513,7.3419495,8.086975,8.5202055,8.707283,8.681026,9.488411,10.925949,11.890873,12.442257,13.8075905,12.711386,9.91836,8.044309,7.6274877,7.125334,6.8562055,7.1187696,7.328821,7.3780518,7.6603084,6.6592827,5.8880005,5.277539,4.962462,5.280821,5.07077,5.175795,6.3474874,7.499488,5.7074876,3.5446157,2.3269746,2.0053334,2.550154,3.9680004,3.5511796,2.9636924,2.5961027,2.5600002,2.6715899,2.806154,3.1770258,3.4592824,3.5610259,3.6463592,2.8914874,3.1409233,3.1277952,2.7864618,3.249231,2.3958976,1.6508719,1.2800001,1.3686155,1.8313848,4.2863593,6.0225644,6.1341543,5.1265645,4.9427695,5.687795,5.6287184,5.2414365,4.31918,1.9396925,1.585231,2.3663592,4.348718,6.889026,8.621949,6.813539,6.0685134,6.422975,7.062975,6.3179493,4.1091285,2.9407182,2.0808206,1.4178462,1.463795,2.5042052,2.4976413,2.8553848,4.240411,6.560821,7.39118,6.7282057,5.3202057,4.0369234,3.892513,4.5128207,4.073026,3.7743592,5.113436,9.888822,10.607591,11.940104,13.108514,12.872206,9.55077,7.062975,6.4295387,7.3353853,9.281642,11.611898,12.33395,11.680821,10.269539,8.690872,7.509334,9.363693,10.138257,9.984001,9.074872,7.5979495,7.1844106,7.5552826,8.044309,8.707283,10.328616,10.453334,9.055181,7.565129,6.550975,5.720616,5.917539,7.1647186,7.456821,6.042257,3.4166157,2.6486156,3.501949,5.149539,6.091488,4.1517954,4.2601027,3.8564105,3.5282054,3.515077,3.7218463,4.2830772,4.7917953,4.7983594,3.9909747,2.1956925,1.9528207,2.5042052,2.7076926,2.041436,0.6268718,0.636718,1.0535386,1.4145643,1.5458462,1.5721027,2.1202054,3.95159,4.420923,3.245949,2.5009232,2.7208207,3.3444104,3.7218463,3.186872,1.0371283,0.512,0.4266667,0.7515898,1.8543591,4.516103,6.1046157,6.8562055,7.3025646,7.450257,6.7905645,5.605744,6.160411,7.8637953,8.845129,5.9503593,2.6190772,3.5052311,5.4186673,5.83877,2.9472823,1.5425643,1.4834872,2.9833848,5.333334,6.8955903,6.675693,6.941539,6.173539,4.535795,3.876103,2.556718,1.6344616,1.3161026,1.910154,3.8137438,4.841026,5.142975,4.768821,3.69559,1.8149745,1.0699488,0.54482055,0.23958977,0.12471796,0.13784617,0.23630771,0.8992821,1.4933335,1.7690258,1.8937438,1.2931283,0.48574364,0.026256412,0.013128206,0.06235898,0.24287182,0.33476925,0.48246157,0.7450257,1.0994873,1.270154,1.467077,1.5524104,1.4572309,1.1749744,0.9321026,0.47589746,0.128,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.036102567,0.14112821,0.33476925,0.22646156,0.22646156,0.17066668,0.049230773,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.02297436,0.04594872,0.3511795,0.6465641,1.3128207,2.3302567,3.2951798,1.9396925,2.0676925,2.5009232,2.4943593,1.723077,1.6278975,2.4549747,3.7907696,5.346462,6.957949,5.2742567,3.882667,3.6496413,4.2962055,4.394667,3.0162053,2.0841026,1.4572309,1.1684103,1.4506668,1.2537436,0.7844103,0.30851284,0.02297436,0.04594872,0.032820515,0.013128206,0.0,0.006564103,0.029538464,0.055794876,0.04266667,0.036102567,0.03938462,0.016410258,0.026256412,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.009846155,0.0,0.0,0.013128206,0.016410258,0.02297436,0.029538464,0.029538464,0.04266667,0.04594872,0.04594872,0.04594872,0.04594872,0.059076928,0.068923086,0.07548718,0.07876924,0.09189744,0.07876924,0.07548718,0.08861539,0.11158975,0.13784617,0.19692309,0.27897438,0.3249231,0.33476925,0.33476925,0.3708718,0.3708718,0.34789747,0.31507695,0.28882053,0.37415388,0.48902568,0.574359,0.636718,0.74830776,0.5513847,0.5940513,0.7220513,0.8402052,0.8992821,0.98461545,0.99774367,0.9682052,0.9353847,0.9616411,1.0108719,1.1323078,1.339077,1.6672822,2.166154,2.412308,3.4527183,4.6112823,5.0674877,3.8465643,3.8695388,3.5544617,3.2918978,3.3641028,3.9384618,5.2315903,6.7807183,8.208411,9.508103,11.047385,12.232206,12.087796,12.074668,11.625027,8.132924,9.281642,13.5318985,16.357744,15.645539,11.703795,8.94359,7.522462,5.8880005,3.7842054,2.2580514,1.4408206,0.90584624,0.5940513,0.446359,0.39712822,1.1060513,2.409026,3.5478978,4.70318,6.9743595,9.196308,9.888822,10.473026,11.493745,12.6063595,15.560206,20.38154,25.898668,30.86113,33.94954,37.51713,41.987286,45.764927,48.76472,52.414364,62.47385,76.38647,91.90073,107.1918,120.86483,119.972115,114.254776,105.21601,93.81088,80.443085,76.672005,76.186264,73.54749,67.26237,59.76616,49.207798,40.854977,35.721848,33.06995,30.395079,27.122873,23.952412,20.883694,17.926565,15.107284,12.504617,10.023385,7.857231,6.0783596,4.637539,3.3312824,2.2383592,1.3817437,0.7811283,0.4266667,0.26912823,0.14769232,0.07876924,0.0951795,0.2297436,0.49887183,0.58420515,0.57764107,0.49887183,0.28882053,0.13128206,0.04594872,0.032820515,0.098461546,0.24287182,3.0654361,6.688821,10.71918,14.483693,17.060104,17.316103,12.517745,7.2336416,4.388103,5.280821,6.0356927,4.8147697,3.0096412,1.6804104,1.5721027,2.097231,1.9331284,1.5622566,1.2242053,0.9321026,0.4660513,0.21333335,0.108307704,0.07548718,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.92225647,0.54482055,0.7811283,0.761436,0.45620516,0.6826667,0.27569234,0.5481026,0.4955898,0.0951795,0.3249231,0.7056411,0.45620516,0.256,0.4660513,1.1126155,0.6662565,0.3052308,0.35446155,0.65312827,0.53825647,0.19692309,0.24943592,0.34133336,0.508718,1.1881026,0.6826667,1.1454359,1.8215386,2.0873847,1.4375386,1.3522053,1.4703591,1.6278975,2.0217438,3.2295387,3.3050258,2.3958976,2.0217438,2.3433847,2.172718,0.90256417,0.53825647,0.7089231,0.9321026,0.6235898,0.72861546,0.77128214,0.5481026,0.20348719,0.2297436,0.50543594,0.62030774,0.6071795,0.51856416,0.4201026,0.2855385,0.24287182,0.24615386,0.23958977,0.16410258,0.118153855,0.06564103,0.036102567,0.032820515,0.052512825,0.18379489,0.49230772,0.5316923,0.3052308,0.27569234,0.5152821,0.46276927,0.29538465,0.18379489,0.27897438,0.5677949,0.3052308,0.08861539,0.13456412,0.256,0.42338464,0.81066674,1.9429746,3.4855387,4.2207184,2.937436,2.5665643,2.5796926,2.6322052,2.550154,2.294154,2.4352822,2.28759,2.1202054,3.1671798,6.265436,5.8814363,5.5958977,6.560821,7.496206,4.020513,3.4691284,3.7940516,3.7874875,3.0916924,2.5993848,2.2482052,1.9331284,1.6344616,1.4276924,1.3095386,1.1848207,1.4112822,2.0086155,2.665026,3.2131286,4.013949,4.97559,5.543385,4.709744,3.7185643,3.2918978,3.1737437,3.0030773,2.3236926,1.7165129,1.3423591,1.1388719,1.148718,1.5195899,1.8871796,2.5074873,3.2656412,4.132103,5.1265645,5.0477953,4.713026,4.384821,4.2207184,4.263385,4.525949,5.106872,5.4843082,5.4974365,5.356308,5.504,5.586052,6.235898,6.9842057,6.2490263,6.3474874,5.927385,5.6451287,5.85518,6.5969234,6.816821,6.9645133,6.8693337,6.6527185,6.705231,7.069539,7.565129,7.4108725,6.957949,7.680001,7.3550773,6.9152827,6.885744,7.076103,6.564103,6.052103,6.114462,6.363898,6.4557953,6.0717955,5.287385,4.7360005,5.1331286,6.048821,5.927385,5.5236926,5.175795,6.157129,7.50277,5.9995904,4.3552823,3.1442053,2.556718,2.6190772,3.186872,2.4976413,2.2514873,2.3958976,2.9111798,3.7809234,3.5544617,3.639795,3.8498464,4.1222568,4.4996924,3.4724104,3.2656412,3.3411283,3.620103,4.4964104,3.5249233,2.2153847,1.3686155,1.2373334,1.5261539,2.4352822,4.2305646,5.077334,4.4800005,3.2722054,3.751385,5.21518,5.835488,5.2447186,4.525949,3.751385,2.5665643,2.1136413,2.6880002,3.7251284,4.020513,4.1156926,4.240411,4.2207184,3.4855387,3.754667,4.2207184,4.3749747,4.31918,4.7491283,6.1374364,7.062975,7.427283,7.6701546,8.759795,10.456616,9.777231,7.9294367,5.914257,4.5390773,3.5872824,2.865231,3.2295387,5.5105643,10.499283,10.253129,9.02236,7.463385,5.940513,4.535795,4.007385,4.578462,5.2414365,6.0225644,7.962257,10.322052,9.334154,7.204103,5.4482055,4.857436,5.72718,6.117744,6.2194877,6.265436,6.5378466,7.3321033,7.325539,7.5913854,8.651488,10.502565,11.736616,10.564924,9.248821,8.726975,8.63836,8.28718,8.579283,8.267488,6.928411,4.969026,3.9548721,3.7120004,4.017231,4.6867695,5.579488,4.84759,4.2371287,4.535795,5.290667,4.785231,3.636513,3.2689233,3.2525132,3.0030773,1.7952822,1.2570257,1.7066668,1.7558975,1.0601027,0.30851284,0.39712822,0.58420515,0.7384616,0.81066674,0.81394875,1.079795,1.6246156,1.5130258,0.83035904,0.67282057,0.95835906,1.4441026,1.6771283,1.591795,1.5130258,1.5261539,1.6246156,3.2295387,6.1505647,8.618668,10.919386,11.411694,10.883283,9.511385,6.8496413,5.5893335,5.3924108,5.477744,5.024821,3.1540515,2.3335385,2.6486156,2.9604106,2.7175386,1.9429746,1.654154,2.2908719,3.8695388,5.58277,5.799385,5.8912826,5.2611284,4.266667,3.3542566,3.045744,2.487795,2.1136413,2.3335385,3.2000003,4.4012313,4.352,3.3903592,2.4549747,1.7985642,0.9747693,0.45292312,0.26256412,0.16738462,0.09189744,0.11158975,0.7089231,1.5425643,1.9922053,1.975795,1.9396925,1.3817437,0.5907693,0.09189744,0.0032820515,0.02297436,0.08205129,0.118153855,0.18707694,0.29210258,0.39056414,0.48246157,0.7581539,1.0765129,1.2373334,0.955077,0.4660513,0.16410258,0.026256412,0.0,0.0,0.03938462,0.026256412,0.006564103,0.0032820515,0.013128206,0.013128206,0.04266667,0.18707694,0.380718,0.41025645,0.2100513,0.0951795,0.032820515,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.068923086,0.13784617,0.36102566,0.8566154,1.6836925,1.6377437,1.5819489,1.529436,1.4933335,1.467077,0.77456415,1.0043077,1.8248206,3.0490258,4.650667,3.9909747,3.0162053,3.255795,4.4438977,4.5423594,3.9909747,2.9604106,1.9035898,1.1848207,1.083077,1.2209232,0.61374366,0.14112821,0.118153855,0.28882053,0.318359,0.2100513,0.0951795,0.055794876,0.128,0.0951795,0.07548718,0.072205134,0.08205129,0.07548718,0.029538464,0.052512825,0.068923086,0.049230773,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0,0.013128206,0.016410258,0.016410258,0.02297436,0.04266667,0.026256412,0.029538464,0.032820515,0.036102567,0.04594872,0.059076928,0.06235898,0.06564103,0.06564103,0.07876924,0.07548718,0.07548718,0.08861539,0.11158975,0.13784617,0.19692309,0.2855385,0.33476925,0.34789747,0.39712822,0.45292312,0.44964105,0.43651286,0.4266667,0.4135385,0.4004103,0.4135385,0.446359,0.47917953,0.49230772,0.46276927,0.4955898,0.56451285,0.6498462,0.7417436,0.86646163,0.9747693,1.0633847,1.1126155,1.1093334,1.0601027,1.0896411,1.2406155,1.5064616,1.847795,2.2219489,3.4691284,5.1200004,6.2129235,5.284103,3.892513,3.620103,3.6332312,3.6430771,3.9253337,4.818052,5.35959,5.930667,6.8332314,8.3134365,10.620719,11.247591,10.929232,9.7673855,7.253334,7.6307697,9.521232,11.149129,11.746463,11.546257,12.163283,11.625027,9.504821,6.2588725,3.1967182,2.048,1.0732309,0.46276927,0.21989745,0.14112821,0.28225642,0.60061544,1.0108719,1.5688206,2.481231,3.501949,4.4800005,5.661539,7.0498466,8.4053335,10.666668,14.375385,19.669334,25.961027,31.947489,37.31036,42.72903,47.17949,50.06113,51.180313,52.480003,55.40103,62.07672,73.117546,87.59139,102.76431,116.44391,119.801445,113.32924,106.84719,98.93416,91.44452,84.42749,77.87652,71.71939,66.42216,58.033234,51.715286,47.986874,42.676517,37.48103,32.958363,28.98708,25.488413,22.406567,19.649643,16.850052,14.053744,11.369026,8.973129,6.99077,5.2742567,3.820308,2.5961027,1.5392822,0.90912825,0.53825647,0.3446154,0.27897438,0.31507695,0.47589746,0.49887183,0.42338464,0.30194873,0.19364104,0.09189744,0.059076928,0.068923086,0.14769232,0.35446155,2.6157951,6.1538467,9.616411,11.572514,10.505847,9.091283,5.917539,3.1934361,2.231795,3.4724104,4.7950773,4.2371287,2.6256413,1.0765129,0.98461545,2.1169233,2.2678976,1.6246156,0.7089231,0.35774362,0.16738462,0.068923086,0.029538464,0.016410258,0.0032820515,0.0,0.006564103,0.013128206,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.24943592,0.34133336,0.6695385,0.58092314,0.2297436,0.5677949,0.6104616,0.7778462,0.6859488,0.56451285,1.2307693,0.8205129,0.39384618,0.17066668,0.36102566,1.1782565,0.47589746,0.15753847,0.33805132,0.8533334,1.2471796,0.36102566,0.128,0.28225642,0.5874872,0.84348726,0.6235898,0.9944616,1.2603078,1.2537436,1.3259488,1.1552821,1.7099489,1.7263591,1.4539489,2.6617439,2.2153847,1.5524104,2.044718,3.1081028,2.1924105,0.6268718,1.1027694,2.048,2.2777438,0.99774367,3.3772311,3.4330258,2.0644104,0.50543594,0.30194873,0.38400003,0.41025645,0.44307697,0.47589746,0.42994875,0.3117949,0.2100513,0.16082053,0.14112821,0.098461546,0.06235898,0.026256412,0.006564103,0.013128206,0.029538464,0.101743594,0.29538465,0.4135385,0.42338464,0.47261542,0.44964105,0.3708718,0.36102566,0.56451285,1.1585642,2.103795,1.9364104,1.6311796,1.7296412,2.3269746,2.4648206,2.409026,2.9210258,3.889231,4.315898,3.5938463,2.5042052,1.9331284,2.1989746,3.045744,3.2754874,3.817026,4.3749747,4.8836927,5.5138464,6.294975,4.9099493,4.0533338,4.4406157,4.824616,3.3772311,3.31159,3.3017437,2.7437952,1.7493335,1.4145643,1.020718,0.6498462,0.41682056,0.46276927,0.6629744,0.52512825,0.512,0.7581539,1.0633847,1.3226668,2.1202054,3.6529233,5.4974365,6.6133337,5.861744,5.408821,5.100308,4.6080003,3.43959,2.6256413,2.0020514,1.4867693,1.1224617,1.0535386,1.3226668,1.6508719,2.028308,2.4484105,2.9078977,2.9210258,2.9472823,3.058872,3.2229745,3.31159,3.3378465,3.4002054,3.31159,3.0293336,2.6617439,2.7569232,2.9210258,3.4592824,4.1550775,4.2535386,4.841026,4.647385,4.585026,5.1167183,6.232616,6.3573337,6.160411,5.677949,5.1659493,5.093744,5.481026,5.4416413,5.093744,4.644103,4.391385,4.571898,5.431795,6.2194877,6.6592827,6.9349747,5.901129,5.0510774,4.6933336,4.6834874,4.414359,4.713026,4.788513,5.72718,7.1876926,7.4141545,6.774154,6.304821,7.0104623,8.083693,6.8955903,6.1374364,5.2414365,4.352,3.7776413,3.9778464,3.9844105,3.9581542,3.5905645,2.9702566,2.5764105,2.4713848,2.9702566,3.383795,3.6004105,4.073026,5.1298466,5.175795,4.7491283,4.5029745,5.1987696,4.522667,3.2722054,2.7634873,2.9735386,2.556718,2.6223593,3.4494362,4.1780515,4.1485133,2.917744,3.2295387,5.0051284,5.989744,5.8978467,6.3901544,5.2414365,3.314872,2.1956925,2.4516926,3.6562054,4.2896414,4.6867695,5.024821,5.169231,4.663795,5.208616,6.0783596,5.9536414,5.034667,5.0477953,5.7698464,6.117744,6.2720003,6.419693,6.764308,7.712821,7.4240007,6.4656415,5.156103,3.5741541,2.2908719,1.522872,1.7887181,3.442872,6.669129,6.6560006,5.674667,4.44718,3.436308,2.8225644,2.7437952,3.31159,3.7382567,4.0008206,4.8344617,6.242462,5.2348723,3.9122055,3.4560003,4.1124105,5.504,5.7698464,5.4843082,5.4613338,6.7577443,7.6143594,7.88677,8.214975,8.726975,9.032206,9.888822,9.856001,9.760821,9.852718,9.826463,9.557334,8.704,7.6767187,6.73477,5.986462,4.33559,3.2196925,3.1770258,4.06318,5.037949,3.6004105,3.3280003,4.128821,4.9296412,3.6594875,3.0523078,2.6518977,2.2711797,1.7985642,1.1913847,0.75487185,0.9714873,1.079795,0.8172308,0.42994875,0.3708718,0.46933338,0.7515898,1.1158975,1.3226668,1.2077949,1.5753847,1.4867693,0.92553854,0.79097444,0.764718,1.1191796,1.7165129,2.809436,5.028103,4.663795,3.8038976,5.0182567,8.408616,11.602052,14.381949,13.426873,10.518975,7.515898,6.3540516,5.277539,4.5095387,3.7054362,2.7602053,1.8051283,2.044718,2.546872,2.806154,2.7175386,2.5829747,2.3433847,2.3236926,2.7142565,3.3214362,3.564308,4.240411,3.5183592,2.6912823,2.428718,2.7733335,2.3204105,1.9561027,1.8773335,2.1070771,2.4976413,2.2022567,1.4703591,0.892718,0.636718,0.46933338,0.23958977,0.17723078,0.13456412,0.08861539,0.14441027,1.1552821,1.847795,2.1858463,2.3269746,2.6223593,1.5589745,0.6432821,0.13456412,0.016410258,0.016410258,0.032820515,0.1148718,0.19364104,0.22646156,0.20348719,0.2855385,0.48246157,0.64000005,0.636718,0.3708718,0.14112821,0.032820515,0.0,0.006564103,0.026256412,0.03938462,0.026256412,0.009846155,0.07548718,0.3708718,0.24615386,0.11158975,0.101743594,0.20020515,0.22646156,0.26912823,0.118153855,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.052512825,0.20348719,0.5218462,0.65641034,0.65312827,0.57764107,0.54482055,0.7187693,0.67938465,0.6629744,0.86974365,1.4473847,2.481231,2.5337439,2.0184617,1.9462565,2.5238976,3.1409233,3.5610259,3.0227695,1.8051283,0.5973334,0.52512825,0.5546667,0.2986667,0.14769232,0.21661541,0.3511795,0.45292312,0.3249231,0.30851284,0.39056414,0.190359,0.118153855,0.06564103,0.06564103,0.101743594,0.108307704,0.032820515,0.06564103,0.072205134,0.02297436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.016410258,0.016410258,0.016410258,0.01969231,0.02297436,0.029538464,0.032820515,0.03938462,0.04594872,0.049230773,0.055794876,0.055794876,0.055794876,0.06564103,0.07548718,0.08205129,0.09189744,0.10502565,0.13784617,0.18379489,0.24615386,0.29538465,0.34133336,0.42994875,0.48246157,0.4955898,0.5021539,0.508718,0.49887183,0.46933338,0.44307697,0.43323082,0.43323082,0.4266667,0.43323082,0.45620516,0.4955898,0.5481026,0.60061544,0.6695385,0.74830776,0.8533334,0.9616411,1.0075898,1.014154,1.0601027,1.1684103,1.3522053,1.6147693,2.0841026,3.1967182,4.9394875,6.426257,5.901129,5.622154,5.5696416,5.2545643,4.84759,5.1954875,6.1046157,6.51159,6.5805135,6.698667,7.4830775,9.45559,10.371283,11.083488,11.30995,9.626257,8.182155,7.9458466,8.004924,8.044309,8.3364105,9.232411,9.055181,7.824411,5.7764106,3.3608208,2.1431797,1.086359,0.4004103,0.10502565,0.049230773,0.049230773,0.08861539,0.190359,0.36102566,0.5973334,0.9156924,2.034872,3.7382567,5.5138464,6.547693,6.951385,7.9261546,10.31877,14.158771,18.668308,23.666874,29.216824,34.487797,38.656002,40.90421,42.085747,42.433643,44.402874,49.352207,57.537647,68.992004,80.74503,91.241035,101.80924,116.65396,121.35057,118.173546,110.165344,100.67693,93.344826,87.04329,76.54729,66.737236,59.58893,54.166977,48.475903,43.0999,38.288414,34.18585,30.831593,27.464207,24.73354,21.779694,18.484514,15.465027,12.612924,10.020103,7.7718983,5.8486156,4.141949,2.8389745,1.9003079,1.2931283,0.9682052,0.8467693,0.8369231,0.69579494,0.47589746,0.25271797,0.12143591,0.04266667,0.02297436,0.04266667,0.11158975,0.27241027,1.2832822,2.9440002,4.6933336,5.7632823,5.1856413,4.4438977,3.05559,2.2121027,2.5238976,4.0467696,5.146257,3.8367183,2.0217438,0.827077,0.6104616,1.1290257,1.1815386,0.8041026,0.28225642,0.11158975,0.04266667,0.013128206,0.0032820515,0.0,0.0,0.006564103,0.029538464,0.032820515,0.026256412,0.06564103,0.06564103,0.029538464,0.013128206,0.016410258,0.009846155,0.0,0.75487185,0.90584624,0.5415385,0.11158975,0.4266667,1.4966155,1.2012309,0.6498462,0.58092314,1.3587693,0.64000005,0.26256412,0.14441027,0.27569234,0.71548724,0.2100513,0.032820515,0.17723078,0.574359,1.1093334,0.4201026,0.098461546,0.15753847,0.38400003,0.34789747,0.4201026,0.8369231,0.827077,0.5481026,1.0633847,1.0732309,2.5140514,2.4516926,1.1881026,2.2580514,1.4244103,1.0535386,1.7001027,2.5731285,1.5458462,0.5513847,1.3062565,2.156308,2.2022567,1.2800001,3.8596926,3.5282054,2.03159,0.6662565,0.28225642,0.29210258,0.82379496,1.5885129,1.8281027,0.3249231,0.27569234,0.17066668,0.09189744,0.06235898,0.036102567,0.026256412,0.128,0.13456412,0.036102567,0.01969231,0.08533334,1.1585642,1.3357949,0.67610264,1.1979488,1.1881026,1.211077,1.1716924,1.1913847,1.591795,2.7241027,3.0818465,3.4560003,4.0041027,4.2568207,3.2656412,2.6256413,2.7142565,3.367385,3.892513,3.6069746,2.802872,3.0162053,4.493129,6.163693,5.2381544,5.3792825,5.868308,6.193231,6.045539,5.85518,4.562052,3.367385,2.7766156,2.5961027,2.2777438,2.2482052,2.0742567,1.5786668,0.8467693,0.63343596,0.36430773,0.15425642,0.08205129,0.20676924,0.36758977,0.2231795,0.118153855,0.15753847,0.20020515,0.2100513,0.56451285,1.6278975,3.436308,5.6976414,6.1997952,6.3573337,6.2851286,5.901129,4.923077,4.269949,3.4855387,2.6223593,1.8248206,1.3259488,1.4211283,1.4309745,1.4441026,1.5163078,1.6705642,1.7558975,1.9856411,2.2908719,2.556718,2.6322052,2.7241027,2.674872,2.4713848,2.1464617,1.7624617,1.7723079,1.7427694,1.8871796,2.3204105,3.0687182,3.945026,3.817026,3.757949,4.3585644,5.720616,5.9667697,5.5729237,5.0609236,4.7261543,4.630975,5.221744,5.2676926,5.0642056,4.6834874,3.9581542,4.460308,5.681231,6.688821,6.994052,6.547693,4.57518,3.2098465,2.789744,3.1113849,3.4560003,5.32677,6.0160003,6.770872,7.8112826,8.326565,8.4053335,7.6307697,7.466667,7.53559,5.602462,5.32677,5.228308,4.95918,4.7327185,5.333334,5.989744,5.5105643,4.138667,2.5140514,1.6607181,1.9954873,2.789744,3.3444104,3.5052311,3.6726158,6.5312824,6.885744,6.1440005,5.4383593,5.602462,4.6605134,3.8596926,4.2535386,5.3005133,4.8640003,4.135385,3.889231,4.1813335,4.460308,3.5577438,3.8038976,4.709744,5.4449234,5.8814363,6.6034875,5.533539,3.5872824,2.4188719,2.7536411,4.414359,5.077334,5.431795,5.5696416,5.425231,4.7983594,5.2020516,5.970052,5.5532312,4.132103,3.6332312,3.626667,3.259077,3.0949745,3.3247182,3.7284105,3.8629746,3.751385,3.4855387,2.9440002,1.8084104,0.9714873,0.4955898,0.5546667,1.2176411,2.4516926,2.6683078,2.5206156,2.3466668,2.2022567,1.8510771,1.6836925,2.03159,2.3663592,2.5271797,2.740513,3.4133337,3.058872,2.9505644,3.5446157,4.466872,5.0477953,5.1364107,5.287385,5.904411,7.240206,7.4797955,7.834257,8.457847,9.275078,9.96759,9.977437,10.597744,11.1294365,11.241027,10.975181,10.157949,8.500513,7.240206,6.7807183,6.6822567,4.453744,3.1770258,3.1573336,3.820308,3.6890259,2.359795,2.2088206,2.8356924,3.4034874,2.6289232,2.356513,1.913436,1.3817437,0.90912825,0.69579494,0.65641034,0.6892308,0.7220513,0.7318975,0.761436,0.81394875,0.90912825,1.1388719,1.4572309,1.6804104,2.0512822,2.8192823,3.058872,2.868513,3.3903592,2.7273848,2.537026,2.993231,4.096,5.7009234,4.95918,4.056616,4.9920006,7.8014364,10.55836,12.970668,12.42913,10.226872,7.975385,7.6110773,6.7282057,5.3005133,3.6069746,2.0906668,1.3423591,1.8281027,2.409026,2.8192823,2.9604106,2.9046156,2.9111798,2.7634873,2.2777438,1.7591796,2.03159,3.114667,2.6584618,2.0151796,1.8609232,2.1825643,1.9035898,1.6114873,1.2931283,1.017436,0.9517949,0.7778462,0.48246157,0.26584616,0.19692309,0.20020515,0.14769232,0.13128206,0.10502565,0.10502565,0.24615386,1.6410258,2.409026,2.733949,2.7995899,2.806154,1.3259488,0.5284103,0.16410258,0.052512825,0.068923086,0.30851284,0.51856416,0.71548724,0.84348726,0.77128214,0.67610264,0.60389745,0.45292312,0.21989745,0.026256412,0.016410258,0.118153855,0.13128206,0.03938462,0.026256412,0.32820517,0.17723078,0.08533334,0.23958977,0.512,0.35774362,0.27569234,0.23630771,0.21989745,0.22646156,0.43651286,0.24943592,0.052512825,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.0,0.006564103,0.016410258,0.01969231,0.016410258,0.032820515,0.072205134,0.06564103,0.068923086,0.27897438,0.49887183,0.4135385,0.34133336,0.5218462,1.1257436,1.591795,1.5360001,1.2964103,1.2209232,1.657436,2.1202054,1.9659488,1.1946667,0.3117949,0.3249231,0.17066668,0.17394873,0.25271797,0.34133336,0.3708718,0.4955898,0.42338464,0.43651286,0.48902568,0.17723078,0.0951795,0.059076928,0.055794876,0.072205134,0.07876924,0.02297436,0.04266667,0.03938462,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.013128206,0.013128206,0.013128206,0.006564103,0.01969231,0.029538464,0.032820515,0.03938462,0.03938462,0.055794876,0.055794876,0.052512825,0.049230773,0.06564103,0.068923086,0.07876924,0.09189744,0.10502565,0.13784617,0.17723078,0.2231795,0.27241027,0.33476925,0.43651286,0.47917953,0.5152821,0.54482055,0.56451285,0.55794877,0.5349744,0.4955898,0.46276927,0.43651286,0.4266667,0.43323082,0.45292312,0.47589746,0.49887183,0.508718,0.51856416,0.54482055,0.61374366,0.7253334,0.8369231,0.92553854,1.017436,1.1126155,1.2471796,1.4933335,2.0873847,3.131077,4.8705645,6.698667,7.13518,7.27959,7.64718,7.778462,7.643898,7.6603084,7.8145647,8.211693,8.628513,9.163487,10.240001,11.516719,11.559385,11.835078,12.140308,10.633847,9.18318,8.887795,9.084719,9.012513,7.781744,7.240206,6.7971287,6.226052,5.211898,3.367385,1.9364104,0.9156924,0.31507695,0.072205134,0.02297436,0.02297436,0.03938462,0.052512825,0.06235898,0.072205134,0.101743594,0.81066674,2.0053334,3.2295387,3.7415388,3.3378465,3.006359,3.4034874,4.7228723,6.698667,9.7673855,13.725539,18.20554,22.662565,26.41395,30.119387,32.439796,34.149746,35.96472,38.547695,43.45108,49.35549,59.01785,73.898674,94.20145,108.72452,118.70196,124.6195,126.75939,125.2234,115.551186,101.73703,86.4197,72.66134,63.914673,58.945644,54.980927,51.01621,46.690464,42.27939,37.293953,33.72308,30.368822,26.95877,24.146053,20.473438,17.027283,13.909334,11.149129,8.687591,6.616616,4.965744,3.7842054,3.0490258,2.6551797,2.297436,1.7952822,1.2274873,0.6826667,0.256,0.06235898,0.009846155,0.016410258,0.049230773,0.118153855,0.28882053,0.56123084,1.0535386,1.6607181,2.0545642,2.1431797,1.9035898,2.1891284,3.3411283,5.1889234,6.042257,3.8006158,1.6278975,0.761436,0.5316923,0.47589746,0.3708718,0.2297436,0.108307704,0.07548718,0.036102567,0.013128206,0.0032820515,0.0,0.0,0.006564103,0.029538464,0.032820515,0.026256412,0.06564103,0.06564103,0.029538464,0.049230773,0.128,0.20348719,0.0,1.2635899,1.2865642,0.65969235,0.098461546,0.44964105,2.2219489,1.654154,0.63343596,0.25271797,0.8369231,0.3249231,0.13128206,0.16082053,0.2231795,0.02297436,0.006564103,0.07548718,0.108307704,0.12471796,0.28225642,0.2855385,0.1148718,0.0,0.006564103,0.036102567,0.24943592,0.7975385,0.7581539,0.28225642,0.6104616,1.3915899,3.5577438,3.5314875,1.7526156,2.678154,1.8609232,1.1815386,0.8008206,0.6498462,0.44964105,0.33805132,0.8041026,0.955077,0.79097444,1.1913847,1.719795,0.90256417,0.40369233,0.58092314,0.4955898,0.508718,1.6246156,3.131077,3.4691284,0.2297436,0.20348719,0.13456412,0.06564103,0.02297436,0.0,0.013128206,0.27241027,0.34789747,0.20020515,0.21333335,0.28882053,2.0184617,2.1202054,0.7975385,1.7493335,2.0841026,2.284308,2.0709746,1.5556924,1.2373334,1.8937438,2.809436,4.2896414,5.7009234,5.464616,3.3903592,2.789744,2.937436,3.2886157,3.495385,3.2623591,3.7251284,5.6320004,8.267488,9.465437,6.3967185,5.8945646,5.865026,5.421949,4.896821,5.687795,5.0084105,3.6332312,2.4188719,2.284308,2.1070771,1.8609232,1.7624617,1.6246156,0.8598975,0.4004103,0.15097436,0.04266667,0.013128206,0.013128206,0.013128206,0.013128206,0.006564103,0.0,0.0,0.0,0.013128206,0.14441027,0.7318975,2.3729234,3.9417439,4.8016415,5.284103,5.5171285,5.412103,5.1856413,4.4865646,3.6004105,2.8258464,2.4484105,2.4943593,2.2153847,1.9790771,1.9331284,2.0086155,1.8707694,1.9462565,2.0709746,2.1300514,2.034872,2.1792822,2.3302567,2.3072822,2.0841026,1.8084104,1.5031796,1.2603078,1.211077,1.4966155,2.284308,3.239385,3.121231,2.9702566,3.4494362,4.844308,5.169231,4.9821544,4.900103,5.1167183,5.428513,5.8092313,6.2916927,6.2720003,5.6418467,4.781949,5.4186673,6.452513,7.3649235,7.325539,5.175795,2.6026669,1.4375386,1.4703591,2.284308,3.2754874,6.564103,7.834257,7.9163084,7.6603084,7.939283,9.291488,8.303591,7.128616,5.9470773,2.9604106,2.7437952,3.4658465,4.332308,5.1331286,6.245744,6.8562055,5.579488,3.6135387,2.0939488,2.0676925,2.7963078,3.6332312,4.4012313,4.850872,4.6539493,6.8988724,7.1909747,6.5870776,5.87159,5.540103,4.1485133,3.817026,4.8049235,6.245744,6.160411,4.9099493,4.2174363,4.3060517,4.7556925,4.519385,4.70318,4.269949,4.33559,4.9887185,5.3234878,4.6080003,3.0785644,1.9954873,2.1234872,3.7349746,4.4307694,4.637539,4.33559,3.623385,2.7306669,3.1573336,3.623385,3.31159,2.3040001,1.6246156,1.3915899,0.86317956,0.50543594,0.6268718,1.3784616,1.3062565,1.1027694,0.90256417,0.6859488,0.25271797,0.049230773,0.0,0.01969231,0.06235898,0.128,0.2231795,0.43651286,0.8369231,1.2077949,1.0469744,0.93866676,1.2012309,1.5031796,1.7296412,2.0020514,2.8816411,3.3969233,3.9844105,4.640821,4.900103,3.7743592,3.761231,4.9329233,6.557539,7.0793853,6.5444107,6.626462,7.6012316,9.472001,11.976206,11.54954,12.143591,12.645744,12.635899,12.379898,10.627283,8.707283,7.397744,6.889026,6.7774363,4.391385,3.6890259,3.9581542,4.128821,2.7798977,2.2514873,2.1300514,2.172718,2.2646155,2.4155898,1.5983591,1.0371283,0.83035904,0.8763078,0.8598975,1.2209232,1.2274873,1.1323078,1.1520001,1.4769232,1.8281027,1.785436,1.6738462,1.657436,1.7591796,3.1343591,4.5095387,5.3727183,5.868308,6.813539,5.172513,4.1550775,3.9154875,3.9023592,2.8947694,2.225231,2.3794873,3.6069746,5.5532312,7.276308,9.110975,10.755282,11.451077,10.893129,9.252103,8.536616,6.7872825,4.8114877,3.2065644,2.3827693,2.487795,2.609231,2.7044106,2.7602053,2.7963078,3.1277952,3.4724104,3.006359,1.9790771,1.7329233,2.6157951,2.4516926,1.9692309,1.5524104,1.2537436,1.394872,1.3554872,1.1257436,0.83035904,0.7581539,0.6826667,0.4955898,0.32164106,0.19692309,0.07876924,0.07548718,0.098461546,0.098461546,0.128,0.3511795,1.910154,2.9997952,3.3608208,2.9833848,2.1431797,0.77128214,0.33476925,0.24287182,0.23630771,0.38728207,0.8763078,1.1454359,1.4473847,1.719795,1.5885129,1.214359,0.88615394,0.5349744,0.22646156,0.16410258,0.14769232,0.3249231,0.3446154,0.17394873,0.08533334,0.7220513,0.45620516,0.27897438,0.4201026,0.34789747,0.27569234,0.39056414,0.4594872,0.4135385,0.34133336,0.49887183,0.30851284,0.0951795,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.0032820515,0.013128206,0.02297436,0.02297436,0.013128206,0.0032820515,0.006564103,0.009846155,0.052512825,0.25271797,0.098461546,0.029538464,0.016410258,0.13784617,0.574359,1.2340513,1.6377437,1.6607181,1.3587693,0.94523084,0.73517954,0.6826667,0.6170257,0.508718,0.4397949,0.2297436,0.24943592,0.39384618,0.5152821,0.446359,0.47917953,0.49230772,0.45292312,0.3446154,0.15425642,0.07876924,0.07876924,0.059076928,0.01969231,0.02297436,0.0032820515,0.013128206,0.016410258,0.0032820515,0.0,0.016410258,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.0032820515,0.006564103,0.016410258,0.016410258,0.016410258,0.02297436,0.029538464,0.032820515,0.036102567,0.068923086,0.06235898,0.052512825,0.059076928,0.07548718,0.06564103,0.072205134,0.08861539,0.108307704,0.13456412,0.18379489,0.22646156,0.27569234,0.33805132,0.4135385,0.45292312,0.508718,0.55794877,0.58420515,0.5874872,0.5677949,0.52512825,0.48902568,0.46276927,0.4397949,0.44307697,0.4594872,0.47261542,0.47261542,0.45620516,0.446359,0.446359,0.48246157,0.56451285,0.69907695,0.827077,0.955077,1.0601027,1.1979488,1.4933335,2.2580514,3.387077,5.1298466,7.273026,9.160206,8.776206,9.645949,10.857026,11.510155,10.71918,9.724719,10.509129,12.20595,14.080001,15.510976,15.346873,13.5778475,12.117334,11.286975,9.819899,11.244308,12.973949,14.569027,14.8709755,12.018872,9.83959,8.477539,7.384616,5.979898,3.636513,1.7427694,0.7089231,0.24287182,0.08533334,0.01969231,0.01969231,0.026256412,0.029538464,0.029538464,0.04266667,0.04266667,0.055794876,0.108307704,0.19364104,0.2855385,0.3446154,0.48246157,0.69251287,0.96492314,1.2898463,2.1202054,3.5282054,5.756718,8.828718,12.57354,17.539284,22.472206,26.397541,28.921438,30.227695,33.217644,36.995285,41.104412,46.125954,53.67467,66.714264,86.87591,110.1916,131.02934,142.12924,136.60555,126.0636,110.80534,93.46954,79.02524,72.22154,68.24042,65.01088,61.292313,56.66134,50.418877,45.31857,40.815594,36.90339,34.12021,29.988106,26.09231,22.373745,18.825848,15.491283,12.6063595,10.200616,8.326565,6.9710774,6.0750775,5.225026,4.2305646,3.1376412,2.0250258,0.98461545,0.4594872,0.19692309,0.08205129,0.032820515,0.02297436,0.052512825,0.101743594,0.256,0.53825647,0.9124103,1.1257436,1.2176411,1.8445129,3.239385,5.2020516,6.160411,3.7710772,1.6377437,0.9944616,0.72861546,0.62030774,0.45620516,0.3446154,0.30194873,0.25271797,0.24287182,0.3249231,0.24943592,0.059076928,0.06235898,0.04266667,0.04266667,0.07548718,0.1148718,0.08533334,0.049230773,0.029538464,0.098461546,0.24943592,0.4201026,0.0,1.0502565,1.4867693,0.9616411,0.18051283,0.8992821,1.1191796,1.6607181,1.404718,0.6892308,1.3128207,0.81066674,0.5316923,0.43323082,0.37743592,0.12143591,0.036102567,0.3708718,0.4135385,0.12143591,0.12143591,0.29210258,0.13456412,0.0,0.036102567,0.18379489,0.6104616,0.63343596,0.50543594,0.45292312,0.67282057,2.6256413,3.4789746,2.9833848,1.8970258,1.9823592,1.1651284,0.38400003,0.3249231,0.8992821,1.2668719,0.47261542,0.5021539,0.43651286,0.128,0.21333335,0.27569234,0.19692309,0.13784617,0.45620516,1.7394873,1.5195899,1.6016412,1.7132308,1.4605129,0.3511795,0.2297436,0.13456412,0.06564103,0.02297436,0.0,0.013128206,0.17066668,0.4397949,0.761436,1.0666667,1.1520001,0.6432821,0.31507695,0.380718,0.5021539,0.9189744,1.1224617,1.0075898,0.6859488,0.5021539,0.47917953,1.1060513,2.8192823,5.208616,7.003898,6.9776416,8.182155,8.303591,6.6560006,4.164923,3.6890259,4.824616,6.514872,7.4765134,6.196513,3.7776413,4.2830772,5.208616,5.3858466,4.95918,4.3618464,2.681436,1.3095386,1.0272821,2.028308,4.263385,4.6211286,4.588308,4.082872,1.4342566,0.446359,0.08861539,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.06564103,0.19692309,0.380718,0.8566154,1.6147693,2.5304618,3.373949,3.2754874,2.9571285,2.809436,3.1442053,4.1813335,4.6572313,4.273231,3.876103,3.764513,3.692308,2.9604106,2.5862565,2.412308,2.2908719,2.0611284,2.097231,2.2055387,2.231795,2.103795,1.847795,1.4933335,1.1552821,0.92553854,1.014154,1.7690258,2.550154,2.1989746,1.8051283,1.9265642,2.546872,2.9997952,4.056616,4.8311796,5.428513,6.941539,5.7698464,6.311385,6.482052,5.4547696,3.6463592,4.1485133,5.1232824,5.7632823,5.5171285,4.089436,2.8914874,2.1464617,1.913436,2.2613335,3.249231,6.8988724,9.104411,8.730257,6.7544622,6.242462,7.5946674,7.5585647,6.6428723,5.2053337,3.4494362,3.5938463,4.06318,4.824616,5.5762057,5.720616,5.3070774,4.086154,3.2000003,3.045744,3.2656412,3.7776413,4.9394875,6.6133337,8.155898,8.438154,5.9963083,5.677949,5.421949,4.6834874,4.4406157,4.1222568,3.8071797,3.5610259,3.1343591,1.9396925,1.4867693,1.5753847,2.228513,3.3608208,4.775385,4.716308,3.8498464,3.190154,3.2000003,3.7842054,2.9407182,2.2088206,1.5327181,1.0502565,1.0994873,1.014154,1.2307693,1.467077,1.5097437,1.204513,1.1815386,1.0469744,0.764718,0.37743592,0.0,0.20676924,0.10502565,0.0,0.0,0.0,0.12143591,0.06235898,0.0,0.02297436,0.108307704,0.02297436,0.0,0.04266667,0.128,0.21333335,0.34789747,0.56451285,1.0043077,1.5458462,1.8149745,2.3040001,2.3335385,2.3696413,2.5632823,2.7470772,3.442872,3.761231,3.7743592,3.754667,4.1813335,4.1682053,4.6867695,5.5236926,6.1046157,5.4941545,4.578462,4.578462,5.664821,7.325539,8.362667,8.618668,9.5146675,10.86359,12.235488,12.954257,11.611898,9.83959,7.463385,5.3727183,5.5072823,3.629949,3.8071797,5.028103,5.6976414,3.6463592,3.6824617,4.525949,4.640821,3.626667,2.1956925,1.024,1.0075898,1.591795,2.2514873,2.4713848,2.7536411,2.9243078,3.1540515,3.3575387,3.1737437,3.367385,2.6584618,2.2121027,2.3827693,2.7011285,3.9581542,5.910975,7.9983597,9.035488,7.2172313,4.1780515,2.7044106,2.156308,1.8806155,1.2209232,1.0502565,1.6672822,2.917744,4.955898,8.241231,11.168821,13.587693,13.072412,9.741129,6.226052,5.8092313,5.2315903,5.5007186,6.449231,6.7282057,5.543385,4.699898,4.0041027,3.6004105,3.9680004,3.2361028,2.9702566,3.0227695,2.930872,1.8904617,1.5622566,1.5064616,1.4342566,1.204513,0.8402052,1.2406155,1.2800001,1.1191796,0.96492314,1.0371283,0.7187693,0.5677949,0.34789747,0.07876924,0.029538464,0.10502565,0.17723078,0.17723078,0.15425642,0.28882053,1.3883078,2.5796926,2.858667,2.1070771,1.0666667,0.5546667,0.36430773,0.4660513,0.81394875,1.3259488,1.4736412,1.4375386,1.5524104,1.723077,1.4178462,1.0043077,0.8730257,0.7253334,0.5546667,0.64000005,0.60389745,0.4397949,0.4201026,0.52512825,0.4266667,0.53825647,0.636718,0.60061544,0.43323082,0.27569234,0.21333335,0.08861539,0.068923086,0.12143591,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.02297436,0.04594872,0.059076928,0.04266667,0.029538464,0.049230773,0.12143591,0.892718,1.7887181,2.1792822,1.8970258,1.2504616,1.1290257,1.273436,1.1257436,0.63343596,0.24287182,0.12143591,0.23958977,0.512,0.7515898,0.64000005,0.4201026,0.45620516,0.512,0.4594872,0.28882053,0.20348719,0.118153855,0.059076928,0.032820515,0.04594872,0.009846155,0.072205134,0.07876924,0.013128206,0.0,0.036102567,0.036102567,0.01969231,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.016410258,0.016410258,0.016410258,0.016410258,0.026256412,0.049230773,0.06235898,0.072205134,0.07548718,0.08205129,0.08861539,0.07548718,0.07548718,0.07548718,0.08205129,0.098461546,0.12143591,0.17066668,0.2297436,0.28225642,0.32820517,0.36758977,0.40369233,0.4660513,0.5152821,0.5415385,0.56451285,0.5513847,0.5218462,0.5021539,0.49887183,0.48902568,0.46276927,0.45620516,0.446359,0.41682056,0.380718,0.380718,0.4004103,0.45620516,0.5415385,0.6268718,0.7220513,0.86646163,1.0075898,1.1979488,1.6016412,2.5435898,3.7120004,5.3398976,7.6603084,10.893129,11.700514,12.934566,14.204719,14.713437,13.259488,12.675283,15.530668,19.11795,21.090464,19.456001,15.254975,11.835078,10.509129,10.896411,10.893129,17.329231,21.379284,22.636309,21.589334,19.623386,17.23077,14.332719,11.264001,8.044309,4.394667,1.9528207,0.81066674,0.32820517,0.1148718,0.029538464,0.029538464,0.029538464,0.02297436,0.01969231,0.029538464,0.029538464,0.029538464,0.04266667,0.06564103,0.09189744,0.09189744,0.118153855,0.16738462,0.23958977,0.3511795,0.5349744,0.88287187,1.4933335,2.540308,4.273231,7.4240007,11.680821,16.049232,20.096,23.942566,27.664412,30.893951,33.98236,36.877132,39.125336,41.859283,48.07549,57.852722,72.19529,93.019905,115.01621,129.09293,134.30154,129.77232,114.68144,96.141136,81.56226,73.72144,71.89662,71.88349,68.06319,62.483696,55.78831,49.014156,43.59221,39.72267,36.276516,32.771286,28.94113,24.71713,20.995283,17.795284,15.05477,12.763899,10.971898,9.6525135,8.260923,6.636308,4.7950773,2.9144619,1.7920002,0.90584624,0.3511795,0.12143591,0.12143591,0.15753847,0.23958977,0.30851284,0.3511795,0.4135385,0.49887183,0.53825647,0.7187693,1.2832822,2.5173335,3.8859491,2.8455386,2.0086155,1.9265642,1.083077,1.1684103,0.9878975,0.8960001,0.92553854,0.7778462,0.92553854,1.4834872,1.214359,0.29210258,0.3052308,0.20676924,0.17394873,0.32164106,0.52512825,0.4266667,0.24287182,0.15097436,0.12143591,0.128,0.15097436,0.0,0.2100513,0.2986667,0.19364104,0.12471796,0.6301539,1.4769232,2.0118976,1.719795,0.8205129,0.26256412,1.020718,0.7417436,0.34133336,0.23302566,0.32820517,0.32164106,0.25271797,0.13456412,0.02297436,0.02297436,0.098461546,0.04594872,0.0,0.006564103,0.036102567,0.37743592,0.62030774,0.67610264,0.62030774,0.6826667,0.9288206,0.99774367,0.8763078,0.7450257,0.95835906,0.7253334,0.4201026,0.29210258,0.34789747,0.36430773,0.18379489,0.23630771,0.27897438,0.2231795,0.15097436,0.7417436,0.8336411,0.5415385,0.21333335,0.4201026,0.41682056,0.5513847,0.636718,0.5546667,0.25271797,0.20020515,0.13784617,0.08861539,0.101743594,0.24287182,0.098461546,0.059076928,0.190359,0.43323082,0.5907693,0.45292312,0.3117949,0.6235898,1.6246156,3.3476925,2.3171284,1.7591796,1.2603078,0.8566154,1.017436,1.1684103,1.2373334,2.3794873,4.3684106,5.5762057,6.8004107,6.925129,6.0750775,4.841026,4.263385,4.5095387,4.266667,3.9844105,3.7218463,3.1442053,2.3860514,2.4320002,2.5009232,2.297436,2.0184617,1.8674873,1.3292309,0.88615394,0.86646163,1.4080001,2.809436,3.698872,3.889231,3.1540515,1.2406155,0.4955898,0.16082053,0.03938462,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.052512825,0.13784617,0.0951795,0.18707694,0.36758977,0.5973334,0.8467693,0.8172308,0.72861546,0.7417436,0.9682052,1.4605129,1.8773335,2.172718,2.5731285,2.986667,3.0227695,3.1277952,3.0884104,3.0326157,2.9538465,2.681436,2.7011285,2.612513,2.3663592,2.028308,1.8084104,1.6016412,1.3259488,1.0896411,0.9682052,1.014154,1.2176411,1.0929232,1.0436924,1.2242053,1.5360001,2.3368206,2.917744,3.242667,3.8728209,5.940513,6.0685134,6.370462,5.8945646,4.775385,4.20759,4.4045134,4.2141542,4.457026,5.093744,5.2480006,4.9887185,4.8640003,4.824616,5.1331286,6.373744,8.969847,9.987283,8.917334,6.813539,6.2884107,7.3616414,7.1581545,6.23918,5.3136415,5.2545643,4.9132314,5.1331286,5.398975,5.3727183,4.903385,4.0992823,3.511795,3.373949,3.626667,3.9253337,4.818052,6.4722056,8.352821,9.4457445,8.241231,5.917539,6.091488,6.235898,5.4974365,4.6966157,3.1770258,2.166154,1.7099489,1.5655385,1.1815386,1.2176411,2.1234872,3.436308,4.493129,4.4340515,3.3476925,2.3729234,1.6836925,1.3784616,1.463795,1.910154,1.8084104,1.1913847,0.45620516,0.37743592,0.23302566,0.38400003,0.6268718,0.7515898,0.5349744,0.4397949,0.33476925,0.2100513,0.08533334,0.0,0.04266667,0.01969231,0.0,0.0,0.0,0.02297436,0.013128206,0.0,0.0032820515,0.02297436,0.0032820515,0.0,0.009846155,0.055794876,0.190359,0.19692309,0.36758977,0.7318975,1.2176411,1.6311796,2.03159,2.0578463,2.0086155,2.3302567,3.5872824,4.9887185,5.353026,4.568616,3.5478978,4.2305646,3.6791797,3.5741541,3.7316926,4.017231,4.332308,4.962462,6.298257,7.351795,7.9261546,8.641642,9.954462,10.807796,10.709334,9.90195,9.340718,9.347282,8.992821,8.320001,7.450257,6.6067696,4.7655387,4.568616,5.037949,4.9460516,2.8160002,2.806154,2.930872,2.674872,2.0151796,1.4276924,2.2186668,3.4592824,3.9942567,3.4855387,2.4352822,2.6387694,3.1638978,3.2689233,3.0260515,3.3214362,2.5895386,1.6082052,1.9232821,3.4691284,4.568616,6.567385,7.1023593,6.6428723,5.5269747,3.9712822,2.4352822,1.6968206,1.3718976,1.1323078,0.7089231,1.1520001,3.4297438,7.88677,13.039591,15.599591,18.110361,17.046976,13.66318,10.082462,9.301334,12.196103,10.131693,7.8736415,7.322257,7.4863596,6.7314878,5.83877,5.1626673,4.906667,5.1265645,4.7458467,3.9089234,3.117949,2.556718,2.0742567,1.4145643,1.1585642,1.079795,1.0732309,1.1552821,1.0994873,1.1979488,1.2242053,1.1552821,1.1585642,0.71548724,0.36102566,0.15097436,0.07548718,0.06564103,0.13128206,0.21661541,0.21989745,0.256,0.6432821,1.2931283,1.595077,1.5097437,1.1716924,0.8960001,0.65641034,0.51856416,0.57764107,0.8598975,1.3161026,1.8707694,2.2219489,2.3204105,2.1792822,1.8838975,1.2340513,0.67610264,0.46276927,0.508718,0.41025645,0.6170257,0.5874872,0.8369231,1.204513,0.84348726,0.67938465,0.41682056,0.23630771,0.15425642,0.055794876,0.04266667,0.016410258,0.013128206,0.02297436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.02297436,0.036102567,0.052512825,0.06235898,0.049230773,0.26256412,0.6170257,0.86974365,0.8795898,0.60389745,0.6498462,0.78769237,0.71548724,0.4135385,0.15753847,0.13456412,0.3052308,0.48246157,0.52512825,0.34789747,0.17723078,0.15097436,0.15753847,0.14769232,0.14441027,0.108307704,0.068923086,0.03938462,0.016410258,0.009846155,0.0032820515,0.013128206,0.04594872,0.068923086,0.036102567,0.013128206,0.013128206,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.013128206,0.016410258,0.02297436,0.036102567,0.049230773,0.08205129,0.101743594,0.1148718,0.11158975,0.101743594,0.101743594,0.09189744,0.0951795,0.108307704,0.12143591,0.13128206,0.18051283,0.2297436,0.27241027,0.32820517,0.37743592,0.4201026,0.4397949,0.446359,0.47917953,0.48574364,0.50543594,0.5218462,0.52512825,0.512,0.48902568,0.48246157,0.46933338,0.446359,0.41682056,0.4266667,0.4397949,0.45620516,0.47589746,0.5021539,0.571077,0.69907695,0.9189744,1.2898463,1.9068719,2.8947694,4.1124105,5.901129,8.598975,12.566976,16.489027,24.392206,29.039593,27.342772,20.352001,24.365952,25.51467,23.210669,18.579693,14.464001,13.223386,11.428103,9.892103,9.035488,8.881231,12.022155,14.221129,15.451899,15.911386,15.996719,14.562463,11.378873,8.067283,5.4974365,3.7710772,1.9659488,0.88615394,0.32164106,0.08533334,0.01969231,0.029538464,0.029538464,0.02297436,0.013128206,0.006564103,0.016410258,0.032820515,0.06564103,0.12143591,0.21333335,0.26256412,0.24943592,0.2231795,0.21989745,0.28882053,0.35446155,0.5284103,0.9124103,1.4998976,2.1497438,3.2853336,5.172513,7.4732313,10.082462,13.124924,16.850052,20.371695,23.958977,27.762875,31.8359,34.500927,38.4558,43.464207,49.598362,57.24226,67.695595,79.89826,93.9159,107.894165,118.07837,117.71734,110.14565,99.28534,88.23139,79.24513,72.90421,69.018265,65.5918,61.57457,56.83857,51.797337,47.44862,43.77272,40.438156,36.791798,31.661951,27.40513,23.811283,20.79836,18.41559,16.367592,14.037334,11.716924,9.475283,7.174565,5.1232824,3.442872,2.1366155,1.1881026,0.574359,0.6301539,0.7318975,0.8172308,0.8960001,1.0338463,1.1881026,1.1881026,1.1979488,1.4276924,2.103795,3.1081028,3.318154,3.511795,3.5577438,2.4024618,2.028308,1.6902566,1.4900514,1.4309745,1.401436,2.3368206,1.9429746,1.1881026,0.6629744,0.5973334,0.5481026,0.6826667,1.1454359,1.8149745,2.294154,1.5458462,1.0699488,0.90912825,0.92553854,0.82379496,0.0,0.0,0.0,0.0,0.04594872,0.23630771,1.339077,2.7437952,2.5238976,0.8533334,0.0,0.42994875,0.50543594,0.34789747,0.14441027,0.15097436,0.18051283,0.101743594,0.026256412,0.0,0.0,0.01969231,0.009846155,0.0,0.0,0.0,0.16410258,0.4397949,0.53825647,0.42994875,0.36758977,0.21989745,0.16082053,0.15097436,0.18379489,0.28225642,0.29210258,0.20348719,0.128,0.0951795,0.072205134,0.06235898,0.09189744,0.12143591,0.12471796,0.072205134,0.79425645,0.7253334,0.380718,0.108307704,0.09189744,0.12471796,0.19364104,0.22646156,0.20348719,0.16410258,0.15097436,0.128,0.118153855,0.14441027,0.23302566,0.072205134,0.013128206,0.059076928,0.3117949,0.97805136,0.96492314,2.2022567,3.3805132,3.9056413,3.9122055,3.626667,3.6857438,4.06318,4.3290257,3.6430771,2.937436,2.1858463,2.6715899,4.1878977,5.044513,5.4843082,5.284103,5.287385,5.924103,7.1909747,7.1548724,5.4941545,3.820308,2.793026,2.1431797,1.4769232,1.2471796,1.1158975,0.98133343,0.9714873,1.3292309,1.1126155,0.72861546,0.47589746,0.53825647,1.0075898,1.404718,1.5031796,1.2012309,0.5218462,0.26256412,0.108307704,0.029538464,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.026256412,0.049230773,0.009846155,0.006564103,0.02297436,0.04594872,0.08533334,0.08205129,0.068923086,0.09189744,0.17066668,0.3117949,0.47261542,0.6662565,1.0699488,1.5885129,1.8543591,2.231795,2.5698464,2.733949,2.865231,3.370667,3.3969233,3.0720003,2.6322052,2.2744617,2.176,2.2088206,2.097231,1.7001027,1.1060513,0.64000005,0.6071795,0.62030774,0.73517954,0.99774367,1.463795,1.8871796,2.3236926,2.934154,3.889231,5.3792825,5.737026,6.196513,5.72718,4.5554876,4.1747694,4.414359,4.2863593,4.204308,4.414359,4.962462,5.0477953,5.7796926,6.8299494,7.817847,8.310155,10.312206,12.258463,11.82195,9.31118,7.6668725,7.8834877,7.9097443,7.3682055,6.5805135,6.567385,5.467898,5.077334,4.8804107,4.594872,4.1682053,3.8728209,4.1485133,4.7556925,5.402257,5.717334,5.5072823,6.692103,7.962257,8.480822,7.8736415,7.525744,8.3823595,7.962257,5.874872,3.8071797,3.0523078,2.300718,1.9429746,1.8576412,1.394872,1.5885129,2.425436,3.1934361,3.4494362,2.9833848,2.2777438,1.7132308,1.2242053,0.86646163,0.83035904,1.2832822,1.4473847,1.3292309,0.9714873,0.43651286,0.12471796,0.15425642,0.27241027,0.3052308,0.14769232,0.23302566,0.128,0.029538464,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.049230773,0.23958977,0.13456412,0.2231795,0.42338464,0.69251287,1.020718,1.5589745,1.9987694,2.100513,2.284308,3.626667,4.4767184,4.3618464,3.9647183,3.5938463,3.190154,3.436308,4.394667,5.5762057,6.363898,6.012718,5.904411,7.3419495,8.487385,8.805744,9.061745,9.31118,9.019077,7.821129,6.2030773,5.5007186,6.436103,7.4797955,7.532308,6.5772314,5.720616,4.7589746,4.161641,3.751385,3.2065644,2.0611284,1.9331284,1.8937438,1.8838975,1.9922053,2.4713848,3.6890259,4.128821,3.8498464,3.367385,3.6726158,4.1189747,4.1485133,3.570872,2.7536411,2.6420515,1.4145643,1.2471796,1.9364104,3.0851285,4.1025643,6.163693,5.83877,4.788513,3.9122055,3.3608208,2.5238976,2.1464617,1.785436,1.3292309,1.0010257,2.294154,5.481026,9.892103,13.925745,15.07118,16.347898,14.933334,12.73436,11.812103,14.372104,15.0777445,11.195078,7.9852314,7.4174366,8.15918,7.8802056,8.277334,8.083693,6.954667,5.4547696,4.8672824,4.0336413,3.190154,2.5042052,2.0644104,1.5195899,2.8225644,2.8947694,1.6246156,1.8871796,1.5622566,1.3653334,1.1257436,0.8336411,0.6695385,0.43323082,0.26256412,0.27241027,0.40697438,0.4135385,0.21989745,0.31507695,0.5218462,0.7778462,1.1355898,1.4309745,1.4998976,1.5130258,1.4703591,1.2012309,0.98133343,1.3587693,1.7526156,2.0873847,2.8127182,3.1737437,2.7503593,2.281026,1.9790771,1.5327181,0.98461545,0.65969235,0.6629744,0.9124103,1.1388719,1.0699488,0.77456415,0.71548724,0.86646163,0.7253334,0.5316923,0.23958977,0.06235898,0.032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.009846155,0.009846155,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.02297436,0.026256412,0.013128206,0.04266667,0.128,0.21661541,0.25271797,0.18707694,0.2855385,0.40369233,0.39056414,0.25271797,0.128,0.28882053,0.43651286,0.49230772,0.42994875,0.26584616,0.15097436,0.17723078,0.2297436,0.21333335,0.06235898,0.059076928,0.04594872,0.02297436,0.0032820515,0.0,0.0,0.0,0.013128206,0.036102567,0.036102567,0.006564103,0.0032820515,0.0032820515,0.0,0.0,0.0,0.006564103,0.013128206,0.04266667,0.13784617,0.049230773,0.03938462,0.052512825,0.06564103,0.072205134,0.032820515,0.02297436,0.029538464,0.04266667,0.055794876,0.098461546,0.10502565,0.108307704,0.1148718,0.1148718,0.1148718,0.108307704,0.101743594,0.11158975,0.13128206,0.13784617,0.17066668,0.20348719,0.23958977,0.29210258,0.33476925,0.3708718,0.39712822,0.40697438,0.42994875,0.44307697,0.47261542,0.50543594,0.5284103,0.53825647,0.5284103,0.52512825,0.51856416,0.50543594,0.48246157,0.48574364,0.49887183,0.508718,0.51856416,0.53825647,0.5907693,0.7318975,1.0010257,1.463795,2.1956925,3.1376412,4.8738465,6.7840004,9.051898,12.681848,24.553028,37.48103,40.733543,32.92226,22.016,22.14072,20.693335,17.880617,14.454155,11.69395,11.047385,10.381129,9.337437,8.247795,8.113232,8.687591,8.490667,8.15918,8.073847,8.372514,7.8703594,6.7610264,5.61559,4.640821,3.6890259,2.2547693,1.079795,0.36102566,0.09189744,0.052512825,0.049230773,0.03938462,0.029538464,0.02297436,0.009846155,0.013128206,0.02297436,0.052512825,0.12471796,0.26256412,0.446359,0.5349744,0.5349744,0.5021539,0.5481026,0.46933338,0.512,0.7187693,1.0305642,1.3161026,1.7165129,2.422154,3.3345644,4.4964104,6.117744,9.015796,11.920411,14.844719,18.064411,22.130873,25.88554,29.942156,34.07426,38.1998,42.407387,48.351185,55.240208,63.91139,74.732315,87.627495,100.13539,107.881035,110.332726,107.4314,99.577446,89.29478,80.88944,74.19077,69.05437,65.35877,61.95857,58.354877,54.495182,50.65518,47.43549,43.506874,39.266464,34.330257,29.394054,26.240002,24.743387,22.14072,18.802874,15.360002,12.708103,10.125129,7.7456417,5.720616,4.076308,2.7273848,2.1956925,2.028308,2.0217438,2.038154,2.0053334,2.4910772,2.7109745,2.7306669,2.7602053,3.1507695,4.023795,4.588308,4.8114877,4.4898467,3.2722054,2.9078977,2.7076926,2.4320002,2.1398976,2.1956925,3.0162053,2.6847181,2.2514873,1.9200002,1.0666667,0.79425645,0.8336411,1.1290257,1.6344616,2.294154,2.15959,1.6771283,1.4572309,1.5261539,1.3489232,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.77456415,1.9593848,1.8313848,0.52512825,0.036102567,0.38400003,0.52512825,0.37415388,0.07548718,0.0,0.02297436,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.036102567,0.19364104,0.24943592,0.16410258,0.09189744,0.01969231,0.009846155,0.02297436,0.052512825,0.14769232,0.3117949,0.15097436,0.016410258,0.016410258,0.02297436,0.01969231,0.026256412,0.032820515,0.032820515,0.02297436,0.45620516,0.34133336,0.14112821,0.06564103,0.072205134,0.098461546,0.10502565,0.101743594,0.0951795,0.09189744,0.09189744,0.08533334,0.098461546,0.4266667,1.6180514,0.74830776,0.27897438,0.7187693,1.7362052,2.1431797,3.876103,4.8311796,5.1889234,5.4383593,6.370462,6.9710774,6.0783596,6.3179493,7.506052,6.633026,5.3070774,4.266667,4.141949,4.8114877,5.412103,4.6244106,4.0369234,4.5423594,5.989744,7.171283,6.4557953,4.601436,2.930872,1.9265642,1.2438976,0.7122052,0.60389745,0.5316923,0.41682056,0.47589746,0.84348726,0.7253334,0.4201026,0.14769232,0.036102567,0.029538464,0.016410258,0.016410258,0.029538464,0.04594872,0.059076928,0.036102567,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.26584616,0.79097444,1.3554872,1.5163078,1.8445129,2.1333334,2.4155898,2.9801028,3.117949,3.0949745,2.7963078,2.3893335,2.3171284,2.481231,2.5698464,2.231795,1.4966155,0.76800007,0.6235898,0.64000005,0.7581539,0.9682052,1.3423591,1.5064616,2.0939488,3.0785644,4.2305646,5.1364107,5.428513,6.1407185,6.0324106,5.041231,4.2535386,4.342154,4.571898,4.6244106,4.630975,5.182359,5.4974365,6.803693,8.92718,11.073642,11.844924,13.538463,15.169642,14.099693,10.597744,7.817847,7.177847,7.3025646,7.4404106,7.2664623,6.8955903,5.333334,4.4734364,4.007385,3.6857438,3.3444104,3.4100516,4.092718,5.2348723,6.3343596,6.554257,5.4974365,5.7829747,6.8988724,7.896616,7.384616,8.674462,8.923898,7.6734366,5.395693,3.4855387,3.8564105,3.8104618,3.515077,3.0260515,2.3105643,2.1234872,2.3663592,2.4681027,2.231795,1.8116925,1.6443079,1.522872,1.4473847,1.4572309,1.6344616,1.8543591,1.975795,1.9626669,1.6410258,0.69251287,0.26912823,0.2231795,0.24943592,0.18707694,0.01969231,0.15425642,0.07548718,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.032820515,0.14769232,0.39056414,0.15425642,0.19692309,0.3446154,0.5284103,0.761436,1.2865642,1.9298463,2.3466668,2.6518977,3.4166157,4.204308,4.7950773,5.4186673,5.586052,4.092718,5.037949,6.491898,7.460103,7.427283,6.377026,6.5345645,7.680001,8.3364105,8.234667,8.316719,7.2861543,6.619898,5.910975,5.1232824,4.588308,4.9493337,5.8256416,5.8453336,4.8672824,3.9745643,4.164923,4.128821,3.9089234,3.43959,2.553436,2.8225644,2.7667694,2.8291285,3.1770258,3.6857438,4.056616,3.7185643,4.073026,5.2644105,6.193231,6.419693,5.733744,4.352,2.937436,2.605949,1.5786668,1.5524104,1.9626669,2.4385643,2.7963078,4.210872,4.1813335,4.2272825,4.6572313,4.5817437,3.879385,3.817026,2.9636924,1.6180514,1.8051283,4.598154,7.653744,9.872411,10.722463,10.230155,10.003693,10.607591,11.257437,12.097642,14.191591,14.7790785,11.85477,10.075898,10.325335,9.711591,10.236719,11.290257,11.933539,11.191795,8.090257,6.1013336,4.348718,3.131077,2.5271797,2.3827693,2.6190772,4.3684106,4.535795,2.9669745,2.4648206,1.8576412,1.3850257,0.99774367,0.71548724,0.6071795,0.38728207,0.37415388,0.4397949,0.5677949,0.8172308,0.636718,0.8795898,1.2307693,1.467077,1.4572309,2.041436,2.5042052,2.9636924,3.318154,3.239385,3.0949745,3.436308,3.5544617,3.4067695,3.620103,3.626667,3.1770258,2.612513,1.9692309,0.9714873,0.90256417,0.73517954,0.764718,1.0732309,1.5589745,1.148718,0.88287187,0.75487185,0.67610264,0.47589746,0.27241027,0.09189744,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.009846155,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.07876924,0.14112821,0.15097436,0.1148718,0.098461546,0.30851284,0.4135385,0.446359,0.41025645,0.30851284,0.20676924,0.24615386,0.2986667,0.26584616,0.072205134,0.108307704,0.0951795,0.06564103,0.03938462,0.02297436,0.01969231,0.009846155,0.006564103,0.009846155,0.01969231,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.006564103,0.013128206,0.04266667,0.13784617,0.059076928,0.07876924,0.0951795,0.09189744,0.14769232,0.052512825,0.02297436,0.03938462,0.06564103,0.049230773,0.072205134,0.09189744,0.0951795,0.0951795,0.10502565,0.118153855,0.12143591,0.118153855,0.12143591,0.13784617,0.15425642,0.17394873,0.19364104,0.2231795,0.29210258,0.32820517,0.36102566,0.39384618,0.41682056,0.42338464,0.4266667,0.4397949,0.46276927,0.48902568,0.51856416,0.5349744,0.5415385,0.5481026,0.5546667,0.5481026,0.5546667,0.574359,0.60389745,0.636718,0.67282057,0.76800007,0.9353847,1.2832822,1.8674873,2.674872,4.2830772,6.7840004,8.982975,11.503591,16.777847,28.077951,36.772106,36.276516,27.51672,18.950565,16.86318,15.376411,14.168616,12.865642,11.040821,9.544206,9.147078,9.153642,9.143796,8.973129,8.3823595,7.1483083,5.7042055,4.673641,4.903385,4.778667,4.716308,4.857436,4.9460516,4.3290257,2.605949,1.1618463,0.36102566,0.18379489,0.2297436,0.15753847,0.08533334,0.04266667,0.026256412,0.016410258,0.016410258,0.016410258,0.029538464,0.07548718,0.17723078,0.3446154,0.4397949,0.46276927,0.4594872,0.52512825,0.4594872,0.4201026,0.47261542,0.62030774,0.79097444,0.9747693,1.2209232,1.4900514,1.8609232,2.5238976,4.2568207,6.009436,7.9524107,10.368001,13.653335,17.178257,21.202053,25.600002,30.175182,34.6519,39.811287,44.28144,48.370876,53.169235,60.557133,72.7237,86.009445,98.33026,107.15898,109.5516,102.649445,93.63693,84.8279,77.78134,73.31119,69.76,66.16616,62.57231,59.313236,57.01908,54.13416,51.14421,46.588722,40.68103,35.27877,32.850056,30.309746,26.945642,22.994053,19.652925,16.239592,13.138052,10.509129,8.306872,6.2752824,5.0543594,4.322462,3.9548721,3.7152824,3.249231,3.7940516,4.269949,4.5029745,4.522667,4.588308,5.037949,5.425231,5.5171285,5.228308,4.6211286,4.516103,4.2568207,3.692308,3.05559,2.9735386,3.3476925,3.3312824,3.1770258,2.7864618,1.6935385,1.2996924,1.2012309,1.273436,1.4834872,1.8970258,2.356513,2.156308,1.8576412,1.7099489,1.654154,0.0,0.0,0.0,0.0,0.0,0.0,0.128,0.108307704,0.049230773,0.02297436,0.072205134,0.7811283,0.73517954,0.42994875,0.15753847,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.006564103,0.0032820515,0.0032820515,0.006564103,0.013128206,0.02297436,0.049230773,0.108307704,0.09189744,0.055794876,0.04594872,0.1148718,0.3249231,0.6629744,0.4660513,0.17723078,0.029538464,0.04594872,0.009846155,0.016410258,0.02297436,0.013128206,0.013128206,0.013128206,0.029538464,0.03938462,0.03938462,0.04266667,0.06235898,0.06235898,0.055794876,0.049230773,0.059076928,0.12143591,0.13784617,0.22646156,0.90584624,3.1081028,1.6410258,0.955077,2.166154,4.1550775,3.5544617,7.1515903,6.5247183,4.9460516,5.0051284,8.579283,9.386667,7.2205133,6.5805135,7.8539495,7.315693,6.5378466,5.8190775,5.21518,5.0116925,5.7107697,4.1780515,2.993231,2.9735386,3.6824617,3.4297438,2.412308,1.5819489,0.98133343,0.5513847,0.12471796,0.10502565,0.28882053,0.29210258,0.0951795,0.036102567,0.026256412,0.016410258,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.03938462,0.23302566,0.65641034,1.3095386,1.1782565,1.1815386,1.4244103,1.7460514,1.6804104,1.9823592,2.605949,3.0654361,3.0358977,2.356513,2.0250258,2.1366155,2.100513,1.6968206,1.0469744,0.9353847,0.96492314,1.0469744,1.0896411,1.0010257,1.1618463,1.9528207,3.117949,4.332308,5.211898,5.028103,5.546667,5.7140517,5.149539,4.1813335,4.1550775,4.5423594,4.95918,5.395693,6.2063594,6.87918,8.362667,11.434668,15.24513,17.299694,18.632206,17.900309,14.562463,9.82318,6.636308,5.3366156,5.097026,5.7042055,6.413129,5.937231,4.4800005,3.5413337,3.0523078,2.802872,2.4516926,2.4484105,2.9243078,4.0369234,5.2676926,5.421949,4.630975,4.352,5.730462,7.765334,7.315693,8.5891285,7.5520005,6.0619493,4.962462,4.082872,4.9099493,5.546667,5.467898,4.7294364,3.9548721,2.8422565,2.2711797,2.0250258,1.8937438,1.6771283,1.6869745,1.785436,2.0250258,2.3729234,2.7011285,2.8488207,2.7470772,2.3794873,1.7394873,0.79425645,0.4004103,0.3511795,0.36102566,0.2855385,0.1148718,0.098461546,0.04266667,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.09189744,0.29210258,0.5349744,0.25928208,0.27241027,0.49887183,0.892718,1.404718,1.6640002,2.1070771,2.986667,4.023795,4.4110775,5.2053337,6.7117953,8.264206,8.900924,7.3682055,8.385642,9.580308,9.045334,7.020308,5.8880005,7.276308,7.9163084,7.79159,7.4043083,7.765334,6.1078978,5.8420515,6.4557953,7.0859494,6.498462,5.041231,4.378257,3.9975388,3.515077,2.674872,3.751385,4.6900516,5.293949,5.297231,4.3651285,5.362872,5.3070774,4.9920006,4.8804107,5.097026,4.4800005,3.9680004,5.6287184,8.52677,8.726975,7.939283,6.6034875,4.785231,3.1573336,2.993231,2.6486156,2.044718,1.8412309,2.0118976,1.8248206,2.3171284,3.1770258,4.716308,6.2555904,6.1374364,5.543385,5.3858466,3.9844105,2.1956925,3.4166157,7.171283,8.986258,8.41518,6.301539,4.778667,4.059898,7.2172313,10.121847,10.902975,9.95118,13.184001,13.072412,13.177437,13.705847,11.510155,13.83713,14.546052,15.1466675,14.923489,10.912822,7.4108725,4.594872,3.2164104,3.2853336,4.086154,5.4580517,5.3103595,4.706462,3.9351797,2.5009232,1.910154,1.5556924,1.3489232,1.2603078,1.3259488,0.88287187,0.78769237,0.65641034,0.58420515,1.1552821,1.404718,2.0545642,2.665026,2.9472823,2.7602053,4.1911798,5.353026,6.3868723,7.0990777,6.954667,6.5444107,6.0291286,5.208616,4.210872,3.4855387,3.370667,3.5905645,3.3509746,2.3762052,0.90584624,1.2668719,0.9878975,0.7778462,0.9353847,1.3718976,0.82379496,0.7975385,0.86317956,0.72861546,0.256,0.052512825,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.013128206,0.006564103,0.009846155,0.049230773,0.14769232,0.21661541,0.28882053,0.34133336,0.318359,0.23302566,0.23302566,0.2231795,0.18051283,0.1148718,0.17066668,0.14769232,0.108307704,0.07876924,0.049230773,0.03938462,0.02297436,0.013128206,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.02297436,0.101743594,0.12143591,0.098461546,0.18379489,0.11158975,0.098461546,0.12143591,0.128,0.03938462,0.09189744,0.15753847,0.15097436,0.08533334,0.08861539,0.12143591,0.13456412,0.13784617,0.13784617,0.14441027,0.16410258,0.17723078,0.190359,0.2231795,0.3117949,0.34789747,0.37743592,0.40697438,0.42994875,0.4266667,0.4201026,0.41025645,0.4135385,0.42994875,0.4594872,0.4955898,0.51856416,0.5415385,0.5677949,0.5973334,0.62030774,0.6695385,0.7318975,0.7975385,0.8533334,1.0305642,1.273436,1.7526156,2.4943593,3.3608208,5.8978467,8.992821,11.762873,15.415796,23.263182,26.072617,24.84513,21.572926,18.146463,16.357744,15.254975,14.785643,14.434463,13.617231,11.67754,9.426052,8.891078,9.865847,11.451077,12.048411,11.336206,9.885539,7.781744,6.048821,6.665847,6.675693,5.8912826,5.5105643,5.5958977,5.0904617,2.6223593,0.9878975,0.27569234,0.256,0.3708718,0.24943592,0.128,0.052512825,0.026256412,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.026256412,0.036102567,0.04266667,0.052512825,0.08861539,0.17723078,0.23958977,0.17394873,0.13456412,0.17394873,0.25271797,0.3314872,0.44307697,0.5973334,0.827077,1.2242053,1.9790771,2.5961027,3.6332312,5.3169236,7.568411,9.728001,12.806565,17.027283,22.022566,26.847181,32.082054,37.569645,42.436928,46.37539,49.631184,53.35303,60.491493,71.3879,84.854164,98.18585,101.983185,100.60144,95.86216,89.26852,81.99221,75.91385,71.74236,68.864006,66.79959,65.21764,62.66421,61.06585,58.29252,53.395695,46.63139,41.81662,38.649437,35.656208,32.07549,27.85149,23.522463,19.639797,16.308514,13.4629755,10.8537445,9.117539,7.8670774,7.1122055,6.4590774,5.106872,5.211898,5.7403083,6.235898,6.370462,5.933949,5.717334,5.674667,5.7665644,5.98318,6.3540516,6.432821,5.920821,5.0510774,4.1911798,3.8367183,3.8400004,3.9089234,3.7185643,3.2295387,2.7044106,2.3827693,2.1497438,2.028308,2.0053334,2.041436,2.5074873,2.612513,2.3138463,1.9232821,2.100513,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.072205134,0.30194873,0.6071795,0.6892308,0.029538464,0.006564103,0.0,0.0,0.0,0.0,0.0,0.026256412,0.032820515,0.016410258,0.016410258,0.03938462,0.06564103,0.11158975,0.24287182,0.5481026,0.45292312,0.27241027,0.101743594,0.032820515,0.16738462,0.6301539,1.142154,0.86646163,0.08205129,0.16738462,0.032820515,0.04594872,0.04594872,0.0,0.0,0.013128206,0.016410258,0.016410258,0.01969231,0.029538464,0.029538464,0.03938462,0.026256412,0.02297436,0.108307704,0.42338464,0.57764107,0.9419488,1.2274873,0.4594872,0.94523084,1.9922053,3.7087183,5.1298466,4.2272825,5.5072823,5.408821,3.8498464,1.9626669,2.0611284,2.8291285,4.5029745,5.041231,3.9089234,2.0906668,3.629949,3.2065644,2.2908719,2.1825643,4.013949,2.4615386,0.98461545,0.24615386,0.21989745,0.18379489,0.21989745,0.35774362,0.40697438,0.29538465,0.07548718,0.026256412,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02297436,0.19692309,0.21333335,0.08861539,0.13784617,0.3708718,0.2986667,0.40369233,0.7417436,0.9616411,1.2898463,1.9495386,4.07959,5.9930263,3.1737437,0.8795898,0.46933338,0.6465641,0.72861546,0.65641034,0.98461545,1.3522053,1.585231,1.5392822,1.0994873,0.9288206,1.5261539,2.7536411,4.309334,5.737026,3.636513,2.7634873,2.4910772,2.484513,2.7175386,3.6069746,3.892513,4.1091285,4.827898,6.6822567,7.8441033,9.396514,14.024206,20.266668,22.537848,22.951385,19.557745,14.168616,8.956718,6.4557953,4.5390773,3.318154,3.255795,3.8400004,3.570872,2.7634873,2.1136413,1.8149745,1.7920002,1.6935385,1.6804104,1.6771283,1.719795,1.9068719,2.3958976,2.9210258,3.4166157,4.138667,5.618872,8.681026,7.8769236,7.565129,7.4371285,6.803693,4.6080003,4.7425647,5.5991797,6.6494365,7.250052,6.6527185,4.2601027,2.9013336,2.425436,2.5206156,2.7175386,2.7634873,2.8422565,2.674872,2.2744617,1.9068719,1.9200002,1.6213335,1.1618463,0.7450257,0.6104616,0.40369233,0.37743592,0.37743592,0.36102566,0.39712822,0.26256412,0.108307704,0.01969231,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.12143591,0.3249231,0.4135385,0.4594872,0.35446155,0.6235898,1.5622566,3.2361028,3.1606157,3.2886157,4.8082056,7.3386674,8.92718,7.240206,6.2162056,7.6996927,10.587898,10.834052,11.687386,13.74195,13.259488,10.476309,9.596719,9.852718,9.258667,9.370257,10.440206,11.428103,9.632821,8.674462,8.697436,8.963283,7.827693,4.9362054,3.314872,2.7109745,2.8225644,3.31159,4.4964104,4.7622566,4.7524104,5.097026,6.439385,7.574975,7.6931286,6.7544622,6.0849237,8.392206,8.635077,7.634052,7.5388722,8.507077,8.726975,6.2490263,4.2929235,2.9440002,2.1891284,1.9068719,2.028308,1.785436,1.5360001,1.5556924,2.044718,2.2022567,2.865231,3.9942567,5.221744,5.8453336,6.1505647,4.450462,3.4494362,4.322462,6.7150774,8.093539,7.7423596,5.7632823,3.3017437,2.5337439,4.3651285,7.6964107,10.125129,10.978462,11.306667,13.748514,13.341539,11.109744,9.291488,11.352616,17.51631,18.07754,15.448617,11.290257,6.5312824,4.210872,3.2656412,4.1025643,6.3310776,8.772923,10.801231,6.803693,3.1540515,2.097231,1.7558975,2.3269746,2.8914874,3.0030773,2.6945643,2.487795,2.0217438,1.5786668,1.1881026,1.0338463,1.4506668,2.3040001,3.7349746,5.3234878,6.7150774,7.643898,9.757539,11.30995,12.724514,13.252924,10.971898,8.822155,7.131898,5.5926156,4.3749747,4.1189747,4.4242053,3.9876926,3.3772311,2.809436,2.1530259,1.9922053,1.6607181,1.2832822,1.0568206,1.2504616,0.8467693,0.4266667,0.16410258,0.072205134,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.02297436,0.036102567,0.06235898,0.13456412,0.17066668,0.15753847,0.10502565,0.029538464,0.01969231,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.013128206,0.08861539,0.19364104,0.256,0.18379489,0.318359,0.45292312,0.4397949,0.27241027,0.07548718,0.380718,0.5021539,0.3708718,0.12471796,0.13784617,0.15097436,0.14441027,0.13784617,0.14441027,0.16738462,0.16738462,0.17723078,0.19692309,0.22646156,0.27569234,0.3117949,0.34789747,0.3708718,0.37743592,0.36758977,0.37743592,0.380718,0.38728207,0.4004103,0.4135385,0.43651286,0.47917953,0.5218462,0.56123084,0.6104616,0.67282057,0.761436,0.8566154,0.9517949,1.0371283,1.2340513,1.6836925,2.356513,3.1770258,4.0434875,6.0816417,9.009232,12.652308,17.243898,23.42072,24.385643,22.30154,21.464617,22.81354,23.926155,19.872822,15.041642,12.363488,12.140308,12.0549755,11.296822,11.464206,12.2157955,14.01436,18.12677,16.955078,13.128206,8.825437,6.2490263,7.6307697,8.717129,7.3583593,6.052103,5.4941545,4.578462,1.7099489,0.47917953,0.0951795,0.029538464,0.029538464,0.04266667,0.036102567,0.02297436,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.02297436,0.029538464,0.029538464,0.029538464,0.04266667,0.04594872,0.04594872,0.04594872,0.04594872,0.04594872,0.072205134,0.12143591,0.2100513,0.380718,0.88287187,1.1093334,1.2537436,1.6114873,2.5632823,5.0543594,7.250052,10.407386,14.578873,18.632206,22.344208,27.024412,32.298668,37.789543,43.136,48.42339,51.997543,54.291695,57.75754,66.852104,79.92452,92.93457,100.76883,100.191185,89.82647,82.29744,79.645546,77.44657,74.14154,71.03016,69.73375,67.32472,64.84677,62.9038,61.643494,55.84739,49.618053,44.90503,41.46544,36.850876,32.626873,27.969643,23.332104,19.193438,16.065641,14.027489,12.977232,12.422565,11.369026,8.329846,7.574975,7.706257,8.211693,8.385642,7.325539,6.7872825,6.2687182,6.2063594,6.672411,7.3550773,7.1220517,6.6625648,6.1013336,5.5696416,5.2020516,5.1167183,4.857436,4.585026,4.4373336,4.5456414,4.315898,3.817026,3.2984617,2.993231,3.1277952,3.0654361,3.062154,3.1343591,3.2820516,3.4789746,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.118153855,0.5973334,0.74830776,0.58092314,0.42338464,0.32820517,0.07876924,0.016410258,0.02297436,0.098461546,0.17723078,0.098461546,0.01969231,0.006564103,0.006564103,0.0032820515,0.0032820515,0.63343596,0.36102566,0.059076928,0.049230773,0.108307704,0.09189744,0.055794876,0.01969231,0.006564103,0.032820515,0.128,0.2297436,0.25271797,0.26584616,0.49887183,0.42994875,0.24943592,0.08205129,0.0,0.0,0.0032820515,0.0032820515,0.17066668,0.33476925,0.006564103,0.25928208,0.13456412,0.47917953,0.955077,0.032820515,0.34133336,1.332513,1.4276924,0.62030774,0.4955898,1.5983591,3.0982566,4.4242053,5.218462,5.349744,6.5444107,5.080616,3.5183592,2.7437952,1.9626669,2.097231,2.2350771,1.9331284,1.2800001,0.90584624,1.3128207,0.95835906,0.54482055,0.47261542,0.8402052,0.51856416,0.2297436,0.08205129,0.06564103,0.049230773,0.04594872,0.072205134,0.09189744,0.08205129,0.026256412,0.006564103,0.009846155,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.04594872,0.06564103,0.08533334,0.2231795,0.6498462,1.0010257,1.1881026,1.1552821,0.88943595,0.8467693,0.9288206,1.3554872,1.8248206,1.5261539,0.5021539,0.190359,0.17066668,0.20020515,0.20348719,0.8566154,1.4276924,1.5031796,1.1684103,1.0010257,0.8402052,1.1782565,2.1398976,3.3476925,3.9056413,2.8717952,1.8838975,1.3981539,1.4736412,1.7624617,2.3236926,2.878359,3.5183592,4.394667,5.730462,7.13518,9.196308,12.937847,16.794258,16.603899,15.908104,12.859077,9.787078,8.041026,7.9786673,6.8463597,5.2053337,3.8104618,3.058872,2.9965131,2.7273848,2.4976413,2.4516926,2.4352822,1.9856411,1.5458462,1.2800001,1.0896411,1.0404103,1.3817437,1.9462565,2.4320002,3.5478978,6.009436,10.538668,11.382154,10.390975,8.795898,6.882462,4.023795,3.308308,4.309334,5.910975,7.026872,6.6034875,4.6112823,3.9909747,4.417641,5.0215387,4.388103,2.993231,2.1070771,1.4966155,1.0436924,0.73517954,0.6301539,0.6170257,0.57764107,0.47589746,0.34133336,0.35774362,0.33805132,0.31507695,0.3052308,0.3117949,0.21661541,0.08861539,0.009846155,0.0032820515,0.013128206,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.052512825,0.18707694,0.4004103,0.15425642,0.15097436,0.5481026,1.6213335,3.7710772,4.0992823,4.8607183,5.654975,6.5870776,8.2904625,9.291488,9.186462,9.238976,10.056206,11.579078,13.154463,14.234258,12.813129,10.308924,11.539693,11.687386,11.782565,12.317539,12.320822,9.366975,8.470975,7.381334,5.907693,4.414359,3.8367183,3.8137438,4.1846156,4.519385,4.4865646,3.8596926,4.4767184,4.962462,5.152821,5.7042055,8.109949,9.120821,8.490667,7.968821,8.070564,8.064001,6.482052,6.6428723,6.9776416,6.6002054,5.297231,4.4307694,3.4264617,2.5042052,2.0873847,2.8225644,2.7208207,2.156308,1.910154,2.1825643,2.5928206,2.9571285,3.56759,3.8629746,4.073026,5.2348723,6.0258465,4.926359,4.670359,5.6352825,5.8092313,6.5345645,5.405539,3.3312824,2.540308,6.5870776,9.82318,10.459898,8.884514,6.918565,7.8145647,13.29559,14.539488,13.5778475,11.546257,8.726975,9.396514,9.688616,8.976411,7.253334,5.139693,4.20759,4.2141542,4.7589746,5.356308,5.4547696,7.890052,6.157129,3.9417439,2.9243078,2.7667694,2.8127182,2.7798977,2.7175386,2.605949,2.3401027,2.0808206,1.8838975,2.484513,3.9581542,5.720616,6.770872,9.042052,11.766154,14.102976,15.140103,16.548103,16.190361,14.211283,11.35918,8.969847,7.768616,6.042257,4.529231,3.5347695,2.937436,3.8465643,3.4297438,2.5074873,1.6377437,1.1257436,1.0075898,0.9911796,0.7975385,0.508718,0.5677949,0.36102566,0.16410258,0.049230773,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.006564103,0.013128206,0.026256412,0.04266667,0.052512825,0.049230773,0.006564103,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.02297436,0.06235898,0.036102567,0.006564103,0.0,0.0032820515,0.0,0.0,0.0,0.006564103,0.036102567,0.108307704,0.15425642,0.2231795,0.29538465,0.28225642,0.11158975,0.44964105,0.446359,0.055794876,0.016410258,0.07548718,0.1148718,0.14769232,0.16410258,0.13784617,0.15097436,0.15753847,0.15753847,0.15097436,0.15425642,0.15425642,0.16410258,0.17394873,0.18707694,0.22646156,0.27241027,0.3117949,0.3446154,0.36758977,0.36758977,0.34789747,0.36102566,0.38400003,0.40697438,0.4004103,0.44307697,0.48246157,0.512,0.5316923,0.56123084,0.6826667,0.81394875,0.9616411,1.1191796,1.2931283,1.6738462,2.297436,3.0851285,4.1222568,5.6418467,8.247795,12.888617,19.498669,26.74872,32.07549,27.736618,21.838772,18.399181,17.703386,16.28554,14.017642,12.498053,12.166565,12.632616,12.665437,13.2562065,14.185027,16.088617,19.075283,22.728207,24.224823,21.700924,16.879591,12.57354,12.681848,14.053744,12.156719,9.947898,8.362667,6.3343596,2.0217438,0.47589746,0.128,0.06564103,0.01969231,0.009846155,0.006564103,0.009846155,0.016410258,0.016410258,0.016410258,0.006564103,0.0032820515,0.006564103,0.016410258,0.006564103,0.013128206,0.01969231,0.01969231,0.01969231,0.01969231,0.029538464,0.032820515,0.032820515,0.032820515,0.032820515,0.04594872,0.06564103,0.10502565,0.19692309,0.56123084,0.77456415,0.98133343,1.2996924,1.8313848,3.4231799,5.1889234,7.5946674,10.679795,14.076719,16.843489,19.652925,23.138464,27.615181,33.089645,38.728207,43.605335,47.241848,50.11693,53.664825,59.805542,69.034676,79.34032,88.65806,94.84473,94.20801,89.00924,83.02277,78.43118,75.82523,74.719185,73.1438,71.47652,69.90113,68.42093,66.3237,62.80534,58.9719,55.03672,50.326977,44.862362,38.915283,32.423386,26.213745,22.025848,20.6999,19.570873,18.20554,16.128002,12.822975,11.293539,10.735591,10.617436,10.489437,9.974154,8.946873,8.100103,7.8408213,8.297027,9.330873,9.636104,9.7214365,9.82318,9.91836,9.708308,9.094564,8.740103,8.480822,8.283898,8.257642,8.231385,7.9885135,7.7948723,7.768616,7.9130263,7.8112826,7.643898,7.456821,7.259898,7.00718,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.098461546,0.2986667,0.49887183,1.214359,1.1946667,0.8566154,0.55794877,0.6301539,0.18379489,0.42338464,0.5349744,0.3117949,0.18707694,0.5513847,0.3052308,0.06564103,0.029538464,0.009846155,0.31507695,0.17394873,0.03938462,0.052512825,0.04594872,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.03938462,0.12471796,0.23302566,0.21333335,0.118153855,0.036102567,0.0,0.0,0.013128206,0.13784617,0.26584616,0.29538465,0.13784617,0.23630771,0.2231795,0.4955898,0.75487185,0.016410258,0.28225642,1.5688206,2.1398976,1.5524104,0.65969235,1.0075898,1.913436,3.5478978,5.5204105,6.8562055,11.332924,7.141744,3.692308,3.5216413,2.284308,1.0962052,0.8041026,0.5973334,0.2986667,0.3446154,0.32164106,0.16738462,0.049230773,0.01969231,0.01969231,0.013128206,0.016410258,0.016410258,0.009846155,0.006564103,0.0,0.0,0.0032820515,0.009846155,0.006564103,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.009846155,0.01969231,0.026256412,0.04266667,0.098461546,0.34789747,0.8041026,1.086359,1.014154,0.5874872,0.48902568,0.77128214,1.3193847,2.1267693,3.2918978,0.9944616,0.18379489,0.118153855,0.2100513,0.036102567,0.32820517,0.57764107,0.6104616,0.52512825,0.6826667,0.8533334,1.142154,1.6377437,2.1956925,2.4516926,1.9167181,1.1946667,0.8172308,0.92553854,1.2603078,1.9429746,2.6551797,3.2623591,3.820308,4.5587697,6.1407185,7.936001,10.505847,12.691693,11.61518,10.505847,8.51036,6.432821,5.159385,5.6418467,6.564103,6.2063594,5.467898,4.9427695,4.923077,4.6276927,4.1747694,4.096,4.1517954,3.3509746,2.0676925,1.3522053,0.9517949,0.8008206,1.0108719,1.5031796,2.2219489,3.892513,6.633026,9.96759,10.236719,8.339693,6.042257,4.1124105,2.3368206,2.5009232,3.7152824,5.031385,5.61559,4.768821,3.764513,3.5807183,3.9089234,4.128821,3.3247182,2.3269746,1.6836925,1.1749744,0.7515898,0.52512825,0.47917953,0.6301539,0.65969235,0.5021539,0.33805132,0.40369233,0.37743592,0.30194873,0.2231795,0.21661541,0.20348719,0.16082053,0.12143591,0.10502565,0.1148718,0.108307704,0.04266667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.07548718,0.2231795,0.26584616,0.58420515,1.1651284,2.4188719,5.179077,6.229334,7.200821,7.325539,7.506052,10.328616,13.459693,13.24636,12.530872,12.166565,11.024411,11.762873,12.84595,12.484924,11.2672825,12.153437,12.22236,13.236514,13.702565,12.570257,9.235693,8.694155,8.454565,6.882462,4.8016415,5.474462,6.2720003,6.1013336,5.737026,5.3891287,4.71959,5.152821,5.8486156,6.6133337,7.768616,10.151385,10.656821,9.580308,8.484103,8.057437,8.109949,7.066257,7.0859494,6.616616,5.218462,3.570872,3.4724104,3.2820516,2.9078977,2.6322052,3.1081028,2.9768207,2.1989746,1.785436,2.0906668,2.806154,3.0818465,3.05559,3.1474874,3.7448208,5.1922054,5.353026,5.3924108,5.805949,6.2129235,5.3727183,4.962462,4.0533338,4.082872,6.0028725,10.262975,12.950975,11.969642,8.103385,4.4767184,6.5312824,8.132924,8.874667,9.229129,8.887795,6.7807183,5.3037953,5.3005133,5.5958977,5.4941545,4.781949,3.8301542,3.1770258,2.8816411,2.934154,3.249231,5.0871797,4.709744,3.9154875,3.6726158,4.1091285,4.20759,3.8104618,3.6627696,3.8662567,3.8695388,3.7054362,4.391385,6.498462,9.462154,11.569232,13.466257,16.183796,18.274464,18.894772,17.818258,15.911386,13.909334,11.556104,9.045334,7.030154,5.8256416,4.598154,3.5511796,2.9210258,2.9702566,3.1442053,2.6223593,2.169436,1.8116925,0.81394875,0.49230772,0.5513847,0.48574364,0.2297436,0.15753847,0.0951795,0.03938462,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.013128206,0.0,0.0,0.0,0.006564103,0.013128206,0.0,0.006564103,0.026256412,0.02297436,0.0032820515,0.013128206,0.032820515,0.01969231,0.0032820515,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.026256412,0.11158975,0.13456412,0.17723078,0.21661541,0.12143591,0.02297436,0.18379489,0.18707694,0.006564103,0.0,0.006564103,0.02297436,0.06235898,0.10502565,0.09189744,0.11158975,0.14112821,0.15097436,0.14112821,0.13456412,0.14112821,0.14769232,0.15097436,0.15425642,0.17723078,0.21989745,0.256,0.29210258,0.3249231,0.33805132,0.32164106,0.3314872,0.36430773,0.40697438,0.42338464,0.47261542,0.512,0.53825647,0.5513847,0.57764107,0.702359,0.85005134,1.0436924,1.332513,1.7985642,2.605949,3.367385,4.519385,6.298257,8.717129,13.02318,18.609232,24.201847,28.665438,31.028515,23.443693,16.439796,13.380924,14.14236,15.123693,14.198155,14.158771,15.172924,16.777847,17.880617,17.253744,17.191385,18.107079,20.020514,22.534565,26.476309,27.733335,25.32431,20.736002,17.929848,17.575386,15.75713,11.9860525,7.3682055,4.578462,1.2865642,0.6826667,0.574359,0.15425642,0.006564103,0.0,0.0,0.0032820515,0.006564103,0.006564103,0.006564103,0.0032820515,0.0,0.0,0.006564103,0.0,0.009846155,0.013128206,0.006564103,0.016410258,0.016410258,0.01969231,0.02297436,0.02297436,0.02297436,0.02297436,0.029538464,0.04266667,0.059076928,0.08861539,0.256,0.49887183,0.8763078,1.3292309,1.6836925,2.8324106,4.5456414,6.6822567,9.074872,11.556104,13.682873,15.67836,17.893745,20.617847,24.080412,29.321848,35.37067,41.06175,45.551594,48.32821,50.530464,55.000618,61.886364,70.79057,80.77457,88.32001,91.28042,90.94565,88.274055,83.89252,80.52185,78.27036,76.29457,74.233444,72.17231,70.74462,69.008415,67.42647,66.067696,64.597336,60.639183,55.315697,47.166363,37.392414,29.830566,28.691694,27.588924,25.498259,22.226053,18.395899,16.564514,15.097437,14.063591,13.266052,12.2387705,11.067078,10.151385,9.645949,9.636104,10.128411,10.801231,11.526565,12.658873,14.043899,15.0088215,15.192616,15.652103,16.219898,16.695797,16.840206,16.987898,16.347898,15.287796,14.152206,13.275898,12.819694,12.534155,12.2157955,11.733335,11.0375395,0.0,0.0,0.0,0.0,0.055794876,0.2855385,0.16082053,0.13784617,0.2855385,0.50543594,0.5546667,1.1060513,1.394872,1.1126155,0.5677949,0.67610264,0.22646156,0.47917953,0.5316923,0.22646156,0.13784617,0.5513847,0.31507695,0.068923086,0.032820515,0.02297436,0.009846155,0.0032820515,0.02297436,0.052512825,0.04594872,0.009846155,0.0,0.0,0.0,0.0,0.0,0.006564103,0.02297436,0.052512825,0.09189744,0.101743594,0.04266667,0.016410258,0.032820515,0.0,0.013128206,0.13784617,0.2231795,0.25928208,0.4004103,0.5349744,0.81394875,0.8598975,0.5481026,0.009846155,0.15425642,2.665026,3.7776413,2.5271797,0.7450257,1.5819489,1.2603078,2.0545642,4.6244106,8.004924,13.804309,7.8769236,2.9078977,2.7109745,2.231795,0.6235898,0.2986667,0.2297436,0.055794876,0.101743594,0.026256412,0.009846155,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.059076928,0.059076928,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.009846155,0.02297436,0.029538464,0.04266667,0.108307704,0.128,0.36102566,0.6859488,0.8730257,0.5677949,0.5677949,1.0075898,1.591795,2.281026,3.2820516,0.955077,0.19364104,0.14112821,0.20020515,0.04266667,0.009846155,0.0,0.01969231,0.098461546,0.3052308,0.6826667,1.1618463,1.5163078,1.6377437,1.5655385,1.332513,0.9747693,0.7089231,0.6892308,0.98461545,1.6672822,2.1530259,2.5042052,2.858667,3.4166157,5.9470773,7.9425645,9.288206,9.793642,9.186462,8.815591,7.778462,6.166975,4.6900516,4.6966157,5.9536414,6.5345645,6.636308,6.560821,6.7183595,6.2884107,5.7074876,5.648411,5.756718,4.644103,2.7142565,1.5819489,1.0404103,0.8960001,0.9747693,1.148718,1.7394873,3.249231,5.346462,6.8594875,6.157129,4.601436,3.1671798,2.297436,1.9035898,2.6354873,3.2754874,3.7907696,3.9089234,3.1409233,3.0654361,3.239385,3.3542566,3.2098465,2.7076926,2.5074873,2.0086155,1.3489232,0.75487185,0.5677949,0.6432821,0.75487185,0.7089231,0.512,0.380718,0.44307697,0.42994875,0.3511795,0.24943592,0.2231795,0.23630771,0.22646156,0.21333335,0.21661541,0.26912823,0.24287182,0.13784617,0.04266667,0.0032820515,0.013128206,0.026256412,0.013128206,0.0,0.0,0.0,0.16082053,0.08205129,0.0,0.08861539,0.43651286,0.8205129,1.8149745,2.6190772,3.7809234,7.1876926,9.826463,9.833026,8.746667,8.402052,10.935796,14.854566,15.31077,14.634667,13.479385,10.834052,11.040821,11.618463,11.54954,10.902975,10.8537445,10.072617,10.450052,10.755282,10.604308,10.466462,9.908514,9.193027,7.755488,6.3934364,7.256616,7.6077952,6.688821,5.3727183,4.5029745,4.9296412,5.175795,6.038975,7.430565,9.009232,10.174359,10.545232,10.112,9.074872,7.975385,7.6701546,6.547693,5.9470773,5.113436,3.948308,3.0326157,3.3903592,3.570872,3.3247182,2.9636924,3.3805132,3.0818465,2.4746668,2.3368206,3.0391798,4.562052,4.3290257,3.754667,3.8400004,4.571898,4.923077,4.312616,4.709744,5.218462,5.287385,4.71959,4.0303593,3.69559,5.1987696,8.539898,12.228924,15.698052,13.078976,8.333129,5.4547696,8.470975,7.8408213,7.030154,6.2720003,5.6385646,5.028103,3.43959,3.69559,4.3684106,4.9985647,6.1013336,4.1714873,2.9801028,2.5074873,2.7175386,3.5478978,4.519385,4.466872,4.457026,4.9985647,6.0324106,6.262154,5.618872,5.225026,5.435077,5.835488,6.685539,8.211693,11.021129,14.401642,16.298668,18.504206,20.470156,20.804924,19.006361,15.445334,12.06154,9.803488,8.077128,6.5969234,5.3760004,4.699898,3.7874875,2.8980515,2.4188719,2.8849232,2.5862565,1.7493335,1.394872,1.4178462,0.5874872,0.23630771,0.24287182,0.2297436,0.09189744,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.013128206,0.0,0.032820515,0.03938462,0.02297436,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.01969231,0.0032820515,0.013128206,0.08205129,0.19692309,0.32164106,0.51856416,0.512,0.3314872,0.0951795,0.006564103,0.006564103,0.013128206,0.016410258,0.013128206,0.013128206,0.013128206,0.016410258,0.029538464,0.04266667,0.049230773,0.07876924,0.118153855,0.13456412,0.12471796,0.1148718,0.118153855,0.12143591,0.12471796,0.128,0.14769232,0.18379489,0.21661541,0.24615386,0.26912823,0.28882053,0.28225642,0.29210258,0.3314872,0.38400003,0.42994875,0.49887183,0.55794877,0.60061544,0.6235898,0.636718,0.764718,0.8730257,1.2570257,1.8806155,2.3401027,2.9636924,4.4767184,6.3343596,8.467693,11.283693,15.875283,20.427488,23.446976,24.25436,22.997335,16.561232,11.293539,9.563898,11.523283,15.113848,14.749539,14.326155,15.346873,17.841232,20.358566,19.748104,19.5479,19.620104,20.059898,21.192207,23.322258,24.86154,23.860516,20.608002,17.64759,17.34236,15.356719,10.66995,4.850872,2.044718,0.702359,0.60389745,0.51856416,0.12471796,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.006564103,0.0032820515,0.009846155,0.009846155,0.009846155,0.013128206,0.013128206,0.009846155,0.013128206,0.01969231,0.029538464,0.03938462,0.04594872,0.09189744,0.28225642,0.6465641,1.0962052,1.4112822,2.3368206,4.092718,6.265436,8.461129,10.305642,11.733335,13.210258,14.588719,15.855591,17.115898,20.886976,25.924925,31.842464,37.858463,42.79139,46.5559,49.906876,53.300518,57.570465,63.917953,73.30134,82.34011,88.90421,91.77929,90.66011,87.75221,84.78852,81.86093,78.97929,76.06155,73.87241,72.126366,70.93826,70.45908,70.87919,70.65929,69.851906,64.79426,55.105644,43.664413,39.21067,36.850876,33.26359,28.054977,23.75549,21.48759,19.495386,17.746052,16.242872,15.0088215,13.896206,12.852514,11.96636,11.369026,11.227899,11.792411,12.583385,13.751796,15.169642,16.406975,17.19795,18.323694,19.442873,20.352001,20.978874,22.038977,21.809233,20.617847,19.026052,17.834667,17.765745,17.408,16.636719,15.573335,14.585437,0.0,0.0,0.0,0.0,0.1148718,0.574359,0.32164106,0.27897438,0.45292312,0.78769237,1.1684103,0.9353847,1.1684103,0.98461545,0.39056414,0.28225642,0.128,0.13128206,0.0951795,0.0,0.0,0.02297436,0.01969231,0.006564103,0.0032820515,0.02297436,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.049230773,0.10502565,0.18379489,0.21333335,0.108307704,0.055794876,0.068923086,0.0,0.0,0.0,0.07876924,0.26256412,0.52512825,0.8566154,1.3784616,1.2865642,0.574359,0.04594872,0.30851284,3.8728209,4.969026,2.6584618,0.8402052,3.4527183,1.9232821,1.1290257,3.3345644,8.185436,11.273847,5.9470773,1.404718,0.8598975,1.5163078,0.5973334,0.3314872,0.190359,0.009846155,0.0,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.118153855,0.118153855,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016410258,0.032820515,0.08205129,0.23302566,0.15097436,0.06235898,0.3511795,0.8205129,0.69907695,0.88615394,1.2209232,1.2865642,1.1618463,1.3850257,0.38400003,0.17066668,0.25271797,0.3511795,0.39384618,0.13128206,0.026256412,0.0,0.0032820515,0.02297436,0.30851284,0.9156924,1.3522053,1.3784616,1.0043077,1.017436,0.98461545,0.8369231,0.69579494,0.88615394,1.2931283,1.2800001,1.3062565,1.6410258,2.3696413,6.009436,8.766359,9.452309,8.684308,8.884514,9.517949,8.848411,7.6143594,6.416411,5.720616,5.504,5.933949,6.242462,6.3212314,6.7216415,6.3901544,5.979898,5.9503593,5.979898,4.969026,3.006359,1.7099489,1.1126155,0.99774367,0.90584624,0.69251287,0.8172308,1.5064616,2.4352822,2.7437952,1.8313848,2.034872,2.5698464,2.930872,2.868513,2.8947694,2.4615386,2.2678976,2.4451284,2.553436,3.1507695,3.511795,3.515077,3.2984617,3.239385,3.318154,2.5632823,1.5458462,0.74830776,0.574359,0.7581539,0.7318975,0.6432821,0.53825647,0.38400003,0.42338464,0.47261542,0.45620516,0.37415388,0.3117949,0.27569234,0.25928208,0.26584616,0.30851284,0.42338464,0.4135385,0.30194873,0.15753847,0.04594872,0.03938462,0.06235898,0.032820515,0.009846155,0.013128206,0.02297436,0.36102566,0.21661541,0.08533334,0.3249231,1.142154,1.6771283,3.0293336,3.7349746,4.4964104,8.178872,12.225642,10.935796,8.651488,8.169026,10.748719,13.633642,14.54277,13.824001,12.209231,10.817642,11.063796,10.384411,9.442462,8.661334,8.195283,6.6592827,5.7501545,6.193231,8.333129,12.12718,11.349334,9.07159,7.6767187,7.6767187,7.7259493,7.0957956,6.340924,4.969026,3.7448208,4.699898,4.857436,5.5204105,6.9382567,8.43159,8.372514,8.94359,9.626257,9.350565,7.9852314,6.340924,4.6276927,3.7710772,3.4822567,3.4855387,3.508513,3.8432825,3.9417439,3.5544617,3.1048207,3.6594875,3.2918978,3.570872,4.2962055,5.7501545,8.674462,7.6077952,6.49518,5.9602056,5.605744,4.013949,3.3411283,3.5413337,3.879385,4.197744,4.919795,5.5236926,5.1626673,6.170257,8.992821,12.173129,15.91795,12.484924,8.707283,8.231385,11.533129,12.064821,9.642668,6.3212314,3.8596926,3.692308,2.8882053,3.6463592,4.276513,5.0838976,8.3593855,5.179077,3.8367183,3.7382567,4.352,5.182359,6.0717955,6.11118,6.3606157,7.1909747,8.293744,8.576,7.965539,7.1089234,6.675693,7.3583593,9.895386,12.163283,14.890668,17.706669,19.157335,20.12554,19.748104,17.80513,14.404924,10.006975,7.857231,6.49518,5.362872,4.391385,3.9942567,4.3060517,3.3969233,2.349949,1.8379488,2.1267693,1.9232821,0.9124103,0.2855385,0.29210258,0.24287182,0.098461546,0.03938462,0.02297436,0.01969231,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.049230773,0.02297436,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.036102567,0.006564103,0.029538464,0.15753847,0.37743592,0.6268718,0.9156924,0.88615394,0.49230772,0.0032820515,0.016410258,0.016410258,0.01969231,0.02297436,0.026256412,0.032820515,0.01969231,0.013128206,0.016410258,0.029538464,0.036102567,0.072205134,0.101743594,0.11158975,0.10502565,0.108307704,0.098461546,0.098461546,0.10502565,0.108307704,0.13128206,0.16410258,0.19364104,0.2100513,0.2231795,0.23958977,0.23958977,0.256,0.28882053,0.33476925,0.39384618,0.48574364,0.58092314,0.7515898,0.9353847,0.9124103,0.97805136,0.96492314,1.6344616,2.7536411,3.1081028,3.1540515,5.5696416,7.9983597,9.885539,12.4685135,15.849027,18.130053,18.786463,17.362053,13.449847,10.771693,8.41518,7.6012316,8.94359,12.435693,12.491488,11.861334,13.049437,16.472616,20.489847,20.74913,19.961437,19.275488,19.288616,20.033642,18.212105,16.879591,15.507693,14.148924,13.453129,13.748514,10.893129,6.5247183,2.412308,0.4397949,0.5316923,0.2231795,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.013128206,0.0032820515,0.016410258,0.01969231,0.026256412,0.036102567,0.052512825,0.07548718,0.15097436,0.4266667,0.8336411,1.0765129,1.6738462,3.2361028,5.408821,7.7456417,9.741129,10.65354,11.572514,12.294565,12.658873,12.553847,14.060308,16.44636,20.499695,26.289232,33.158566,41.16677,46.98585,50.41231,52.194466,54.019287,58.525543,66.50093,75.697235,84.178055,90.29252,91.82524,90.240005,87.67673,85.008415,81.83467,78.50011,75.346054,72.42503,70.18996,69.490875,71.614365,75.60862,76.78359,72.56616,62.49026,53.805954,47.763695,40.71385,32.817234,28.071386,25.27836,23.095797,21.001848,19.055592,17.870771,16.827078,15.606155,14.395078,13.4400015,13.019898,13.170873,13.650052,14.053744,14.25395,14.404924,14.943181,16.006565,16.95836,17.732924,18.822565,21.090464,21.897848,21.444925,20.348719,19.626669,20.52595,20.338873,19.26236,17.85436,17.033848,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.006564103,0.41025645,1.2800001,2.3040001,2.0709746,1.2635899,0.8533334,0.9156924,0.6104616,0.14769232,0.013128206,0.0,0.0,0.0,0.013128206,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.049230773,0.12471796,0.101743594,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.36758977,0.4397949,0.19364104,0.2297436,1.5360001,2.3368206,2.300718,1.6804104,1.3259488,4.4767184,2.6354873,2.1858463,4.6933336,6.928411,4.450462,2.3762052,1.1355898,0.6629744,0.380718,0.08861539,0.016410258,0.009846155,0.0,0.0,0.013128206,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.02297436,0.036102567,0.06235898,0.049230773,0.036102567,0.23302566,0.4660513,0.19692309,0.69907695,1.0436924,1.020718,1.1290257,2.5928206,0.71548724,0.28225642,0.81066674,1.5655385,1.5425643,0.56451285,0.128,0.0,0.0,0.0,0.0,0.009846155,0.02297436,0.03938462,0.07548718,0.18707694,0.47917953,0.764718,0.95835906,1.0666667,1.2012309,0.9156924,0.6301539,0.67610264,1.2964103,4.1550775,7.194257,8.766359,8.687591,8.224821,7.9327188,6.8332314,5.979898,5.504,4.6244106,3.9286156,3.6791797,3.7284105,3.95159,4.2568207,4.4406157,4.210872,3.7710772,3.442872,3.6627696,2.550154,1.5327181,0.95835906,0.74830776,0.380718,0.19692309,0.19692309,0.36430773,0.6071795,0.7778462,0.8992821,3.1638978,5.0674877,5.1889234,3.1737437,1.3423591,0.74830776,0.8336411,1.4178462,2.7011285,3.9351797,3.9318976,3.4658465,3.0949745,3.1442053,2.5928206,1.8510771,1.1815386,0.7581539,0.67282057,0.90256417,0.9419488,1.0043077,0.9714873,0.39712822,0.34789747,0.5284103,0.5874872,0.45620516,0.33476925,0.24943592,0.3117949,0.36102566,0.38728207,0.5349744,0.6695385,0.53825647,0.35446155,0.2100513,0.07548718,0.03938462,0.049230773,0.055794876,0.06235898,0.12143591,0.19692309,0.27897438,0.42994875,0.8730257,1.9823592,2.5206156,2.4352822,2.0086155,2.3072822,5.1889234,7.788308,7.3386674,5.5893335,6.2818465,15.16636,14.995693,12.343796,9.596719,8.254359,8.92718,8.4512825,6.774154,5.786257,5.861744,5.874872,6.2162056,6.961231,8.224821,10.151385,12.908309,11.894155,9.728001,8.805744,9.363693,9.458873,8.008205,8.2215395,8.612103,7.9819493,5.431795,6.163693,5.6254363,5.4974365,6.3245134,7.506052,7.8112826,8.064001,7.7325134,6.488616,4.1813335,4.5456414,4.6572313,5.097026,5.622154,5.156103,4.1452312,3.9548721,4.0336413,3.9384618,3.3411283,3.8432825,6.0816417,7.962257,9.908514,14.87754,12.947693,10.515693,7.574975,4.57518,2.425436,3.121231,4.3684106,5.3694363,6.3967185,8.789334,12.340514,10.089026,8.812308,10.197334,10.817642,7.3780518,6.7183595,6.9382567,7.748924,10.482873,10.505847,7.2894363,4.391385,3.3509746,3.692308,3.620103,3.892513,4.2240005,5.428513,9.4457445,5.661539,3.3608208,2.7569232,3.4494362,4.4242053,7.3682055,9.019077,9.842873,10.161232,10.161232,10.587898,10.742155,9.337437,7.3321033,7.9195905,11.286975,14.76595,17.96595,20.368412,21.330053,18.694565,14.427898,10.200616,7.1154876,5.723898,4.7950773,3.9023592,3.2754874,2.9210258,2.6387694,2.7864618,1.9889232,1.2209232,0.90584624,0.9321026,0.39384618,0.12143591,0.01969231,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.0032820515,0.0,0.0,0.0032820515,0.016410258,0.026256412,0.03938462,0.052512825,0.059076928,0.04594872,0.02297436,0.032820515,0.059076928,0.072205134,0.06235898,0.08533334,0.09189744,0.09189744,0.0951795,0.108307704,0.108307704,0.098461546,0.09189744,0.0951795,0.108307704,0.13128206,0.15425642,0.17394873,0.190359,0.21333335,0.21333335,0.2231795,0.23958977,0.27241027,0.32164106,0.39384618,0.512,1.1060513,1.8642052,1.7558975,1.5458462,1.3128207,2.0644104,3.629949,4.670359,5.0477953,6.944821,8.795898,10.308924,12.481642,15.556924,17.024002,16.656412,14.450873,10.604308,8.408616,6.6592827,5.6451287,5.221744,4.8082056,6.73477,10.200616,15.035078,20.719591,26.397541,23.834259,16.768002,13.026463,14.6871805,18.080822,18.435284,17.736206,16.613745,15.428925,14.283488,9.508103,5.0215387,2.1103592,0.9156924,0.4266667,0.108307704,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.016410258,0.016410258,0.026256412,0.03938462,0.04594872,0.052512825,0.07548718,0.101743594,0.15097436,0.77456415,1.6377437,1.5425643,1.2471796,2.0250258,3.6496413,6.0783596,9.458873,10.8996935,11.306667,11.099898,10.614155,10.102155,9.429334,10.663385,12.770463,15.556924,19.669334,26.456617,33.65744,42.003696,50.07754,54.275288,54.09149,56.50052,61.23652,67.843285,75.67098,82.98011,87.611084,90.18093,90.9555,89.84288,85.474464,81.12247,77.0396,73.31119,69.8716,66.21867,66.067696,68.844315,73.80678,80.02954,74.35488,61.31529,47.323902,36.55549,30.976002,28.2519,25.521233,23.312412,21.461334,19.104822,17.893745,16.768002,15.77354,15.044924,14.8020525,14.887385,15.750566,16.324924,16.01641,14.710155,14.332719,14.483693,14.752822,15.123693,15.990155,18.103796,18.724104,18.248207,17.171694,16.098463,17.184822,17.814976,17.942976,17.85436,18.15631,0.0,0.0,0.0,0.0,0.0,0.0,0.06235898,0.86646163,1.8346668,2.231795,1.1684103,1.083077,0.6859488,0.42338464,0.44307697,0.5874872,0.15097436,0.016410258,0.0,0.0,0.0,0.0032820515,0.0,0.0,0.006564103,0.036102567,0.07548718,0.072205134,0.108307704,0.17394873,0.13456412,0.026256412,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.026256412,0.01969231,0.0,0.0,0.0,0.2855385,0.2855385,0.0032820515,0.02297436,0.92225647,3.3312824,2.9833848,0.2986667,0.37415388,0.95835906,1.0765129,1.6869745,3.383795,6.36718,6.1013336,3.1507695,1.7690258,2.612513,2.7273848,1.7362052,1.4441026,1.6410258,1.7362052,0.77128214,0.21661541,0.032820515,0.0032820515,0.0,0.0,0.013128206,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.013128206,0.049230773,0.07548718,0.41682056,0.51856416,0.4397949,0.8467693,0.56451285,0.9485129,1.4309745,1.7066668,1.7165129,0.8598975,0.47917953,0.47261542,0.6662565,0.7975385,0.5021539,0.18051283,0.006564103,0.0,0.0,0.0,0.0032820515,0.0032820515,0.009846155,0.026256412,0.049230773,0.12143591,0.32164106,0.55794877,0.58092314,0.8205129,0.7450257,0.54482055,0.43651286,0.6498462,1.6607181,2.868513,4.2436924,5.3037953,5.113436,4.076308,3.121231,2.5895386,2.4385643,2.2416413,1.9856411,1.9823592,2.1070771,2.176,1.9265642,1.7952822,2.1333334,2.5928206,2.9078977,2.8914874,2.9144619,1.9659488,0.9714873,0.40369233,0.27241027,0.23630771,0.32164106,0.54482055,0.79425645,0.827077,0.8205129,1.4506668,1.9035898,1.8576412,1.463795,1.4211283,1.9987694,2.6847181,3.0490258,2.737231,2.553436,2.1825643,1.7493335,1.3981539,1.2996924,1.0732309,0.955077,0.7844103,0.571077,0.47589746,0.6104616,0.764718,1.4900514,2.3696413,2.0217438,0.8960001,0.58092314,0.5415385,0.46933338,0.2986667,0.29210258,0.41682056,0.44964105,0.39056414,0.44964105,0.67938465,0.7187693,0.60061544,0.39712822,0.23630771,0.17066668,0.068923086,0.009846155,0.013128206,0.02297436,0.29210258,0.48246157,0.74830776,1.4966155,3.387077,4.8705645,5.3891287,5.0510774,4.6080003,5.4580517,7.1876926,8.740103,9.435898,10.066052,12.898462,10.870154,7.643898,5.1856413,4.535795,5.8125134,7.397744,8.881231,9.984001,10.125129,8.438154,8.507077,8.2904625,7.384616,6.547693,7.683283,7.9786673,7.3714876,6.7610264,6.6133337,6.944821,7.171283,7.322257,7.250052,7.4929237,9.278359,10.840616,9.83959,7.788308,6.038975,5.786257,6.2096415,6.8332314,6.820103,6.0258465,4.9985647,4.709744,5.169231,5.3694363,4.903385,3.9614363,6.36718,7.9458466,7.9524107,6.941539,6.770872,6.5969234,5.674667,4.8705645,5.2742567,8.201847,8.185436,6.422975,4.7983594,4.57518,6.380308,6.813539,5.8157954,4.450462,3.9122055,5.5532312,6.186667,9.15036,13.292309,16.305231,14.762668,13.351386,11.411694,8.139488,5.3760004,7.6012316,9.238976,7.3091288,4.640821,2.9965131,3.0949745,3.1081028,3.6036925,4.8016415,6.764308,9.383386,8.608821,7.5946674,7.0925136,7.328821,8.01477,10.57477,12.137027,11.664412,9.882257,9.29477,11.090053,14.411489,18.379488,22.793848,28.146873,30.273643,29.45313,26.991592,23.663591,19.695591,13.866668,9.271795,6.3212314,4.9821544,4.781949,4.1189747,3.2918978,2.5895386,2.1366155,1.8937438,1.6804104,1.2537436,1.1454359,1.2931283,1.0666667,0.32164106,0.059076928,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.049230773,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.01969231,0.016410258,0.016410258,0.026256412,0.026256412,0.03938462,0.04594872,0.052512825,0.059076928,0.059076928,0.052512825,0.049230773,0.052512825,0.06235898,0.06235898,0.07548718,0.08533334,0.09189744,0.08861539,0.08205129,0.08205129,0.08205129,0.07876924,0.07876924,0.08205129,0.108307704,0.13128206,0.15425642,0.17394873,0.190359,0.21989745,0.23630771,0.25271797,0.27569234,0.29538465,0.36102566,0.45292312,0.7253334,1.0732309,1.1684103,1.0502565,1.2176411,1.7952822,2.612513,3.1803079,3.1474874,4.8836927,8.139488,12.22236,15.996719,19.2,18.425438,16.49231,14.116103,9.908514,7.683283,5.4153852,4.089436,4.1485133,5.4908724,6.6002054,8.293744,13.131488,20.276514,25.494976,24.365952,18.537027,15.369847,16.938667,20.010668,20.207592,19.954874,18.704412,15.727591,10.108719,5.4514875,3.131077,2.1858463,1.5753847,0.15753847,0.0951795,0.032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.006564103,0.0,0.0,0.0,0.0,0.006564103,0.016410258,0.016410258,0.026256412,0.03938462,0.055794876,0.07548718,0.101743594,0.14441027,0.2100513,0.4004103,0.6662565,0.77128214,0.9288206,1.5195899,2.609231,4.204308,6.23918,8.694155,10.7158985,11.69395,11.290257,9.429334,7.5881033,7.1876926,8.027898,10.010257,13.138052,17.700104,23.11877,29.584412,36.696617,43.483902,48.301952,53.277542,57.724724,61.49908,64.9879,71.15816,76.681854,80.896,83.75139,85.8158,85.45806,83.82359,80.70893,76.80329,73.70175,70.74462,68.75242,66.7799,65.253746,65.96924,67.59057,67.68903,63.245132,54.56739,45.31857,37.41867,32.02626,29.049438,27.680822,26.377848,23.814566,21.014977,18.710976,17.24718,16.584206,16.41354,16.994463,18.087385,18.944002,18.310566,17.45395,16.518566,15.563488,14.808617,14.647796,16.02954,17.132309,17.463797,17.161848,16.978052,18.628925,19.554462,19.442873,19.042463,20.148514,0.0,0.0,0.0,0.0,0.0,0.0,0.26256412,0.8008206,1.3161026,1.4112822,0.60061544,0.7220513,0.73517954,0.7056411,0.80738467,1.3489232,0.47589746,0.33476925,0.2297436,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.01969231,0.03938462,0.036102567,0.055794876,0.08533334,0.06564103,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14441027,0.14441027,0.0032820515,0.013128206,0.46276927,5.225026,5.8157954,2.0939488,2.28759,2.0118976,1.404718,1.7165129,3.698872,7.6307697,6.1341543,4.1058464,3.0490258,2.9801028,2.4549747,0.955077,0.67282057,0.9124103,1.024,0.39384618,0.19692309,0.059076928,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.026256412,0.049230773,0.24615386,0.2986667,0.27897438,0.6301539,0.48574364,0.7187693,1.2832822,1.9429746,2.300718,1.276718,0.7975385,0.60061544,0.53825647,0.5546667,1.1224617,1.2012309,0.92553854,0.5021539,0.20020515,0.10502565,0.049230773,0.016410258,0.0,0.006564103,0.006564103,0.013128206,0.10502565,0.26584616,0.37415388,0.42338464,0.5546667,0.77456415,0.96492314,0.8533334,0.9353847,1.5786668,2.7569232,3.7710772,3.2525132,2.553436,2.1202054,2.156308,2.609231,3.186872,2.740513,2.5829747,2.5895386,2.481231,1.8281027,1.5392822,1.5819489,1.6869745,1.7132308,1.6475899,1.975795,1.7690258,1.3193847,0.88615394,0.7122052,0.6662565,0.6629744,0.72861546,0.77456415,0.5907693,0.57764107,0.7318975,1.0436924,1.5753847,2.4648206,3.2262566,3.6168208,3.501949,2.8488207,1.7033848,1.2176411,0.88287187,0.63343596,0.4660513,0.41682056,0.37415388,0.40369233,0.3708718,0.27569234,0.23630771,0.36758977,0.54482055,1.2931283,2.297436,2.3991797,1.6672822,0.9682052,0.56123084,0.42338464,0.25271797,0.23630771,0.318359,0.3511795,0.2986667,0.26256412,0.571077,0.7975385,0.84348726,0.7089231,0.48574364,0.2231795,0.08533334,0.04266667,0.06235898,0.09189744,0.31507695,0.48902568,0.7384616,1.719795,4.634257,6.678975,7.171283,7.0990777,7.3747697,8.828718,11.162257,12.156719,12.035283,11.52,11.835078,10.112,6.6067696,4.1911798,3.9122055,4.9887185,6.5312824,7.4207187,8.132924,8.323282,6.816821,6.3212314,5.7665644,5.172513,4.772103,5.0051284,4.71959,4.4767184,4.4898467,5.024821,6.3901544,7.4830775,7.7259493,7.75877,8.375795,10.512411,10.512411,8.953437,7.463385,6.6034875,5.868308,5.8223596,6.452513,6.75118,6.173539,4.6539493,5.2480006,6.436103,6.6395903,5.658257,4.6769233,7.827693,9.055181,8.362667,6.9349747,7.145026,7.2992826,7.5881033,7.27959,6.5870776,6.669129,5.7403083,4.9985647,5.1659493,6.4000006,8.293744,11.23118,11.421539,9.481847,6.997334,6.5411286,6.163693,10.197334,14.792206,16.49559,12.268309,13.692719,11.441232,7.9950776,6.0028725,8.264206,8.832001,6.5378466,3.9844105,2.6026669,2.6617439,3.2918978,4.706462,6.7216415,8.78277,9.990565,10.8307705,11.080206,10.788103,10.223591,9.882257,11.45436,13.794462,15.228719,15.862155,17.575386,22.426258,27.654566,33.043694,37.635284,39.702976,37.792824,33.30626,27.14913,20.59159,15.258258,10.725744,7.5487185,5.6320004,4.604718,3.82359,3.4166157,2.550154,1.8215386,1.4506668,1.270154,1.2800001,1.5261539,1.4473847,0.9714873,0.4955898,0.14112821,0.01969231,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.02297436,0.013128206,0.013128206,0.013128206,0.009846155,0.009846155,0.009846155,0.0032820515,0.0032820515,0.009846155,0.009846155,0.01969231,0.02297436,0.029538464,0.03938462,0.03938462,0.036102567,0.04266667,0.049230773,0.052512825,0.052512825,0.052512825,0.049230773,0.052512825,0.06235898,0.06235898,0.06564103,0.08205129,0.08861539,0.08205129,0.07548718,0.068923086,0.072205134,0.07548718,0.07548718,0.07548718,0.09189744,0.12143591,0.15425642,0.18051283,0.20020515,0.2231795,0.24287182,0.26584616,0.29210258,0.3249231,0.3511795,0.4201026,0.5907693,0.8369231,1.0502565,1.2077949,1.2438976,1.3456411,1.6640002,2.3138463,3.117949,5.169231,8.1755905,11.858052,15.95077,17.266872,15.832617,13.495796,10.817642,7.069539,5.4514875,5.4547696,5.8092313,6.189949,7.2172313,7.7259493,7.827693,9.842873,13.889642,17.906874,17.316103,14.739694,14.037334,15.91795,17.910154,17.555695,17.06995,14.444309,9.869129,5.730462,3.6102567,1.9790771,1.0994873,0.7122052,0.036102567,0.06564103,0.03938462,0.009846155,0.0,0.0,0.0,0.0,0.009846155,0.026256412,0.01969231,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.006564103,0.016410258,0.016410258,0.026256412,0.03938462,0.06235898,0.0951795,0.13456412,0.190359,0.27569234,0.38400003,0.51856416,0.7089231,1.014154,1.5327181,2.2153847,3.006359,3.8301542,5.280821,6.9677954,8.306872,8.667898,7.384616,5.7632823,5.110154,5.691077,7.4240007,9.856001,13.157744,16.99118,21.54995,26.965336,33.316105,39.266464,45.252926,50.996517,56.159184,60.320824,63.9639,67.78749,71.8277,75.75303,78.8677,80.48903,80.00001,78.56575,76.5998,73.77396,71.21724,69.0839,66.64206,63.789955,61.042877,60.845955,61.774773,61.824005,59.73662,55.000618,47.829338,41.284927,36.47344,33.522873,31.576618,29.184002,26.200617,23.394463,21.280823,20.132105,19.373951,19.557745,20.361847,21.113438,20.795078,19.744822,19.035898,17.920002,16.433231,15.402668,15.799796,16.416822,17.152,18.336823,20.739285,23.141745,22.912003,21.221745,19.626669,20.069746,0.0,0.0,0.0,0.0,0.03938462,0.190359,0.39056414,0.6826667,0.90256417,0.8960001,0.508718,0.47917953,0.5481026,0.761436,1.0765129,1.3554872,0.46276927,0.5349744,0.57764107,0.27897438,0.006564103,0.006564103,0.009846155,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.052512825,0.256,3.0194874,5.933949,5.280821,2.3138463,3.2722054,2.5337439,1.7066668,1.6508719,2.9111798,5.7009234,4.9854364,3.7776413,2.9111798,2.553436,2.2186668,0.6432821,0.23630771,0.24615386,0.23958977,0.08205129,0.13456412,0.08533334,0.026256412,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.016410258,0.049230773,0.08205129,0.13456412,0.25928208,0.3117949,0.42338464,0.8369231,1.5327181,2.1924105,1.4080001,1.0404103,0.86646163,0.75487185,0.6892308,1.2373334,1.4933335,1.3193847,0.85005134,0.50543594,0.4397949,0.5218462,0.49230772,0.31507695,0.18379489,0.04594872,0.0032820515,0.032820515,0.18051283,0.5874872,0.44307697,0.508718,0.90256417,1.4769232,1.8018463,1.529436,1.6836925,2.169436,2.5928206,2.2777438,2.3663592,2.5206156,2.7798977,3.18359,3.7842054,3.1671798,2.740513,2.5009232,2.297436,1.8084104,1.6672822,1.7526156,1.5885129,1.1848207,1.0568206,1.3095386,1.5130258,1.5786668,1.463795,1.1749744,0.92225647,0.7253334,0.61374366,0.5284103,0.3052308,0.53825647,1.1093334,1.8182565,2.5665643,3.370667,3.4166157,3.18359,2.5862565,1.6902566,0.7089231,0.39384618,0.20676924,0.118153855,0.0951795,0.11158975,0.108307704,0.12143591,0.108307704,0.07548718,0.06564103,0.17066668,0.34789747,0.81066674,1.4178462,1.6738462,1.6771283,1.2800001,0.79097444,0.40697438,0.2297436,0.25928208,0.27897438,0.28225642,0.24615386,0.14769232,0.48246157,0.764718,0.9124103,0.90584624,0.79097444,0.39384618,0.15753847,0.10502565,0.19692309,0.318359,0.36430773,0.5481026,0.94523084,2.3236926,6.1308722,8.231385,7.3583593,6.806975,8.004924,10.489437,13.584412,13.482668,12.117334,10.925949,10.84718,9.931488,7.5881033,6.055385,5.7107697,5.093744,5.832206,5.677949,5.937231,6.5345645,6.012718,5.6254363,4.1878977,3.3903592,3.5183592,3.436308,2.9636924,2.8553848,3.383795,4.6178465,6.4032826,7.4863596,7.781744,8.146052,9.042052,10.561642,9.074872,7.529026,7.2631803,7.890052,7.3025646,6.1341543,6.088206,6.485334,6.564103,5.4974365,6.2129235,7.3682055,7.200821,6.0356927,6.294975,8.004924,8.513641,7.9425645,7.076103,7.3583593,8.280616,10.834052,11.848206,10.71918,9.403078,6.3901544,5.9634876,6.921847,8.300308,9.357129,12.800001,12.947693,10.978462,8.569437,7.8703594,7.768616,12.009027,15.908104,16.000002,10.069334,10.492719,8.789334,7.069539,6.6527185,8.070564,7.2631803,5.225026,3.6496413,3.1967182,3.515077,4.1550775,5.940513,8.146052,10.151385,11.467488,12.268309,12.757335,12.813129,12.596514,12.544001,13.371078,15.75713,18.707693,21.848618,25.422771,30.742977,34.97354,38.029133,39.223797,37.293953,33.57867,28.514463,22.708515,17.017437,12.553847,9.685334,7.529026,5.940513,4.6900516,3.4625645,2.9046156,2.0906668,1.4802053,1.2340513,1.1913847,1.3423591,1.5031796,1.2504616,0.61374366,0.072205134,0.026256412,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.01969231,0.02297436,0.02297436,0.032820515,0.02297436,0.013128206,0.009846155,0.016410258,0.02297436,0.02297436,0.02297436,0.029538464,0.03938462,0.04594872,0.03938462,0.04594872,0.049230773,0.04594872,0.04594872,0.04594872,0.04594872,0.049230773,0.055794876,0.06235898,0.06564103,0.07876924,0.08205129,0.07548718,0.07548718,0.06564103,0.068923086,0.07548718,0.07876924,0.08205129,0.08861539,0.11158975,0.14112821,0.17394873,0.20676924,0.2297436,0.25271797,0.28225642,0.38728207,0.7056411,0.6301539,0.6268718,0.80738467,1.083077,1.1848207,1.3128207,1.9068719,2.0020514,1.6640002,1.9790771,3.2098465,5.76,8.349539,10.538668,12.747488,13.082257,12.087796,10.128411,7.5946674,4.886975,4.896821,6.373744,7.4469748,7.634052,7.827693,8.779488,9.383386,10.656821,12.970668,16.032822,14.316309,12.232206,11.769437,12.921437,13.705847,13.558155,12.822975,9.849437,5.504,3.1671798,2.4976413,1.1520001,0.22646156,0.013128206,0.0,0.049230773,0.055794876,0.036102567,0.013128206,0.04266667,0.03938462,0.013128206,0.009846155,0.026256412,0.01969231,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.016410258,0.02297436,0.032820515,0.059076928,0.098461546,0.14769232,0.21661541,0.32164106,0.45292312,0.6235898,0.8533334,1.1848207,1.6508719,2.1202054,2.5107694,2.806154,3.3017437,4.027077,4.8049235,5.2545643,4.7917953,4.027077,3.9811285,4.893539,6.675693,8.897642,11.648001,14.450873,17.657436,21.54995,26.358156,31.389542,36.26667,41.892105,48.23303,54.3278,58.21375,61.75836,65.414566,68.87057,71.04329,73.12739,73.51467,73.275085,72.39549,69.77641,67.91878,66.43529,64.89272,62.897236,60.09108,57.682056,56.336414,56.241234,56.608826,55.680004,52.04021,47.51098,43.30667,39.922874,37.14298,34.323696,31.077745,28.107489,25.80677,24.25108,23.305847,23.3879,23.85395,23.798155,22.04554,20.535797,19.889233,19.055592,17.736206,16.410257,16.554668,16.987898,18.402462,21.490873,26.935797,29.699284,27.710361,23.972105,20.801643,19.849848,0.0,0.0,0.0,0.0,0.07548718,0.37743592,0.37743592,0.65641034,0.92553854,0.9517949,0.56123084,0.2986667,0.108307704,0.3708718,0.8041026,0.49887183,0.16410258,0.5021539,0.8402052,0.77128214,0.13128206,0.07876924,0.04266667,0.02297436,0.006564103,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.01969231,0.0032820515,0.0,0.0,0.27241027,1.3554872,6.692103,4.926359,1.8609232,0.7778462,2.4484105,2.2482052,1.9495386,1.7788719,1.9462565,2.665026,3.2787695,2.162872,1.1552821,0.90912825,0.90256417,0.24615386,0.11158975,0.08861539,0.032820515,0.072205134,0.072205134,0.08205129,0.052512825,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0,0.013128206,0.03938462,0.06235898,0.06564103,0.0951795,0.20348719,0.43323082,0.7515898,1.0601027,1.1257436,1.148718,1.1191796,1.0666667,1.0371283,0.8730257,0.9616411,0.955077,0.81394875,0.78769237,0.81066674,1.1355898,1.2438976,1.0929232,1.1191796,0.46276927,0.118153855,0.01969231,0.19692309,0.79425645,0.6170257,0.48246157,0.7450257,1.4966155,2.5698464,2.2678976,2.034872,1.8116925,1.7723079,2.3302567,2.937436,3.1737437,3.0720003,2.8291285,2.802872,2.353231,1.8543591,1.4769232,1.3128207,1.3620514,1.4408206,1.8937438,1.8642052,1.339077,1.1651284,1.276718,1.2931283,1.3718976,1.4276924,1.1257436,0.7122052,0.4266667,0.27569234,0.2100513,0.128,0.6301539,1.7263591,2.6518977,2.993231,2.7208207,1.5491283,0.9878975,0.6859488,0.446359,0.2100513,0.13128206,0.052512825,0.029538464,0.052512825,0.072205134,0.026256412,0.02297436,0.029538464,0.029538464,0.006564103,0.04266667,0.19364104,0.36430773,0.508718,0.6235898,0.98133343,1.2242053,0.9878975,0.44307697,0.26912823,0.4004103,0.37415388,0.3117949,0.256,0.17723078,0.4266667,0.6432821,0.8205129,0.9747693,1.1224617,0.7253334,0.3314872,0.21333335,0.380718,0.5973334,0.56123084,0.80738467,1.463795,3.2787695,7.634052,10.266257,7.7456417,6.3540516,8.132924,10.889847,13.334975,12.232206,10.417232,9.40636,9.40636,9.18318,8.763078,8.27077,7.322257,4.9985647,5.3234878,5.024821,5.330052,6.3310776,7.0137444,7.020308,5.0642056,3.6890259,3.5610259,3.4625645,3.186872,3.3312824,3.9909747,5.0477953,6.166975,7.39118,7.506052,7.6668725,8.556309,10.377847,8.815591,7.499488,7.637334,8.67118,8.27077,6.173539,5.5007186,6.235898,7.6964107,8.5202055,8.507077,8.641642,7.75877,6.7117953,8.372514,7.9917955,8.572719,9.088,9.127385,8.900924,10.804514,13.778052,15.081027,14.139078,12.550565,9.238976,9.429334,10.213744,10.276103,9.908514,11.844924,10.138257,8.050873,7.3747697,8.438154,9.242257,13.53518,16.866463,16.275694,10.266257,6.8299494,5.874872,5.973334,6.2227697,6.2555904,5.2644105,4.7392826,4.8114877,5.284103,5.6287184,5.5663595,6.810257,8.582564,10.555078,12.816411,12.763899,12.872206,13.436719,14.437745,15.553642,16.055796,17.155283,19.373951,22.478771,25.488413,28.09108,29.351387,28.977234,27.06708,24.086977,21.704206,18.796309,16.137848,13.784616,11.090053,8.963283,7.1187696,5.5696416,4.345436,3.495385,2.7766156,2.2186668,1.8084104,1.585231,1.6311796,1.4900514,0.9156924,0.5316923,0.40697438,0.03938462,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.016410258,0.02297436,0.036102567,0.052512825,0.032820515,0.01969231,0.013128206,0.016410258,0.026256412,0.026256412,0.01969231,0.01969231,0.029538464,0.03938462,0.03938462,0.049230773,0.049230773,0.04266667,0.04266667,0.04266667,0.04266667,0.04266667,0.04594872,0.059076928,0.068923086,0.072205134,0.07548718,0.07548718,0.07548718,0.06235898,0.06564103,0.072205134,0.07548718,0.08205129,0.08861539,0.098461546,0.118153855,0.14441027,0.19364104,0.2297436,0.256,0.29210258,0.47917953,1.0666667,0.92553854,0.94523084,1.3620514,1.847795,1.5064616,1.2898463,2.8455386,3.4067695,2.5698464,2.294154,3.2787695,6.363898,9.002667,9.911796,9.097847,9.435898,8.999385,7.574975,5.5893335,4.1189747,5.8912826,7.39118,8.001641,7.88677,7.9983597,11.142565,14.076719,16.95836,19.636515,21.635284,16.242872,11.703795,9.80677,10.240001,10.59118,10.709334,9.544206,7.312411,4.6539493,2.6420515,1.4506668,0.48574364,0.02297436,0.0,0.0032820515,0.04266667,0.06564103,0.052512825,0.032820515,0.0951795,0.098461546,0.055794876,0.02297436,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.013128206,0.02297436,0.04594872,0.08205129,0.12471796,0.20676924,0.31507695,0.45620516,0.65312827,0.9156924,1.2438976,1.6508719,2.0873847,2.5107694,2.9078977,3.239385,3.2918978,3.2032824,3.0687182,2.9472823,2.986667,3.6496413,4.965744,6.8529234,9.110975,11.500309,13.955283,16.57436,19.492104,22.889027,26.633848,29.535181,33.22421,38.38031,44.734364,51.30503,56.68103,60.914875,63.88513,65.28657,67.11795,68.23714,68.174774,66.724106,63.94093,62.516518,61.4958,60.45867,59.38216,58.61416,56.963287,55.135185,53.11344,51.27221,50.349953,49.486774,48.26585,46.749542,44.872208,42.453335,39.03344,35.49867,32.610462,30.441029,28.3799,27.782566,28.681849,29.193848,27.697233,22.820105,20.102566,18.71754,18.064411,17.526155,16.475899,16.968206,17.719797,19.787489,23.998362,30.926771,33.473644,31.054771,27.201643,24.159182,22.89231,0.0,0.0,0.0,0.0,0.0,0.0,0.32820517,0.16410258,0.0,0.036102567,0.18379489,0.574359,0.27897438,0.016410258,0.032820515,0.108307704,0.3511795,0.4201026,0.7253334,1.0601027,0.5940513,0.3249231,0.12143591,0.036102567,0.03938462,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01969231,0.09189744,0.01969231,0.0,0.0,0.84348726,4.210872,3.259077,1.2537436,0.15425642,0.3708718,0.761436,2.740513,3.7185643,3.3969233,2.359795,2.0906668,1.847795,1.0075898,0.5021539,0.45292312,0.18379489,0.12143591,0.068923086,0.026256412,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.016410258,0.016410258,0.0032820515,0.0,0.0,0.006564103,0.029538464,0.06564103,0.29538465,0.4660513,0.48574364,0.4135385,0.75487185,1.1881026,1.4145643,1.404718,1.404718,1.270154,1.1093334,0.81394875,0.58092314,0.88615394,0.71548724,0.94523084,1.4572309,2.3171284,3.767795,1.8510771,0.5481026,0.0,0.0,0.0,0.0,0.055794876,0.34133336,0.8598975,1.4342566,1.2406155,1.9790771,2.4976413,2.806154,4.089436,4.089436,3.0818465,2.15959,1.7165129,1.4342566,1.4966155,1.463795,1.4342566,1.4703591,1.6180514,1.3718976,1.2931283,1.1158975,0.88615394,0.94523084,1.0075898,0.7187693,0.36102566,0.101743594,0.016410258,0.03938462,0.09189744,0.14112821,0.16410258,0.15097436,0.3117949,0.75487185,1.0469744,0.9517949,0.4266667,0.08533334,0.009846155,0.016410258,0.016410258,0.016410258,0.052512825,0.032820515,0.032820515,0.06235898,0.06235898,0.02297436,0.016410258,0.026256412,0.04266667,0.029538464,0.01969231,0.068923086,0.21661541,0.4397949,0.67282057,0.65969235,0.6104616,0.53825647,0.46276927,0.4266667,0.5481026,0.50543594,0.36102566,0.23958977,0.33476925,0.26256412,0.46276927,0.77456415,1.1093334,1.463795,1.086359,0.6268718,0.44307697,0.574359,0.7318975,1.0371283,1.332513,1.9429746,3.764513,8.27077,13.945437,12.33395,11.437949,13.6467705,15.747283,14.306462,11.556104,9.682052,8.930462,7.5979495,8.392206,8.113232,6.4000006,4.204308,3.8137438,5.097026,4.9132314,4.450462,4.7655387,6.806975,5.720616,6.6002054,7.5421543,7.7357955,7.4929237,5.464616,5.7468724,6.0225644,5.605744,5.4482055,9.07159,8.549745,6.8430777,6.6560006,10.453334,10.404103,8.1755905,6.764308,6.6100516,5.586052,4.522667,5.0543594,7.4896417,10.948924,13.367796,13.879796,12.688411,11.424822,10.889847,11.047385,10.499283,12.501334,13.912617,13.479385,11.85477,15.064616,14.158771,13.344822,12.931283,9.291488,11.720206,15.927796,17.079796,14.060308,9.4457445,12.583385,10.722463,8.388924,8.011488,9.90195,11.588924,13.88636,15.540514,14.979283,10.315488,6.8004107,5.5630774,5.3694363,5.4875903,5.7074876,6.3179493,7.578257,8.621949,8.828718,7.827693,7.2664623,7.5913854,8.897642,10.679795,11.841642,12.06154,12.983796,14.211283,15.248411,15.51754,15.579899,14.460719,13.587693,13.2562065,12.635899,12.465232,12.2387705,12.501334,12.809847,11.733335,10.610872,9.386667,8.077128,6.7085133,5.3398976,4.571898,3.8564105,3.3641028,3.0916924,2.8849232,3.2000003,3.1442053,2.7766156,2.3171284,2.1202054,1.204513,0.51856416,0.14769232,0.03938462,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01969231,0.029538464,0.026256412,0.016410258,0.016410258,0.006564103,0.006564103,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.02297436,0.029538464,0.029538464,0.029538464,0.029538464,0.029538464,0.029538464,0.032820515,0.04594872,0.04594872,0.055794876,0.06564103,0.07548718,0.07548718,0.052512825,0.04594872,0.052512825,0.059076928,0.04594872,0.068923086,0.0951795,0.11158975,0.13128206,0.16738462,0.20348719,0.2231795,0.26584616,0.33476925,0.39712822,0.4201026,0.88615394,2.1431797,3.2787695,2.1070771,1.7033848,2.8389745,3.5446157,3.4166157,3.6004105,4.7622566,8.411898,11.365745,11.953232,10.023385,8.595693,7.351795,5.7403083,4.069744,3.508513,4.9854364,7.351795,8.815591,9.462154,11.244308,18.91118,23.581541,26.01354,26.686361,25.833027,13.1872835,7.653744,7.90318,11.1294365,13.046155,10.9456415,8.178872,5.609026,3.7185643,2.5928206,0.64000005,0.068923086,0.009846155,0.0032820515,0.016410258,0.016410258,0.016410258,0.02297436,0.032820515,0.04594872,0.108307704,0.14112821,0.12143591,0.06235898,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.0032820515,0.009846155,0.026256412,0.052512825,0.07548718,0.15097436,0.23302566,0.36102566,0.5481026,0.79425645,1.1093334,1.5097437,1.9987694,2.5435898,3.0654361,3.4100516,3.5938463,3.6627696,3.6562054,3.629949,3.7776413,4.263385,5.4482055,7.243488,9.124104,10.564924,13.223386,15.8654375,18.202257,20.873848,24.513643,27.638157,29.797747,31.524105,34.33354,41.206158,47.894978,54.400005,60.43898,65.44411,67.373955,68.05662,67.28206,64.941956,61.036312,58.069336,56.26421,54.751183,53.392414,52.78195,52.877132,52.9198,52.48657,51.328003,49.362057,46.50667,44.465233,43.47077,43.405132,43.808823,42.587902,40.415184,38.12431,35.7678,32.594055,32.384003,35.885952,36.936207,32.915695,24.74995,19.64636,16.94195,15.924514,15.671796,15.061335,15.281232,15.977027,17.362053,19.817028,23.896618,25.83631,27.346054,29.24636,31.671797,34.087387,0.0,0.0,0.0,0.0,0.0,0.0,0.06564103,1.4178462,1.4080001,0.11158975,0.318359,0.5907693,0.36758977,0.13128206,0.08861539,0.18051283,0.2100513,0.16738462,0.36102566,0.67610264,0.58420515,0.33476925,0.18707694,0.108307704,0.068923086,0.016410258,0.0032820515,0.013128206,0.01969231,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.01969231,0.0032820515,0.0,0.009846155,0.20676924,0.93866676,0.69251287,0.26912823,0.052512825,0.28225642,1.0436924,3.3641028,3.8564105,3.0358977,1.9528207,2.2121027,1.7132308,0.9944616,1.0436924,1.6377437,1.3292309,0.6629744,0.24943592,0.049230773,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.026256412,0.02297436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.016410258,0.0032820515,0.0,0.0,0.0,0.006564103,0.02297436,0.09189744,0.15097436,0.17066668,0.15425642,0.36102566,0.67282057,0.96492314,1.211077,1.463795,1.8576412,2.100513,2.1333334,1.8543591,1.1060513,0.6498462,0.45292312,0.46276927,0.6268718,0.88943595,0.40697438,0.1148718,0.0,0.0,0.0,0.0,0.1148718,0.4594872,0.79425645,0.51856416,0.35446155,0.99774367,2.0808206,3.0326157,3.0654361,2.0775387,1.5622566,1.6443079,2.1431797,2.605949,2.6584618,2.4484105,2.3269746,2.3433847,2.2777438,1.7985642,1.654154,1.5885129,1.4933335,1.3981539,2.0151796,1.6246156,0.9616411,0.4660513,0.27241027,0.13128206,0.10502565,0.108307704,0.098461546,0.06564103,0.098461546,0.5546667,1.4572309,2.0742567,0.90256417,0.20020515,0.01969231,0.016410258,0.016410258,0.016410258,0.04266667,0.04266667,0.04266667,0.04266667,0.013128206,0.013128206,0.016410258,0.016410258,0.01969231,0.01969231,0.006564103,0.049230773,0.16410258,0.3314872,0.52512825,0.5907693,0.53825647,0.45620516,0.38400003,0.318359,0.51856416,0.53825647,0.47917953,0.3708718,0.17723078,0.2100513,0.39712822,0.6301539,0.8598975,1.086359,1.0108719,0.77128214,0.48574364,0.34789747,0.6235898,0.6629744,1.2242053,2.162872,3.8334363,7.0859494,10.732308,11.0145645,11.85477,13.512206,12.57354,10.390975,9.288206,8.448001,7.4896417,6.452513,5.799385,5.431795,5.333334,5.2709746,4.8049235,5.2447186,5.0576415,5.2414365,6.3868723,8.648206,7.171283,6.8562055,7.7423596,8.576,6.806975,5.6320004,5.5236926,5.609026,5.2709746,4.164923,6.9021544,9.908514,9.179898,5.937231,6.619898,7.322257,8.211693,8.267488,7.716103,8.0377445,8.585847,9.301334,10.476309,11.480617,10.755282,9.626257,8.320001,8.277334,9.360411,9.852718,10.755282,11.828514,11.611898,10.30236,9.744411,11.989334,14.536206,16.354464,15.983591,11.526565,12.822975,15.061335,14.759386,11.539693,8.12636,9.780514,9.750975,8.674462,7.637334,8.182155,8.041026,12.534155,15.113848,13.364513,8.982975,7.030154,6.485334,6.452513,7.0137444,9.235693,11.963078,13.10195,13.111795,12.3306675,10.978462,10.748719,11.113027,11.32636,11.414975,12.182976,12.842668,12.924719,12.612924,12.219078,12.173129,11.989334,11.191795,10.30236,9.442462,8.3134365,7.574975,7.1581545,6.954667,6.8233852,6.557539,6.432821,5.4580517,4.0467696,2.7142565,2.0676925,1.8084104,1.7033848,1.7558975,1.8838975,1.9331284,2.0742567,1.657436,1.3193847,1.148718,0.67938465,0.32164106,0.118153855,0.029538464,0.006564103,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.01969231,0.01969231,0.026256412,0.026256412,0.01969231,0.013128206,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.01969231,0.01969231,0.029538464,0.029538464,0.02297436,0.02297436,0.029538464,0.032820515,0.032820515,0.04266667,0.055794876,0.06564103,0.06564103,0.049230773,0.04594872,0.04594872,0.04594872,0.032820515,0.059076928,0.08205129,0.10502565,0.128,0.15425642,0.21333335,0.256,0.29538465,0.42994875,0.8598975,1.6180514,1.9561027,2.609231,3.4330258,3.4231799,2.1136413,1.7920002,2.28759,3.5216413,5.4941545,9.094564,12.422565,13.492514,12.0549755,9.596719,7.194257,6.8693337,6.813539,6.314667,5.7435904,6.2227697,8.612103,11.1064625,13.443283,16.886156,23.59467,28.760618,27.969643,21.395695,13.784616,11.264001,9.025641,8.14277,8.585847,9.212719,10.033232,6.99077,3.8400004,2.0676925,0.8960001,0.4004103,0.11158975,0.006564103,0.013128206,0.016410258,0.016410258,0.016410258,0.21333335,0.67938465,1.3653334,1.6016412,1.7526156,1.719795,1.3489232,0.4266667,0.10502565,0.016410258,0.013128206,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.0032820515,0.0032820515,0.006564103,0.013128206,0.026256412,0.06235898,0.11158975,0.190359,0.3052308,0.45292312,0.6826667,0.955077,1.3357949,1.8051283,2.2613335,2.7798977,3.170462,3.3608208,3.4166157,3.5577438,3.9876926,4.6900516,5.605744,6.8266673,8.598975,10.459898,12.35036,13.968411,15.258258,16.420103,19.157335,22.967796,26.83077,29.604105,29.997952,32.341335,36.660515,42.640415,49.713234,57.071594,62.93662,66.56657,67.885956,67.06216,64.51529,61.12821,58.325336,55.10893,51.616825,49.14216,47.921234,47.599594,47.668518,47.757133,47.62913,46.385235,44.356926,42.38113,40.950157,40.231388,40.37908,40.224823,39.565132,38.501747,37.425232,39.141747,43.21149,42.919388,36.099285,25.140514,20.358566,17.979078,17.060104,16.46277,14.815181,14.372104,14.329437,14.8020525,16.052513,18.500925,19.639797,22.304823,25.481848,27.749746,27.27713,0.0,0.0,0.0,0.0,0.0,0.0,0.06564103,0.80738467,0.8369231,0.16410258,0.18707694,0.45292312,0.702359,0.5874872,0.20348719,0.08861539,0.3052308,0.17066668,0.118153855,0.25271797,0.3314872,0.75487185,0.63343596,0.512,0.5284103,0.41025645,0.190359,0.06235898,0.013128206,0.016410258,0.026256412,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.01969231,0.049230773,0.01969231,0.009846155,0.03938462,0.23958977,0.83035904,2.9046156,3.4691284,3.0326157,2.231795,1.8412309,1.1323078,0.97805136,2.3335385,3.9220517,2.2219489,0.76800007,0.18379489,0.02297436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.06235898,0.12471796,0.14769232,0.072205134,0.013128206,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.032820515,0.052512825,0.072205134,0.2297436,0.380718,0.58092314,0.86317956,1.2242053,1.6738462,1.9889232,2.1792822,2.231795,2.0841026,1.7001027,1.2964103,0.88943595,0.508718,0.19692309,0.21333335,0.2297436,0.14441027,0.0,0.0,0.0,0.052512825,0.20020515,0.318359,0.1148718,0.07548718,0.35446155,0.86317956,1.3193847,1.2406155,0.83035904,0.7975385,1.2570257,2.041436,2.7241027,2.7963078,2.6518977,2.7175386,2.9801028,2.989949,2.5337439,2.4582565,2.5862565,2.6486156,2.281026,2.166154,1.657436,1.2012309,1.1257436,1.654154,1.2012309,0.90912825,0.81066674,0.77128214,0.5218462,0.25928208,0.29210258,0.702359,1.0535386,0.4266667,0.108307704,0.049230773,0.052512825,0.049230773,0.07876924,0.059076928,0.03938462,0.02297436,0.013128206,0.0,0.0032820515,0.006564103,0.006564103,0.006564103,0.006564103,0.0,0.02297436,0.10502565,0.24287182,0.39712822,0.47589746,0.45292312,0.39056414,0.3511795,0.41682056,0.446359,0.52512825,0.56451285,0.5218462,0.39384618,0.41682056,0.46933338,0.50543594,0.571077,0.77128214,0.78769237,0.5907693,0.34133336,0.38728207,1.273436,1.972513,4.125539,5.8190775,6.764308,8.2904625,10.499283,10.807796,10.663385,10.072617,7.604513,7.8080006,7.906462,7.1844106,5.7731285,4.663795,4.8804107,4.841026,4.7360005,4.6080003,4.3552823,4.821334,5.504,6.5247183,7.7292314,8.677744,7.4765134,6.8496413,7.069539,7.174565,4.9427695,4.007385,3.6135387,3.636513,4.0336413,4.844308,6.514872,8.582564,9.32759,8.536616,7.509334,8.41518,9.120821,8.953437,8.228104,8.247795,8.966565,10.315488,10.889847,10.630565,10.824206,9.580308,8.320001,8.612103,9.931488,9.662359,8.89436,8.930462,10.535385,13.466257,16.449642,18.560001,18.62236,16.902565,13.909334,10.374565,10.735591,12.872206,13.443283,11.369026,7.8145647,7.433847,7.8769236,7.899898,7.4765134,7.824411,9.005949,12.645744,14.329437,12.829539,10.115283,8.392206,7.4141545,7.0400004,7.6603084,10.20718,12.550565,13.00677,12.2617445,11.126155,10.528821,10.427077,10.55836,10.725744,10.880001,11.132719,11.536411,11.398565,11.001437,10.594462,10.374565,10.358154,9.872411,9.042052,8.01477,6.948103,6.298257,5.7534366,5.1298466,4.4340515,3.892513,3.882667,3.18359,2.2219489,1.3915899,1.0666667,1.0568206,1.148718,1.2931283,1.4211283,1.4375386,1.1027694,0.6629744,0.4135385,0.3446154,0.128,0.03938462,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.006564103,0.0,0.0,0.0,0.009846155,0.016410258,0.01969231,0.029538464,0.02297436,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.006564103,0.013128206,0.016410258,0.016410258,0.02297436,0.02297436,0.016410258,0.016410258,0.02297436,0.02297436,0.029538464,0.03938462,0.049230773,0.052512825,0.06235898,0.049230773,0.03938462,0.04266667,0.052512825,0.03938462,0.072205134,0.098461546,0.11158975,0.118153855,0.13456412,0.48246157,0.7089231,0.8992821,1.086359,1.2603078,2.1924105,2.1924105,2.156308,2.425436,2.7634873,1.8937438,1.5491283,2.0676925,3.7152824,6.688821,11.999181,12.219078,10.5780525,8.982975,7.9983597,7.282872,7.6110773,8.5661545,9.517949,9.626257,10.325335,10.758565,12.048411,15.783386,24.034464,28.65231,30.720003,27.109745,19.10154,12.393026,13.08554,11.972924,10.04636,8.352821,7.9983597,7.512616,5.0576415,2.7864618,1.4178462,0.23630771,0.15097436,0.059076928,0.016410258,0.02297436,0.02297436,0.016410258,0.108307704,0.40697438,1.1355898,2.6289232,3.9614363,4.2962055,3.9056413,2.740513,0.43323082,0.12471796,0.02297436,0.006564103,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.0,0.0,0.0,0.0,0.006564103,0.02297436,0.04266667,0.07548718,0.13456412,0.2297436,0.3708718,0.54482055,0.8041026,1.1355898,1.4276924,1.9396925,2.3072822,2.546872,2.7175386,2.9440002,3.4166157,4.0500517,4.778667,5.733744,7.250052,9.032206,10.752001,12.179693,13.092104,13.272616,14.674052,17.335796,21.162668,25.133951,27.313232,28.009027,30.024208,33.476925,38.31467,44.310978,51.072002,57.75754,61.9717,63.20903,62.87426,62.40821,61.47939,59.821953,57.216003,53.49744,49.601646,47.169643,45.613953,44.78031,44.934566,44.737644,43.83508,42.505848,40.96985,39.381336,38.912003,39.187695,39.424004,39.279594,38.85621,40.66462,43.85149,42.77498,36.260105,27.592207,23.61436,21.13313,19.643078,18.566566,17.253744,15.954053,15.27795,15.40595,16.54154,18.907898,21.766565,24.953438,26.272823,24.533335,19.551182,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0,0.072205134,0.12143591,0.14112821,0.13128206,0.101743594,0.2297436,0.6301539,0.6301539,0.23958977,0.15097436,0.508718,0.4135385,0.18707694,0.03938462,0.101743594,0.62030774,0.5546667,0.46276927,0.50543594,0.4135385,0.21333335,0.08533334,0.026256412,0.013128206,0.026256412,0.029538464,0.02297436,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.055794876,0.016410258,0.009846155,0.13784617,0.42994875,0.8533334,2.4155898,3.9680004,3.889231,2.422154,1.657436,1.3554872,2.0775387,3.3345644,3.8596926,1.6114873,0.4594872,0.068923086,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02297436,0.02297436,0.0,0.0,0.0,0.059076928,0.13456412,0.190359,0.190359,0.03938462,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.036102567,0.17723078,0.20020515,0.28225642,0.51856416,0.9124103,1.2570257,1.6082052,1.9396925,2.2646155,2.6387694,2.546872,2.2613335,1.8215386,1.2996924,0.8008206,0.65641034,0.55794877,0.380718,0.17394873,0.15753847,0.07548718,0.026256412,0.006564103,0.006564103,0.0,0.02297436,0.055794876,0.072205134,0.09189744,0.17394873,0.3117949,0.46276927,0.9419488,1.8281027,2.9440002,3.1803079,2.9407182,2.8389745,3.0162053,3.1113849,2.9801028,3.0523078,3.1967182,3.190154,2.7241027,1.9462565,1.4506668,1.2996924,1.5622566,2.3138463,2.048,1.6180514,1.270154,1.0371283,0.73517954,0.40697438,0.3314872,0.512,0.6662565,0.21333335,0.08533334,0.118153855,0.17066668,0.17723078,0.128,0.12471796,0.055794876,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.072205134,0.20020515,0.32820517,0.36430773,0.36102566,0.32820517,0.32164106,0.42994875,0.3708718,0.47261542,0.5677949,0.6170257,0.7187693,0.764718,0.6892308,0.5316923,0.42338464,0.60061544,0.60061544,0.47261542,0.3708718,0.83035904,2.7437952,5.681231,7.0432825,8.372514,9.849437,10.299078,11.139283,11.08677,10.423796,9.153642,7.000616,7.6176414,7.8703594,7.328821,6.3179493,5.920821,7.1515903,6.925129,6.1078978,5.3398976,5.037949,4.634257,5.0904617,6.547693,8.474257,9.642668,8.487385,7.1187696,6.518154,6.2916927,4.6933336,3.0851285,2.294154,2.1858463,2.9965131,5.3202057,7.0400004,7.785026,8.595693,9.366975,8.822155,10.19077,10.791386,10.499283,9.524513,8.41518,9.321027,10.217027,10.226872,9.777231,10.581334,10.33518,9.494975,10.098872,11.467488,10.194052,8.113232,8.621949,13.869949,22.534565,29.850258,28.983797,22.967796,15.894976,10.41395,7.719385,7.785026,10.174359,11.946668,11.336206,7.722667,6.4689236,6.3474874,6.626462,7.0334363,7.75877,9.403078,11.254155,12.189539,11.956513,11.191795,9.458873,7.893334,7.1154876,7.581539,9.586872,10.873437,10.683078,9.803488,9.061745,9.314463,9.088,9.334154,9.688616,10.003693,10.345026,10.627283,10.102155,9.4916935,9.117539,8.904206,9.179898,8.966565,8.260923,7.2960005,6.547693,6.0783596,5.412103,4.6211286,3.767795,2.8947694,3.0194874,2.9013336,2.5042052,1.9922053,1.7394873,1.4900514,1.273436,1.0633847,0.88287187,0.79097444,0.43651286,0.190359,0.07548718,0.055794876,0.04266667,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.006564103,0.0,0.0,0.0,0.009846155,0.016410258,0.016410258,0.02297436,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.013128206,0.009846155,0.009846155,0.009846155,0.006564103,0.013128206,0.016410258,0.016410258,0.016410258,0.016410258,0.013128206,0.013128206,0.016410258,0.016410258,0.02297436,0.036102567,0.04266667,0.04266667,0.055794876,0.052512825,0.04266667,0.04594872,0.059076928,0.052512825,0.07548718,0.10502565,0.128,0.16410258,0.27569234,0.9353847,0.92553854,0.95835906,1.276718,1.6508719,2.0611284,1.7033848,1.2964103,1.214359,1.4769232,1.5130258,1.654154,2.2219489,3.4330258,5.3891287,9.366975,8.707283,7.2205133,6.6494365,6.6560006,7.0104623,7.6209235,8.89436,10.55836,11.644719,12.95754,12.484924,13.551591,17.897026,25.659079,28.278156,27.457644,22.777437,16.384,12.967385,12.960821,10.857026,8.625232,7.2303596,6.633026,5.218462,3.4560003,2.1169233,1.2307693,0.068923086,0.026256412,0.016410258,0.02297436,0.032820515,0.04266667,0.059076928,0.26256412,0.7056411,1.5163078,2.8914874,4.059898,4.352,3.9548721,2.8455386,0.78769237,0.3511795,0.098461546,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.009846155,0.01969231,0.04594872,0.0951795,0.16738462,0.26912823,0.42994875,0.6301539,0.8008206,1.2012309,1.847795,2.1891284,2.1956925,2.3663592,2.6420515,3.1507695,3.761231,4.4996924,5.546667,7.056411,8.651488,10.134975,11.185231,11.329642,11.746463,12.76718,15.238565,18.986668,22.826668,23.942566,24.874668,26.354874,28.819695,32.423386,37.97662,45.075695,50.61252,53.474464,54.53457,56.631798,58.95549,60.90503,61.71898,60.45539,56.90093,53.727184,50.84226,48.433235,46.959595,45.50236,44.402874,43.411697,42.35816,41.153645,40.060722,39.581543,39.552002,39.53559,38.81354,39.95241,41.665646,40.677746,36.404514,30.946465,27.999182,25.580309,23.542156,21.779694,20.243694,18.756924,17.634462,17.411283,18.471386,21.064207,24.602259,26.906258,25.911797,21.35959,14.788924,0.0,0.0,0.0,0.009846155,0.029538464,0.04594872,0.06235898,0.06235898,0.049230773,0.049230773,0.108307704,0.072205134,0.21989745,0.25271797,0.18379489,0.3249231,0.6498462,0.67282057,0.47917953,0.21989745,0.108307704,0.02297436,0.0032820515,0.009846155,0.016410258,0.02297436,0.04266667,0.06235898,0.04594872,0.036102567,0.17066668,0.1148718,0.06235898,0.02297436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02297436,0.11158975,0.032820515,0.026256412,0.26584616,0.7187693,1.1355898,1.9593848,4.388103,4.522667,2.3762052,1.8838975,2.3269746,3.43959,3.18359,1.4572309,0.07548718,0.026256412,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.04266667,0.04266667,0.0,0.0,0.0,0.0,0.01969231,0.08533334,0.23302566,0.04594872,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.108307704,0.108307704,0.118153855,0.24615386,0.58092314,0.82379496,1.2537436,1.7362052,2.166154,2.4976413,2.7076926,2.740513,2.6157951,2.3466668,1.9364104,1.4539489,1.0929232,0.8008206,0.571077,0.46933338,0.2100513,0.068923086,0.009846155,0.0,0.0,0.0,0.0,0.0,0.02297436,0.12143591,0.24943592,0.29210258,0.61374366,1.4966155,3.1671798,3.5774362,3.117949,2.6157951,2.4516926,2.546872,2.7700515,2.993231,2.989949,2.7437952,2.4484105,1.6804104,1.2832822,1.2209232,1.4080001,1.6869745,2.0184617,1.7066668,1.1290257,0.6301539,0.50543594,0.446359,0.79097444,1.4342566,1.8281027,0.9616411,0.42338464,0.2855385,0.30851284,0.30194873,0.11158975,0.16082053,0.068923086,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.098461546,0.29210258,0.46933338,0.39056414,0.33476925,0.29538465,0.27569234,0.3117949,0.35446155,0.46276927,0.53825647,0.6301539,0.9353847,1.1257436,1.017436,0.7778462,0.67938465,1.1224617,1.6902566,1.4112822,1.0896411,1.657436,4.1550775,9.242257,8.78277,9.275078,11.762873,11.83836,11.864616,11.510155,11.680821,12.202667,11.818667,10.272821,9.747693,9.524513,9.380103,9.577026,9.990565,9.091283,8.109949,7.5913854,7.3682055,6.0849237,5.5926156,6.816821,9.409642,11.753027,9.941334,7.5191803,6.4590774,6.616616,5.7468724,3.6069746,2.6847181,2.4910772,3.0949745,5.139693,7.1647186,7.6077952,7.3386674,7.177847,7.890052,9.91836,11.625027,11.851488,10.512411,8.576,10.069334,10.066052,9.603283,9.186462,8.789334,9.537642,10.000411,11.474052,12.813129,10.443488,9.40636,12.0549755,19.554462,29.873234,37.789543,32.101746,22.603489,14.053744,8.887795,7.210667,7.6274877,9.6,10.912822,10.217027,7.0400004,6.2162056,5.3858466,5.579488,6.8430777,8.2445135,8.769642,9.032206,9.90195,11.332924,12.386462,11.011283,9.028924,7.6143594,7.394462,8.4512825,9.074872,8.726975,8.231385,8.086975,8.477539,8.152616,8.809027,9.216001,9.291488,10.098872,10.443488,9.429334,8.264206,7.5552826,7.3058467,7.8834877,7.8670774,7.2303596,6.3507695,6.0225644,5.6418467,4.906667,4.276513,3.8367183,3.2853336,3.4756925,4.0533338,3.9548721,3.1803079,2.789744,2.1234872,1.3259488,0.636718,0.19692309,0.06235898,0.101743594,0.08205129,0.08533334,0.1148718,0.08533334,0.016410258,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.013128206,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.006564103,0.0032820515,0.0032820515,0.0032820515,0.013128206,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.006564103,0.006564103,0.016410258,0.016410258,0.016410258,0.036102567,0.03938462,0.036102567,0.04594872,0.06235898,0.059076928,0.059076928,0.06564103,0.072205134,0.08205129,0.12143591,0.17066668,0.25271797,0.45620516,1.1388719,0.7089231,0.42994875,0.80738467,1.6180514,1.3259488,0.88615394,0.56123084,0.44307697,0.47589746,1.2209232,1.6836925,2.3794873,3.1474874,3.1507695,4.069744,5.3037953,6.6527185,7.5618467,7.1187696,6.567385,6.8299494,7.584821,8.746667,10.456616,12.032001,12.20595,13.6467705,16.643284,19.111385,20.345438,19.121233,15.858873,12.120616,10.624001,9.042052,5.8945646,4.667077,5.4153852,4.7589746,3.9089234,2.6322052,1.6311796,0.96492314,0.059076928,0.02297436,0.013128206,0.02297436,0.04266667,0.06564103,0.1148718,0.34133336,0.8205129,1.4408206,1.8871796,1.7755898,1.8379488,1.8182565,1.6114873,1.2537436,0.63343596,0.19364104,0.0032820515,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.02297436,0.055794876,0.11158975,0.19692309,0.3052308,0.4201026,0.67282057,1.6114873,2.03159,1.8084104,1.8773335,2.03159,2.428718,2.934154,3.4756925,4.0434875,5.1659493,6.4065647,7.817847,9.18318,10.033232,10.289231,10.31877,11.132719,13.200411,16.423386,18.566566,19.748104,20.762259,22.042257,23.657028,27.07036,31.90154,36.676926,40.231388,41.678772,44.399593,49.092926,54.272003,59.011288,62.92021,63.91139,63.681644,62.447594,60.16985,56.546467,51.823593,48.44308,46.148926,44.816414,44.468517,43.585644,42.27939,41.38339,40.795902,39.46667,39.525745,39.686565,39.286156,37.714054,34.422157,32.305233,30.260515,28.110771,25.764105,23.200823,21.904411,20.54236,19.761232,20.187899,22.455797,24.507078,24.776207,22.46236,18.103796,13.568001,0.0,0.0,0.0,0.02297436,0.0951795,0.2297436,0.26584616,0.24615386,0.15425642,0.036102567,0.0,0.19692309,0.26256412,0.21333335,0.14441027,0.2297436,0.5218462,0.4955898,0.65312827,0.90256417,0.5481026,0.12143591,0.02297436,0.02297436,0.013128206,0.0,0.0,0.0,0.006564103,0.18379489,0.8533334,0.32820517,0.07876924,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.0032820515,0.036102567,0.26256412,0.6465641,0.97805136,0.6104616,1.4178462,2.2777438,2.5895386,2.2744617,2.6880002,2.225231,1.1979488,0.18707694,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.072205134,0.072205134,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.15425642,0.16082053,0.029538464,0.09189744,0.2855385,0.6826667,1.2274873,1.8116925,2.28759,2.5206156,2.7241027,2.9078977,3.0227695,2.9768207,2.6584618,2.1497438,1.6049232,1.1290257,0.761436,0.2986667,0.08205129,0.009846155,0.0,0.0,0.0,0.0,0.0,0.013128206,0.06235898,0.108307704,0.07548718,0.13128206,0.6170257,2.044718,2.2416413,1.9232821,1.6607181,1.657436,1.7558975,1.7920002,2.048,2.0118976,1.7165129,1.7394873,1.5195899,1.0896411,0.6859488,0.4660513,0.5021539,0.9911796,1.0404103,0.6432821,0.14112821,0.21333335,0.5546667,1.5458462,2.8160002,3.623385,2.8521028,1.4375386,0.6629744,0.31507695,0.17394873,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.22646156,0.6662565,1.0666667,0.761436,0.5218462,0.3446154,0.24943592,0.27569234,0.4955898,0.6235898,0.6104616,0.5940513,0.8992821,1.3522053,1.3554872,1.270154,1.6738462,3.3575387,6.3343596,5.0116925,3.1737437,2.7241027,3.6758976,6.8627696,9.947898,11.963078,12.547283,11.946668,13.203693,12.045129,12.973949,16.275694,18.021746,15.602873,14.201437,13.610668,12.944411,10.650257,6.62318,5.5696416,6.5837955,8.477539,9.796924,11.149129,11.736616,12.091078,12.435693,12.678565,9.481847,7.1909747,6.62318,6.747898,4.6834874,4.588308,4.7458467,4.916513,5.10359,5.5532312,5.1265645,5.037949,4.9460516,4.568616,3.6791797,5.618872,8.549745,9.248821,7.6110773,6.62318,8.379078,9.862565,9.747693,8.021334,5.98318,5.858462,9.380103,12.57354,12.786873,8.697436,11.579078,16.692514,20.292925,20.65067,18.051283,11.37559,11.040821,11.933539,12.3995905,14.267078,15.218873,15.61272,12.822975,7.7718983,4.9296412,4.4274874,4.210872,5.6385646,8.477539,10.893129,11.273847,10.305642,10.880001,13.558155,16.587488,16.06236,13.4859495,10.41395,8.205129,8.011488,8.644924,8.960001,8.818872,8.257642,7.4765134,7.6603084,8.310155,8.707283,8.815591,9.291488,9.156924,8.464411,7.574975,6.695385,5.8912826,6.8299494,6.882462,6.0324106,4.9952826,5.2020516,4.972308,4.4110775,4.1911798,4.5554876,5.32677,4.4701543,5.182359,4.785231,3.058872,2.228513,1.8248206,0.73517954,0.06564103,0.036102567,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.026256412,0.03938462,0.04594872,0.04594872,0.04594872,0.08205129,0.09189744,0.08533334,0.08533334,0.12143591,0.15753847,0.2231795,0.26584616,0.27241027,0.25928208,0.30851284,0.32820517,0.33476925,0.3249231,0.27569234,0.27569234,0.42994875,0.508718,0.4266667,0.24287182,1.0371283,1.2635899,2.4713848,4.381539,4.8836927,5.970052,7.9327188,10.748719,12.832822,11.063796,8.205129,7.069539,6.308103,5.8420515,6.8660517,7.709539,8.073847,6.4656415,4.342154,6.1341543,6.3901544,8.03118,8.756514,7.4732313,4.2896414,3.31159,3.1573336,4.7392826,6.5017443,4.4406157,3.2820516,2.422154,1.270154,0.0951795,0.04594872,0.009846155,0.009846155,0.032820515,0.06564103,0.09189744,0.09189744,0.09189744,0.07876924,0.055794876,0.029538464,0.01969231,0.02297436,0.12143591,0.32820517,0.5940513,0.37415388,0.13784617,0.016410258,0.016410258,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.013128206,0.016410258,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.032820515,0.06564103,0.10502565,0.15097436,0.23958977,0.38728207,0.5940513,0.827077,1.024,1.7427694,1.9593848,2.2646155,2.8225644,3.370667,3.8498464,4.535795,5.5532312,6.885744,8.362667,9.449026,10.085744,10.548513,10.965334,11.306667,12.99036,14.851283,16.265848,17.017437,17.273438,19.006361,21.556515,24.815592,28.130465,30.290054,32.229748,35.37067,39.742363,45.331696,52.09272,59.821953,67.72185,74.079185,76.859085,73.69846,66.04472,59.214775,53.251286,48.84021,47.300926,47.13026,46.749542,45.938877,44.691696,43.2279,41.409645,40.119797,39.75549,39.54872,37.58277,35.554462,33.86749,32.15426,30.027489,27.083488,24.946875,23.46995,22.09149,21.19877,22.12431,21.832207,20.17477,17.746052,15.179488,13.154463,0.0,0.0,0.0,0.0032820515,0.02297436,0.068923086,0.7122052,0.83035904,0.56451285,0.16738462,0.02297436,0.072205134,0.08205129,0.055794876,0.029538464,0.04594872,0.1148718,0.37415388,0.80738467,0.9944616,0.13456412,0.029538464,0.01969231,0.032820515,0.055794876,0.12143591,0.02297436,0.0,0.016410258,0.101743594,0.35446155,0.18051283,0.055794876,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.029538464,0.07548718,0.07548718,0.016410258,0.013128206,2.2383592,5.8847184,7.1909747,3.9023592,3.7316926,4.2338467,4.125539,3.2623591,2.1234872,1.0896411,0.37743592,0.04594872,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01969231,0.03938462,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.029538464,0.032820515,0.009846155,0.029538464,0.108307704,0.33805132,0.7056411,1.1651284,1.6410258,2.0020514,2.2580514,2.4418464,2.550154,2.5600002,2.3893335,2.1136413,1.785436,1.4309745,1.0568206,0.65969235,0.33476925,0.11158975,0.0,0.0,0.0,0.0,0.0,0.006564103,0.036102567,0.04594872,0.032820515,0.04266667,0.14769232,0.43323082,0.6498462,0.9878975,1.2242053,1.2340513,1.0108719,0.9189744,0.9911796,1.017436,0.9321026,0.8008206,0.6301539,0.47589746,0.37743592,0.34133336,0.30851284,0.39712822,0.41682056,0.26912823,0.055794876,0.09189744,0.18051283,0.40369233,0.77456415,1.2832822,1.9003079,1.0404103,0.53825647,0.27897438,0.17066668,0.13784617,0.28225642,0.19364104,0.06564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.10502565,0.36758977,0.8008206,1.1684103,1.2931283,1.083077,0.6695385,0.4201026,0.39712822,0.30851284,0.24943592,0.24287182,0.26584616,0.40369233,1.3915899,2.9472823,5.169231,8.54318,10.8996935,8.260923,5.139693,3.8498464,4.519385,7.2861543,12.859077,15.796514,15.812924,17.782156,17.778873,14.299898,13.098668,15.14995,16.640001,12.691693,10.410667,9.051898,8.4283085,8.904206,10.873437,12.3306675,14.211283,15.849027,14.972719,14.569027,13.564719,13.377642,13.46954,11.362462,8.457847,9.504821,11.749744,12.681848,10.043077,7.0367184,7.059693,7.778462,7.637334,5.87159,5.277539,7.7259493,11.08677,13.105232,11.405129,9.271795,7.509334,6.6822567,7.017026,8.392206,8.470975,8.595693,8.900924,9.701744,11.510155,15.264822,19.682463,21.53354,20.138668,17.375181,18.28431,20.555489,19.508514,14.6871805,9.8592825,13.239796,13.344822,12.872206,13.896206,17.844515,13.220103,9.025641,6.1505647,4.7294364,4.1714873,4.6276927,6.6067696,8.4972315,9.95118,11.871181,13.206975,12.133744,11.257437,12.356924,16.390566,17.683693,16.505438,13.712411,10.696206,9.3768215,9.035488,9.554052,9.993847,9.90195,9.29477,8.989539,8.858257,8.786052,8.65477,8.339693,7.50277,6.363898,5.4482055,4.8705645,4.3290257,4.4077954,4.069744,3.5774362,3.1573336,2.993231,3.239385,3.2098465,3.2525132,3.4100516,3.3969233,2.3269746,1.8707694,1.4244103,1.079795,1.6180514,1.020718,0.35774362,0.016410258,0.016410258,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0032820515,0.0032820515,0.0032820515,0.0032820515,0.0032820515,0.013128206,0.016410258,0.016410258,0.013128206,0.0032820515,0.0032820515,0.009846155,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.01969231,0.026256412,0.026256412,0.03938462,0.04594872,0.04594872,0.04594872,0.04594872,0.06235898,0.11158975,0.15425642,0.16738462,0.13456412,0.12143591,0.15097436,0.18379489,0.23302566,0.35774362,0.25928208,0.18707694,0.19692309,0.25928208,0.24943592,0.23958977,0.256,0.26584616,0.25928208,0.23302566,0.39056414,0.5152821,1.2603078,2.861949,5.139693,7.906462,12.173129,13.124924,10.482873,8.500513,5.7796926,5.0871797,5.937231,6.521436,3.7284105,3.9187696,4.57518,4.4373336,3.7054362,4.0336413,5.8912826,6.7314878,6.518154,5.602462,4.70318,5.395693,4.525949,4.4898467,4.893539,2.546872,1.6705642,1.148718,0.64000005,0.14769232,0.02297436,0.013128206,0.006564103,0.013128206,0.026256412,0.029538464,0.03938462,0.04266667,0.03938462,0.036102567,0.029538464,0.01969231,0.016410258,0.036102567,0.07876924,0.14441027,0.098461546,0.052512825,0.026256412,0.026256412,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.013128206,0.006564103,0.18379489,0.46276927,0.512,0.13128206,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.029538464,0.049230773,0.06564103,0.1148718,0.17394873,0.24943592,0.3446154,0.47261542,0.764718,1.0568206,1.4506668,2.0020514,2.737231,3.2918978,3.8728209,4.5128207,5.2545643,6.163693,7.240206,8.109949,8.92718,9.711591,10.368001,11.073642,12.068104,13.039591,13.718975,13.866668,13.892924,15.015386,16.971489,19.51836,22.452515,23.952412,25.32759,27.510157,31.34031,37.56636,44.60308,51.59057,59.152416,67.551186,76.701546,80.30852,77.312004,69.74688,60.0878,51.245953,49.568825,48.60062,48.19036,47.95077,47.268105,46.444313,45.32513,44.18298,43.073643,41.829746,38.193233,36.12554,35.203285,34.31713,31.635695,29.305439,27.375591,25.878977,24.756516,23.857233,22.600206,19.872822,16.932104,14.480412,12.678565,0.0,0.0,0.006564103,0.006564103,0.0032820515,0.013128206,0.3446154,0.39712822,0.27569234,0.118153855,0.08533334,0.318359,0.44307697,0.33805132,0.08861539,0.0,0.013128206,0.14112821,0.33805132,0.40697438,0.013128206,0.0032820515,0.006564103,0.01969231,0.032820515,0.06235898,0.013128206,0.0,0.006564103,0.032820515,0.09189744,0.055794876,0.01969231,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.032820515,0.072205134,0.08861539,0.04594872,0.4397949,0.9944616,2.7175386,4.7917953,4.568616,2.4352822,2.8553848,3.6332312,3.5544617,2.3827693,1.332513,0.5316923,0.11158975,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.01969231,0.0,0.0,0.0,0.0,0.036102567,0.17394873,0.23958977,0.14112821,0.03938462,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.026256412,0.12143591,0.318359,0.6235898,1.0502565,1.4539489,1.7427694,1.9200002,2.0118976,2.034872,1.9528207,1.8215386,1.6443079,1.4244103,1.148718,0.8566154,0.5513847,0.27897438,0.08861539,0.009846155,0.0032820515,0.0,0.0032820515,0.009846155,0.013128206,0.01969231,0.016410258,0.04266667,0.07548718,0.03938462,0.11158975,0.40369233,0.73517954,1.2373334,2.353231,2.537026,1.847795,1.1979488,0.9747693,1.020718,0.9353847,0.86974365,0.90256417,0.97805136,0.8992821,0.7056411,0.49887183,0.27897438,0.12471796,0.21661541,0.22646156,0.20676924,0.24287182,0.44964105,0.95835906,0.69251287,0.5284103,0.49887183,0.5349744,0.46933338,0.5152821,0.39712822,0.20020515,0.029538464,0.0,0.013128206,0.02297436,0.026256412,0.032820515,0.055794876,0.06235898,0.052512825,0.06564103,0.13784617,0.32820517,0.53825647,0.64000005,0.6432821,0.57764107,0.5021539,0.36758977,0.24615386,0.15425642,0.0951795,0.06235898,0.128,0.7384616,1.9954873,3.817026,5.904411,6.3245134,4.768821,3.2065644,2.7470772,3.623385,6.012718,9.7903595,12.432411,14.381949,19.02277,21.047796,18.471386,16.584206,17.050259,17.906874,14.129231,12.163283,11.270565,11.690667,14.611693,18.838976,18.477951,16.879591,15.58318,14.316309,14.257232,15.415796,16.249437,15.96718,14.529642,11.053949,11.290257,14.250668,17.30954,16.226463,11.684103,10.755282,10.410667,9.357129,8.011488,8.891078,10.233437,10.95877,10.71918,9.885539,8.297027,7.4043083,7.4075904,8.149334,9.117539,7.4863596,6.678975,7.3649235,9.55077,12.563693,15.809642,18.33354,20.276514,21.02154,19.2,16.662975,15.963899,13.929027,10.325335,7.8506675,11.605334,12.100924,11.85477,12.297847,13.774771,9.764103,6.918565,5.792821,5.910975,5.7764106,6.0192823,7.4929237,9.009232,10.131693,11.162257,12.041847,10.79795,9.117539,8.572719,10.594462,12.763899,13.318565,12.176412,10.390975,10.131693,10.226872,10.870154,11.464206,11.651283,11.32636,10.033232,9.045334,8.3593855,7.7718983,6.885744,5.5729237,5.031385,4.6211286,4.197744,4.1091285,3.4198978,3.18359,3.0818465,2.989949,2.9801028,2.7602053,2.4155898,2.353231,2.5173335,2.3729234,1.2800001,0.6235898,0.28882053,0.26584616,0.64000005,0.39712822,0.14441027,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.013128206,0.016410258,0.016410258,0.013128206,0.009846155,0.009846155,0.013128206,0.016410258,0.016410258,0.02297436,0.016410258,0.016410258,0.026256412,0.04266667,0.049230773,0.052512825,0.049230773,0.04594872,0.049230773,0.06564103,0.09189744,0.1148718,0.13128206,0.13784617,0.118153855,0.12471796,0.13456412,0.15097436,0.18379489,0.25271797,0.20020515,0.15097436,0.15753847,0.21333335,0.23630771,0.25271797,0.24287182,0.24943592,0.25928208,0.21989745,0.23302566,0.27897438,0.65641034,1.7788719,4.1517954,8.887795,12.599796,13.364513,11.080206,7.4469748,6.189949,5.7009234,5.7009234,5.3005133,3.0096412,4.519385,5.034667,4.844308,4.571898,5.156103,7.2336416,6.705231,5.618872,4.775385,3.7349746,3.498667,2.7273848,2.4943593,2.5304618,1.2406155,0.62030774,0.45620516,0.31507695,0.09189744,0.02297436,0.02297436,0.016410258,0.013128206,0.013128206,0.006564103,0.009846155,0.013128206,0.016410258,0.01969231,0.013128206,0.006564103,0.013128206,0.013128206,0.006564103,0.013128206,0.01969231,0.02297436,0.02297436,0.01969231,0.016410258,0.009846155,0.009846155,0.009846155,0.006564103,0.0,0.0032820515,0.006564103,0.12143591,0.38728207,0.76800007,0.6235898,0.45292312,0.21989745,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.02297436,0.032820515,0.04594872,0.068923086,0.0951795,0.118153855,0.14769232,0.20676924,0.318359,0.58420515,0.8960001,1.3193847,2.0939488,2.6322052,3.1540515,3.6332312,4.161641,4.97559,5.8157954,6.5411286,7.3550773,8.237949,8.933744,9.38995,10.092308,10.771693,11.244308,11.405129,10.86359,10.834052,11.460924,12.964104,15.648822,17.545847,19.452719,21.267694,23.207386,25.80677,31.232002,37.858463,45.59426,54.15713,63.071186,70.91529,76.18298,78.66093,77.52206,71.32555,63.78339,57.206158,52.8279,50.898056,50.688004,50.41231,49.942978,49.24062,48.39385,47.62585,44.865646,42.28267,40.034466,37.933952,35.439594,34.070976,32.856617,31.22872,29.213541,27.441233,26.128412,22.95795,20.079592,18.235079,16.761436,0.0,0.009846155,0.026256412,0.02297436,0.0032820515,0.0,0.02297436,0.059076928,0.08205129,0.12471796,0.2855385,0.48574364,0.50543594,0.34789747,0.12471796,0.08533334,0.04266667,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.013128206,0.032820515,0.072205134,0.08533334,0.06235898,0.026256412,0.6859488,2.4976413,3.0424619,1.9954873,1.1454359,0.7450257,1.2964103,1.8412309,1.8051283,1.017436,0.62030774,0.27897438,0.08861539,0.036102567,0.0,0.0,0.013128206,0.013128206,0.0,0.0,0.013128206,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.036102567,0.17394873,0.23958977,0.14112821,0.03938462,0.009846155,0.04266667,0.055794876,0.02297436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03938462,0.16410258,0.38400003,0.67610264,0.9517949,1.2242053,1.4178462,1.5097437,1.529436,1.4605129,1.3718976,1.2635899,1.1323078,0.96492314,0.78769237,0.574359,0.3511795,0.15097436,0.026256412,0.006564103,0.0,0.0032820515,0.009846155,0.013128206,0.009846155,0.009846155,0.036102567,0.068923086,0.032820515,0.013128206,0.101743594,0.28882053,0.8041026,2.1202054,2.7306669,2.28759,1.7624617,1.5655385,1.5425643,1.3292309,1.1060513,1.0765129,1.1815386,1.1093334,0.90256417,0.761436,0.574359,0.45292312,0.7220513,0.8730257,0.6629744,0.4266667,0.34133336,0.4201026,0.4201026,0.4594872,0.56451285,0.6629744,0.5874872,0.6892308,0.6826667,0.44964105,0.12143591,0.06564103,0.08533334,0.08205129,0.108307704,0.17066668,0.23302566,0.14769232,0.1148718,0.09189744,0.07876924,0.10502565,0.09189744,0.13128206,0.2855385,0.512,0.65641034,0.58420515,0.41682056,0.21661541,0.07876924,0.128,0.25928208,0.41682056,0.9419488,1.7558975,2.3466668,1.9035898,1.7066668,1.6213335,1.7362052,2.3663592,4.1485133,5.989744,8.576,12.580104,18.668308,20.434053,18.46154,15.960617,14.647796,14.752822,13.699283,13.761642,14.437745,15.711181,18.048002,19.698874,18.271181,16.505438,15.51754,14.79877,15.451899,16.692514,17.040411,16.41354,16.128002,12.534155,10.788103,12.550565,15.91795,15.415796,12.553847,11.523283,10.699488,9.885539,10.312206,9.91836,8.684308,7.4797955,7.2237954,8.891078,10.601027,11.808822,11.825232,10.81436,9.819899,7.64718,7.6242056,9.019077,10.925949,12.265027,12.340514,12.117334,13.974976,16.876308,16.38072,12.665437,11.116308,9.83959,8.474257,8.172308,9.409642,9.77395,10.029949,10.262975,9.856001,7.702975,6.741334,6.76759,7.174565,6.961231,6.928411,7.3353853,7.890052,8.388924,8.710565,9.110975,8.576,7.4896417,6.4656415,6.370462,8.119796,9.718155,10.256411,9.961026,10.180923,10.167795,10.541949,11.001437,11.218052,10.843898,9.051898,7.6603084,6.7117953,6.009436,5.113436,4.027077,3.882667,3.8432825,3.6430771,3.5872824,2.8127182,2.7700515,2.8947694,2.9013336,2.7569232,2.176,1.7394873,1.5327181,1.467077,1.2865642,0.58092314,0.20348719,0.055794876,0.032820515,0.055794876,0.068923086,0.03938462,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.009846155,0.009846155,0.009846155,0.009846155,0.009846155,0.009846155,0.013128206,0.016410258,0.02297436,0.02297436,0.016410258,0.02297436,0.036102567,0.049230773,0.055794876,0.049230773,0.04266667,0.03938462,0.04266667,0.059076928,0.0951795,0.108307704,0.11158975,0.11158975,0.11158975,0.13128206,0.14112821,0.15097436,0.16082053,0.16738462,0.16738462,0.16082053,0.17066668,0.19364104,0.21661541,0.24943592,0.24615386,0.24615386,0.24287182,0.19692309,0.20348719,0.20676924,0.39056414,1.1290257,2.9735386,8.464411,11.638155,13.033027,12.507898,9.252103,8.303591,7.1089234,6.0849237,5.4843082,5.395693,5.9634876,5.8157954,5.0543594,4.4800005,5.609026,6.370462,5.477744,4.128821,2.92759,1.8609232,1.4539489,1.3489232,1.2504616,0.96492314,0.4135385,0.118153855,0.13784617,0.13784617,0.036102567,0.02297436,0.032820515,0.02297436,0.016410258,0.013128206,0.0,0.0,0.0,0.0032820515,0.006564103,0.0,0.0,0.006564103,0.006564103,0.0,0.0,0.02297436,0.01969231,0.013128206,0.009846155,0.009846155,0.013128206,0.016410258,0.016410258,0.013128206,0.0,0.0,0.006564103,0.029538464,0.15425642,0.512,0.55794877,0.446359,0.21989745,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.006564103,0.006564103,0.006564103,0.016410258,0.026256412,0.03938462,0.09189744,0.20020515,0.28882053,0.36758977,0.512,0.45620516,0.571077,0.73517954,0.9616411,1.4112822,1.8970258,2.409026,2.9013336,3.4166157,4.076308,4.713026,5.3005133,5.9569235,6.698667,7.450257,7.64718,8.146052,8.65477,8.887795,8.579283,8.628513,8.211693,8.021334,8.55959,10.138257,11.923694,14.188309,16.633438,18.868515,20.434053,23.066257,27.152412,32.961643,39.955696,46.798775,54.9678,63.970467,72.71057,79.32719,81.16842,77.2759,71.59795,65.48677,60.064827,56.25108,54.068516,52.90339,52.063183,51.28862,50.737236,49.772312,48.098465,45.748516,42.909542,39.94913,39.184414,38.34749,36.466873,33.929848,32.495594,31.182772,27.976208,26.105438,26.25313,26.548515,0.0,0.01969231,0.03938462,0.049230773,0.04266667,0.02297436,0.03938462,0.13128206,0.17066668,0.20348719,0.4594872,0.40697438,0.17394873,0.036102567,0.072205134,0.17066668,0.072205134,0.01969231,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.036102567,0.06235898,0.06564103,0.07548718,0.08533334,0.10502565,0.17723078,0.380718,1.2603078,3.9384618,3.4166157,0.17066668,0.16410258,0.42994875,0.35446155,0.20676924,0.12143591,0.1148718,0.18379489,0.16410258,0.11158975,0.059076928,0.0,0.0,0.03938462,0.03938462,0.0,0.0,0.029538464,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01969231,0.0951795,0.118153855,0.049230773,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03938462,0.15425642,0.3249231,0.446359,0.5152821,0.7450257,0.9714873,1.1093334,1.142154,1.0568206,0.9517949,0.8369231,0.7220513,0.60389745,0.512,0.40697438,0.27569234,0.13456412,0.03938462,0.013128206,0.0032820515,0.006564103,0.01969231,0.04594872,0.036102567,0.036102567,0.04594872,0.049230773,0.036102567,0.016410258,0.009846155,0.0032820515,0.03938462,0.19692309,0.9485129,1.4572309,1.7558975,1.8412309,1.6836925,1.1815386,0.7515898,0.5940513,0.65312827,0.6235898,0.5940513,0.7384616,0.77128214,0.79097444,1.2800001,1.6804104,1.3128207,0.85005134,0.5874872,0.47589746,0.47917953,0.58420515,0.69251287,0.7515898,0.761436,1.2635899,1.4703591,1.2274873,0.7417436,0.58420515,0.58420515,0.51856416,0.5284103,0.6104616,0.63343596,0.32820517,0.27241027,0.3446154,0.4397949,0.46933338,0.3249231,0.26912823,0.34133336,0.5218462,0.7187693,0.7581539,0.5415385,0.26912823,0.13456412,0.3249231,0.5940513,0.6826667,0.7417436,0.81066674,0.82379496,0.86646163,1.2635899,1.5163078,1.4966155,1.4539489,2.5238976,4.0303593,7.1056414,11.756309,16.876308,15.737437,13.180719,10.331899,8.4053335,8.710565,12.012309,14.171899,15.287796,15.474873,14.8709755,12.928001,13.095386,14.795488,16.79754,17.237335,18.100513,16.90913,15.58318,14.897232,14.496821,11.319796,8.763078,9.045334,11.011283,10.118565,10.089026,9.626257,9.281642,9.485129,10.532104,7.532308,5.648411,5.861744,8.169026,11.588924,15.455181,16.70236,15.356719,12.452104,10.010257,9.301334,10.883283,12.504617,12.977232,12.153437,8.887795,6.7971287,7.857231,10.883283,11.516719,9.544206,8.999385,8.753231,8.5202055,8.835282,9.5146675,11.431385,12.58995,12.081232,10.102155,7.6307697,6.557539,6.419693,6.669129,6.672411,6.701949,6.5903597,6.196513,5.730462,5.723898,6.1997952,6.9710774,7.328821,7.0104623,6.2194877,6.7774363,8.28718,9.573745,9.990565,9.449026,8.4972315,8.254359,8.306872,8.192,7.4108725,5.924103,4.7524104,4.007385,3.5840003,3.1803079,2.937436,2.7766156,2.789744,2.8127182,2.4352822,2.1497438,2.176,2.2678976,2.1825643,1.6640002,1.204513,1.0535386,0.8041026,0.40697438,0.18379489,0.06235898,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.02297436,0.029538464,0.01969231,0.01969231,0.032820515,0.04266667,0.04594872,0.049230773,0.036102567,0.032820515,0.032820515,0.029538464,0.032820515,0.06235898,0.0951795,0.108307704,0.11158975,0.1148718,0.128,0.14441027,0.16410258,0.18707694,0.19692309,0.20348719,0.21333335,0.21661541,0.21661541,0.20020515,0.21661541,0.2100513,0.19364104,0.17394873,0.16738462,0.14769232,0.13456412,0.256,0.7778462,2.1136413,6.5247183,10.226872,12.737642,13.8075905,13.4400015,11.201642,9.065026,7.706257,7.581539,8.923898,6.6592827,5.730462,4.8738465,4.164923,5.0182567,3.6562054,3.045744,1.9331284,0.4660513,0.19364104,0.83035904,1.3128207,1.214359,0.5973334,0.0032820515,0.013128206,0.029538464,0.032820515,0.02297436,0.013128206,0.032820515,0.02297436,0.013128206,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.006564103,0.016410258,0.04594872,0.036102567,0.01969231,0.009846155,0.0,0.009846155,0.016410258,0.016410258,0.013128206,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.009846155,0.016410258,0.026256412,0.026256412,0.026256412,0.026256412,0.049230773,0.1148718,0.23958977,0.5546667,0.88943595,1.1684103,1.4178462,1.7591796,1.5589745,1.522872,1.5261539,1.4802053,1.3554872,1.6344616,1.9889232,2.4615386,2.986667,3.3936412,3.95159,4.4996924,4.9460516,5.395693,6.1374364,5.8781543,6.0783596,6.419693,6.419693,5.4449234,6.2194877,6.1374364,5.989744,6.091488,6.2851286,7.1483083,8.677744,11.451077,15.212309,18.888206,19.80718,20.647387,23.122053,27.749746,33.847797,40.64821,47.734158,55.32226,63.583183,72.65478,79.75057,82.01847,79.625854,73.728004,66.44842,60.911594,57.219288,54.580517,52.640823,51.475697,51.360825,51.282055,50.30072,48.078773,44.868927,44.084515,42.902977,40.86154,38.73149,38.528004,37.00841,34.225235,35.236107,40.077133,43.75303,0.0,0.0,0.0,0.072205134,0.16738462,0.108307704,0.0951795,0.13784617,0.16082053,0.15425642,0.16738462,0.19364104,0.08861539,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.055794876,0.15097436,0.23630771,0.19692309,0.052512825,0.02297436,0.24287182,0.7975385,1.723077,3.7743592,4.6080003,2.8914874,0.01969231,0.09189744,0.14112821,0.1148718,0.055794876,0.04266667,0.21333335,0.1148718,0.118153855,0.08205129,0.0,0.0,0.0,0.055794876,0.055794876,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.04594872,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.009846155,0.006564103,0.029538464,0.14112821,0.34133336,0.5973334,0.8369231,0.94523084,0.90912825,0.80738467,0.65641034,0.48246157,0.33476925,0.26256412,0.19692309,0.12471796,0.052512825,0.016410258,0.026256412,0.02297436,0.032820515,0.068923086,0.108307704,0.15425642,0.18707694,0.19692309,0.18379489,0.12143591,0.072205134,0.04266667,0.01969231,0.0,0.0,0.0,0.0,0.072205134,0.34133336,0.97805136,0.36758977,0.12143591,0.04266667,0.013128206,0.0,0.0,0.036102567,0.20020515,0.54482055,1.083077,1.5721027,1.529436,1.3522053,1.2209232,1.0994873,1.3554872,1.585231,1.7296412,1.8215386,1.9692309,3.1770258,3.5413337,3.3247182,2.793026,2.2416413,2.1956925,2.0086155,1.8313848,1.6738462,1.404718,0.8041026,0.7581539,1.1355898,1.6180514,1.6771283,1.0075898,0.47261542,0.20348719,0.18379489,0.24287182,0.14769232,0.07548718,0.08205129,0.21661541,0.5349744,0.98461545,1.024,0.78769237,0.46933338,0.33476925,0.36102566,0.64000005,0.92225647,1.0371283,0.9156924,1.6836925,3.7907696,7.072821,10.259693,10.955488,9.114257,6.564103,5.405539,6.5870776,9.91836,16.521847,17.046976,13.147899,7.962257,6.121026,8.316719,11.474052,13.226667,13.856822,16.295385,16.856617,15.681643,15.199181,15.107284,12.360206,8.979693,8.507077,10.095591,12.317539,13.184001,11.18195,9.895386,9.563898,9.055181,5.8453336,6.124308,10.121847,13.607386,14.834873,14.54277,13.466257,10.463181,8.477539,8.129642,7.6898465,10.935796,11.82195,11.224616,10.637129,12.176412,8.648206,7.0990777,7.200821,7.939283,7.5979495,7.8441033,7.381334,7.4075904,8.310155,9.688616,14.693745,24.769644,28.75077,23.663591,14.739694,7.90318,5.0510774,4.4340515,4.841026,5.586052,5.681231,5.6976414,5.330052,4.772103,4.699898,5.5663595,6.698667,7.522462,7.8670774,7.965539,7.965539,8.385642,8.897642,8.973129,7.8736415,6.5444107,5.7698464,5.028103,4.0533338,2.868513,2.1234872,1.6443079,1.2800001,1.0568206,1.1913847,1.7887181,2.0217438,2.0578463,1.9593848,1.6771283,1.6180514,1.5753847,1.3620514,1.017436,0.80738467,0.6629744,0.3708718,0.118153855,0.02297436,0.12143591,0.15753847,0.06564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.02297436,0.036102567,0.04266667,0.029538464,0.029538464,0.029538464,0.036102567,0.049230773,0.06235898,0.049230773,0.04594872,0.03938462,0.032820515,0.04594872,0.04594872,0.055794876,0.06235898,0.06564103,0.09189744,0.10502565,0.13456412,0.190359,0.25928208,0.32164106,0.3446154,0.3511795,0.3314872,0.2855385,0.21333335,0.190359,0.17394873,0.15425642,0.14441027,0.16738462,0.118153855,0.068923086,0.108307704,0.4660513,1.5425643,3.3247182,7.8080006,12.12718,15.199181,17.700104,14.171899,12.87877,11.316514,9.301334,8.973129,6.9809237,6.0258465,6.550975,7.5421543,6.5312824,3.8334363,1.8773335,0.7056411,0.27897438,0.47261542,0.92553854,0.86317956,0.79097444,0.6859488,0.016410258,0.016410258,0.016410258,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01969231,0.029538464,0.03938462,0.07548718,0.07548718,0.06564103,0.06235898,0.049230773,0.0,0.0,0.01969231,0.02297436,0.016410258,0.016410258,0.016410258,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.026256412,0.049230773,0.06235898,0.06564103,0.07548718,0.07548718,0.11158975,0.2297436,0.50543594,1.0666667,2.2153847,2.934154,3.498667,4.017231,4.394667,4.322462,4.420923,4.2568207,3.7710772,3.2951798,2.8914874,2.5632823,2.605949,3.0162053,3.4789746,4.027077,4.4406157,4.6539493,4.7589746,4.9887185,4.4274874,4.3716927,4.3585644,4.089436,3.4166157,2.989949,3.387077,4.2863593,5.0149746,4.562052,4.4406157,4.7589746,5.802667,8.096821,12.406155,17.496616,20.059898,20.273232,19.86954,22.14072,27.181952,33.48021,40.658054,48.301952,55.955696,63.120415,69.90113,76.530876,81.87734,83.46585,77.177444,69.983185,63.504414,58.459904,54.688824,52.355286,51.478977,50.504208,49.092926,48.141132,47.678364,46.19816,44.629337,43.897438,44.93785,43.33621,41.764107,49.030567,63.005543,70.64616,0.08533334,0.06564103,0.02297436,0.013128206,0.032820515,0.02297436,0.01969231,0.026256412,0.04266667,0.068923086,0.13128206,0.118153855,0.15097436,0.27897438,0.446359,0.47589746,0.318359,0.128,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.032820515,0.06235898,0.07548718,0.08861539,0.049230773,0.04266667,0.9189744,2.5665643,3.8859491,2.428718,1.404718,0.5940513,0.072205134,0.21333335,0.06564103,0.029538464,0.052512825,0.08205129,0.06564103,0.5546667,0.4135385,0.14112821,0.0,0.0,0.0,0.009846155,0.026256412,0.055794876,0.13456412,0.026256412,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.072205134,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.006564103,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0,0.006564103,0.03938462,0.12471796,0.26912823,0.44964105,0.6170257,0.6859488,0.69251287,0.6104616,0.45292312,0.2855385,0.19364104,0.14112821,0.0951795,0.055794876,0.03938462,0.072205134,0.09189744,0.10502565,0.10502565,0.08205129,0.072205134,0.059076928,0.14441027,0.29210258,0.318359,0.12143591,0.09189744,0.07548718,0.032820515,0.013128206,0.013128206,0.013128206,0.02297436,0.072205134,0.20676924,0.0951795,0.032820515,0.009846155,0.0032820515,0.0,0.0,0.006564103,0.03938462,0.14441027,0.4004103,0.7417436,1.2570257,1.3259488,0.99774367,0.96492314,1.2898463,1.8576412,2.097231,1.9265642,1.7624617,3.0949745,3.9712822,4.2469745,4.1583595,4.2830772,4.778667,5.287385,5.3234878,4.8836927,4.417641,3.4494362,3.1015387,3.314872,3.8038976,4.069744,3.7120004,2.4648206,1.5064616,1.2832822,1.4998976,1.1290257,1.0502565,1.014154,1.0568206,1.5097437,4.138667,6.0291286,5.8420515,3.7842054,1.5688206,0.7811283,0.4201026,0.34133336,0.58420515,1.3784616,3.1737437,5.3891287,7.817847,9.800206,10.223591,9.065026,8.297027,8.884514,11.464206,16.338053,14.985847,9.301334,5.435077,5.2676926,6.422975,9.02236,10.729027,12.07795,13.216822,13.892924,15.29436,16.97477,16.666258,13.919181,10.138257,12.675283,14.342566,14.372104,13.51877,14.063591,12.274873,9.69518,7.768616,6.4754877,4.3290257,8.234667,11.080206,11.634872,10.312206,9.170052,8.214975,6.636308,6.491898,8.910769,14.086565,13.673027,10.676514,7.6898465,6.3540516,7.3550773,7.529026,8.749949,9.573745,9.350565,8.208411,7.6635904,6.997334,7.181129,8.198565,9.042052,16.177233,28.160002,31.291079,22.54113,9.563898,6.0192823,4.634257,4.3585644,4.3749747,4.096,4.1747694,4.7622566,5.113436,5.228308,5.858462,6.8233852,7.9885135,8.851693,8.884514,7.5388722,6.738052,5.98318,5.8289237,6.048821,5.651693,5.044513,4.2240005,3.1442053,2.0545642,1.5261539,1.3587693,1.5786668,1.5458462,1.4112822,2.1300514,2.4451284,2.2678976,1.7920002,1.2800001,1.0666667,0.65641034,0.47261542,0.35774362,0.25271797,0.2100513,0.14112821,0.07548718,0.02297436,0.04266667,0.20676924,0.128,0.08533334,0.04266667,0.013128206,0.072205134,0.09189744,0.03938462,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.016410258,0.12471796,0.48246157,0.18051283,0.07548718,0.06235898,0.072205134,0.08533334,0.06235898,0.049230773,0.049230773,0.052512825,0.04594872,0.036102567,0.049230773,0.06564103,0.08533334,0.14112821,0.14441027,0.16410258,0.2100513,0.25928208,0.27241027,0.23630771,0.23630771,0.24287182,0.23958977,0.22646156,0.190359,0.17394873,0.15097436,0.12471796,0.13128206,0.12143591,0.098461546,0.108307704,0.27241027,0.761436,2.3860514,5.87159,9.780514,13.223386,15.832617,12.842668,13.952001,12.36677,7.719385,6.091488,5.2348723,5.7632823,5.7698464,5.0051284,4.8705645,2.2613335,0.8402052,0.2986667,0.41682056,1.0699488,1.404718,0.8533334,0.3314872,0.15097436,0.016410258,0.016410258,0.016410258,0.013128206,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.049230773,0.11158975,0.19692309,0.23630771,0.2297436,0.18707694,0.118153855,0.049230773,0.049230773,0.03938462,0.01969231,0.0032820515,0.0032820515,0.0032820515,0.009846155,0.04594872,0.21661541,0.69579494,0.38400003,0.128,0.032820515,0.18707694,0.69907695,1.1618463,1.3686155,1.404718,1.3522053,1.2832822,1.5983591,2.1300514,2.7963078,3.6168208,4.706462,6.741334,8.096821,8.828718,9.357129,10.499283,10.610872,10.171078,9.268514,7.9917955,6.419693,6.1046157,5.7107697,5.175795,4.601436,4.2371287,3.7710772,4.0533338,4.3060517,4.315898,4.4406157,4.082872,3.95159,3.764513,3.3345644,2.5764105,2.7142565,2.8291285,3.2361028,3.7185643,3.501949,3.4166157,3.2328207,3.5577438,4.6539493,6.422975,9.337437,13.019898,16.89272,19.88595,20.407797,20.545643,22.86277,26.93908,32.278976,38.304825,46.690464,56.10667,64.9879,71.35508,72.78606,74.68308,77.72226,78.23754,74.93908,68.9198,63.570057,60.212517,57.711594,55.141747,51.7678,49.125748,47.422363,46.742977,47.169643,48.78113,48.160824,49.85108,62.336006,79.24513,79.32719,0.28882053,0.18379489,0.06235898,0.0,0.0,0.0,0.036102567,0.036102567,0.02297436,0.01969231,0.049230773,0.03938462,0.06564103,0.14769232,0.24615386,0.27569234,0.190359,0.07876924,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.01969231,0.029538464,0.0,0.0,0.0,0.0,0.0032820515,0.01969231,0.009846155,0.04266667,0.04266667,0.04266667,0.17066668,0.28225642,0.702359,2.4713848,4.338872,2.7667694,1.079795,0.2855385,0.032820515,0.04266667,0.098461546,0.01969231,0.0032820515,0.01969231,0.036102567,0.013128206,0.27241027,0.2855385,0.19692309,0.21661541,0.60389745,0.128,0.009846155,0.013128206,0.029538464,0.06564103,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.036102567,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.032820515,0.16410258,0.032820515,0.0032820515,0.06564103,0.12471796,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.032820515,0.09189744,0.18379489,0.31507695,0.4397949,0.50543594,0.48902568,0.42994875,0.4135385,0.24943592,0.14769232,0.08205129,0.03938462,0.026256412,0.09189744,0.128,0.13456412,0.10502565,0.03938462,0.029538464,0.013128206,0.052512825,0.128,0.14769232,0.052512825,0.09189744,0.12143591,0.098461546,0.06235898,0.04594872,0.036102567,0.029538464,0.026256412,0.02297436,0.052512825,0.06235898,0.049230773,0.02297436,0.0,0.0,0.0,0.0,0.01969231,0.09189744,0.2297436,0.52512825,0.5907693,0.42994875,0.446359,0.69251287,1.0732309,1.1749744,0.9682052,0.81066674,1.585231,2.3729234,2.8750772,3.0194874,2.9604106,2.7733335,3.045744,3.2951798,3.3772311,3.4888208,2.733949,2.3630772,2.5107694,2.9702566,3.1770258,3.2623591,3.2787695,3.4297438,3.7284105,4.020513,3.9056413,3.4592824,2.8389745,2.5600002,3.495385,7.069539,9.005949,9.094564,7.5881033,5.1922054,2.9144619,1.2242053,0.76800007,1.6443079,3.4100516,3.9220517,5.4186673,7.4797955,9.147078,8.914052,8.320001,9.078155,9.997129,10.262975,9.43918,7.0990777,5.034667,4.768821,6.2687182,7.936001,11.126155,11.634872,11.861334,12.422565,12.163283,14.011078,16.09518,15.547078,12.356924,9.363693,11.431385,14.267078,15.474873,14.523078,12.754052,13.026463,11.815386,9.140513,6.042257,4.565334,7.450257,8.73354,9.02236,8.759795,8.241231,10.108719,10.883283,10.35159,9.498257,10.505847,9.019077,6.705231,4.893539,4.2240005,4.6572313,5.2644105,6.3540516,7.3747697,8.03118,8.27077,8.067283,8.146052,8.612103,9.222565,9.366975,12.265027,16.62031,16.610462,11.480617,5.533539,4.342154,3.7874875,3.564308,3.4789746,3.43959,3.8728209,4.8082056,5.297231,5.290667,5.664821,6.47877,6.436103,6.426257,6.5050263,5.8945646,5.221744,4.1682053,3.508513,3.3772311,3.2754874,2.92759,2.409026,1.6344616,0.9156924,0.9517949,1.1257436,1.0338463,0.9419488,1.0535386,1.4966155,1.5261539,1.1618463,0.73517954,0.446359,0.37415388,0.16738462,0.07876924,0.04266667,0.02297436,0.02297436,0.0032820515,0.0,0.0,0.01969231,0.09189744,0.049230773,0.036102567,0.02297436,0.013128206,0.06564103,0.08205129,0.032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016410258,0.101743594,0.34789747,0.3052308,0.17723078,0.098461546,0.101743594,0.101743594,0.10502565,0.108307704,0.108307704,0.10502565,0.101743594,0.101743594,0.10502565,0.09189744,0.072205134,0.098461546,0.11158975,0.12471796,0.15425642,0.20348719,0.23302566,0.21989745,0.21989745,0.23302566,0.24943592,0.256,0.22646156,0.2231795,0.20348719,0.17066668,0.15097436,0.14112821,0.12143591,0.45292312,1.1815386,2.0217438,4.2502565,8.201847,12.740924,16.515284,17.96595,13.689437,12.3536415,10.742155,8.146052,6.3606157,5.5663595,5.0149746,4.3060517,3.5413337,3.3476925,1.9889232,0.8960001,0.27569234,0.18051283,0.48902568,0.6170257,0.3511795,0.0951795,0.016410258,0.016410258,0.006564103,0.006564103,0.006564103,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.01969231,0.052512825,0.09189744,0.118153855,0.12471796,0.101743594,0.06235898,0.032820515,0.026256412,0.016410258,0.006564103,0.0,0.0,0.16082053,0.5907693,0.9517949,1.1716924,1.4112822,1.1585642,1.0305642,1.2274873,1.6640002,1.9692309,2.1169233,2.3466668,2.5895386,2.8521028,3.2065644,3.9351797,4.70318,5.5171285,6.3245134,7.0334363,9.101129,10.676514,11.69395,12.452104,13.59754,14.063591,13.945437,13.354668,12.225642,10.325335,8.704,8.103385,7.450257,6.416411,5.4416413,4.699898,4.516103,4.4077954,4.2207184,4.1189747,3.9384618,3.698872,3.18359,2.412308,1.6607181,1.6836925,1.8379488,2.1136413,2.4188719,2.5665643,2.428718,2.225231,2.3466668,2.9013336,3.7185643,5.093744,7.3714876,10.482873,13.7386675,15.845745,17.864206,19.045746,20.657232,23.072823,25.750977,30.634668,37.69108,46.372105,55.259903,62.08657,68.841034,73.51795,75.02113,73.68862,71.299286,69.42852,67.36739,65.243904,62.608414,58.466465,54.747902,51.856415,50.067696,49.631184,50.76021,51.03262,52.558773,59.55939,68.355286,67.364105,0.44964105,0.2986667,0.118153855,0.013128206,0.0,0.0,0.036102567,0.036102567,0.016410258,0.0951795,0.48246157,0.39056414,0.48902568,0.52512825,0.40697438,0.23302566,0.13128206,0.059076928,0.049230773,0.09189744,0.1148718,0.14112821,0.098461546,0.04266667,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.01969231,0.032820515,0.01969231,0.01969231,0.006564103,0.009846155,0.029538464,0.049230773,0.052512825,0.15097436,0.23630771,0.32820517,0.5907693,1.0371283,1.1126155,2.1234872,3.1376412,1.0043077,0.256,0.055794876,0.03938462,0.01969231,0.01969231,0.0032820515,0.0,0.0,0.013128206,0.06235898,0.04266667,0.118153855,0.15097436,0.23630771,0.702359,0.18707694,0.03938462,0.016410258,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.032820515,0.16410258,0.032820515,0.0,0.08533334,0.17394873,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.016410258,0.04594872,0.11158975,0.21661541,0.2855385,0.32164106,0.35446155,0.44964105,0.28882053,0.17066668,0.09189744,0.049230773,0.02297436,0.072205134,0.09189744,0.08861539,0.059076928,0.009846155,0.03938462,0.04266667,0.052512825,0.06235898,0.036102567,0.016410258,0.06235898,0.0951795,0.08861539,0.055794876,0.04594872,0.04594872,0.03938462,0.032820515,0.02297436,0.04594872,0.06564103,0.059076928,0.026256412,0.0,0.0,0.0,0.0,0.0,0.0,0.06235898,0.07548718,0.06564103,0.06235898,0.072205134,0.19692309,0.31507695,0.34133336,0.32820517,0.46276927,0.42338464,0.7450257,1.1191796,1.3062565,1.1651284,0.71548724,0.7450257,0.93866676,1.1848207,1.5458462,1.3161026,1.014154,1.0108719,1.276718,1.401436,1.7460514,2.5698464,3.3444104,3.7973337,3.9187696,3.95159,3.7120004,3.2918978,3.1507695,4.1124105,7.13518,8.418462,8.530052,7.7981544,6.314667,4.096,2.2646155,1.6738462,2.4418464,3.9581542,4.2863593,5.366154,6.6428723,7.3747697,6.633026,6.3179493,7.066257,7.5552826,6.7840004,4.066462,4.3618464,5.3005133,6.3474874,7.259898,8.067283,10.925949,10.771693,10.098872,9.783795,9.074872,10.620719,13.594257,14.158771,11.513436,7.90318,8.569437,11.956513,15.02195,15.744001,13.138052,13.305437,13.289026,10.6469755,6.2851286,4.457026,7.0367184,9.163487,10.161232,10.000411,9.288206,11.21477,11.805539,10.295795,7.4075904,5.3398976,4.516103,3.9253337,3.8629746,4.2436924,4.6145644,4.391385,4.57518,5.4186673,6.701949,7.7456417,7.781744,8.408616,9.03877,9.094564,8.024616,7.328821,6.432821,5.169231,3.948308,3.7809234,3.7218463,3.5478978,3.3476925,3.259077,3.4691284,3.7251284,4.201026,4.2994876,4.013949,3.948308,4.352,3.9187696,3.5905645,3.6660516,3.7874875,3.5052311,2.878359,2.2088206,1.7296412,1.5786668,1.4178462,1.017436,0.6301539,0.45292312,0.63343596,0.69251287,0.48902568,0.4135385,0.5415385,0.64000005,0.5152821,0.23958977,0.04266667,0.0032820515,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.026256412,0.036102567,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02297436,0.08205129,0.17066668,0.4660513,0.6268718,0.58092314,0.36430773,0.11158975,0.11158975,0.118153855,0.1148718,0.108307704,0.11158975,0.13128206,0.128,0.11158975,0.0951795,0.108307704,0.14441027,0.16082053,0.18051283,0.2100513,0.24287182,0.24615386,0.25928208,0.2855385,0.31507695,0.318359,0.2986667,0.2986667,0.28225642,0.23302566,0.16082053,0.16082053,0.33805132,0.8172308,1.7755898,3.4592824,6.262154,11.457642,16.420103,19.016207,17.631182,12.908309,9.5146675,7.6701546,6.8693337,5.8945646,5.277539,3.9023592,2.7273848,2.1202054,1.8346668,1.3850257,0.79097444,0.32820517,0.0951795,0.006564103,0.009846155,0.009846155,0.013128206,0.013128206,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.013128206,0.013128206,0.009846155,0.009846155,0.0032820515,0.0,0.0032820515,0.0032820515,0.0,0.18707694,0.7253334,1.2373334,1.5163078,1.5491283,1.5491283,1.6804104,2.2022567,3.0752823,3.945026,4.332308,4.076308,3.7973337,3.8334363,4.2568207,4.7950773,5.5269747,6.3573337,7.128616,7.6012316,9.009232,10.213744,11.057232,11.674257,12.488206,12.754052,12.511181,11.949949,11.10318,9.8363085,8.188719,7.7948723,7.5191803,6.803693,5.677949,4.821334,4.4274874,4.2338467,4.076308,3.889231,3.6693337,3.3378465,2.6354873,1.6836925,0.9878975,0.892718,1.0469744,1.2406155,1.4080001,1.6508719,1.6443079,1.6180514,1.7001027,1.975795,2.5009232,3.1540515,4.197744,5.674667,7.653744,10.230155,13.650052,15.205745,16.357744,17.578669,18.346668,20.118977,23.666874,29.476105,37.218464,45.75836,54.626465,60.800003,64.78442,67.216415,68.87057,69.57621,69.07406,67.98769,66.4517,64.101746,61.25949,58.11857,55.230362,53.287388,53.116722,53.192207,53.044518,53.937237,55.542156,55.922874,1.0404103,0.9124103,0.4004103,0.068923086,0.04266667,0.0,0.0,0.0,0.0,0.19364104,0.9682052,0.7778462,0.98133343,1.0338463,0.77456415,0.4004103,0.24287182,0.15425642,0.21661541,0.37743592,0.4660513,0.380718,0.2297436,0.09189744,0.016410258,0.032820515,0.059076928,0.052512825,0.036102567,0.02297436,0.032820515,0.04594872,0.04594872,0.026256412,0.006564103,0.036102567,0.049230773,0.049230773,0.06564103,0.11158975,0.18051283,0.4004103,0.6268718,0.76800007,0.8598975,1.0699488,1.7591796,1.083077,0.3446154,0.07876924,0.032820515,0.03938462,0.04266667,0.03938462,0.036102567,0.03938462,0.006564103,0.0,0.0,0.032820515,0.15097436,0.08533334,0.055794876,0.03938462,0.059076928,0.20020515,0.13456412,0.101743594,0.059076928,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.08861539,0.17394873,0.12143591,0.02297436,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.02297436,0.052512825,0.10502565,0.16082053,0.2231795,0.318359,0.256,0.17723078,0.118153855,0.07876924,0.032820515,0.032820515,0.01969231,0.006564103,0.0,0.0,0.059076928,0.09189744,0.12143591,0.13456412,0.108307704,0.098461546,0.072205134,0.03938462,0.013128206,0.013128206,0.02297436,0.052512825,0.055794876,0.03938462,0.04594872,0.02297436,0.02297436,0.02297436,0.013128206,0.0,0.0032820515,0.0,0.0,0.0,0.0,0.098461546,0.049230773,0.013128206,0.02297436,0.013128206,0.032820515,0.026256412,0.08533334,0.28225642,0.67282057,0.13456412,0.009846155,0.07548718,0.18707694,0.27569234,0.25271797,0.29210258,0.24943592,0.16738462,0.26912823,0.49230772,0.28225642,0.0951795,0.10502565,0.21333335,0.52512825,0.9878975,1.3259488,1.4112822,1.2570257,1.2274873,1.6180514,2.0250258,2.3663592,2.878359,4.266667,4.8016415,4.667077,4.194462,3.8695388,3.242667,2.6256413,2.28759,2.28759,2.4976413,3.754667,4.7261543,5.0510774,4.6900516,3.9318976,3.6168208,3.2820516,3.3378465,3.9844105,5.1922054,7.778462,7.834257,6.9809237,6.232616,5.9930263,8.008205,8.385642,7.8736415,6.957949,5.85518,6.7938466,10.870154,12.865642,10.768411,5.7632823,6.2884107,10.177642,14.155488,16.003283,14.572309,12.291283,12.393026,11.044104,7.755488,5.3858466,8.500513,12.176412,13.10195,11.113027,9.196308,8.5202055,7.2205133,5.4482055,3.7316926,2.9440002,3.2951798,3.498667,4.092718,5.034667,5.7107697,4.827898,4.562052,4.962462,5.7501545,6.308103,6.193231,6.803693,7.315693,6.9645133,5.0642056,4.0434875,3.6135387,3.5282054,3.6562054,3.9581542,3.8859491,3.6758976,3.4527183,3.3312824,3.4198978,3.1081028,2.6945643,2.284308,1.9429746,1.7132308,1.7493335,1.9626669,2.0873847,2.0808206,2.1464617,2.0512822,1.9626669,1.6049232,1.0568206,0.73517954,0.74830776,0.3117949,0.14112821,0.318359,0.318359,0.10502565,0.18051283,0.2297436,0.17394873,0.18379489,0.06564103,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.016410258,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.04594872,0.11158975,0.17723078,0.53825647,1.020718,1.1651284,0.85005134,0.28225642,0.15425642,0.098461546,0.07548718,0.06564103,0.07876924,0.15097436,0.15425642,0.15097436,0.16738462,0.20020515,0.24943592,0.27897438,0.29538465,0.30194873,0.31507695,0.3117949,0.33476925,0.3708718,0.40697438,0.39712822,0.39056414,0.38400003,0.3511795,0.29538465,0.24943592,0.3052308,0.77128214,1.2307693,2.1858463,5.0871797,8.595693,14.316309,18.927591,19.482258,13.420309,9.209436,6.4590774,4.95918,4.3749747,4.2436924,3.9220517,2.7503593,1.529436,0.761436,0.65312827,0.35446155,0.30851284,0.3052308,0.21333335,0.013128206,0.0032820515,0.0,0.0032820515,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.0032820515,0.055794876,0.28882053,0.63343596,0.96492314,1.083077,1.3357949,1.782154,2.5698464,3.7743592,5.3891287,6.2785645,5.5007186,4.394667,3.7152824,3.6529233,3.4691284,3.9023592,4.640821,5.428513,6.042257,6.564103,7.0957956,7.4174366,7.5946674,7.9983597,7.6701546,6.957949,6.0816417,5.3169236,5.0084105,4.7261543,4.772103,4.9394875,4.896821,4.1550775,3.3378465,3.117949,3.2032824,3.3476925,3.3542566,3.062154,2.6551797,1.9823592,1.1684103,0.6432821,0.6301539,0.67610264,0.7450257,0.8172308,0.88943595,1.1093334,1.2373334,1.3029745,1.4145643,1.7558975,2.300718,3.0884104,3.8006158,4.529231,5.796103,7.9819493,9.984001,11.904001,13.541744,14.391796,15.333745,16.54154,18.615797,22.022566,27.096617,35.19344,43.54626,51.492107,58.15139,62.421337,64.05252,65.17498,65.8839,66.41888,67.16062,66.18913,63.94421,61.08226,58.39754,56.815594,55.440414,53.609028,52.08616,51.695595,53.30708,3.190154,3.0916924,1.3193847,0.19692309,0.20676924,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.0032820515,0.0,0.0,0.009846155,0.04594872,0.19364104,0.34789747,0.6301539,0.97805136,1.1749744,0.5021539,0.16082053,0.026256412,0.032820515,0.16738462,0.28882053,0.26584616,0.18051283,0.118153855,0.16738462,0.2297436,0.22646156,0.128,0.0,0.0,0.06235898,0.16738462,0.2297436,0.30194873,0.5940513,1.595077,1.9364104,1.7657437,1.3161026,0.8992821,1.0699488,1.1126155,0.8467693,0.37415388,0.108307704,0.08205129,0.08533334,0.07876924,0.052512825,0.016410258,0.0032820515,0.0,0.006564103,0.04266667,0.15097436,0.055794876,0.013128206,0.049230773,0.10502565,0.029538464,0.07876924,0.2100513,0.18051283,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06564103,0.19364104,0.37743592,0.6104616,0.12143591,0.009846155,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.036102567,0.06564103,0.08533334,0.12143591,0.15753847,0.15097436,0.118153855,0.08205129,0.04594872,0.04594872,0.01969231,0.0,0.0,0.0,0.0,0.06564103,0.07548718,0.059076928,0.16738462,0.31507695,0.23302566,0.09189744,0.013128206,0.06235898,0.072205134,0.12143591,0.14112821,0.13128206,0.16738462,0.04594872,0.016410258,0.016410258,0.013128206,0.0,0.013128206,0.006564103,0.0,0.0,0.0,0.0,0.009846155,0.009846155,0.013128206,0.06235898,0.013128206,0.026256412,0.026256412,0.0,0.0,0.0,0.009846155,0.02297436,0.055794876,0.15097436,0.14112821,0.072205134,0.029538464,0.036102567,0.06235898,0.20676924,0.1148718,0.029538464,0.055794876,0.15097436,0.24943592,0.18379489,0.14112821,0.14769232,0.06235898,0.15753847,0.37415388,0.60061544,0.8402052,1.204513,0.9747693,0.761436,0.5481026,0.4266667,0.6104616,0.84348726,1.2406155,1.5688206,1.5819489,1.0075898,0.94523084,0.9944616,1.591795,2.4057438,2.3204105,1.9298463,1.6016412,2.0841026,4.007385,7.890052,7.8408213,7.059693,5.0871797,2.8553848,2.6847181,5.2381544,8.392206,9.813334,8.94359,7.003898,8.274052,10.148104,10.098872,7.79159,5.080616,5.6418467,10.771693,13.545027,12.547283,11.88759,8.480822,8.664616,10.902975,13.026463,12.22236,11.588924,11.300103,9.524513,6.422975,4.164923,3.9712822,4.1878977,3.8334363,3.1540515,3.6168208,4.1058464,3.7316926,3.5249233,3.8432825,4.378257,3.879385,3.9187696,3.7054362,3.242667,3.3411283,3.3542566,3.767795,3.8071797,3.4034874,3.2196925,3.4034874,3.879385,4.3618464,4.568616,4.2272825,3.4198978,2.6715899,2.0906668,1.7985642,1.9068719,1.8084104,1.4276924,1.148718,1.0896411,1.1126155,1.4441026,1.7460514,2.044718,2.231795,2.0611284,1.6935385,1.1913847,0.76800007,0.49230772,0.25928208,0.17394873,0.12471796,0.06564103,0.0,0.0,0.20676924,0.10502565,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.026256412,0.016410258,0.016410258,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.036102567,0.10502565,0.190359,0.27569234,0.22646156,0.26912823,0.7515898,1.3226668,0.9321026,0.42994875,0.18707694,0.08861539,0.06564103,0.09189744,0.36102566,0.3446154,0.27241027,0.24943592,0.27569234,0.3117949,0.34789747,0.37743592,0.4004103,0.4135385,0.44964105,0.45620516,0.45620516,0.45620516,0.45620516,0.46933338,0.45620516,0.39384618,0.38400003,0.64000005,0.8598975,1.2832822,2.0808206,4.086154,8.772923,14.25395,17.473642,21.07077,21.48759,8.986258,3.8104618,3.8006158,5.0149746,5.3202057,4.378257,3.3050258,2.1202054,1.1191796,0.54482055,0.58092314,0.36102566,0.26912823,0.21333335,0.13456412,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.03938462,0.036102567,0.108307704,0.28882053,0.5349744,0.86317956,1.7690258,2.930872,3.8137438,3.692308,3.4494362,3.4067695,2.9472823,2.0775387,1.4178462,0.8336411,0.7417436,1.0272821,1.5392822,2.0742567,2.2449234,2.537026,2.8160002,2.993231,3.006359,2.7241027,2.7273848,2.3729234,1.6377437,1.1126155,1.1749744,0.9517949,0.7253334,0.64000005,0.702359,0.65312827,0.64000005,0.8730257,1.3522053,1.8773335,2.0250258,1.4998976,0.90912825,0.55794877,0.47261542,0.49887183,0.5316923,0.56123084,0.5940513,0.65641034,0.72861546,0.8566154,0.99774367,1.1323078,1.2668719,1.6935385,2.1398976,2.858667,3.9286156,5.2348723,6.491898,7.456821,8.464411,9.547488,10.436924,11.474052,12.320822,13.61395,15.635694,18.297438,21.910976,26.292515,32.141132,39.240208,46.480415,53.267696,59.231186,63.898262,67.06216,68.77211,67.87939,66.17272,64.70236,63.491287,61.538467,58.1317,55.696415,53.999596,53.41867,54.931698,1.1126155,0.8402052,0.34789747,0.06564103,0.052512825,0.0,0.0,0.0,0.0032820515,0.009846155,0.0032820515,0.07876924,0.03938462,0.0,0.0032820515,0.009846155,0.03938462,0.068923086,0.12471796,0.19692309,0.23630771,0.14112821,0.07548718,0.032820515,0.01969231,0.04594872,0.068923086,0.07876924,0.07876924,0.068923086,0.068923086,0.052512825,0.059076928,0.16082053,0.28225642,0.19692309,1.0469744,0.9485129,0.571077,0.5152821,1.3161026,1.9856411,1.3259488,0.60389745,0.3511795,0.37415388,0.3708718,0.39056414,0.47917953,0.508718,0.18051283,0.07876924,0.098461546,0.17394873,0.21661541,0.101743594,0.049230773,0.029538464,0.016410258,0.009846155,0.029538464,0.009846155,0.02297436,0.04266667,0.04594872,0.029538464,0.08861539,0.17066668,0.17394873,0.108307704,0.098461546,0.01969231,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07876924,0.10502565,0.07548718,0.12143591,0.14112821,0.24943592,0.19364104,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.013128206,0.016410258,0.02297436,0.06235898,0.0951795,0.1148718,0.108307704,0.068923086,0.059076928,0.03938462,0.01969231,0.009846155,0.0,0.0,0.013128206,0.04594872,0.068923086,0.032820515,0.072205134,0.06564103,0.032820515,0.0032820515,0.013128206,0.013128206,0.02297436,0.029538464,0.029538464,0.04594872,0.013128206,0.07548718,0.101743594,0.052512825,0.0,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0032820515,0.013128206,0.0032820515,0.006564103,0.006564103,0.0,0.0,0.009846155,0.049230773,0.14441027,0.23958977,0.190359,0.08861539,0.04266667,0.026256412,0.02297436,0.049230773,0.15753847,0.26584616,0.22646156,0.108307704,0.22646156,0.26584616,0.23302566,0.16082053,0.08205129,0.02297436,0.032820515,0.07548718,0.12471796,0.17723078,0.23958977,0.19364104,0.15097436,0.13456412,0.17394873,0.318359,0.3249231,0.4004103,0.47589746,0.50543594,0.45620516,0.39712822,0.380718,0.43651286,0.58420515,0.83035904,1.3292309,2.1333334,2.5009232,3.1540515,6.2523084,4.5817437,3.8662567,3.4527183,2.806154,1.4998976,2.2547693,4.2240005,7.2205133,9.954462,10.006975,8.598975,7.1844106,5.8978467,4.516103,2.4320002,3.5413337,7.578257,10.758565,11.913847,12.484924,9.458873,9.590155,11.053949,11.71036,9.097847,7.0465646,5.924103,5.07077,4.0992823,2.8947694,2.740513,2.674872,2.5928206,2.8455386,4.2272825,3.7382567,2.930872,2.4320002,2.3433847,2.2547693,2.1267693,2.103795,2.097231,2.1103592,2.2678976,2.7864618,3.0720003,2.9440002,2.556718,2.4024618,2.7602053,2.861949,2.740513,2.3794873,1.723077,1.3193847,1.4375386,1.4473847,1.3193847,1.6147693,1.3883078,0.9911796,0.75487185,0.8369231,1.211077,1.7263591,1.9593848,1.9298463,1.6180514,0.9485129,0.61374366,0.41025645,0.26256412,0.14112821,0.06564103,0.036102567,0.055794876,0.09189744,0.108307704,0.06235898,0.18051283,0.08533334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.032820515,0.049230773,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.016410258,0.0032820515,0.013128206,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.026256412,0.06564103,0.128,0.21333335,0.21333335,0.4135385,0.73517954,0.95835906,0.7220513,0.8467693,0.90584624,0.80738467,0.5349744,0.14112821,0.5349744,0.8369231,0.6826667,0.256,0.2986667,0.31507695,0.34789747,0.38400003,0.4201026,0.4594872,0.46933338,0.46933338,0.48574364,0.508718,0.51856416,0.512,0.49230772,0.6465641,1.0929232,1.8871796,2.172718,2.612513,3.5971284,5.32677,7.7981544,13.797745,18.822565,20.342155,16.505438,6.157129,3.5971284,4.6276927,5.6352825,5.169231,3.9154875,3.308308,2.0742567,0.9911796,0.41025645,0.24943592,0.15753847,0.10502565,0.06564103,0.026256412,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.006564103,0.055794876,0.16082053,0.27897438,0.55794877,1.2471796,2.0151796,2.5796926,2.6912823,2.6912823,2.5107694,2.1530259,1.6508719,1.0896411,0.56123084,0.4266667,0.3708718,0.318359,0.4266667,0.46276927,0.5284103,0.5874872,0.6268718,0.6498462,0.9944616,1.4966155,1.719795,1.4867693,0.892718,0.446359,0.28225642,0.2297436,0.21661541,0.23958977,0.23958977,0.25928208,0.33476925,0.4594872,0.58420515,0.6498462,0.571077,0.47261542,0.42338464,0.42338464,0.4594872,0.47917953,0.50543594,0.5415385,0.58420515,0.6268718,0.74830776,0.9616411,1.276718,1.6935385,2.0053334,2.353231,3.0162053,3.9745643,4.9296412,5.756718,6.340924,6.8233852,7.2861543,7.788308,8.41518,9.173334,9.95118,10.95877,12.740924,15.182771,18.343386,22.163694,26.59118,31.573336,35.862976,41.091286,47.44862,54.596928,61.666466,66.67487,69.04452,69.333336,67.83344,64.54154,60.626057,57.764107,56.077133,55.391182,55.2238,1.4572309,2.6387694,1.6672822,0.72861546,0.48902568,0.118153855,0.17066668,0.24287182,0.23958977,0.15425642,0.09189744,0.15097436,0.27569234,0.2100513,0.0032820515,0.01969231,0.0032820515,0.006564103,0.026256412,0.07876924,0.17394873,0.38400003,0.73517954,0.574359,0.029538464,0.006564103,0.17394873,0.77456415,1.3226668,1.6278975,1.785436,1.4998976,1.2996924,0.81394875,0.20348719,0.15097436,0.58092314,0.5284103,0.30851284,0.24287182,0.63343596,1.0305642,0.88287187,0.67938465,0.5152821,0.108307704,0.07876924,0.08533334,0.17394873,0.30851284,0.36430773,0.75487185,0.56451285,0.3117949,0.26584616,0.4594872,0.44964105,0.23630771,0.13456412,0.15425642,0.0,0.0,0.009846155,0.016410258,0.013128206,0.013128206,0.036102567,0.068923086,0.07876924,0.06235898,0.059076928,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.10502565,0.10502565,0.0,0.0,0.059076928,0.3511795,0.34133336,0.04266667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.032820515,0.052512825,0.06564103,0.06564103,0.055794876,0.032820515,0.02297436,0.01969231,0.0,0.0,0.0,0.013128206,0.029538464,0.0,0.013128206,0.036102567,0.055794876,0.059076928,0.036102567,0.04266667,0.02297436,0.009846155,0.009846155,0.006564103,0.009846155,0.03938462,0.049230773,0.036102567,0.055794876,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016410258,0.016410258,0.0,0.0,0.0032820515,0.02297436,0.072205134,0.13128206,0.17066668,0.072205134,0.026256412,0.009846155,0.009846155,0.01969231,0.06564103,0.13784617,0.14769232,0.098461546,0.098461546,0.12143591,0.10502565,0.06564103,0.026256412,0.006564103,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0,0.009846155,0.059076928,0.14769232,0.24287182,0.14441027,0.16082053,0.21333335,0.256,0.28225642,0.18707694,0.16410258,0.11158975,0.06564103,0.2100513,0.7122052,1.1716924,1.2077949,1.270154,2.6322052,2.612513,2.156308,1.9364104,1.8445129,1.0043077,1.2373334,2.3171284,4.263385,6.088206,5.796103,5.024821,4.076308,3.1376412,2.3958976,2.034872,4.020513,6.370462,8.713847,10.364718,10.33518,7.8473854,6.5969234,6.4722056,6.485334,4.7917953,3.242667,2.9046156,2.8521028,2.605949,2.1202054,2.1202054,2.172718,2.097231,2.044718,2.5206156,2.1267693,1.6180514,1.3718976,1.4112822,1.4211283,1.6475899,1.6180514,1.7099489,1.8576412,1.5589745,2.097231,2.487795,2.5173335,2.2121027,1.8313848,1.8149745,1.7165129,1.5392822,1.3653334,1.3259488,0.7515898,0.6629744,0.6629744,0.6301539,0.7089231,0.6432821,0.7056411,0.9517949,1.3095386,1.5753847,1.5130258,1.3751796,1.1355898,0.7975385,0.37743592,0.20348719,0.13456412,0.101743594,0.07548718,0.06235898,0.013128206,0.013128206,0.03938462,0.055794876,0.029538464,0.068923086,0.032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.0032820515,0.0032820515,0.016410258,0.02297436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.009846155,0.029538464,0.02297436,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.068923086,0.16738462,0.20676924,0.24287182,0.4660513,0.7450257,0.9353847,0.90912825,1.5360001,1.6935385,1.785436,2.231795,3.4658465,4.391385,4.0533338,2.6486156,0.9747693,0.4135385,0.30851284,0.3117949,0.34789747,0.39056414,0.446359,0.45292312,0.47261542,0.512,0.56451285,0.6071795,0.60389745,0.7253334,1.1651284,1.8576412,2.5009232,3.6824617,4.5554876,5.4843082,6.514872,7.3616414,9.504821,11.608616,11.923694,9.714872,5.2545643,3.8695388,4.8016415,5.586052,5.1954875,4.0467696,4.6145644,3.876103,2.3663592,0.8172308,0.14112821,0.101743594,0.08533334,0.118153855,0.14769232,0.036102567,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.30851284,0.67282057,0.8960001,0.8369231,0.88615394,1.0568206,1.3062565,1.5753847,1.8182565,1.8445129,1.7362052,1.5261539,1.2012309,0.7220513,0.512,0.42338464,0.24943592,0.02297436,0.016410258,0.016410258,0.01969231,0.026256412,0.032820515,0.04266667,0.24287182,0.5546667,0.7384616,0.67282057,0.36430773,0.14769232,0.09189744,0.09189744,0.098461546,0.10502565,0.12471796,0.15097436,0.27241027,0.47589746,0.65312827,0.52512825,0.40369233,0.35446155,0.37743592,0.40369233,0.42338464,0.446359,0.4660513,0.48902568,0.51856416,0.5546667,0.62030774,0.7318975,0.90256417,1.1520001,1.4834872,1.9003079,2.422154,3.0129232,3.5807183,4.161641,4.5390773,5.169231,6.160411,7.282872,7.177847,7.1187696,7.2664623,7.8112826,8.973129,10.492719,12.616206,15.199181,18.169437,21.540104,24.4119,28.054977,32.856617,38.688824,44.931286,51.64308,57.366978,61.587696,64.085335,64.93539,64.66626,64.53498,64.73518,65.903595,69.10359,1.2176411,2.605949,2.0086155,1.2471796,0.8730257,0.15425642,0.19364104,0.47917953,0.6104616,0.4660513,0.20676924,0.23958977,0.4135385,0.52512825,0.5481026,0.64000005,0.446359,0.40369233,0.6071795,0.97805136,1.2537436,1.0305642,1.2537436,1.020718,0.3117949,0.013128206,0.23302566,0.88615394,1.591795,2.0709746,2.1464617,1.6902566,1.4342566,0.8763078,0.190359,0.23958977,0.36758977,0.35774362,0.24287182,0.12143591,0.15097436,0.44964105,0.6629744,0.7122052,0.5284103,0.052512825,0.28882053,0.79425645,1.2274873,1.3915899,1.2373334,1.3686155,1.024,0.9156924,1.2931283,1.9331284,1.3587693,0.6071795,0.21661541,0.20348719,0.06235898,0.06235898,0.02297436,0.0,0.0,0.006564103,0.0,0.006564103,0.009846155,0.01969231,0.06564103,0.1148718,0.13784617,0.13128206,0.09189744,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.03938462,0.18379489,0.17394873,0.029538464,0.01969231,0.0032820515,0.25928208,0.27897438,0.04266667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.02297436,0.036102567,0.032820515,0.026256412,0.02297436,0.01969231,0.006564103,0.0,0.0032820515,0.0032820515,0.0,0.0,0.013128206,0.032820515,0.068923086,0.1148718,0.14769232,0.10502565,0.068923086,0.049230773,0.03938462,0.01969231,0.01969231,0.013128206,0.0032820515,0.009846155,0.055794876,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.032820515,0.026256412,0.009846155,0.04266667,0.009846155,0.0032820515,0.0032820515,0.02297436,0.108307704,0.052512825,0.026256412,0.013128206,0.006564103,0.006564103,0.009846155,0.013128206,0.03938462,0.055794876,0.0,0.013128206,0.006564103,0.0,0.0,0.0,0.0,0.03938462,0.10502565,0.14441027,0.08533334,0.026256412,0.016410258,0.049230773,0.108307704,0.14769232,0.0951795,0.14441027,0.18051283,0.17723078,0.17394873,0.101743594,0.098461546,0.068923086,0.036102567,0.11158975,0.47261542,0.48902568,0.30851284,0.18051283,0.47589746,1.5195899,1.719795,1.5589745,1.3095386,1.020718,1.3226668,1.785436,2.3204105,2.6157951,2.1202054,2.2088206,2.294154,2.0906668,1.8346668,2.281026,3.9876926,4.768821,5.7534366,6.820103,6.6002054,5.0051284,3.436308,2.5993848,2.3893335,1.9035898,1.2209232,1.3620514,1.5261539,1.4309745,1.3226668,1.3751796,1.6311796,1.6311796,1.332513,1.1060513,1.2964103,1.3128207,1.3653334,1.4966155,1.5688206,1.9331284,1.9528207,1.9626669,1.9200002,1.4080001,1.4112822,1.5327181,1.595077,1.4802053,1.148718,0.90912825,0.764718,0.67938465,0.6892308,0.9321026,0.44307697,0.25928208,0.2986667,0.42338464,0.4397949,0.508718,0.8402052,1.1815386,1.3620514,1.3062565,0.9616411,0.702359,0.47917953,0.27897438,0.14769232,0.08205129,0.055794876,0.049230773,0.055794876,0.055794876,0.009846155,0.0,0.0,0.0,0.0,0.0,0.009846155,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.006564103,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.02297436,0.029538464,0.03938462,0.04594872,0.036102567,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.052512825,0.14769232,0.20676924,0.31507695,0.7089231,0.9944616,1.0436924,0.9878975,1.5261539,1.7723079,2.0709746,3.0720003,5.7435904,7.312411,7.138462,5.3202057,2.7634873,1.1913847,0.6498462,0.4660513,0.4397949,0.4660513,0.53825647,0.6235898,1.0272821,1.1585642,0.95835906,0.9124103,1.1126155,1.3587693,1.9823592,2.8882053,3.5807183,4.706462,5.986462,6.75118,7.000616,7.4043083,7.6242056,7.506052,6.885744,5.933949,5.146257,4.46359,4.900103,5.3858466,5.3727183,4.841026,5.044513,4.378257,2.9407182,1.2668719,0.33476925,0.21989745,0.128,0.12471796,0.15425642,0.049230773,0.072205134,0.04594872,0.06235898,0.101743594,0.04266667,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.5481026,1.1454359,1.4539489,1.270154,1.142154,1.0896411,1.1323078,1.2471796,1.3554872,1.1881026,1.0994873,0.97805136,0.76800007,0.47917953,0.446359,0.38400003,0.2231795,0.032820515,0.016410258,0.016410258,0.016410258,0.01969231,0.02297436,0.02297436,0.02297436,0.08861539,0.16410258,0.19692309,0.12471796,0.08205129,0.07876924,0.08533334,0.09189744,0.098461546,0.118153855,0.16738462,0.34789747,0.6301539,0.8467693,0.6662565,0.47589746,0.3708718,0.36758977,0.39056414,0.40697438,0.4266667,0.44307697,0.45620516,0.47589746,0.5021539,0.5284103,0.5546667,0.5973334,0.6629744,0.90584624,1.2209232,1.5458462,1.8543591,2.156308,2.5009232,2.7175386,3.242667,4.2207184,5.5171285,5.579488,5.654975,5.664821,5.76,6.3540516,7.2336416,8.579283,10.31877,12.347078,14.5263605,16.42995,18.520617,21.215181,24.763079,29.203695,35.219696,41.04862,46.464005,51.406773,55.981953,59.62175,62.87098,67.18031,73.31775,81.3719,0.0,0.15753847,0.7975385,1.1323078,0.8402052,0.08205129,0.04594872,0.46933338,0.74830776,0.6465641,0.28882053,0.26256412,0.31507695,0.65312827,1.1684103,1.4506668,0.96492314,0.8172308,1.1716924,1.847795,2.2908719,1.3850257,1.1093334,1.0305642,0.78769237,0.13456412,0.28225642,0.47917953,0.9156924,1.2964103,0.827077,0.4397949,0.4955898,0.52512825,0.41682056,0.39384618,0.6826667,0.6662565,0.47917953,0.30851284,0.42338464,0.71548724,0.6859488,0.48246157,0.27569234,0.25271797,0.8041026,1.7920002,2.5665643,2.7109745,2.0644104,1.4178462,1.2570257,1.723077,2.6289232,3.4527183,2.15959,0.9321026,0.25928208,0.15425642,0.16082053,0.14441027,0.06235898,0.016410258,0.026256412,0.029538464,0.009846155,0.009846155,0.013128206,0.03938462,0.12143591,0.23630771,0.30194873,0.2986667,0.21333335,0.04266667,0.013128206,0.0032820515,0.0032820515,0.0032820515,0.0,0.009846155,0.006564103,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.02297436,0.098461546,0.23630771,0.21333335,0.055794876,0.036102567,0.006564103,0.06564103,0.09189744,0.07548718,0.108307704,0.06235898,0.01969231,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.01969231,0.01969231,0.013128206,0.013128206,0.0032820515,0.009846155,0.009846155,0.0032820515,0.0,0.009846155,0.013128206,0.04266667,0.11158975,0.21989745,0.12143591,0.098461546,0.09189744,0.07876924,0.04594872,0.032820515,0.02297436,0.013128206,0.006564103,0.009846155,0.006564103,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.036102567,0.03938462,0.026256412,0.029538464,0.101743594,0.02297436,0.009846155,0.006564103,0.006564103,0.03938462,0.036102567,0.036102567,0.026256412,0.013128206,0.013128206,0.0032820515,0.0,0.0032820515,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.08533334,0.2100513,0.28882053,0.18051283,0.059076928,0.026256412,0.02297436,0.02297436,0.006564103,0.07548718,0.13456412,0.10502565,0.029538464,0.04266667,0.04594872,0.049230773,0.036102567,0.06564103,0.26912823,0.5874872,0.5973334,0.446359,0.3314872,0.5152821,0.9321026,1.7460514,1.9462565,1.4966155,1.3193847,1.7001027,1.782154,1.6508719,1.4769232,1.522872,1.5983591,1.9298463,2.2350771,2.4746668,2.858667,3.249231,2.9078977,2.5928206,2.6683078,3.0949745,2.487795,1.8084104,1.3095386,1.0896411,1.1093334,0.86974365,0.7384616,0.69907695,0.71548724,0.7384616,0.7450257,1.0469744,1.1716924,1.0371283,0.9517949,1.5261539,1.785436,1.8642052,1.8642052,1.8642052,2.1398976,2.1956925,2.044718,1.7493335,1.404718,0.82379496,0.46933338,0.3708718,0.42338464,0.4004103,0.26912823,0.190359,0.14441027,0.118153855,0.08533334,0.049230773,0.16738462,0.43323082,0.74830776,0.9124103,0.955077,1.1126155,1.0436924,0.7318975,0.48574364,0.35774362,0.28882053,0.21661541,0.13456412,0.07548718,0.036102567,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.02297436,0.04266667,0.032820515,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0,0.0,0.02297436,0.07548718,0.13456412,0.128,0.08533334,0.04266667,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.055794876,0.18379489,0.3511795,0.90912825,1.2668719,1.2307693,0.9878975,1.0502565,1.3686155,1.7460514,2.7208207,5.5729237,7.3682055,8.083693,6.9842057,4.4767184,2.1202054,1.0765129,0.69907695,0.61374366,0.6235898,0.702359,0.892718,1.7591796,1.9987694,1.5163078,1.4112822,1.9987694,2.3433847,3.0096412,3.9909747,4.6966157,4.772103,6.0160003,6.5739493,6.3901544,7.1876926,8.720411,8.635077,7.207385,5.398975,4.857436,4.8836927,5.2578464,5.8092313,6.2096415,5.970052,4.44718,3.5347695,2.7634873,1.8806155,0.8533334,0.4594872,0.20020515,0.059076928,0.016410258,0.026256412,0.16410258,0.15425642,0.21333335,0.2986667,0.0951795,0.01969231,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.49887183,1.0404103,1.3259488,1.1290257,0.9878975,1.1323078,1.3620514,1.5130258,1.4605129,1.142154,0.90912825,0.7056411,0.51856416,0.37415388,0.29210258,0.21333335,0.12471796,0.04266667,0.02297436,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.02297436,0.10502565,0.21333335,0.20348719,0.08861539,0.07876924,0.08861539,0.0951795,0.10502565,0.118153855,0.190359,0.34789747,0.5415385,0.6465641,0.58420515,0.47917953,0.39056414,0.35446155,0.37415388,0.40369233,0.41682056,0.42994875,0.446359,0.45620516,0.46933338,0.49230772,0.5152821,0.53825647,0.574359,0.63343596,0.69907695,0.8369231,1.0305642,1.214359,1.3292309,1.4145643,1.4933335,1.7296412,2.4155898,3.2000003,4.1124105,4.4077954,4.1846156,4.397949,4.9920006,5.8256416,6.941539,8.267488,9.626257,10.765129,11.867898,13.298873,15.468308,18.848822,23.122053,26.77826,30.486977,34.806156,40.16903,45.650055,51.203285,58.72575,68.80493,80.70565,0.0,0.0,0.15425642,0.31507695,0.32820517,0.04594872,0.009846155,0.0,0.006564103,0.068923086,0.28882053,0.059076928,0.0,0.098461546,0.4004103,1.024,0.4135385,0.11158975,0.06564103,0.23958977,0.65641034,0.26584616,0.15753847,0.5546667,1.0371283,0.5481026,0.7581539,1.1191796,1.6705642,1.8149745,0.3511795,0.27897438,1.0469744,1.3226668,0.7844103,0.13784617,0.35774362,0.45620516,0.4397949,0.48574364,0.9616411,1.0469744,0.9321026,0.8205129,0.8041026,0.8402052,1.1454359,1.0108719,0.72861546,0.574359,0.79425645,0.6465641,1.3062565,1.782154,1.8510771,2.0611284,1.4605129,0.8172308,0.40369233,0.25928208,0.19692309,0.11158975,0.072205134,0.08533334,0.1148718,0.09189744,0.04266667,0.049230773,0.072205134,0.08533334,0.06235898,0.049230773,0.118153855,0.17394873,0.16410258,0.09189744,0.04266667,0.02297436,0.016410258,0.013128206,0.0,0.049230773,0.032820515,0.016410258,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.06235898,0.08533334,0.06564103,0.026256412,0.0,0.0,0.0,0.0,0.13456412,0.37415388,0.5349744,0.31507695,0.10502565,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.006564103,0.006564103,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.036102567,0.06235898,0.059076928,0.04594872,0.032820515,0.029538464,0.029538464,0.032820515,0.04594872,0.032820515,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08533334,0.04266667,0.02297436,0.06564103,0.07548718,0.026256412,0.006564103,0.0,0.0032820515,0.016410258,0.052512825,0.02297436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02297436,0.02297436,0.009846155,0.009846155,0.04594872,0.032820515,0.07548718,0.0951795,0.06564103,0.029538464,0.09189744,0.07876924,0.036102567,0.006564103,0.029538464,0.04266667,0.026256412,0.016410258,0.108307704,0.48902568,0.6104616,0.7417436,0.80738467,0.7975385,0.74830776,0.5415385,0.8369231,1.3062565,1.6475899,1.5885129,1.5885129,1.4867693,1.3653334,1.2898463,1.3259488,1.4145643,1.7099489,2.2580514,3.2000003,4.775385,4.532513,3.436308,2.3072822,1.7755898,2.28759,2.03159,1.3554872,0.90256417,0.8992821,1.1454359,0.9353847,0.81066674,0.9517949,1.2635899,1.3718976,1.4572309,1.4703591,1.3620514,1.2438976,1.404718,1.3423591,1.0699488,0.72861546,0.571077,0.9616411,1.1191796,1.014154,0.8960001,0.8041026,0.5481026,0.37743592,0.28882053,0.18051283,0.059076928,0.04594872,0.02297436,0.006564103,0.006564103,0.013128206,0.0,0.15753847,0.35446155,0.6662565,0.99774367,1.083077,0.9616411,0.6662565,0.29210258,0.032820515,0.16738462,0.118153855,0.098461546,0.06235898,0.016410258,0.016410258,0.016410258,0.016410258,0.009846155,0.0,0.0,0.0,0.0,0.0,0.009846155,0.04594872,0.108307704,0.10502565,0.055794876,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.013128206,0.0,0.0,0.036102567,0.1148718,0.21333335,0.27569234,0.36102566,0.20676924,0.055794876,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02297436,0.12143591,0.18379489,0.318359,0.892718,1.5983591,1.463795,1.5261539,1.7066668,1.9331284,2.5829747,4.4865646,5.3169236,5.717334,5.0674877,3.4527183,1.6311796,0.7056411,0.5546667,0.6235898,0.65312827,0.702359,0.8730257,1.3456411,1.5721027,1.5556924,1.8609232,2.802872,3.367385,4.0434875,4.562052,3.892513,3.6332312,3.9745643,4.279795,4.525949,5.293949,7.686565,7.5520005,5.7632823,3.7710772,3.6004105,4.309334,5.9602056,7.8703594,8.753231,6.7150774,4.673641,4.394667,4.273231,3.4166157,1.6475899,0.69579494,0.3117949,0.128,0.0032820515,0.016410258,0.16082053,0.30851284,0.4594872,0.47261542,0.04594872,0.009846155,0.0,0.0,0.0,0.0,0.0,0.009846155,0.009846155,0.0032820515,0.016410258,0.016410258,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08205129,0.31507695,0.5546667,0.45620516,0.43323082,0.88615394,1.3718976,1.7558975,2.1825643,2.2416413,1.7460514,1.1913847,0.75487185,0.28882053,0.118153855,0.07548718,0.068923086,0.059076928,0.04594872,0.02297436,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.02297436,0.036102567,0.04594872,0.04594872,0.059076928,0.068923086,0.08205129,0.09189744,0.09189744,0.1148718,0.13128206,0.16082053,0.20676924,0.24287182,0.26912823,0.30194873,0.3314872,0.3511795,0.3511795,0.38728207,0.40697438,0.42338464,0.446359,0.45620516,0.46933338,0.49230772,0.508718,0.52512825,0.5481026,0.5973334,0.65641034,0.7220513,0.8008206,0.88615394,0.9714873,1.0469744,1.1027694,1.148718,1.2209232,1.3686155,1.6246156,1.9298463,2.284308,2.7634873,3.5314875,4.07959,4.824616,5.8420515,6.8660517,7.5881033,8.490667,9.53436,10.692924,11.963078,14.342566,18.01518,21.69436,25.153643,29.206976,33.70995,39.525745,42.79467,46.342567,59.648006,0.0,0.0,0.029538464,0.06235898,0.06564103,0.009846155,0.0032820515,0.0,0.0,0.013128206,0.059076928,0.013128206,0.0,0.01969231,0.07876924,0.20348719,0.101743594,0.032820515,0.016410258,0.068923086,0.18051283,0.072205134,0.15425642,0.56123084,0.9878975,0.69579494,0.74830776,0.9747693,1.024,0.7253334,0.118153855,0.34789747,0.7975385,1.2077949,1.1552821,0.03938462,0.18051283,0.22646156,0.17394873,0.14441027,0.38728207,0.73517954,1.0732309,1.1979488,1.2406155,1.6705642,1.1158975,0.764718,0.8992821,1.2603078,1.0502565,0.8041026,0.8172308,1.2996924,1.9167181,1.8051283,1.9167181,1.7394873,1.6836925,1.5753847,0.6268718,0.23630771,0.23302566,0.5677949,0.9156924,0.67610264,0.256,0.128,0.09189744,0.06235898,0.036102567,0.013128206,0.052512825,0.07548718,0.055794876,0.029538464,0.068923086,0.049230773,0.016410258,0.0032820515,0.013128206,0.013128206,0.006564103,0.0032820515,0.0032820515,0.013128206,0.0032820515,0.013128206,0.01969231,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.016410258,0.013128206,0.006564103,0.006564103,0.036102567,0.006564103,0.0,0.055794876,0.15425642,0.20348719,0.08205129,0.01969231,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03938462,0.19692309,0.03938462,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.006564103,0.0,0.0,0.0032820515,0.009846155,0.013128206,0.013128206,0.0,0.009846155,0.0032820515,0.0032820515,0.009846155,0.0,0.0,0.006564103,0.013128206,0.013128206,0.009846155,0.006564103,0.006564103,0.006564103,0.006564103,0.009846155,0.006564103,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.059076928,0.036102567,0.013128206,0.016410258,0.026256412,0.006564103,0.0,0.0,0.006564103,0.026256412,0.055794876,0.052512825,0.032820515,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.02297436,0.08205129,0.26584616,0.20348719,0.118153855,0.068923086,0.055794876,0.01969231,0.08861539,0.1148718,0.24943592,0.4135385,0.3117949,0.15753847,0.09189744,0.06564103,0.0951795,0.26912823,0.4004103,0.5349744,0.702359,0.827077,0.7122052,0.45620516,0.4660513,0.5316923,0.55794877,0.5874872,0.60389745,0.58420515,0.6301539,0.8763078,1.4506668,2.3072822,2.9046156,3.629949,4.4767184,5.044513,4.322462,3.2098465,2.1202054,1.394872,1.3128207,1.1913847,0.8730257,0.6498462,0.6892308,1.0108719,1.339077,1.657436,1.8838975,1.9200002,1.6311796,0.9353847,0.58092314,0.4955898,0.6071795,0.8533334,0.6859488,0.42338464,0.25928208,0.23630771,0.26584616,0.30851284,0.25271797,0.20020515,0.17394873,0.12143591,0.118153855,0.14441027,0.13456412,0.09189744,0.068923086,0.14441027,0.13784617,0.07548718,0.036102567,0.17066668,0.43651286,0.761436,0.9714873,0.92553854,0.5218462,0.30194873,0.19364104,0.118153855,0.072205134,0.118153855,0.049230773,0.02297436,0.013128206,0.0032820515,0.0032820515,0.0032820515,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.013128206,0.068923086,0.09189744,0.101743594,0.08533334,0.049230773,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.013128206,0.013128206,0.0,0.0,0.013128206,0.08533334,0.190359,0.26256412,0.37743592,0.58420515,0.6268718,0.44964105,0.19692309,0.03938462,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.02297436,0.07548718,0.19364104,0.7089231,1.2635899,0.8041026,1.4998976,3.0720003,3.9909747,4.0041027,4.1189747,3.9351797,3.6693337,3.1507695,2.4188719,1.7427694,1.3817437,1.2209232,0.98461545,0.65969235,0.4955898,1.0371283,1.6311796,2.2121027,2.6584618,2.789744,3.6693337,4.3290257,4.8705645,5.0838976,4.453744,3.7185643,3.4822567,3.5577438,3.7382567,3.7940516,4.1747694,4.5554876,4.3684106,3.9253337,4.417641,5.5072823,5.8978467,6.445949,6.954667,6.1768208,4.138667,3.2853336,2.8849232,2.3860514,1.4145643,0.88287187,0.44964105,0.26256412,0.38400003,0.7975385,0.48246157,0.508718,0.5349744,0.508718,0.65641034,1.2931283,0.6235898,0.04266667,0.0,0.0,0.0,0.009846155,0.013128206,0.009846155,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.006564103,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016410258,0.08861539,0.22646156,0.4201026,0.36758977,0.4594872,0.7975385,1.1979488,1.204513,1.529436,1.4342566,1.1684103,0.86974365,0.58420515,0.17723078,0.068923086,0.059076928,0.04594872,0.032820515,0.01969231,0.006564103,0.0032820515,0.0032820515,0.0032820515,0.013128206,0.016410258,0.013128206,0.013128206,0.02297436,0.032820515,0.052512825,0.068923086,0.07876924,0.07876924,0.1148718,0.13784617,0.17394873,0.21661541,0.24287182,0.28882053,0.3117949,0.3314872,0.35774362,0.38728207,0.39384618,0.39712822,0.41682056,0.44307697,0.446359,0.4660513,0.49230772,0.508718,0.5218462,0.53825647,0.57764107,0.6170257,0.6695385,0.7318975,0.78769237,0.8533334,0.90912825,0.9616411,1.0075898,1.0633847,1.1881026,1.3587693,1.5425643,1.7427694,2.0053334,2.5304618,3.0752823,3.748103,4.588308,5.586052,6.304821,7.604513,8.569437,8.89436,8.874667,10.738873,13.092104,15.248411,17.355488,20.391386,24.477541,27.72349,30.893951,36.10585,46.85457,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.0032820515,0.0032820515,0.009846155,0.02297436,0.009846155,0.06235898,0.2297436,0.4004103,0.3117949,0.30851284,0.39056414,0.36102566,0.24287182,0.26256412,0.44307697,0.48574364,0.5481026,0.5218462,0.006564103,0.08533334,0.10502565,0.06564103,0.0951795,0.446359,0.8467693,1.0075898,1.020718,1.0502565,1.3554872,1.4736412,1.2800001,1.3423591,1.595077,1.3522053,1.6311796,1.3456411,1.3226668,1.7657437,2.2416413,2.156308,1.913436,1.8379488,1.7132308,0.7975385,0.6826667,0.60389745,0.9189744,1.3850257,1.1815386,0.6695385,0.2986667,0.098461546,0.029538464,0.02297436,0.013128206,0.02297436,0.055794876,0.07548718,0.04266667,0.08205129,0.10502565,0.08533334,0.03938462,0.006564103,0.0,0.0,0.0,0.0,0.006564103,0.016410258,0.01969231,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.01969231,0.0032820515,0.18051283,0.24615386,0.14112821,0.049230773,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01969231,0.098461546,0.01969231,0.0,0.0032820515,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0,0.009846155,0.013128206,0.0032820515,0.0,0.0032820515,0.0032820515,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.01969231,0.013128206,0.0032820515,0.0032820515,0.016410258,0.032820515,0.029538464,0.029538464,0.032820515,0.013128206,0.072205134,0.08205129,0.049230773,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.036102567,0.101743594,0.18379489,0.16082053,0.16082053,0.19692309,0.24943592,0.23630771,0.22646156,0.28882053,0.35446155,0.35446155,0.19692309,0.11158975,0.09189744,0.08533334,0.09189744,0.15097436,0.22646156,0.27897438,0.3446154,0.40369233,0.36430773,0.26912823,0.24615386,0.2297436,0.21333335,0.21661541,0.23302566,0.2986667,0.42338464,0.7187693,1.3883078,2.300718,2.665026,2.993231,3.3641028,3.4166157,2.7208207,2.0545642,1.6213335,1.4933335,1.5983591,1.585231,1.401436,1.1979488,1.142154,1.3981539,1.5327181,1.2406155,1.0272821,1.0108719,0.8960001,0.57764107,0.5415385,0.56123084,0.5481026,0.5513847,1.0666667,0.7778462,0.5021539,0.44964105,0.2297436,0.0951795,0.036102567,0.01969231,0.016410258,0.016410258,0.12471796,0.25928208,0.28882053,0.19692309,0.08533334,0.13128206,0.14769232,0.15425642,0.18707694,0.31507695,0.7318975,0.76800007,0.65641034,0.5218462,0.4004103,0.20020515,0.08861539,0.059076928,0.068923086,0.04266667,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.029538464,0.036102567,0.03938462,0.03938462,0.02297436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.013128206,0.0032820515,0.0,0.0,0.0032820515,0.029538464,0.07548718,0.11158975,0.16082053,0.27897438,0.32820517,0.27569234,0.20676924,0.23958977,0.38400003,0.36758977,0.16082053,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01969231,0.07548718,0.3052308,0.5907693,0.5677949,1.0108719,2.5829747,3.7251284,4.1682053,4.9427695,2.4451284,2.0578463,2.3269746,2.5895386,2.9604106,2.0808206,1.5491283,1.3423591,1.1618463,0.40697438,1.1946667,1.7493335,2.2547693,2.8192823,3.4691284,3.8104618,4.7950773,6.23918,7.0498466,5.2348723,3.7415388,3.2656412,3.2098465,3.5413337,4.772103,5.5532312,5.2709746,5.044513,5.287385,5.7042055,7.781744,7.453539,6.4000006,5.6287184,5.504,4.7294364,3.8400004,3.3378465,2.9243078,1.467077,0.7318975,0.36430773,0.2297436,0.46933338,1.4867693,1.6508719,1.7165129,1.5721027,1.463795,1.9889232,2.5238976,1.5458462,0.5152821,0.06564103,0.0,0.0,0.009846155,0.016410258,0.013128206,0.009846155,0.009846155,0.013128206,0.01969231,0.01969231,0.01969231,0.01969231,0.016410258,0.013128206,0.009846155,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.07548718,0.256,0.4135385,0.54482055,0.8763078,1.3489232,1.6114873,1.6935385,1.339077,0.8992821,0.56123084,0.30851284,0.101743594,0.04594872,0.03938462,0.032820515,0.02297436,0.016410258,0.013128206,0.006564103,0.0,0.0,0.0032820515,0.013128206,0.009846155,0.0032820515,0.016410258,0.01969231,0.032820515,0.049230773,0.06235898,0.07548718,0.11158975,0.14112821,0.17066668,0.20676924,0.25271797,0.29538465,0.3249231,0.3511795,0.37743592,0.40697438,0.4135385,0.4135385,0.4266667,0.44307697,0.45292312,0.46276927,0.47261542,0.48246157,0.49230772,0.49887183,0.52512825,0.5546667,0.5940513,0.64000005,0.67938465,0.7122052,0.7581539,0.8041026,0.8533334,0.892718,0.97805136,1.1093334,1.2668719,1.4441026,1.6607181,2.0053334,2.3696413,2.8488207,3.4658465,4.1747694,4.886975,6.0160003,6.87918,7.2894363,7.525744,8.835282,10.226872,11.247591,12.232206,14.296617,19.170464,22.28513,25.77395,32.15426,44.35036,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.01969231,0.009846155,0.013128206,0.01969231,0.06235898,0.23958977,0.29538465,0.190359,0.07876924,0.029538464,0.006564103,0.036102567,0.055794876,0.06235898,0.12143591,0.38400003,0.60061544,0.571077,0.512,0.5349744,0.65312827,1.2832822,1.270154,1.1979488,1.3357949,1.6377437,2.8192823,2.6683078,2.1891284,2.0118976,2.409026,2.284308,2.041436,1.7657437,1.4506668,0.99774367,1.3357949,1.3095386,1.3456411,1.5031796,1.467077,1.1782565,0.7581539,0.40697438,0.21661541,0.16082053,0.18051283,0.108307704,0.06564103,0.072205134,0.049230773,0.06235898,0.16082053,0.23958977,0.23302566,0.098461546,0.052512825,0.036102567,0.036102567,0.03938462,0.02297436,0.01969231,0.013128206,0.032820515,0.052512825,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.18051283,0.23302566,0.12471796,0.10502565,0.13456412,0.27569234,0.21989745,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.029538464,0.029538464,0.032820515,0.049230773,0.06564103,0.128,0.101743594,0.04266667,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.029538464,0.07548718,0.09189744,0.1148718,0.2231795,0.36430773,0.49887183,0.571077,0.5152821,0.47589746,0.39384618,0.26584616,0.15097436,0.118153855,0.12143591,0.15097436,0.190359,0.19364104,0.14441027,0.15753847,0.16738462,0.15425642,0.14441027,0.18379489,0.22646156,0.24943592,0.23630771,0.18707694,0.18707694,0.23958977,0.33476925,0.5546667,1.083077,1.847795,2.1891284,2.2646155,2.1825643,2.0086155,1.4441026,1.1158975,1.0666667,1.3193847,1.8740515,1.6180514,1.5622566,1.4900514,1.4408206,1.7165129,1.9823592,1.7099489,1.1093334,0.56451285,0.65312827,1.0568206,1.2340513,1.1552821,0.88287187,0.56451285,1.0699488,0.9321026,0.6859488,0.51856416,0.23958977,0.14112821,0.06235898,0.06235898,0.12471796,0.16738462,0.33476925,0.36102566,0.2855385,0.17723078,0.128,0.16082053,0.24287182,0.2855385,0.30194873,0.40697438,0.69251287,0.5152821,0.27241027,0.18707694,0.30851284,0.2100513,0.098461546,0.04266667,0.036102567,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.006564103,0.006564103,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.0,0.0,0.0,0.0,0.0,0.009846155,0.04594872,0.049230773,0.013128206,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.009846155,0.009846155,0.01969231,0.052512825,0.12143591,0.29538465,0.4955898,0.5546667,0.39056414,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02297436,0.068923086,0.17723078,0.4135385,0.892718,2.1891284,3.131077,3.6135387,4.585026,1.8609232,1.7296412,2.5862565,3.387077,3.6562054,2.7175386,2.0512822,1.8871796,1.8576412,0.98461545,1.8116925,2.1234872,2.3105643,2.6551797,3.3542566,3.757949,4.6834874,6.1407185,7.181129,5.904411,4.886975,4.2830772,3.7874875,4.0467696,6.6527185,7.6603084,7.8145647,7.1680007,6.4032826,6.813539,7.755488,8.27077,7.568411,5.904411,4.604718,5.9667697,5.9569235,5.208616,3.948308,1.9856411,0.8402052,0.38400003,0.37415388,0.69251287,1.332513,1.591795,1.8510771,2.4188719,2.917744,2.2646155,2.3204105,1.5031796,0.79425645,0.508718,0.256,0.08533334,0.02297436,0.009846155,0.009846155,0.016410258,0.016410258,0.029538464,0.036102567,0.036102567,0.036102567,0.04266667,0.03938462,0.03938462,0.03938462,0.03938462,0.016410258,0.013128206,0.009846155,0.006564103,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01969231,0.09189744,0.27569234,0.47261542,0.8205129,1.3128207,1.7952822,1.8576412,1.3686155,0.77128214,0.318359,0.052512825,0.029538464,0.029538464,0.029538464,0.026256412,0.009846155,0.013128206,0.016410258,0.009846155,0.0,0.0,0.0,0.006564103,0.006564103,0.006564103,0.009846155,0.013128206,0.02297436,0.03938462,0.055794876,0.07548718,0.108307704,0.13128206,0.15425642,0.190359,0.24615386,0.28225642,0.32164106,0.35446155,0.380718,0.40697438,0.4135385,0.42338464,0.42994875,0.4397949,0.446359,0.446359,0.44964105,0.45292312,0.45620516,0.4660513,0.48246157,0.49230772,0.512,0.54482055,0.58420515,0.60061544,0.63343596,0.67938465,0.72861546,0.761436,0.8172308,0.92553854,1.079795,1.2570257,1.4539489,1.6771283,1.8970258,2.1989746,2.5928206,3.0096412,3.5905645,4.3749747,5.1889234,5.937231,6.629744,7.7456417,8.795898,9.403078,9.898667,11.32636,15.281232,18.491077,24.329847,37.215183,62.62811,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.016410258,0.01969231,0.02297436,0.052512825,0.1148718,0.17394873,0.13784617,0.052512825,0.029538464,0.072205134,0.2297436,0.5940513,0.6662565,0.5940513,0.53825647,0.79425645,1.8018463,3.43959,3.817026,3.495385,3.0162053,2.9144619,2.6715899,2.7569232,2.6157951,2.2449234,2.1891284,2.412308,2.2514873,1.847795,1.5655385,1.972513,2.0709746,1.8970258,1.4473847,0.88943595,0.56451285,0.5218462,0.34133336,0.16082053,0.072205134,0.101743594,0.11158975,0.23630771,0.38728207,0.446359,0.23630771,0.128,0.08205129,0.07548718,0.07876924,0.049230773,0.009846155,0.0,0.052512825,0.108307704,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.04266667,0.20676924,0.26584616,0.55794877,0.45620516,0.016410258,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.009846155,0.013128206,0.013128206,0.016410258,0.03938462,0.032820515,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.03938462,0.14769232,0.16082053,0.08861539,0.02297436,0.0,0.0032820515,0.013128206,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.049230773,0.14112821,0.21989745,0.40369233,0.63343596,0.86317956,1.0633847,1.0633847,0.8992821,0.71548724,0.5874872,0.52512825,0.4594872,0.4135385,0.40697438,0.40369233,0.34133336,0.18051283,0.21661541,0.28882053,0.30194873,0.22646156,0.41025645,0.6235898,0.74830776,0.69251287,0.39384618,0.34133336,0.29538465,0.27897438,0.36102566,0.65312827,1.214359,1.7296412,1.9068719,1.8215386,1.9331284,1.3193847,0.9517949,0.827077,0.9878975,1.5130258,0.9485129,1.0010257,1.0994873,1.1454359,1.5031796,2.2678976,2.858667,2.4057438,1.3062565,1.2209232,1.913436,1.9954873,1.7985642,1.5031796,1.1388719,0.9419488,0.9156924,0.7253334,0.36758977,0.13784617,0.21989745,0.128,0.15097436,0.31507695,0.37743592,0.49230772,0.30851284,0.1148718,0.068923086,0.190359,0.25271797,0.3708718,0.36758977,0.27897438,0.36430773,0.32820517,0.18707694,0.07876924,0.059076928,0.128,0.13456412,0.08533334,0.029538464,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.009846155,0.013128206,0.013128206,0.013128206,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.0032820515,0.0,0.0,0.0032820515,0.016410258,0.0032820515,0.0032820515,0.006564103,0.013128206,0.016410258,0.036102567,0.101743594,0.10502565,0.036102567,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.02297436,0.15753847,0.24615386,0.42994875,0.5349744,0.06564103,0.072205134,0.029538464,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02297436,0.06564103,0.13784617,0.2855385,1.0469744,2.2646155,2.8980515,2.8947694,3.1934361,2.3991797,2.540308,3.3214362,4.0008206,3.3608208,3.0162053,2.6354873,2.5435898,2.546872,1.9364104,2.4352822,2.4418464,2.349949,2.3860514,2.605949,3.4330258,3.945026,4.571898,5.353026,5.943795,6.0685134,5.579488,4.97559,5.3136415,8.214975,8.917334,10.440206,9.622975,7.1581545,7.565129,6.449231,8.342975,9.403078,8.123077,5.3202057,7.8506675,9.120821,7.7948723,4.7261543,2.9440002,1.4080001,0.7089231,0.73517954,1.020718,0.7384616,0.60061544,0.955077,2.5009232,3.8465643,1.4802053,1.5753847,1.0896411,0.9714873,1.2996924,1.2964103,0.65641034,0.24287182,0.04594872,0.006564103,0.013128206,0.016410258,0.036102567,0.049230773,0.049230773,0.04594872,0.06564103,0.07876924,0.08533334,0.08205129,0.07876924,0.049230773,0.036102567,0.026256412,0.016410258,0.016410258,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.072205134,0.35446155,0.71548724,1.0699488,1.3686155,1.6213335,1.3456411,0.81066674,0.28882053,0.02297436,0.032820515,0.07876924,0.14112821,0.17723078,0.10502565,0.049230773,0.02297436,0.006564103,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.0032820515,0.009846155,0.02297436,0.04266667,0.06235898,0.072205134,0.098461546,0.11158975,0.13456412,0.17394873,0.21989745,0.256,0.29210258,0.32820517,0.36102566,0.38400003,0.38728207,0.41025645,0.4266667,0.4266667,0.42338464,0.42338464,0.43323082,0.43323082,0.42994875,0.45292312,0.45292312,0.446359,0.45620516,0.48246157,0.512,0.5349744,0.55794877,0.5940513,0.64000005,0.6695385,0.7187693,0.81066674,0.9419488,1.0929232,1.2471796,1.401436,1.5786668,1.7788719,1.9987694,2.2350771,2.5862565,3.1015387,3.8859491,4.850872,5.7107697,6.9809237,8.14277,8.907488,9.478565,10.564924,12.068104,15.097437,24.33313,45.49908,85.36616,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.01969231,0.029538464,0.055794876,0.052512825,0.17394873,0.35774362,0.32164106,0.08861539,0.059076928,0.24615386,0.8992821,2.487795,0.79097444,0.24615386,0.35774362,0.8467693,1.6771283,1.9593848,3.0818465,4.1091285,4.8672824,5.9667697,3.9154875,4.6211286,5.7731285,6.229334,5.9963083,4.4832826,3.1245131,2.2153847,2.2022567,3.692308,3.9975388,4.3290257,3.761231,2.3827693,1.2964103,0.892718,0.702359,0.4955898,0.29538465,0.380718,0.44307697,0.39384618,0.3314872,0.28225642,0.19692309,0.101743594,0.059076928,0.026256412,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.036102567,0.07876924,0.08533334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.029538464,0.04266667,0.026256412,0.032820515,0.08861539,0.19692309,0.16082053,0.06235898,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.06235898,0.036102567,0.013128206,0.0,0.0032820515,0.016410258,0.016410258,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.029538464,0.128,0.33476925,0.58092314,0.8795898,1.2504616,1.6344616,1.8904617,2.0873847,2.1267693,1.9856411,1.7460514,1.585231,1.4998976,1.3423591,1.0568206,0.69579494,0.4266667,0.3052308,0.36758977,0.5316923,0.65312827,0.51856416,1.2012309,1.8018463,2.1989746,2.0775387,0.9321026,0.7220513,0.6432821,0.508718,0.34789747,0.39712822,0.46933338,0.571077,0.9124103,1.7362052,3.31159,2.297436,1.522872,1.394872,1.4900514,0.5481026,0.512,0.40369233,0.26256412,0.2100513,0.44307697,1.0896411,2.1103592,2.7536411,2.6354873,1.7690258,1.5753847,1.6180514,1.9298463,2.3827693,2.7011285,2.6026669,1.9823592,1.214359,0.56451285,0.19692309,0.2231795,0.14769232,0.23958977,0.4266667,0.3052308,0.14769232,0.098461546,0.108307704,0.15097436,0.21333335,0.2855385,0.23302566,0.14112821,0.068923086,0.04594872,0.02297436,0.016410258,0.02297436,0.029538464,0.029538464,0.01969231,0.006564103,0.0,0.0,0.0,0.0,0.0,0.006564103,0.016410258,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.01969231,0.029538464,0.01969231,0.006564103,0.0,0.0032820515,0.016410258,0.0032820515,0.009846155,0.032820515,0.06564103,0.07548718,0.08861539,0.101743594,0.08205129,0.036102567,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02297436,0.13128206,0.27897438,0.380718,0.32164106,0.3708718,0.15097436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.03938462,0.14112821,0.39712822,0.43323082,1.6246156,2.3991797,2.5928206,3.4494362,3.4855387,3.3214362,3.3312824,3.370667,2.7634873,2.5042052,2.6256413,2.9965131,3.117949,2.1070771,1.6771283,1.6344616,1.7165129,1.8379488,2.1070771,2.1431797,2.546872,3.5282054,4.6145644,4.637539,3.9318976,4.276513,5.58277,7.3353853,8.605539,10.315488,11.539693,10.804514,8.772923,8.224821,9.284924,10.010257,10.9686165,11.83836,11.398565,10.873437,12.389745,10.138257,4.9099493,4.1058464,2.2383592,1.394872,1.0338463,0.94523084,1.2504616,1.3489232,1.2176411,1.8281027,2.6026669,1.4178462,3.4560003,2.7766156,1.8379488,2.0775387,3.9220517,2.4320002,1.0436924,0.23302566,0.02297436,0.0,0.02297436,0.049230773,0.06235898,0.059076928,0.04594872,0.0951795,0.1148718,0.1148718,0.10502565,0.09189744,0.09189744,0.06564103,0.03938462,0.026256412,0.016410258,0.016410258,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.36758977,1.079795,1.5195899,1.4802053,1.1749744,1.0666667,0.98133343,0.6892308,0.256,0.06235898,0.098461546,0.28882053,0.5874872,0.78769237,0.51856416,0.20020515,0.049230773,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.0032820515,0.01969231,0.036102567,0.049230773,0.06235898,0.08533334,0.101743594,0.118153855,0.14769232,0.18379489,0.21989745,0.256,0.29210258,0.3249231,0.33476925,0.34789747,0.38728207,0.41682056,0.42338464,0.4135385,0.4135385,0.4201026,0.4201026,0.4135385,0.4266667,0.4397949,0.44307697,0.45620516,0.47589746,0.48902568,0.49887183,0.512,0.5316923,0.55794877,0.5940513,0.6432821,0.702359,0.78769237,0.90584624,1.0535386,1.1881026,1.3292309,1.4769232,1.6246156,1.7690258,1.9659488,2.3630772,3.0391798,3.9876926,5.110154,6.442667,7.5913854,8.4512825,9.101129,9.796924,10.5780525,14.336001,24.42831,42.686363,69.39898,0.15753847,0.032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.029538464,0.04266667,0.055794876,0.06564103,0.07548718,0.08533334,0.08861539,0.06235898,0.10502565,0.17066668,0.30851284,0.6432821,0.49887183,0.50543594,0.69251287,0.955077,1.0436924,1.1684103,1.2996924,2.048,3.249231,3.9778464,3.820308,4.128821,4.571898,4.9788723,5.3136415,4.46359,4.20759,4.516103,4.7950773,3.8990772,3.5511796,4.020513,4.2207184,3.6102567,2.1989746,2.7142565,2.9636924,2.5271797,1.5327181,0.6498462,0.8369231,1.0108719,1.0962052,1.014154,0.67282057,0.4397949,0.25928208,0.15097436,0.098461546,0.06235898,0.013128206,0.0,0.01969231,0.03938462,0.0,0.0,0.013128206,0.01969231,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02297436,0.09189744,0.13784617,0.0,0.0,0.006564103,0.016410258,0.016410258,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.08533334,0.0951795,0.07876924,0.07876924,0.15097436,0.14112821,0.098461546,0.118153855,0.17066668,0.12143591,0.02297436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.006564103,0.0032820515,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.04266667,0.15097436,0.5152821,0.9878975,1.4408206,1.785436,2.0020514,2.0808206,2.0906668,2.0184617,1.910154,1.8806155,1.8248206,1.7755898,1.6968206,1.595077,1.4998976,1.214359,0.99774367,0.85005134,0.76800007,0.7515898,1.1224617,1.595077,1.785436,1.6278975,1.3686155,1.2012309,0.90584624,0.6301539,0.45620516,0.41025645,0.43323082,0.5284103,0.53825647,0.75487185,1.9200002,2.3433847,1.5458462,1.3292309,1.8248206,1.4998976,1.3292309,0.76800007,0.3708718,0.3052308,0.3314872,0.636718,1.0535386,1.3193847,1.2931283,0.9517949,0.9124103,1.1257436,1.847795,2.7109745,2.7241027,2.1891284,1.7165129,1.2406155,0.7844103,0.4660513,0.40369233,0.29210258,0.2100513,0.18379489,0.15753847,0.16738462,0.16738462,0.15753847,0.14441027,0.128,0.0951795,0.06235898,0.036102567,0.013128206,0.009846155,0.0032820515,0.0032820515,0.0032820515,0.006564103,0.006564103,0.0032820515,0.0,0.0032820515,0.013128206,0.013128206,0.0032820515,0.0,0.0,0.006564103,0.016410258,0.02297436,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.036102567,0.1148718,0.04594872,0.01969231,0.006564103,0.0032820515,0.016410258,0.013128206,0.013128206,0.02297436,0.04594872,0.08861539,0.072205134,0.09189744,0.08861539,0.049230773,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.026256412,0.08861539,0.17723078,0.2231795,0.2231795,0.24943592,0.16082053,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.013128206,0.036102567,0.0951795,0.21333335,0.14441027,0.4201026,0.83035904,1.3226668,2.0217438,3.6890259,4.017231,3.8695388,3.4921029,2.5304618,3.308308,5.398975,6.12759,4.6900516,2.1431797,1.4309745,1.5163078,1.9823592,2.5435898,3.045744,2.553436,2.665026,3.2131286,4.086154,5.211898,4.857436,5.031385,5.431795,5.83877,6.1538467,8.0377445,8.940309,8.946873,8.684308,9.298052,10.916103,10.315488,9.573745,9.737847,10.811078,11.421539,14.516514,13.308719,7.584821,3.7021542,2.0873847,1.273436,1.0699488,1.1782565,1.1913847,1.0338463,1.1093334,1.7657437,2.546872,2.2121027,5.159385,5.5171285,4.9099493,4.6145644,5.5696416,5.4482055,4.342154,3.4625645,2.6420515,0.34133336,0.39712822,0.20676924,0.08205129,0.0951795,0.08205129,0.08205129,0.08533334,0.07876924,0.068923086,0.06564103,0.08533334,0.09189744,0.07548718,0.036102567,0.016410258,0.026256412,0.026256412,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.60061544,1.1323078,1.5327181,1.657436,1.273436,1.0371283,0.7318975,0.41025645,0.14441027,0.036102567,0.11158975,0.6071795,1.0535386,1.2012309,1.020718,0.79097444,0.5874872,0.35774362,0.128,0.013128206,0.0032820515,0.0,0.0,0.0,0.0032820515,0.0,0.009846155,0.02297436,0.03938462,0.06235898,0.08533334,0.101743594,0.1148718,0.13128206,0.15753847,0.20348719,0.23630771,0.26256412,0.2855385,0.2986667,0.32164106,0.34789747,0.37415388,0.39384618,0.4135385,0.4135385,0.4201026,0.4201026,0.4135385,0.4135385,0.43651286,0.44964105,0.45620516,0.46276927,0.46276927,0.47589746,0.4955898,0.508718,0.51856416,0.5349744,0.5940513,0.64000005,0.69579494,0.7778462,0.892718,0.99774367,1.0929232,1.1881026,1.3029745,1.4408206,1.6246156,1.9035898,2.3466668,3.1343591,4.5489235,6.3606157,7.6110773,8.375795,8.950154,9.882257,10.604308,13.833847,22.327797,33.33908,38.623184,0.3446154,0.4266667,0.6071795,0.48574364,0.118153855,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.01969231,0.02297436,0.049230773,0.10502565,0.15097436,0.10502565,0.049230773,0.072205134,0.118153855,0.19364104,0.35774362,0.571077,0.53825647,0.4660513,0.4594872,0.5021539,0.702359,1.1060513,1.9265642,2.9669745,3.6168208,4.013949,3.8137438,3.3280003,3.0162053,3.4756925,3.8400004,4.2929235,4.4340515,4.164923,3.6758976,4.585026,4.384821,4.9493337,5.586052,3.0227695,2.7995899,3.3444104,3.446154,2.934154,2.7044106,1.9331284,1.3718976,1.404718,1.9232821,2.3401027,1.6607181,1.404718,1.0994873,0.7187693,0.69907695,0.5874872,0.4004103,0.2297436,0.128,0.108307704,0.06564103,0.03938462,0.11158975,0.21661541,0.14769232,0.052512825,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.04594872,0.068923086,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03938462,0.04594872,0.036102567,0.029538464,0.055794876,0.098461546,0.09189744,0.10502565,0.128,0.08861539,0.03938462,0.032820515,0.059076928,0.072205134,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01969231,0.098461546,0.6498462,1.0994873,1.0994873,0.8598975,1.142154,1.4900514,1.6082052,1.7066668,1.8642052,2.0184617,2.0053334,1.9922053,2.0217438,2.0709746,2.044718,1.8116925,1.8182565,1.8806155,1.8806155,1.8051283,1.9462565,2.1989746,2.2482052,2.0578463,1.8838975,1.7099489,1.404718,1.0929232,0.84348726,0.6695385,0.52512825,0.45620516,0.61374366,1.0633847,1.7723079,1.9987694,1.4998976,1.2603078,1.3522053,0.9714873,0.98133343,0.702359,0.47261542,0.43323082,0.52512825,0.5481026,0.93866676,1.2373334,1.2274873,0.9321026,0.9321026,1.1158975,1.5491283,2.0118976,2.0086155,1.6836925,1.4375386,1.2668719,1.142154,1.0272821,0.86317956,0.6498462,0.44307697,0.2986667,0.26912823,0.28225642,0.23302566,0.15753847,0.08205129,0.06235898,0.029538464,0.013128206,0.0032820515,0.006564103,0.026256412,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.006564103,0.0,0.0,0.0,0.0,0.006564103,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.04266667,0.20020515,0.57764107,0.6071795,0.26256412,0.01969231,0.02297436,0.07876924,0.12471796,0.128,0.118153855,0.101743594,0.101743594,0.04594872,0.055794876,0.0951795,0.11158975,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.026256412,0.055794876,0.10502565,0.24287182,0.16738462,0.18707694,0.18051283,0.10502565,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.04594872,0.049230773,0.068923086,0.055794876,0.036102567,0.08533334,0.07548718,0.12471796,0.30851284,0.69251287,1.3062565,3.4330258,4.519385,4.571898,3.8564105,2.8914874,3.6758976,5.221744,5.3694363,3.8367183,2.225231,2.484513,3.3641028,3.9876926,4.0434875,3.7842054,4.7425647,4.7294364,4.2469745,4.086154,5.3366156,5.031385,5.832206,7.000616,7.79159,7.460103,6.678975,7.1647186,7.9852314,8.907488,10.381129,12.1928215,11.011283,10.9226675,11.529847,7.975385,12.324103,15.2155905,13.4170265,8.254359,5.6320004,3.3936412,2.0118976,1.4933335,1.4998976,1.3686155,1.8215386,1.8970258,1.8937438,2.1300514,2.9604106,4.9854364,5.4875903,5.8847184,6.5345645,6.741334,6.2720003,5.8190775,6.0225644,6.0947695,3.7973337,1.1618463,0.34133336,0.17394873,0.08533334,0.072205134,0.068923086,0.06235898,0.055794876,0.052512825,0.052512825,0.068923086,0.08861539,0.08533334,0.059076928,0.04266667,0.049230773,0.04266667,0.026256412,0.009846155,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.29210258,0.82379496,1.3653334,1.6902566,1.5819489,1.5031796,1.1191796,0.58092314,0.13456412,0.12143591,0.07548718,0.27897438,0.53825647,0.72861546,0.8041026,0.7581539,0.60061544,0.4004103,0.21333335,0.06235898,0.013128206,0.0,0.0,0.0,0.0,0.006564103,0.013128206,0.026256412,0.04266667,0.06235898,0.08533334,0.101743594,0.12143591,0.14441027,0.16082053,0.19692309,0.21661541,0.23958977,0.26256412,0.28225642,0.3052308,0.3249231,0.34133336,0.36102566,0.38400003,0.4004103,0.4135385,0.42338464,0.42994875,0.42994875,0.4397949,0.45292312,0.45620516,0.4594872,0.4660513,0.47917953,0.4955898,0.5021539,0.50543594,0.508718,0.5546667,0.60061544,0.6498462,0.7089231,0.79097444,0.85005134,0.92225647,1.014154,1.1257436,1.2406155,1.3915899,1.6213335,1.9396925,2.4549747,3.3575387,5.1232824,6.889026,8.208411,9.081436,9.96759,10.397539,11.67754,14.998976,18.770052,18.609232,0.26584616,0.42994875,1.7920002,2.605949,2.1530259,0.761436,0.17723078,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.026256412,0.11158975,0.20348719,0.15753847,0.08205129,0.07548718,0.13128206,0.24615386,0.42338464,0.49887183,0.44964105,0.5316923,0.78769237,1.0666667,1.1093334,1.585231,1.9429746,2.1989746,2.9440002,3.3969233,3.255795,2.5796926,1.8281027,1.8904617,2.425436,2.9407182,3.1803079,3.1770258,3.2853336,4.59159,4.923077,6.226052,7.4929237,4.7917953,3.1343591,3.3280003,3.5413337,3.2164104,3.0949745,2.0709746,1.3686155,1.2307693,1.595077,2.097231,1.5655385,1.4244103,1.1913847,0.9124103,1.1881026,1.2176411,0.86317956,0.60389745,0.6268718,0.8369231,0.33476925,0.13456412,0.74830776,1.4605129,0.33476925,0.108307704,0.01969231,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.006564103,0.013128206,0.18707694,0.21661541,0.2297436,0.25271797,0.18051283,0.16410258,0.08533334,0.059076928,0.072205134,0.0,0.0,0.006564103,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.029538464,0.14769232,0.65969235,1.0962052,0.9485129,0.45292312,0.5874872,0.75487185,0.81394875,0.9517949,1.2438976,1.6738462,1.9856411,1.9954873,1.9331284,2.038154,2.556718,2.3433847,2.1924105,2.3138463,2.540308,2.3368206,2.6223593,2.6420515,2.550154,2.422154,2.2547693,2.028308,1.7001027,1.401436,1.1552821,0.85005134,0.65969235,0.57764107,0.7253334,1.0436924,1.2898463,1.2570257,1.1520001,1.0699488,0.9714873,0.6892308,0.81394875,0.86317956,0.88287187,0.9485129,1.1716924,1.2242053,1.6443079,1.9035898,1.7591796,1.2603078,1.4506668,1.7460514,1.9429746,1.9889232,1.9790771,1.7690258,1.657436,1.5622566,1.467077,1.4080001,1.2176411,0.97805136,0.71548724,0.47589746,0.33476925,0.28882053,0.2100513,0.118153855,0.03938462,0.01969231,0.009846155,0.013128206,0.009846155,0.006564103,0.026256412,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.052512825,0.19364104,0.5415385,0.6268718,0.28225642,0.029538464,0.03938462,0.10502565,0.13784617,0.13784617,0.12143591,0.101743594,0.07548718,0.04594872,0.04266667,0.07548718,0.101743594,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.026256412,0.04266667,0.072205134,0.19692309,0.12143591,0.0951795,0.118153855,0.14441027,0.059076928,0.029538464,0.009846155,0.009846155,0.01969231,0.006564103,0.07876924,0.098461546,0.118153855,0.14441027,0.13784617,0.098461546,0.0951795,0.06235898,0.013128206,0.01969231,0.049230773,0.08533334,0.15097436,0.34789747,0.84348726,2.6322052,3.508513,3.8038976,3.6332312,2.8816411,4.532513,5.464616,4.9296412,3.5183592,3.170462,4.023795,4.9099493,5.543385,5.910975,6.262154,7.7390776,7.3682055,6.2588725,5.671385,7.0334363,7.017026,7.6767187,8.953437,10.354873,10.981745,10.085744,11.158976,11.355898,11.369026,15.415796,13.725539,11.480617,12.481642,14.815181,10.840616,15.067899,18.448412,15.868719,9.412924,8.372514,5.8912826,4.2896414,3.1737437,2.4024618,2.1103592,2.8980515,3.56759,3.1474874,2.4615386,4.132103,5.2480006,5.7009234,5.9470773,6.265436,6.7774363,6.38359,6.987488,7.7981544,7.9917955,6.7249236,3.0030773,1.273436,0.54482055,0.256,0.26256412,0.26584616,0.13456412,0.04594872,0.04594872,0.04594872,0.052512825,0.06564103,0.072205134,0.06564103,0.055794876,0.04594872,0.036102567,0.029538464,0.01969231,0.016410258,0.006564103,0.0032820515,0.0,0.0,0.0,0.029538464,0.380718,0.84348726,1.2570257,1.5064616,1.6935385,1.4834872,0.98461545,0.4135385,0.12143591,0.032820515,0.0032820515,0.068923086,0.2100513,0.34789747,0.39056414,0.318359,0.22646156,0.15097436,0.055794876,0.036102567,0.016410258,0.0032820515,0.0,0.0,0.013128206,0.016410258,0.026256412,0.04266667,0.06235898,0.08533334,0.101743594,0.12143591,0.15097436,0.16082053,0.18707694,0.20348719,0.2231795,0.24287182,0.26256412,0.28225642,0.30194873,0.32164106,0.33805132,0.36758977,0.38728207,0.40369233,0.42338464,0.446359,0.45620516,0.45620516,0.46276927,0.47261542,0.47917953,0.48574364,0.49230772,0.5021539,0.512,0.51856416,0.5218462,0.55794877,0.5973334,0.6432821,0.69907695,0.75487185,0.8041026,0.88287187,0.98461545,1.0896411,1.1716924,1.3095386,1.5327181,1.7887181,2.0906668,2.4910772,3.7349746,5.431795,6.9842057,8.28718,9.741129,10.171078,10.102155,9.764103,9.222565,8.352821,0.0032820515,0.03938462,2.3696413,4.2371287,4.089436,1.591795,0.38400003,0.032820515,0.029538464,0.059076928,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.013128206,0.013128206,0.009846155,0.013128206,0.06235898,0.13128206,0.15097436,0.14441027,0.128,0.18707694,0.3314872,0.49887183,0.54482055,0.7220513,1.2307693,1.9528207,2.4320002,2.0709746,1.9626669,1.4802053,0.9747693,1.782154,1.9987694,2.2777438,2.1431797,1.6640002,1.4736412,1.2996924,1.339077,1.9331284,2.7503593,2.8160002,3.114667,4.71959,6.636308,7.650462,6.3310776,3.9581542,3.3214362,2.9505644,2.3072822,1.785436,1.4572309,1.2209232,0.8763078,0.47589746,0.33805132,0.42338464,0.45292312,0.42338464,0.512,1.0568206,1.2996924,0.955077,0.82379496,1.1684103,1.7460514,1.0043077,0.86974365,1.9429746,2.8849232,0.4135385,0.14769232,0.032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.013128206,0.01969231,0.04266667,0.37743592,0.4135385,0.41682056,0.44307697,0.33476925,0.3052308,0.14769232,0.052512825,0.059076928,0.049230773,0.009846155,0.013128206,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.036102567,0.18707694,0.43651286,0.8369231,0.90912825,0.6432821,0.512,0.19364104,0.08205129,0.11158975,0.3249231,0.88287187,1.4867693,1.5195899,1.394872,1.5688206,2.540308,2.3269746,1.8084104,1.7657437,2.1234872,1.9462565,2.4516926,2.3401027,2.2153847,2.2580514,2.2121027,1.9495386,1.6016412,1.3718976,1.2307693,0.9189744,0.7975385,0.8598975,0.8205129,0.6662565,0.65312827,0.79097444,0.96492314,1.1520001,1.3423591,1.5425643,1.6836925,1.910154,2.1825643,2.4188719,2.4943593,2.8225644,3.1474874,3.1277952,2.6978464,2.0676925,2.4549747,2.7995899,2.878359,2.7175386,2.5928206,2.2580514,2.097231,1.8576412,1.5392822,1.3751796,1.204513,1.017436,0.78769237,0.51856416,0.23302566,0.15425642,0.098461546,0.059076928,0.029538464,0.0,0.0,0.02297436,0.02297436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.029538464,0.032820515,0.026256412,0.049230773,0.08205129,0.055794876,0.032820515,0.036102567,0.06564103,0.04594872,0.029538464,0.029538464,0.03938462,0.029538464,0.055794876,0.04594872,0.032820515,0.02297436,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.032820515,0.06564103,0.06564103,0.03938462,0.04594872,0.08861539,0.108307704,0.068923086,0.029538464,0.026256412,0.049230773,0.032820515,0.2297436,0.31507695,0.38400003,0.41682056,0.30194873,0.190359,0.0951795,0.03938462,0.01969231,0.0032820515,0.006564103,0.029538464,0.055794876,0.15097436,0.45620516,1.4572309,1.4276924,1.7887181,2.674872,2.9440002,5.0642056,5.72718,5.277539,4.519385,4.706462,6.1341543,5.8256416,5.970052,7.3419495,9.284924,9.724719,9.124104,8.1755905,7.817847,9.216001,9.67877,9.869129,10.5780525,12.153437,14.464001,16.177233,17.99877,16.269129,13.735386,19.570873,13.833847,10.84718,12.232206,16.082052,16.94195,18.914463,23.105642,19.72513,11.008,11.195078,8.201847,6.5312824,4.9920006,3.6004105,3.5741541,3.767795,4.827898,4.7360005,3.7776413,4.5423594,5.9634876,7.1680007,6.5247183,4.9427695,5.85518,6.242462,7.312411,7.6931286,7.282872,7.243488,6.4295387,3.6890259,1.7558975,1.4473847,1.6672822,1.1093334,0.4201026,0.055794876,0.055794876,0.052512825,0.04594872,0.04266667,0.049230773,0.052512825,0.04266667,0.01969231,0.016410258,0.02297436,0.029538464,0.01969231,0.01969231,0.009846155,0.0032820515,0.0,0.0032820515,0.0,0.029538464,0.18707694,0.49230772,0.90256417,1.2340513,1.3193847,1.1323078,0.6892308,0.032820515,0.009846155,0.0,0.0,0.0,0.0,0.009846155,0.013128206,0.013128206,0.01969231,0.036102567,0.09189744,0.055794876,0.016410258,0.0032820515,0.0,0.009846155,0.013128206,0.02297436,0.036102567,0.059076928,0.08205129,0.098461546,0.118153855,0.13784617,0.15097436,0.17723078,0.20020515,0.21989745,0.23630771,0.24615386,0.26256412,0.29210258,0.31507695,0.33476925,0.3708718,0.38400003,0.40697438,0.43323082,0.45620516,0.47917953,0.48246157,0.48902568,0.49887183,0.508718,0.508718,0.5152821,0.5218462,0.5349744,0.5481026,0.56123084,0.5973334,0.6268718,0.6695385,0.7253334,0.7778462,0.84348726,0.93866676,1.0404103,1.1355898,1.2176411,1.3620514,1.5688206,1.7723079,1.9593848,2.166154,2.7076926,3.6627696,4.850872,6.3573337,8.549745,9.314463,9.32759,8.51036,7.056411,5.428513,0.016410258,0.0032820515,0.0,0.0,0.068923086,0.33476925,0.15097436,0.04266667,0.14769232,0.29210258,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01969231,0.04266667,0.06235898,0.06235898,0.049230773,0.036102567,0.02297436,0.026256412,0.07548718,0.15097436,0.12143591,0.19692309,0.49887183,1.083077,1.7657437,2.2121027,2.412308,2.5435898,2.9440002,2.409026,1.595077,1.1093334,1.1848207,1.7099489,0.9878975,0.94523084,1.1158975,1.522872,2.6715899,2.8160002,2.294154,1.8609232,1.8510771,2.1825643,1.7657437,2.422154,3.0949745,3.5249233,4.2568207,3.757949,2.6518977,1.657436,1.3456411,2.1530259,2.162872,1.4802053,0.9485129,0.86317956,0.9616411,0.99774367,0.82379496,0.46276927,0.10502565,0.09189744,0.14112821,0.14441027,0.27897438,0.6826667,1.463795,2.3433847,3.3312824,3.2525132,1.9298463,0.18379489,0.15753847,0.06235898,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01969231,0.09189744,0.446359,0.40697438,0.2297436,0.10502565,0.15097436,0.15097436,0.19692309,0.25928208,0.29210258,0.24287182,0.049230773,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.08861539,0.16082053,0.12471796,0.013128206,0.0,0.013128206,0.006564103,0.006564103,0.016410258,0.016410258,0.016410258,0.04266667,0.4397949,0.90256417,0.48902568,0.5481026,0.69251287,0.77128214,0.85005134,1.1913847,1.079795,1.0994873,1.3357949,1.6016412,1.4178462,1.273436,1.1913847,1.142154,1.1126155,1.1126155,0.9419488,1.0108719,1.204513,1.4703591,1.8018463,1.9593848,2.100513,2.3991797,2.9111798,3.570872,3.9745643,4.522667,5.2315903,5.6287184,4.775385,5.2512827,5.5269747,5.1298466,4.315898,4.059898,4.082872,3.6758976,3.121231,2.6322052,2.349949,2.0808206,1.7033848,1.3489232,1.0962052,0.9616411,0.69251287,0.47917953,0.38728207,0.318359,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01969231,0.036102567,0.049230773,0.06235898,0.02297436,0.006564103,0.006564103,0.016410258,0.016410258,0.016410258,0.006564103,0.006564103,0.01969231,0.029538464,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.016410258,0.032820515,0.04594872,0.049230773,0.06235898,0.049230773,0.04594872,0.03938462,0.04594872,0.108307704,0.3511795,0.60389745,0.7450257,0.72861546,0.5940513,0.42338464,0.15097436,0.0,0.0032820515,0.016410258,0.03938462,0.072205134,0.108307704,0.16082053,0.25928208,0.3446154,0.5021539,0.61374366,1.5031796,4.95918,2.7142565,1.8215386,3.1409233,5.4514875,5.4613338,9.770667,7.7357955,6.124308,7.1614366,8.530052,8.041026,8.461129,8.241231,7.433847,7.6898465,8.201847,10.006975,11.808822,13.2562065,14.953027,16.968206,16.902565,13.686155,9.38995,9.232411,8.523488,7.9819493,8.664616,10.7158985,13.351386,20.883694,23.003899,17.700104,10.440206,14.17518,7.8408213,4.900103,3.8498464,4.0500517,5.720616,4.2568207,3.1113849,4.1452312,5.4449234,1.3423591,4.84759,8.861539,9.288206,6.4295387,4.9887185,5.3070774,4.204308,3.6496413,4.2436924,5.218462,11.785847,8.136206,4.7228723,5.1331286,6.0717955,3.239385,1.0666667,0.09189744,0.08861539,0.07548718,0.052512825,0.036102567,0.029538464,0.029538464,0.029538464,0.01969231,0.016410258,0.02297436,0.029538464,0.029538464,0.029538464,0.029538464,0.01969231,0.0032820515,0.016410258,0.0032820515,0.0,0.0,0.013128206,0.06235898,0.15753847,0.256,0.27569234,0.19364104,0.04594872,0.02297436,0.006564103,0.0,0.0,0.0,0.0,0.0,0.029538464,0.098461546,0.18379489,0.21989745,0.128,0.04266667,0.013128206,0.0,0.0,0.009846155,0.02297436,0.032820515,0.04594872,0.068923086,0.0951795,0.11158975,0.128,0.15097436,0.17723078,0.20020515,0.22646156,0.24615386,0.25928208,0.28225642,0.30851284,0.3314872,0.35774362,0.380718,0.40697438,0.4397949,0.46276927,0.47917953,0.5021539,0.5152821,0.51856416,0.51856416,0.5218462,0.5349744,0.55794877,0.56451285,0.571077,0.5874872,0.6104616,0.63343596,0.67610264,0.7187693,0.764718,0.8402052,0.8763078,0.93866676,1.0371283,1.1684103,1.3259488,1.4605129,1.5786668,1.6705642,1.7526156,1.8609232,2.0676925,2.422154,3.0654361,4.059898,5.402257,6.3901544,7.571693,7.686565,6.73477,5.9667697,0.4660513,0.446359,0.32164106,0.14769232,0.01969231,0.09189744,1.1388719,1.8773335,1.6246156,0.636718,0.108307704,0.02297436,0.013128206,0.02297436,0.01969231,0.0,0.009846155,0.0032820515,0.009846155,0.01969231,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.036102567,0.072205134,0.108307704,0.17723078,0.37415388,0.40369233,0.24943592,0.16082053,0.22646156,0.18051283,0.11158975,0.128,0.3511795,0.54482055,0.57764107,0.54482055,0.5316923,0.60061544,0.8763078,1.3489232,1.7591796,1.9035898,1.6475899,1.0633847,0.79097444,0.7384616,0.98461545,1.7920002,2.0841026,3.1967182,3.8137438,3.8564105,4.4898467,3.4691284,2.5600002,2.162872,2.4582565,3.4133337,3.4133337,3.239385,2.7798977,2.0611284,1.2373334,1.083077,0.9419488,1.204513,2.0644104,3.5478978,3.0293336,1.8445129,0.83035904,0.35446155,0.3249231,0.256,0.19364104,0.18051283,0.23302566,0.34133336,0.5481026,0.8467693,0.9616411,0.77128214,0.3052308,0.08533334,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.04266667,0.0951795,0.036102567,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.01969231,0.18707694,0.13128206,0.20676924,0.43651286,0.4955898,0.47589746,0.5218462,0.63343596,0.69907695,0.512,0.2100513,0.17066668,0.118153855,0.0,0.0,0.049230773,0.08205129,0.059076928,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.032820515,0.026256412,0.0032820515,0.0,0.0032820515,0.0,0.006564103,0.013128206,0.0032820515,0.0032820515,0.009846155,0.09189744,0.190359,0.098461546,0.21661541,0.28882053,0.3511795,0.43651286,0.54482055,0.8533334,1.0043077,1.0305642,0.9485129,0.7844103,0.84348726,0.9156924,0.9682052,1.017436,1.1257436,1.2176411,1.3751796,1.5688206,1.8379488,2.2646155,2.8324106,3.1934361,3.4494362,3.692308,4.010667,4.33559,4.7392826,5.037949,5.106872,4.896821,4.699898,4.630975,4.3716927,3.9286156,3.6430771,3.4133337,2.9144619,2.3794873,1.9396925,1.6311796,1.3718976,1.0765129,0.7844103,0.5349744,0.36430773,0.2297436,0.12471796,0.07876924,0.06235898,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.01969231,0.02297436,0.02297436,0.016410258,0.013128206,0.01969231,0.026256412,0.026256412,0.026256412,0.026256412,0.068923086,0.12471796,0.06564103,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.006564103,0.013128206,0.016410258,0.013128206,0.02297436,0.06235898,0.049230773,0.04594872,0.068923086,0.08205129,0.3249231,0.5513847,0.7778462,0.88287187,0.58420515,0.4201026,0.31507695,0.23958977,0.16082053,0.026256412,0.032820515,0.03938462,0.08533334,0.17066668,0.24615386,0.3511795,0.39056414,0.40369233,0.6170257,1.4572309,2.2482052,2.7798977,3.43959,4.1156926,4.204308,5.0477953,6.048821,8.530052,11.477334,11.556104,8.792616,6.695385,5.733744,6.265436,8.533334,9.055181,9.659078,12.2847185,14.700309,10.499283,12.025436,11.516719,11.1983595,11.0375395,8.730257,10.121847,8.500513,7.496206,8.369231,10.020103,12.005745,12.511181,12.530872,13.046155,15.05477,8.874667,7.2336416,6.889026,6.918565,8.736821,8.073847,6.550975,5.9667697,5.927385,3.8564105,5.8289237,10.860309,12.320822,9.337437,6.7840004,4.7950773,3.4494362,3.2656412,3.623385,2.7634873,9.419488,9.278359,5.9930263,3.170462,4.3651285,2.412308,0.9616411,0.2986667,0.22646156,0.08861539,0.318359,0.21989745,0.08205129,0.029538464,0.01969231,0.006564103,0.009846155,0.016410258,0.01969231,0.01969231,0.029538464,0.029538464,0.029538464,0.026256412,0.026256412,0.016410258,0.0032820515,0.0,0.0032820515,0.013128206,0.032820515,0.052512825,0.055794876,0.03938462,0.009846155,0.013128206,0.16738462,0.37743592,0.512,0.4135385,0.33805132,0.30194873,0.380718,0.512,0.49887183,0.26256412,0.08861539,0.009846155,0.0032820515,0.0,0.0,0.009846155,0.016410258,0.02297436,0.032820515,0.068923086,0.08861539,0.0951795,0.10502565,0.128,0.16082053,0.19692309,0.2297436,0.26256412,0.28225642,0.30851284,0.3314872,0.3511795,0.3708718,0.39384618,0.40697438,0.43323082,0.45292312,0.4660513,0.49230772,0.512,0.51856416,0.52512825,0.5349744,0.55794877,0.574359,0.5973334,0.61374366,0.62030774,0.63343596,0.6498462,0.6826667,0.7089231,0.72861546,0.75487185,0.79097444,0.8402052,0.90912825,1.0010257,1.1191796,1.1848207,1.2635899,1.3686155,1.5064616,1.654154,1.7427694,1.8937438,2.162872,2.6026669,3.2525132,4.97559,5.58277,6.2720003,7.2205133,7.6143594,0.955077,1.3784616,1.3193847,0.92225647,0.42338464,0.17723078,1.1815386,1.6443079,1.4769232,0.8763078,0.32164106,0.1148718,0.03938462,0.032820515,0.052512825,0.072205134,0.055794876,0.036102567,0.029538464,0.029538464,0.026256412,0.036102567,0.013128206,0.013128206,0.03938462,0.055794876,0.026256412,0.036102567,0.068923086,0.08533334,0.01969231,0.0032820515,0.029538464,0.101743594,0.16738462,0.12143591,0.30851284,0.636718,0.6465641,0.3314872,0.13784617,0.17066668,0.28882053,0.26256412,0.10502565,0.08533334,0.108307704,0.072205134,0.029538464,0.013128206,0.016410258,0.22646156,0.67282057,1.270154,1.8970258,2.3827693,1.847795,1.0666667,0.58420515,0.5677949,0.81066674,0.9288206,1.972513,3.045744,3.8400004,4.644103,4.850872,3.639795,2.3072822,1.6935385,2.2153847,2.740513,2.9440002,2.5796926,1.8018463,1.1618463,0.702359,0.5677949,0.7417436,1.2996924,2.4188719,1.9068719,1.6607181,1.5261539,1.404718,1.2504616,0.9911796,0.79097444,0.5546667,0.2855385,0.07876924,0.049230773,0.108307704,0.18051283,0.20676924,0.13456412,0.026256412,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02297436,0.049230773,0.01969231,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0,0.049230773,0.02297436,0.22646156,0.61374366,0.8008206,0.67938465,0.60061544,0.6432821,0.7253334,0.6071795,0.42338464,0.512,0.5152821,0.35446155,0.23958977,0.14441027,0.11158975,0.06564103,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.01969231,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0,0.052512825,0.07548718,0.098461546,0.13456412,0.16082053,0.36430773,0.5349744,0.65969235,0.7122052,0.67282057,0.8402052,0.9189744,0.9288206,0.9156924,0.94523084,0.9353847,1.0535386,1.2603078,1.5163078,1.785436,2.0545642,2.4549747,2.665026,2.6617439,2.7470772,3.117949,3.2164104,3.2229745,3.2098465,3.1606157,2.9801028,2.8258464,2.6256413,2.3729234,2.1398976,1.8904617,1.5491283,1.214359,0.9321026,0.7187693,0.5546667,0.4135385,0.27897438,0.15753847,0.08533334,0.04594872,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.009846155,0.016410258,0.02297436,0.032820515,0.04266667,0.04266667,0.013128206,0.013128206,0.02297436,0.029538464,0.02297436,0.013128206,0.016410258,0.059076928,0.098461546,0.03938462,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.0,0.013128206,0.02297436,0.016410258,0.0,0.006564103,0.0,0.0032820515,0.006564103,0.009846155,0.016410258,0.04266667,0.032820515,0.032820515,0.059076928,0.0951795,0.26584616,0.5284103,0.7089231,0.7122052,0.52512825,0.41682056,0.31507695,0.2231795,0.13128206,0.013128206,0.01969231,0.016410258,0.06564103,0.16082053,0.22646156,0.27569234,0.256,0.24615386,0.7844103,2.8488207,2.986667,3.1343591,3.692308,4.9985647,7.3419495,7.213949,7.5454364,8.697436,9.718155,8.333129,7.6734366,9.731283,9.984001,7.8736415,6.820103,9.314463,10.092308,11.168821,12.248616,10.70277,10.187488,10.345026,11.116308,11.428103,9.193027,8.861539,10.026668,10.226872,9.03877,8.077128,13.348104,11.280411,9.810052,11.188514,11.979488,9.02236,9.780514,9.055181,6.3179493,5.681231,14.8709755,12.2847185,8.195283,6.672411,5.5565133,6.8496413,9.442462,10.299078,9.130668,8.375795,5.182359,2.8422565,2.0250258,2.2777438,2.0151796,6.2818465,10.203898,9.035488,4.3651285,4.128821,3.370667,1.4178462,0.23630771,0.20676924,0.13784617,0.256,0.3052308,0.28882053,0.20020515,0.032820515,0.006564103,0.009846155,0.013128206,0.006564103,0.006564103,0.01969231,0.02297436,0.026256412,0.029538464,0.029538464,0.026256412,0.01969231,0.013128206,0.009846155,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0032820515,0.18051283,0.42994875,0.64000005,0.702359,0.7515898,0.6465641,0.5874872,0.5677949,0.37743592,0.13784617,0.032820515,0.0,0.0,0.0,0.0,0.009846155,0.01969231,0.026256412,0.03938462,0.055794876,0.07876924,0.098461546,0.1148718,0.14112821,0.17723078,0.20676924,0.23958977,0.27569234,0.2986667,0.31507695,0.33476925,0.34789747,0.36102566,0.3708718,0.38728207,0.40697438,0.42338464,0.446359,0.46933338,0.48574364,0.5021539,0.5152821,0.5316923,0.56451285,0.5907693,0.62030774,0.64000005,0.6465641,0.6498462,0.65641034,0.67282057,0.6859488,0.6892308,0.6859488,0.7089231,0.73517954,0.764718,0.81066674,0.88615394,0.92553854,0.9878975,1.0732309,1.1749744,1.2537436,1.3095386,1.404718,1.5589745,1.785436,2.0841026,3.0358977,3.5347695,4.266667,5.4875903,7.026872,1.0043077,1.4375386,1.4703591,1.2832822,1.1684103,1.5392822,1.0043077,0.8008206,0.7844103,0.77456415,0.5349744,0.24943592,0.13128206,0.08861539,0.07876924,0.12143591,0.08205129,0.059076928,0.108307704,0.20348719,0.23958977,0.12471796,0.04266667,0.08533334,0.571077,2.0578463,2.2219489,1.8412309,1.3554872,0.8992821,0.3117949,0.072205134,0.06235898,0.23958977,0.46933338,0.5316923,0.47917953,0.5316923,0.446359,0.2100513,0.06564103,0.072205134,0.21333335,0.23958977,0.12143591,0.06564103,0.036102567,0.029538464,0.01969231,0.009846155,0.02297436,0.032820515,0.15753847,0.5021539,1.1093334,1.9561027,1.6082052,0.92225647,0.4660513,0.4266667,0.6170257,0.636718,1.2931283,2.1234872,2.8849232,3.5478978,4.46359,3.7316926,2.4320002,1.467077,1.5425643,2.1366155,2.4057438,2.2449234,1.8084104,1.5097437,1.2209232,1.4080001,1.5031796,1.4145643,1.5360001,1.1290257,1.5458462,2.169436,2.5600002,2.4549747,2.0906668,1.8051283,1.6114873,1.3357949,0.6104616,0.17066668,0.03938462,0.04594872,0.06564103,0.04266667,0.01969231,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.15097436,0.40697438,0.5677949,0.4660513,0.39384618,0.45292312,0.574359,0.49230772,0.53825647,0.71548724,0.764718,0.6170257,0.40369233,0.26256412,0.21333335,0.16082053,0.072205134,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.032820515,0.09189744,0.03938462,0.009846155,0.0,0.0,0.0,0.0,0.04266667,0.04266667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.049230773,0.14769232,0.28225642,0.4004103,0.4266667,0.55794877,0.60061544,0.5907693,0.55794877,0.5546667,0.48246157,0.5349744,0.6662565,0.8172308,0.8992821,0.8960001,1.1257436,1.2340513,1.1618463,1.1552821,1.401436,1.3522053,1.2668719,1.2504616,1.2406155,1.1979488,1.079795,0.9517949,0.8402052,0.7220513,0.5907693,0.4594872,0.33476925,0.22646156,0.13784617,0.07876924,0.049230773,0.02297436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.02297436,0.09189744,0.1148718,0.16082053,0.21661541,0.15753847,0.055794876,0.02297436,0.02297436,0.029538464,0.02297436,0.0032820515,0.006564103,0.02297436,0.03938462,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.0,0.013128206,0.026256412,0.02297436,0.0032820515,0.0,0.0032820515,0.013128206,0.01969231,0.02297436,0.02297436,0.03938462,0.029538464,0.01969231,0.032820515,0.0951795,0.19692309,0.4266667,0.574359,0.5907693,0.574359,0.446359,0.2855385,0.16738462,0.09189744,0.0,0.006564103,0.01969231,0.049230773,0.101743594,0.17723078,0.27569234,0.21333335,0.17066668,0.69579494,2.6978464,2.2646155,2.4943593,3.2229745,4.7327185,7.768616,9.9282055,10.049642,8.795898,7.0925136,6.114462,7.5552826,11.185231,11.700514,8.477539,5.5630774,8.342975,9.701744,10.167795,10.397539,11.16554,10.620719,11.349334,11.651283,11.011283,10.082462,9.429334,10.509129,10.896411,9.737847,7.778462,14.04718,13.879796,13.528616,14.17518,11.910565,9.268514,14.424617,13.249642,6.1472826,8.024616,17.870771,13.607386,7.968821,6.0619493,5.362872,5.684513,6.091488,6.51159,6.9842057,7.6635904,5.6320004,3.9384618,2.9144619,2.4746668,2.1169233,3.2328207,10.5780525,13.420309,9.068309,2.865231,2.7208207,1.1651284,0.14769232,0.14112821,0.13784617,0.128,0.21333335,0.26256412,0.21661541,0.08861539,0.072205134,0.036102567,0.009846155,0.0,0.0,0.006564103,0.009846155,0.016410258,0.02297436,0.02297436,0.02297436,0.02297436,0.01969231,0.016410258,0.016410258,0.006564103,0.006564103,0.0032820515,0.0,0.0,0.0,0.098461546,0.24287182,0.38400003,0.4955898,0.58092314,0.4955898,0.4004103,0.32164106,0.14769232,0.029538464,0.0,0.0032820515,0.006564103,0.006564103,0.006564103,0.016410258,0.026256412,0.03938462,0.052512825,0.055794876,0.07876924,0.101743594,0.12143591,0.14769232,0.16738462,0.19364104,0.21661541,0.24287182,0.26912823,0.2855385,0.2986667,0.31507695,0.32820517,0.3314872,0.3511795,0.36102566,0.37743592,0.4004103,0.4201026,0.44307697,0.4660513,0.48902568,0.508718,0.54482055,0.58420515,0.61374366,0.636718,0.6498462,0.6498462,0.6465641,0.65312827,0.65641034,0.6498462,0.6301539,0.63343596,0.6432821,0.65312827,0.6662565,0.702359,0.72861546,0.77128214,0.8172308,0.8598975,0.8992821,0.9878975,1.083077,1.1815386,1.3029745,1.4572309,1.719795,2.0841026,2.605949,3.623385,5.7829747,0.6629744,0.65641034,0.6826667,1.0305642,1.8937438,3.3805132,1.148718,0.4004103,0.4201026,0.702359,0.94523084,0.6104616,0.48246157,0.38728207,0.26912823,0.190359,0.10502565,0.14112821,0.4594872,0.92553854,1.1027694,0.5021539,0.256,0.43323082,1.723077,5.4514875,5.0510774,4.315898,3.876103,3.4625645,1.8773335,0.62030774,0.21661541,0.4955898,1.0699488,1.3554872,0.827077,0.33476925,0.059076928,0.006564103,0.0,0.02297436,0.03938462,0.052512825,0.072205134,0.108307704,0.049230773,0.052512825,0.04266667,0.013128206,0.02297436,0.0032820515,0.0,0.0032820515,0.10502565,0.4955898,0.48246157,0.4266667,0.4135385,0.5349744,0.90912825,1.0272821,1.5524104,1.8248206,1.8248206,2.1825643,2.809436,2.6912823,2.2088206,1.7427694,1.6836925,1.7591796,1.8773335,2.044718,2.1169233,1.7887181,2.0250258,2.8225644,3.2722054,3.1343591,2.8356924,2.6026669,2.8127182,3.3969233,3.9942567,3.9318976,3.6069746,3.2820516,3.2886157,3.3411283,2.546872,0.8205129,0.190359,0.08205129,0.11158975,0.08533334,0.036102567,0.02297436,0.013128206,0.0,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.006564103,0.0032820515,0.009846155,0.03938462,0.08205129,0.21661541,0.36102566,0.26912823,0.45620516,0.60061544,0.6432821,0.56451285,0.39712822,0.36102566,0.36430773,0.2986667,0.15753847,0.032820515,0.009846155,0.0,0.0,0.0,0.0,0.006564103,0.029538464,0.068923086,0.11158975,0.15097436,0.07548718,0.02297436,0.016410258,0.032820515,0.0,0.0,0.08861539,0.08861539,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.0,0.0,0.0,0.0,0.0,0.009846155,0.013128206,0.01969231,0.02297436,0.013128206,0.02297436,0.03938462,0.059076928,0.08205129,0.12143591,0.12471796,0.13128206,0.13784617,0.14441027,0.13456412,0.12471796,0.1148718,0.108307704,0.108307704,0.108307704,0.108307704,0.101743594,0.07876924,0.059076928,0.098461546,0.08861539,0.032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.006564103,0.0,0.0,0.0,0.0,0.0,0.009846155,0.032820515,0.18379489,0.25271797,0.34789747,0.4201026,0.28225642,0.13784617,0.059076928,0.029538464,0.02297436,0.02297436,0.006564103,0.0032820515,0.0032820515,0.0032820515,0.02297436,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.016410258,0.013128206,0.009846155,0.02297436,0.049230773,0.059076928,0.049230773,0.049230773,0.06564103,0.049230773,0.02297436,0.02297436,0.098461546,0.15097436,0.34133336,0.5349744,0.67282057,0.7581539,0.5349744,0.27897438,0.14112821,0.108307704,0.01969231,0.016410258,0.03938462,0.036102567,0.029538464,0.1148718,0.30851284,0.23302566,0.15753847,0.17394873,0.19692309,0.30194873,1.1913847,1.972513,2.7011285,4.342154,9.248821,10.443488,8.595693,6.3277955,8.205129,9.96759,10.312206,9.639385,8.152616,5.85518,6.616616,7.9917955,9.399796,10.315488,10.262975,11.611898,12.806565,12.173129,10.28595,9.957745,11.250873,9.472001,8.464411,9.212719,9.813334,12.071385,15.067899,18.697847,20.680206,16.587488,9.95118,17.56882,16.984617,8.388924,14.6182575,16.000002,11.369026,8.03118,7.1483083,3.757949,2.92759,2.7700515,3.6594875,5.0116925,5.3136415,6.8529234,6.5247183,5.218462,3.6857438,2.5271797,1.270154,8.644924,14.693745,13.08554,1.148718,0.72861546,0.48574364,0.28225642,0.118153855,0.098461546,0.068923086,0.032820515,0.02297436,0.055794876,0.12471796,0.14112821,0.08205129,0.04594872,0.052512825,0.029538464,0.009846155,0.0,0.006564103,0.013128206,0.013128206,0.013128206,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.009846155,0.0032820515,0.0032820515,0.0032820515,0.0032820515,0.0032820515,0.0032820515,0.0032820515,0.0032820515,0.0032820515,0.0032820515,0.0,0.0032820515,0.0032820515,0.0032820515,0.009846155,0.01969231,0.01969231,0.01969231,0.029538464,0.03938462,0.052512825,0.06235898,0.07548718,0.08533334,0.0951795,0.108307704,0.13128206,0.128,0.14441027,0.16082053,0.17394873,0.19692309,0.21989745,0.23630771,0.25271797,0.27241027,0.28225642,0.29538465,0.30194873,0.3117949,0.3314872,0.3446154,0.38400003,0.4135385,0.4397949,0.4660513,0.49887183,0.5349744,0.571077,0.60389745,0.6235898,0.6301539,0.62030774,0.6235898,0.6235898,0.6104616,0.5874872,0.571077,0.574359,0.57764107,0.57764107,0.5874872,0.5973334,0.6170257,0.6235898,0.636718,0.69251287,0.8172308,0.88943595,0.9288206,0.97805136,1.1126155,1.2898463,1.4539489,1.9462565,3.1507695,5.4875903,0.5021539,0.4660513,0.3117949,0.8008206,1.9790771,3.1737437,1.9790771,1.0929232,1.0436924,1.654154,2.044718,1.5819489,1.401436,1.273436,1.0075898,0.45620516,0.23958977,0.45620516,1.4408206,2.7864618,3.370667,1.5885129,1.0075898,1.4703591,3.2886157,7.2336416,3.2886157,3.511795,6.521436,9.15036,6.452513,2.412308,0.7450257,0.98133343,2.038154,2.1956925,1.6114873,0.86974365,0.30194873,0.036102567,0.0,0.108307704,0.15425642,0.13128206,0.068923086,0.04594872,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.01969231,0.07876924,0.21333335,0.4955898,0.56451285,0.6629744,0.6892308,0.21333335,0.45620516,0.8763078,1.1388719,1.2668719,1.6311796,2.3269746,2.1924105,2.0676925,2.2219489,2.3204105,1.5261539,1.2373334,1.339077,1.5556924,1.4342566,1.6902566,2.477949,3.6791797,5.0576415,6.23918,6.6428723,6.8004107,6.872616,6.7610264,6.1046157,5.8945646,5.431795,5.2414365,5.733744,7.1876926,2.5107694,0.7122052,0.19364104,0.036102567,0.0,0.0,0.06564103,0.06564103,0.0032820515,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01969231,0.036102567,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.04594872,0.0951795,0.068923086,0.06564103,0.108307704,0.18379489,0.14769232,0.108307704,0.12143591,0.20020515,0.33476925,0.41025645,0.3708718,0.26256412,0.13128206,0.04594872,0.02297436,0.006564103,0.0,0.0,0.0,0.036102567,0.15425642,0.26584616,0.25928208,0.016410258,0.026256412,0.013128206,0.08533334,0.17066668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.029538464,0.006564103,0.0,0.0,0.0,0.0,0.0,0.009846155,0.059076928,0.098461546,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.02297436,0.04594872,0.16738462,0.318359,0.36758977,0.29538465,0.19692309,0.19692309,0.13456412,0.055794876,0.0,0.0,0.013128206,0.016410258,0.009846155,0.009846155,0.04594872,0.02297436,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.016410258,0.02297436,0.04594872,0.068923086,0.11158975,0.13128206,0.12143591,0.12143591,0.108307704,0.068923086,0.032820515,0.049230773,0.18379489,0.15753847,0.5907693,0.8795898,0.892718,0.97805136,0.69579494,0.24943592,0.06564103,0.15097436,0.09189744,0.07876924,0.049230773,0.036102567,0.055794876,0.09189744,0.128,0.13784617,0.15097436,0.17394873,0.19692309,0.23630771,0.26256412,0.4955898,1.0338463,1.8773335,3.6463592,4.667077,5.47118,7.6701546,13.932309,15.0777445,12.025436,10.614155,10.84718,6.882462,5.7468724,5.5630774,7.387898,9.849437,9.140513,10.568206,13.331694,13.223386,9.810052,6.4557953,8.467693,7.9819493,6.8430777,7.958975,15.320617,14.244103,9.813334,11.32636,18.710976,22.505028,10.761847,10.118565,12.3766165,13.115078,11.687386,13.909334,13.98154,16.738462,17.64759,2.793026,2.0217438,1.9331284,3.8498464,6.2523084,4.775385,11.113027,8.612103,4.522667,2.5764105,2.989949,1.5392822,1.2471796,4.3552823,7.680001,2.6256413,1.3193847,1.2012309,0.8795898,0.17066668,0.12143591,0.072205134,0.032820515,0.009846155,0.0032820515,0.016410258,0.052512825,0.098461546,0.190359,0.26256412,0.15097436,0.04266667,0.006564103,0.006564103,0.013128206,0.0,0.013128206,0.016410258,0.02297436,0.026256412,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.02297436,0.01969231,0.0032820515,0.016410258,0.016410258,0.02297436,0.029538464,0.029538464,0.029538464,0.04266667,0.04594872,0.052512825,0.06235898,0.06235898,0.08533334,0.09189744,0.09189744,0.0951795,0.108307704,0.0951795,0.101743594,0.108307704,0.11158975,0.13784617,0.15097436,0.16082053,0.17394873,0.18707694,0.19692309,0.2100513,0.2231795,0.23630771,0.24615386,0.25928208,0.30851284,0.34789747,0.37743592,0.40369233,0.4266667,0.45292312,0.48574364,0.5218462,0.5546667,0.58092314,0.5907693,0.5874872,0.58092314,0.574359,0.5481026,0.52512825,0.508718,0.5021539,0.5021539,0.5021539,0.5021539,0.5021539,0.5218462,0.55794877,0.5940513,0.6301539,0.6235898,0.6465641,0.761436,0.9911796,1.1388719,1.4145643,2.681436,5.034667,7.781744,0.101743594,0.09189744,0.15097436,0.5021539,0.9288206,0.76800007,0.57764107,0.5677949,0.88615394,1.5753847,2.5829747,3.620103,3.114667,2.858667,3.0884104,2.4582565,1.1749744,0.60061544,0.9156924,1.7033848,1.9561027,0.827077,0.76800007,2.0578463,4.164923,5.756718,2.8488207,1.7755898,3.4888208,7.706257,12.947693,8.694155,4.273231,1.6705642,1.5031796,3.0391798,4.397949,4.8804107,3.6496413,1.463795,0.6826667,0.6662565,0.7253334,0.61374366,0.50543594,0.99774367,1.7624617,1.3095386,0.64000005,0.28225642,0.29210258,0.83035904,1.3456411,1.7427694,1.8510771,1.4112822,0.6268718,0.32164106,0.21333335,0.15425642,0.1148718,0.21333335,0.45620516,0.86646163,1.1618463,0.764718,0.8467693,0.9944616,1.2209232,1.5458462,2.0151796,1.591795,2.1202054,2.3893335,2.038154,1.5556924,1.3161026,1.3095386,2.0939488,3.3444104,3.8859491,4.2502565,4.900103,5.7829747,6.8299494,7.958975,8.123077,7.1581545,5.874872,4.785231,4.0992823,2.1956925,1.0010257,0.36102566,0.0951795,0.0,0.0,0.026256412,0.08205129,0.13456412,0.13784617,0.026256412,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.032820515,0.06235898,0.75487185,0.37743592,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.016410258,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.009846155,0.01969231,0.013128206,0.013128206,0.02297436,0.036102567,0.049230773,0.11158975,0.10502565,0.049230773,0.10502565,0.22646156,0.3052308,0.29210258,0.19364104,0.068923086,0.016410258,0.009846155,0.016410258,0.032820515,0.072205134,0.14769232,0.101743594,0.08861539,0.12143591,0.052512825,0.036102567,0.04266667,0.04594872,0.032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.029538464,0.06564103,0.036102567,0.026256412,0.009846155,0.0,0.0,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.01969231,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.013128206,0.01969231,0.016410258,0.02297436,0.12471796,0.21661541,0.24287182,0.20676924,0.19692309,0.22646156,0.16410258,0.07876924,0.029538464,0.049230773,0.02297436,0.016410258,0.013128206,0.013128206,0.02297436,0.016410258,0.01969231,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.0032820515,0.0032820515,0.006564103,0.01969231,0.032820515,0.059076928,0.08533334,0.10502565,0.11158975,0.12143591,0.14769232,0.14769232,0.108307704,0.06235898,0.098461546,0.18051283,0.6629744,1.4178462,1.9692309,1.4900514,0.9353847,0.5316923,0.33805132,0.256,0.01969231,0.055794876,0.052512825,0.052512825,0.068923086,0.06564103,0.1148718,0.14769232,0.17066668,0.17723078,0.17394873,0.21989745,0.2297436,0.28882053,0.5349744,1.1323078,1.6049232,1.9889232,2.5993848,3.69559,5.4843082,5.861744,4.9854364,5.2545643,6.6461544,6.7117953,7.1876926,7.860513,9.672206,12.406155,14.706873,11.260718,9.921641,10.94236,12.993642,13.180719,9.472001,9.344001,9.035488,8.625232,12.012309,16.006565,13.732103,11.72677,11.812103,11.1064625,10.581334,13.377642,14.41477,12.800001,11.808822,14.578873,11.0145645,8.333129,7.453539,2.986667,1.9167181,3.7251284,8.1755905,11.096616,4.384821,7.3714876,7.381334,5.7632823,4.273231,5.077334,6.055385,4.4996924,11.503591,21.431797,11.913847,4.338872,1.3161026,0.4201026,0.190359,0.12143591,0.08205129,0.08861539,0.06564103,0.009846155,0.0032820515,0.009846155,0.026256412,0.068923086,0.13128206,0.17723078,0.15425642,0.07548718,0.01969231,0.013128206,0.013128206,0.013128206,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.029538464,0.049230773,0.03938462,0.029538464,0.036102567,0.04594872,0.049230773,0.03938462,0.049230773,0.052512825,0.049230773,0.03938462,0.052512825,0.04266667,0.032820515,0.036102567,0.04266667,0.04266667,0.04594872,0.052512825,0.06564103,0.072205134,0.06235898,0.07548718,0.07876924,0.07876924,0.08205129,0.0951795,0.09189744,0.08533334,0.09189744,0.11158975,0.12471796,0.128,0.13784617,0.14441027,0.15097436,0.16082053,0.17394873,0.18707694,0.20348719,0.22646156,0.24615386,0.26584616,0.29210258,0.318359,0.34133336,0.36758977,0.39056414,0.41682056,0.44964105,0.48574364,0.51856416,0.5415385,0.54482055,0.53825647,0.5284103,0.52512825,0.49887183,0.47917953,0.46276927,0.45620516,0.45620516,0.45620516,0.46933338,0.49230772,0.5152821,0.5218462,0.53825647,0.57764107,0.65312827,0.77456415,0.9189744,0.99774367,1.3718976,2.546872,4.332308,5.8289237,0.036102567,0.108307704,0.33805132,0.702359,0.92553854,0.46933338,0.25271797,0.21989745,0.35774362,0.69907695,1.3259488,2.7109745,3.5774362,4.325744,5.0642056,5.5958977,4.345436,2.4582565,1.1946667,0.8369231,0.67610264,0.41682056,0.7515898,2.9078977,6.7610264,10.824206,5.802667,2.4976413,1.8838975,3.9023592,7.466667,6.409847,4.594872,3.4822567,3.7415388,5.2644105,6.7938466,8.201847,6.0816417,1.5786668,0.37743592,0.446359,0.4660513,0.6301539,0.9517949,1.2373334,2.1333334,1.6082052,0.94523084,0.7253334,0.8336411,0.8960001,1.1782565,1.4375386,1.4900514,1.2406155,0.5940513,0.33476925,0.29538465,0.44964105,0.88943595,0.9485129,0.77456415,0.8008206,0.98133343,0.76800007,0.61374366,0.8205129,1.0765129,1.2865642,1.5622566,1.2996924,1.8445129,2.0841026,1.7624617,1.4966155,1.1290257,1.0765129,1.7099489,2.6223593,2.6190772,2.7963078,2.7798977,3.3411283,4.417641,5.1265645,5.0904617,4.713026,4.2896414,3.9778464,3.8104618,3.2328207,2.422154,1.5360001,0.7056411,0.055794876,0.19364104,0.32820517,0.4660513,0.6104616,0.761436,0.39384618,0.18051283,0.101743594,0.16738462,0.4397949,0.6301539,0.3314872,0.06564103,0.016410258,0.03938462,0.37743592,0.190359,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.01969231,0.026256412,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.04594872,0.03938462,0.0032820515,0.01969231,0.072205134,0.1148718,0.13456412,0.13128206,0.11158975,0.0951795,0.06235898,0.032820515,0.026256412,0.04594872,0.07876924,0.049230773,0.055794876,0.08861539,0.032820515,0.016410258,0.01969231,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.032820515,0.01969231,0.013128206,0.03938462,0.055794876,0.04266667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.029538464,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0,0.013128206,0.036102567,0.03938462,0.01969231,0.006564103,0.08205129,0.17723078,0.22646156,0.23302566,0.28225642,0.27241027,0.20348719,0.118153855,0.059076928,0.06235898,0.06235898,0.06564103,0.07548718,0.07548718,0.052512825,0.029538464,0.02297436,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.009846155,0.013128206,0.01969231,0.026256412,0.029538464,0.03938462,0.06235898,0.08205129,0.10502565,0.14112821,0.21989745,0.26256412,0.20676924,0.09189744,0.06564103,0.15425642,1.1552821,2.6256413,3.6693337,2.934154,2.356513,1.7657437,1.079795,0.40697438,0.04594872,0.049230773,0.036102567,0.036102567,0.059076928,0.098461546,0.17723078,0.17723078,0.16410258,0.15753847,0.15753847,0.18707694,0.18379489,0.24943592,0.4004103,0.571077,0.7187693,0.9747693,1.3817437,2.2416413,4.1222568,3.4921029,4.348718,6.3343596,8.090257,7.253334,8.960001,9.737847,10.361437,11.244308,12.425847,10.545232,8.592411,8.605539,10.354873,11.319796,10.308924,11.9860525,13.193847,12.62277,10.781539,12.199386,14.303181,13.000206,9.409642,9.892103,11.992617,13.873232,12.514462,9.55077,11.273847,14.221129,10.584617,6.816821,5.097026,3.31159,1.9232821,3.9122055,7.1647186,8.805744,5.1954875,5.395693,5.4514875,6.091488,7.2303596,7.972103,10.473026,9.088,13.961847,22.833233,21.018257,8.346257,2.3401027,0.35446155,0.190359,0.0951795,0.08861539,0.12471796,0.12143591,0.06564103,0.009846155,0.016410258,0.02297436,0.029538464,0.049230773,0.08205129,0.14112821,0.108307704,0.08205129,0.08205129,0.06235898,0.032820515,0.013128206,0.009846155,0.016410258,0.016410258,0.016410258,0.01969231,0.036102567,0.052512825,0.055794876,0.049230773,0.052512825,0.06235898,0.068923086,0.06564103,0.07548718,0.07876924,0.07548718,0.07548718,0.08861539,0.08205129,0.07876924,0.07876924,0.08533334,0.09189744,0.098461546,0.10502565,0.11158975,0.12143591,0.1148718,0.12143591,0.13456412,0.13456412,0.12471796,0.128,0.128,0.12471796,0.12471796,0.128,0.14112821,0.14112821,0.14441027,0.14769232,0.15097436,0.16082053,0.16738462,0.17723078,0.190359,0.21333335,0.25271797,0.27897438,0.29538465,0.3117949,0.33805132,0.37743592,0.40369233,0.4266667,0.44964105,0.47261542,0.5021539,0.5284103,0.53825647,0.5415385,0.5349744,0.5284103,0.5021539,0.47917953,0.45292312,0.42994875,0.4135385,0.42338464,0.42994875,0.4397949,0.45292312,0.47589746,0.51856416,0.56123084,0.6170257,0.69251287,0.80738467,1.0371283,1.595077,2.5271797,3.446154,3.5478978,0.10502565,0.34789747,0.446359,0.60061544,0.8992821,1.3193847,1.5360001,1.0962052,0.636718,0.47589746,0.60389745,1.5819489,2.7142565,3.6562054,4.5029745,5.792821,5.8912826,5.431795,4.161641,2.281026,0.45292312,0.60389745,1.4834872,4.972308,9.527796,10.177642,7.6274877,3.3969233,0.9353847,0.99774367,1.6640002,2.4024618,2.993231,3.5446157,4.06318,4.453744,4.9526157,6.088206,4.630975,1.3193847,0.8730257,0.7056411,0.39712822,0.41025645,0.71548724,0.77128214,1.3193847,1.086359,0.94523084,1.1684103,1.4080001,1.1716924,0.81394875,0.72861546,0.9124103,0.9616411,0.5481026,0.4266667,0.4266667,0.53825647,0.92553854,0.9419488,0.85005134,0.88287187,0.9944616,0.86646163,1.1191796,1.5885129,1.8248206,1.7263591,1.5556924,1.2012309,1.2668719,1.3095386,1.2471796,1.3915899,1.4145643,1.3915899,1.7263591,2.2547693,2.2219489,2.3072822,1.723077,2.166154,3.4002054,3.239385,2.7831798,3.3312824,3.6562054,3.3509746,2.8225644,2.6354873,2.2350771,1.591795,0.8402052,0.28225642,0.571077,0.6892308,0.74830776,0.8467693,1.0666667,0.6892308,0.46276927,0.40697438,0.53825647,0.8730257,1.1224617,0.5874872,0.14769232,0.08205129,0.08861539,0.052512825,0.03938462,0.02297436,0.0,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.01969231,0.026256412,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01969231,0.059076928,0.101743594,0.09189744,0.059076928,0.029538464,0.016410258,0.02297436,0.013128206,0.013128206,0.036102567,0.055794876,0.02297436,0.0032820515,0.0032820515,0.01969231,0.04266667,0.072205134,0.068923086,0.029538464,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.032820515,0.055794876,0.04266667,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0,0.006564103,0.006564103,0.0,0.0,0.08861539,0.059076928,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01969231,0.04266667,0.04594872,0.029538464,0.029538464,0.072205134,0.16082053,0.21333335,0.2297436,0.26912823,0.30851284,0.29210258,0.21333335,0.10502565,0.055794876,0.08533334,0.09189744,0.08533334,0.068923086,0.052512825,0.029538464,0.02297436,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016410258,0.02297436,0.026256412,0.029538464,0.029538464,0.036102567,0.049230773,0.068923086,0.10502565,0.15097436,0.26256412,0.34133336,0.29210258,0.14769232,0.055794876,0.14441027,1.2898463,2.7798977,3.7316926,3.0752823,3.0982566,2.5009232,1.463795,0.4266667,0.06564103,0.03938462,0.02297436,0.016410258,0.06235898,0.23958977,0.32164106,0.24615386,0.15753847,0.12471796,0.12143591,0.12471796,0.12471796,0.190359,0.30194873,0.3249231,0.51856416,0.72861546,0.92225647,1.4572309,3.0916924,2.6715899,4.926359,7.6307697,8.953437,7.4371285,10.482873,12.166565,11.720206,10.131693,10.138257,9.796924,8.569437,7.9852314,8.52677,9.659078,9.885539,10.515693,11.506873,12.015591,10.377847,8.841846,11.723488,12.534155,10.8767185,12.4685135,12.747488,14.322873,12.517745,8.395488,8.769642,12.370052,12.137027,9.984001,7.4469748,5.684513,2.7766156,3.2196925,5.4875903,7.4929237,6.567385,5.106872,5.280821,8.086975,12.107488,13.525334,15.451899,13.436719,12.744206,15.202463,19.203283,9.590155,3.4034874,0.65969235,0.29210258,0.16738462,0.101743594,0.118153855,0.14441027,0.13128206,0.026256412,0.036102567,0.06564103,0.059076928,0.02297436,0.02297436,0.0951795,0.10502565,0.1148718,0.13784617,0.14769232,0.098461546,0.049230773,0.02297436,0.02297436,0.026256412,0.026256412,0.036102567,0.04594872,0.055794876,0.072205134,0.072205134,0.07548718,0.08533334,0.09189744,0.08861539,0.101743594,0.10502565,0.108307704,0.118153855,0.12471796,0.13456412,0.13456412,0.13456412,0.14112821,0.15097436,0.16410258,0.17394873,0.18707694,0.19692309,0.19692309,0.190359,0.20348719,0.2100513,0.20020515,0.19692309,0.190359,0.190359,0.18379489,0.17723078,0.190359,0.18379489,0.17723078,0.17394873,0.17723078,0.17394873,0.18379489,0.20020515,0.2297436,0.30851284,0.508718,0.6301539,0.69251287,0.61374366,0.45620516,0.4266667,0.47261542,0.55794877,0.6662565,0.7515898,0.761436,0.827077,0.8467693,0.8369231,0.81394875,0.8041026,0.7384616,0.6465641,0.5349744,0.43651286,0.39712822,0.40369233,0.40697438,0.4135385,0.43323082,0.46933338,0.5218462,0.54482055,0.57764107,0.6826667,0.9419488,1.3883078,1.9429746,2.4648206,2.7044106,2.3269746,0.318359,0.8992821,0.636718,0.28225642,0.49230772,1.8313848,2.7700515,2.225231,1.8674873,2.038154,1.7526156,1.5688206,1.6049232,1.6869745,1.972513,2.9604106,4.5587697,7.131898,7.6635904,5.3891287,1.782154,1.7591796,2.8914874,6.6395903,9.580308,3.4100516,6.2096415,3.4855387,1.148718,1.0502565,0.9616411,1.1618463,2.162872,3.170462,3.5380516,2.7798977,1.8740515,1.463795,1.7001027,2.3958976,3.0260515,2.3433847,1.6640002,0.9321026,0.28882053,0.07548718,0.13456412,0.26584616,0.6465641,1.1913847,1.5556924,1.5360001,0.7056411,0.3708718,0.7450257,0.92553854,0.55794877,0.49230772,0.42338464,0.33476925,0.50543594,0.61374366,0.9714873,1.4080001,1.5425643,0.77456415,1.8806155,2.8422565,2.917744,2.2022567,1.6246156,1.1782565,0.99774367,1.0043077,1.1323078,1.3095386,1.7558975,1.6935385,1.6771283,1.8871796,2.1169233,2.2383592,1.7920002,2.5665643,4.1485133,3.9351797,2.8980515,3.5971284,3.764513,2.6912823,1.270154,1.1257436,0.892718,0.6170257,0.4266667,0.5481026,0.8336411,0.86974365,0.79425645,0.7450257,0.8566154,0.7417436,0.69251287,0.7318975,0.8369231,0.9353847,1.0502565,0.57764107,0.24287182,0.23958977,0.24287182,0.14769232,0.118153855,0.072205134,0.013128206,0.02297436,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.04266667,0.08205129,0.08205129,0.032820515,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.036102567,0.03938462,0.006564103,0.0,0.0032820515,0.013128206,0.02297436,0.0032820515,0.0032820515,0.013128206,0.032820515,0.052512825,0.01969231,0.072205134,0.118153855,0.14441027,0.20020515,0.18707694,0.08533334,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.006564103,0.0,0.0,0.0,0.026256412,0.029538464,0.0032820515,0.0,0.118153855,0.09189744,0.036102567,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.006564103,0.0,0.0,0.04594872,0.02297436,0.0,0.0,0.0,0.0,0.0,0.006564103,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.029538464,0.049230773,0.06564103,0.108307704,0.10502565,0.14112821,0.16738462,0.16738462,0.15425642,0.27897438,0.3249231,0.26256412,0.13128206,0.052512825,0.08205129,0.08533334,0.055794876,0.01969231,0.01969231,0.013128206,0.01969231,0.016410258,0.006564103,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.03938462,0.04594872,0.029538464,0.02297436,0.032820515,0.036102567,0.04266667,0.049230773,0.06564103,0.10502565,0.15097436,0.25928208,0.35774362,0.34789747,0.21989745,0.06564103,0.14112821,0.83035904,1.5819489,1.9692309,1.6869745,2.5042052,2.1891284,1.2800001,0.3708718,0.08533334,0.026256412,0.013128206,0.006564103,0.06564103,0.33476925,0.39056414,0.26256412,0.13456412,0.08861539,0.068923086,0.06235898,0.068923086,0.09189744,0.15097436,0.28882053,0.5218462,0.6892308,0.7811283,0.81066674,0.81394875,1.3751796,3.9942567,6.1768208,6.944821,6.8463597,11.178667,14.87754,14.503386,11.0145645,9.747693,9.626257,9.156924,8.946873,9.485129,11.155693,9.153642,6.196513,4.9952826,6.377026,9.268514,7.604513,7.8736415,9.747693,11.96636,12.340514,10.643693,13.00677,12.721231,8.677744,5.3694363,8.960001,12.822975,13.459693,10.8537445,8.474257,4.0467696,2.349949,4.325744,7.890052,7.9491286,7.13518,8.070564,11.946668,17.122463,19.140924,18.73395,16.006565,10.955488,6.5706673,8.841846,8.572719,5.4613338,2.3171284,0.57764107,0.29210258,0.13128206,0.09189744,0.13128206,0.16082053,0.055794876,0.055794876,0.108307704,0.10502565,0.03938462,0.03938462,0.068923086,0.08205129,0.101743594,0.15425642,0.2855385,0.3314872,0.2297436,0.11158975,0.049230773,0.04594872,0.04594872,0.055794876,0.06235898,0.068923086,0.0951795,0.098461546,0.10502565,0.1148718,0.118153855,0.108307704,0.12143591,0.12471796,0.13456412,0.15097436,0.15097436,0.17066668,0.17066668,0.17394873,0.190359,0.20348719,0.21989745,0.23630771,0.256,0.26584616,0.26584616,0.256,0.25928208,0.26584616,0.27241027,0.26256412,0.24943592,0.24943592,0.24615386,0.23958977,0.24943592,0.23958977,0.21989745,0.21333335,0.21661541,0.19692309,0.23958977,0.40369233,0.574359,0.77128214,1.1585642,1.3522053,1.4408206,1.214359,0.7844103,0.58420515,0.8369231,1.204513,1.595077,1.9068719,2.03159,2.2678976,2.353231,2.3401027,2.28759,2.2744617,2.1530259,1.8904617,1.4473847,0.90584624,0.46276927,0.4201026,0.41025645,0.4266667,0.4594872,0.4955898,0.5316923,0.5481026,0.636718,0.86974365,1.3259488,1.8149745,2.1956925,2.4976413,2.7536411,2.9997952,0.9156924,2.1103592,1.6508719,0.7122052,0.049230773,0.0,0.11158975,0.63343596,3.1638978,6.193231,5.097026,2.6190772,2.484513,2.1103592,1.0568206,1.0075898,1.7263591,3.3542566,5.504,6.774154,4.7589746,4.345436,4.2962055,3.754667,2.7011285,1.9692309,1.8576412,3.058872,4.322462,4.903385,4.562052,4.8311796,6.2162056,7.857231,9.005949,9.019077,7.4174366,4.923077,5.080616,7.2861543,6.774154,5.8945646,5.546667,3.9351797,1.332513,0.07548718,0.026256412,0.016410258,0.016410258,0.128,0.58092314,0.77456415,0.45620516,0.23302566,0.32820517,0.5940513,0.62030774,0.49887183,0.4135385,0.6892308,1.8018463,2.5337439,2.6880002,3.0424619,3.0194874,0.702359,2.4713848,3.7382567,3.0916924,1.1224617,0.4266667,0.4397949,1.3850257,2.15959,2.1530259,1.2373334,1.0272821,1.2340513,1.4276924,1.4473847,1.3718976,1.4834872,1.8412309,2.5107694,3.5216413,4.850872,2.8258464,1.4506668,1.0043077,1.5491283,2.930872,3.1376412,2.0644104,0.92225647,0.36758977,0.48902568,0.40369233,0.67282057,0.80738467,0.6859488,0.56451285,0.61374366,0.6432821,0.60061544,0.48574364,0.3511795,0.32820517,0.32164106,0.3511795,0.40369233,0.4266667,0.23302566,0.19364104,0.14441027,0.06235898,0.06235898,0.049230773,0.01969231,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.21989745,0.41025645,0.4135385,0.16738462,0.032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01969231,0.03938462,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.01969231,0.072205134,0.13784617,0.13784617,0.07548718,0.318359,0.40369233,0.27569234,0.27569234,0.24943592,0.12471796,0.026256412,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06564103,0.068923086,0.013128206,0.0,0.013128206,0.016410258,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.026256412,0.026256412,0.0,0.0,0.23302566,0.1148718,0.0,0.0,0.0,0.0,0.0,0.029538464,0.06235898,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01969231,0.07876924,0.16738462,0.2297436,0.16738462,0.1148718,0.10502565,0.118153855,0.108307704,0.0951795,0.055794876,0.029538464,0.03938462,0.07548718,0.07548718,0.0951795,0.101743594,0.07876924,0.029538464,0.006564103,0.0,0.013128206,0.029538464,0.029538464,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.06564103,0.19692309,0.12471796,0.06235898,0.029538464,0.036102567,0.06235898,0.049230773,0.055794876,0.07876924,0.1148718,0.15097436,0.24943592,0.33805132,0.35774362,0.28225642,0.13784617,0.07548718,0.07876924,0.128,0.25928208,0.56451285,1.1388719,1.1979488,0.9353847,0.5481026,0.24287182,0.049230773,0.0,0.0,0.006564103,0.029538464,0.06564103,0.049230773,0.029538464,0.032820515,0.04594872,0.059076928,0.06235898,0.072205134,0.0951795,0.108307704,0.23958977,0.60389745,0.96492314,1.1191796,0.8992821,0.86317956,1.3128207,2.2646155,3.7316926,5.720616,10.496001,16.338053,17.942976,14.007796,7.2336416,9.905231,9.7214365,9.472001,10.545232,12.924719,11.1294365,6.954667,3.511795,2.7864618,5.6320004,5.802667,6.311385,6.0849237,4.8114877,2.930872,3.5282054,3.761231,3.8695388,4.06318,4.5029745,4.342154,7.4896417,10.699488,11.158976,6.485334,4.1156926,1.9790771,1.3489232,3.3345644,8.864821,12.796719,13.768207,15.491283,18.018463,17.762463,15.136822,15.27795,13.801026,9.7214365,5.4482055,10.06277,11.296822,7.322257,1.0732309,0.24287182,0.17066668,0.12471796,0.101743594,0.09189744,0.09189744,0.09189744,0.072205134,0.06564103,0.07548718,0.07548718,0.07548718,0.07548718,0.068923086,0.15097436,0.51856416,0.9353847,0.73517954,0.3708718,0.108307704,0.04594872,0.04594872,0.055794876,0.06564103,0.08205129,0.108307704,0.118153855,0.12143591,0.1148718,0.108307704,0.12143591,0.13456412,0.128,0.128,0.14112821,0.15097436,0.15097436,0.16082053,0.18051283,0.20348719,0.2297436,0.25271797,0.25928208,0.27241027,0.28882053,0.28882053,0.28882053,0.28225642,0.27569234,0.27569234,0.27569234,0.26256412,0.26912823,0.27569234,0.27569234,0.27569234,0.27569234,0.256,0.24287182,0.24615386,0.25928208,0.3708718,1.0929232,1.719795,2.0250258,2.2580514,2.2449234,2.1136413,1.8346668,1.4375386,1.020718,1.9987694,3.1113849,4.1124105,4.9132314,5.586052,6.232616,6.557539,6.629744,6.5706673,6.5444107,6.436103,5.904411,4.6178465,2.6978464,0.7318975,0.512,0.45620516,0.46933338,0.4955898,0.51856416,0.5546667,0.6826667,0.9714873,1.3653334,1.6935385,1.7427694,2.0578463,3.0523078,4.562052,5.8453336,0.19692309,0.5907693,0.7778462,1.0732309,1.595077,2.2580514,1.4112822,0.7187693,1.079795,2.0939488,2.0676925,1.0666667,1.4769232,2.540308,3.4888208,3.5446157,2.3827693,2.937436,3.4002054,3.5478978,4.7360005,3.2754874,4.9296412,5.211898,3.2525132,1.7985642,3.3969233,6.0324106,6.8955903,5.72718,4.818052,6.619898,8.513641,9.219283,8.356103,6.4557953,5.832206,4.325744,3.3641028,3.2853336,3.3575387,2.8291285,2.5042052,2.8455386,3.1343591,1.4572309,0.5973334,0.76800007,1.4441026,1.9265642,1.3718976,0.9714873,0.65969235,0.508718,0.5021539,0.54482055,0.69907695,0.8041026,0.8402052,1.0601027,1.9954873,2.8160002,3.6463592,4.1222568,3.5511796,0.90912825,1.2635899,2.1333334,2.674872,2.5731285,2.0151796,1.9692309,1.5721027,1.7526156,2.297436,1.8707694,1.4375386,2.481231,3.8465643,4.8377438,5.1954875,3.3903592,2.0808206,1.6640002,1.9626669,2.228513,1.6082052,1.8051283,2.5173335,3.1638978,2.8914874,2.1825643,1.5097437,1.1388719,1.3292309,2.3204105,0.69251287,0.37743592,0.4266667,0.39712822,0.380718,0.48902568,0.5415385,0.5021539,0.38728207,0.25271797,0.21989745,0.32820517,0.47917953,0.55794877,0.4135385,0.17066668,0.12471796,0.29210258,0.58420515,0.8172308,0.24943592,0.32164106,0.60389745,0.74830776,0.47589746,0.13456412,0.06235898,0.06235898,0.04266667,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.04266667,0.07876924,0.0951795,0.08205129,0.032820515,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.009846155,0.02297436,0.029538464,0.026256412,0.026256412,0.016410258,0.072205134,0.098461546,0.07876924,0.07876924,0.055794876,0.055794876,0.09189744,0.12143591,0.02297436,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.013128206,0.0032820515,0.0,0.0032820515,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.02297436,0.016410258,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.006564103,0.0,0.0,0.21333335,0.10502565,0.0,0.0,0.0,0.0,0.0,0.026256412,0.052512825,0.0,0.0,0.0,0.02297436,0.049230773,0.0,0.0,0.0,0.0,0.0,0.0,0.118153855,0.059076928,0.029538464,0.059076928,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.029538464,0.03938462,0.08205129,0.15097436,0.19364104,0.17066668,0.14441027,0.14441027,0.18707694,0.25271797,0.15425642,0.1148718,0.13784617,0.17066668,0.08861539,0.07876924,0.08861539,0.098461546,0.09189744,0.04266667,0.01969231,0.0032820515,0.0032820515,0.009846155,0.01969231,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.013128206,0.04594872,0.098461546,0.17394873,0.17723078,0.118153855,0.059076928,0.032820515,0.049230773,0.036102567,0.04266667,0.06564103,0.108307704,0.16410258,0.24287182,0.318359,0.3511795,0.3249231,0.24615386,0.18707694,0.13784617,0.108307704,0.13784617,0.29538465,0.49887183,0.6432821,0.65969235,0.5415385,0.35446155,0.09189744,0.016410258,0.006564103,0.0,0.006564103,0.02297436,0.02297436,0.013128206,0.006564103,0.009846155,0.029538464,0.072205134,0.108307704,0.13456412,0.15425642,0.21333335,0.4397949,0.8369231,1.2012309,1.1093334,1.0404103,1.0010257,1.2406155,2.1956925,4.4898467,9.028924,11.992617,12.35036,11.10318,11.30995,11.45436,11.648001,11.024411,10.256411,11.58236,13.223386,10.962052,7.282872,4.516103,4.8607183,4.8082056,6.931693,7.1483083,5.8912826,8.093539,6.738052,5.874872,8.293744,12.603078,13.22995,7.9917955,9.196308,12.166565,12.727796,7.194257,3.7120004,2.0250258,1.7493335,2.6223593,4.519385,4.5456414,5.0182567,7.5881033,10.528821,8.726975,10.128411,10.240001,9.344001,7.509334,4.604718,6.5739493,8.129642,7.3353853,4.594872,2.6617439,1.5425643,0.7220513,0.28882053,0.16738462,0.128,0.098461546,0.08205129,0.07876924,0.08205129,0.06564103,0.12143591,0.108307704,0.08205129,0.08861539,0.15097436,0.3052308,0.39056414,0.5481026,0.6695385,0.4135385,0.22646156,0.1148718,0.06564103,0.055794876,0.068923086,0.09189744,0.118153855,0.13784617,0.13784617,0.12143591,0.12471796,0.13128206,0.14112821,0.15097436,0.16410258,0.18379489,0.19692309,0.21333335,0.22646156,0.23958977,0.24615386,0.24615386,0.256,0.26584616,0.26584616,0.27569234,0.29210258,0.2986667,0.30194873,0.3117949,0.2986667,0.28225642,0.26912823,0.26584616,0.2855385,0.27569234,0.27241027,0.27241027,0.33805132,0.56451285,1.7394873,2.4057438,2.8488207,3.1606157,3.2361028,2.8225644,2.422154,2.3171284,2.5271797,2.8160002,3.5872824,4.637539,5.622154,6.416411,7.0990777,7.529026,7.709539,7.5913854,7.3091288,7.1548724,6.4032826,4.8804107,2.9243078,1.1651284,0.53825647,0.49230772,0.50543594,0.5415385,0.58092314,0.6170257,0.7318975,0.90912825,1.1454359,1.4309745,1.7427694,2.6912823,4.699898,7.13518,8.874667,8.310155,0.006564103,0.08533334,0.23958977,0.57764107,1.0601027,1.522872,1.4178462,1.2504616,1.148718,1.0469744,0.69907695,0.32820517,0.5284103,1.3883078,2.4188719,2.5337439,2.0118976,2.4713848,2.8882053,3.0818465,3.7316926,3.1671798,4.900103,4.9854364,3.1376412,2.7175386,4.0303593,7.6701546,7.6603084,4.023795,2.7667694,3.6857438,4.391385,4.4242053,3.9647183,3.817026,3.879385,3.4297438,2.917744,2.5009232,2.0644104,1.6968206,1.8674873,3.0391798,4.8147697,5.9470773,3.639795,2.2022567,1.7066668,1.6607181,1.024,0.5973334,0.39384618,0.28882053,0.22646156,0.21333335,0.2855385,0.37415388,0.44964105,0.7056411,1.5688206,1.9068719,2.3269746,2.422154,1.8609232,0.38400003,0.4004103,0.7089231,1.0404103,1.1749744,0.96492314,0.93866676,0.6498462,0.65969235,0.9353847,0.81066674,0.6170257,1.1158975,1.9265642,2.7602053,3.4297438,3.0293336,2.989949,2.7536411,2.2219489,1.7460514,1.7033848,1.6836925,2.1924105,2.9997952,3.121231,2.5928206,2.2350771,1.8871796,1.5589745,1.4506668,0.58420515,0.45292312,0.4955898,0.42994875,0.24287182,0.31507695,0.35446155,0.39384618,0.41025645,0.3117949,0.44307697,0.40697438,0.38728207,0.40369233,0.32820517,0.15425642,0.15097436,0.42994875,0.84348726,0.9878975,0.5218462,0.6268718,0.7581539,0.6892308,0.48574364,0.21333335,0.12471796,0.09189744,0.049230773,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.02297436,0.016410258,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.006564103,0.0,0.0,0.0,0.0032820515,0.009846155,0.013128206,0.013128206,0.0032820515,0.013128206,0.04266667,0.06235898,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016410258,0.016410258,0.0,0.0,0.006564103,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.009846155,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02297436,0.04266667,0.0,0.08205129,0.04266667,0.0,0.0,0.0,0.04266667,0.02297436,0.009846155,0.01969231,0.0,0.0,0.0,0.013128206,0.02297436,0.0,0.0,0.0,0.0,0.006564103,0.036102567,0.101743594,0.07548718,0.06564103,0.072205134,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.03938462,0.08205129,0.118153855,0.118153855,0.1148718,0.128,0.16410258,0.23302566,0.35446155,0.27569234,0.23630771,0.256,0.29210258,0.24615386,0.16082053,0.11158975,0.08205129,0.06235898,0.026256412,0.016410258,0.006564103,0.0,0.0,0.006564103,0.0,0.0,0.0,0.0032820515,0.009846155,0.03938462,0.036102567,0.052512825,0.098461546,0.16738462,0.17066668,0.108307704,0.049230773,0.036102567,0.055794876,0.04266667,0.03938462,0.04266667,0.07548718,0.15097436,0.23630771,0.2986667,0.34133336,0.36758977,0.35774362,0.30194873,0.2231795,0.14441027,0.108307704,0.15425642,0.23630771,0.28225642,0.30194873,0.27897438,0.18051283,0.059076928,0.02297436,0.009846155,0.0,0.0,0.013128206,0.016410258,0.016410258,0.01969231,0.01969231,0.01969231,0.08205129,0.15097436,0.20020515,0.23302566,0.3052308,0.5513847,0.9714873,1.3686155,1.3522053,1.404718,1.3686155,1.3522053,1.9364104,4.1714873,6.925129,10.026668,11.21477,10.824206,11.815386,12.265027,12.678565,11.69395,9.511385,7.9228725,9.15036,8.320001,6.6494365,5.9667697,8.687591,5.5597954,6.196513,6.2194877,5.648411,8.907488,10.896411,11.588924,12.42913,14.106257,16.564514,13.02318,10.331899,10.994873,12.393026,6.774154,4.092718,4.2272825,4.972308,5.8453336,8.103385,7.4436927,4.827898,3.7054362,4.2436924,3.3017437,4.089436,4.2962055,4.4964104,4.7950773,4.824616,4.0303593,6.1440005,9.173334,10.745437,8.116513,4.8049235,1.8740515,0.35446155,0.17394873,0.15425642,0.12471796,0.098461546,0.08533334,0.08205129,0.07876924,0.1148718,0.1148718,0.10502565,0.09189744,0.07876924,0.10502565,0.17723078,0.32164106,0.4660513,0.42994875,0.41025645,0.30851284,0.21333335,0.16082053,0.1148718,0.11158975,0.1148718,0.12143591,0.12471796,0.12143591,0.128,0.14112821,0.15097436,0.16410258,0.17723078,0.19364104,0.20348719,0.20676924,0.21333335,0.22646156,0.24943592,0.25928208,0.26256412,0.25928208,0.25928208,0.26584616,0.27241027,0.28225642,0.28882053,0.30194873,0.2986667,0.28882053,0.28225642,0.28225642,0.2986667,0.30194873,0.30851284,0.32164106,0.38728207,0.5874872,1.8445129,2.605949,3.1967182,3.7054362,3.9811285,4.201026,4.391385,4.5128207,4.562052,4.565334,5.074052,5.874872,6.62318,7.1515903,7.4765134,7.5191803,7.525744,7.243488,6.5280004,5.3398976,3.5314875,2.2777438,1.3029745,0.61374366,0.49887183,0.50543594,0.5546667,0.6235898,0.6892308,0.7318975,0.8533334,0.98133343,1.1257436,1.3193847,1.654154,2.7831798,4.4701543,6.052103,6.705231,5.428513,0.0,0.0,0.016410258,0.118153855,0.30194873,0.5152821,1.3226668,2.2022567,2.3663592,1.7460514,0.9911796,0.5513847,1.4736412,2.8849232,3.629949,2.2711797,2.359795,3.767795,4.857436,4.778667,3.4756925,4.0041027,6.0225644,6.2194877,4.263385,2.8192823,3.31159,5.5696416,5.0904617,2.0086155,1.1027694,1.0568206,1.024,1.1290257,1.4703591,2.0841026,2.4418464,2.4648206,2.4385643,2.4582565,2.412308,2.6190772,2.3893335,2.681436,3.9778464,6.2720003,4.3651285,2.5206156,1.3883078,0.97805136,0.69907695,0.51856416,0.44964105,0.35446155,0.25271797,0.318359,0.4397949,0.4266667,0.41025645,0.55794877,1.0633847,0.8467693,0.79097444,0.6662565,0.39056414,0.006564103,0.08533334,0.08205129,0.03938462,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.013128206,0.0032820515,0.0,0.14769232,0.508718,1.086359,1.8970258,2.4352822,2.484513,2.2186668,2.1924105,2.5600002,2.2646155,2.100513,2.3433847,2.737231,2.7011285,2.5895386,2.2547693,1.6869745,1.0108719,0.83035904,0.67938465,0.51856416,0.34133336,0.16410258,0.30851284,0.49887183,0.51856416,0.36430773,0.23958977,0.48574364,0.49230772,0.3708718,0.27897438,0.4135385,0.4135385,0.4266667,0.60061544,0.8467693,0.84348726,0.60061544,0.5907693,0.5316923,0.37743592,0.3249231,0.25928208,0.26256412,0.2297436,0.13456412,0.04266667,0.029538464,0.009846155,0.006564103,0.04266667,0.13456412,0.098461546,0.04266667,0.006564103,0.0,0.0,0.0,0.02297436,0.029538464,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.006564103,0.006564103,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.01969231,0.01969231,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.029538464,0.052512825,0.049230773,0.02297436,0.013128206,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.032820515,0.072205134,0.04266667,0.009846155,0.0,0.0,0.0,0.0,0.04266667,0.03938462,0.01969231,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.029538464,0.036102567,0.02297436,0.006564103,0.036102567,0.04266667,0.04594872,0.049230773,0.04266667,0.0,0.0,0.026256412,0.026256412,0.006564103,0.036102567,0.006564103,0.013128206,0.032820515,0.032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.04594872,0.07876924,0.09189744,0.07548718,0.07548718,0.108307704,0.15097436,0.20676924,0.2986667,0.28882053,0.28225642,0.3117949,0.35446155,0.32164106,0.18707694,0.101743594,0.052512825,0.029538464,0.016410258,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.03938462,0.029538464,0.032820515,0.06235898,0.108307704,0.10502565,0.06564103,0.03938462,0.03938462,0.055794876,0.04266667,0.029538464,0.02297436,0.04594872,0.13128206,0.2297436,0.28225642,0.32820517,0.37415388,0.4004103,0.35446155,0.26912823,0.17394873,0.10502565,0.101743594,0.15753847,0.15097436,0.12471796,0.09189744,0.04594872,0.03938462,0.04266667,0.04266667,0.03938462,0.049230773,0.06564103,0.055794876,0.03938462,0.029538464,0.029538464,0.032820515,0.08861539,0.15425642,0.2100513,0.24943592,0.34789747,0.6104616,1.024,1.4375386,1.5721027,1.6213335,1.657436,1.6771283,2.03159,3.4100516,4.841026,7.5979495,9.160206,8.907488,8.119796,8.470975,8.67118,8.441437,7.463385,5.3760004,5.2578464,6.2030773,7.2369237,8.231385,9.878975,6.012718,6.5739493,7.4863596,7.4141545,7.755488,10.709334,12.130463,11.536411,10.65354,13.403898,12.2157955,9.107693,9.252103,10.788103,4.8082056,4.84759,6.340924,7.3616414,8.392206,12.3306675,12.035283,7.653744,3.5052311,1.5556924,1.4211283,1.2668719,1.3587693,1.8313848,2.7634873,4.1780515,2.556718,3.876103,7.020308,9.622975,8.070564,5.8781543,4.3684106,2.6157951,0.827077,0.31507695,0.16738462,0.108307704,0.08205129,0.072205134,0.07876924,0.08533334,0.098461546,0.098461546,0.0951795,0.098461546,0.10502565,0.118153855,0.14769232,0.19692309,0.27241027,0.3511795,0.31507695,0.27241027,0.256,0.21333335,0.15425642,0.13128206,0.12471796,0.128,0.13456412,0.14769232,0.15425642,0.16082053,0.17066668,0.18379489,0.190359,0.20020515,0.2100513,0.21989745,0.23302566,0.26912823,0.2855385,0.29210258,0.28882053,0.28882053,0.28882053,0.28882053,0.29210258,0.30194873,0.30851284,0.30851284,0.36430773,0.45292312,0.52512825,0.48246157,0.36102566,0.34133336,0.3708718,0.53825647,1.086359,2.1398976,3.0358977,3.817026,4.4767184,4.972308,5.874872,6.8233852,7.3583593,7.2664623,6.5870776,6.3606157,6.5969234,6.7938466,6.770872,6.6461544,6.439385,6.1374364,5.4186673,4.2207184,2.733949,1.204513,0.63343596,0.5152821,0.5218462,0.5218462,0.5481026,0.61374366,0.67938465,0.7384616,0.78769237,0.88287187,0.97805136,1.086359,1.2603078,1.5983591,2.3401027,2.9997952,3.3050258,3.062154,2.1398976,0.0,0.0,0.0,0.009846155,0.068923086,0.24287182,1.211077,2.5238976,2.92759,2.3072822,1.6869745,1.0272821,2.8882053,5.110154,5.7009234,2.8225644,2.7437952,4.8836927,6.265436,5.5958977,3.2722054,4.082872,6.3212314,6.9382567,4.9887185,1.6213335,1.654154,1.595077,1.4342566,1.214359,1.0502565,0.9124103,1.086359,1.6114873,2.034872,1.4080001,1.657436,1.6705642,1.7427694,2.172718,3.2525132,4.0041027,2.737231,1.4966155,1.3029745,2.1398976,2.1202054,1.4834872,0.94523084,0.76800007,0.76800007,0.9189744,1.0108719,0.892718,0.6892308,0.7778462,1.1323078,1.2307693,1.1716924,1.0043077,0.7122052,0.26584616,0.06564103,0.0032820515,0.0032820515,0.013128206,0.13784617,0.128,0.059076928,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.02297436,0.0032820515,0.0,0.0,0.04594872,0.23302566,0.827077,0.6235898,0.69579494,1.3718976,2.231795,2.8717952,3.4133337,2.9538465,1.9265642,2.103795,2.297436,2.3433847,2.2908719,2.1924105,2.1136413,1.8773335,1.404718,1.014154,0.8467693,0.8369231,0.86646163,1.1946667,1.1060513,0.5874872,0.3052308,0.5349744,0.79097444,0.74830776,0.65969235,1.3554872,1.5721027,1.1388719,0.79097444,0.73517954,0.6301539,0.5349744,0.41682056,0.28882053,0.20348719,0.21989745,0.34789747,0.49887183,0.54482055,0.48902568,0.4660513,0.318359,0.1148718,0.016410258,0.09189744,0.29210258,0.21333335,0.09189744,0.013128206,0.0,0.0,0.0,0.036102567,0.055794876,0.04266667,0.006564103,0.0,0.0032820515,0.0032820515,0.006564103,0.006564103,0.0,0.0,0.0,0.0,0.0032820515,0.026256412,0.03938462,0.04266667,0.052512825,0.098461546,0.098461546,0.07548718,0.04266667,0.016410258,0.0032820515,0.0,0.0,0.0,0.0032820515,0.02297436,0.055794876,0.055794876,0.032820515,0.009846155,0.04266667,0.12143591,0.13784617,0.101743594,0.04266667,0.013128206,0.0032820515,0.0,0.0032820515,0.009846155,0.026256412,0.01969231,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02297436,0.026256412,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.059076928,0.072205134,0.06235898,0.04594872,0.03938462,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.006564103,0.0,0.0,0.0,0.0,0.009846155,0.009846155,0.0,0.0,0.0,0.0,0.01969231,0.055794876,0.08533334,0.016410258,0.0,0.0,0.0,0.0,0.0,0.036102567,0.036102567,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.059076928,0.072205134,0.059076928,0.032820515,0.0,0.009846155,0.0032820515,0.0032820515,0.009846155,0.0,0.0,0.06235898,0.072205134,0.03938462,0.08205129,0.032820515,0.04594872,0.072205134,0.072205134,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01969231,0.04594872,0.06564103,0.072205134,0.072205134,0.07876924,0.098461546,0.12143591,0.14112821,0.15425642,0.19364104,0.24943592,0.3446154,0.42338464,0.37415388,0.23302566,0.118153855,0.04594872,0.01969231,0.016410258,0.006564103,0.0,0.0,0.0,0.0,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.016410258,0.016410258,0.026256412,0.026256412,0.032820515,0.04266667,0.04266667,0.032820515,0.02297436,0.016410258,0.036102567,0.11158975,0.20020515,0.25271797,0.2986667,0.34133336,0.36430773,0.33476925,0.26912823,0.17723078,0.098461546,0.08205129,0.12471796,0.15753847,0.13456412,0.07548718,0.052512825,0.06564103,0.10502565,0.13128206,0.14112821,0.15753847,0.17066668,0.13128206,0.07548718,0.03938462,0.036102567,0.059076928,0.08533334,0.12143591,0.16082053,0.20676924,0.3117949,0.54482055,0.90912825,1.3259488,1.6311796,1.654154,1.719795,1.9200002,2.1956925,2.3269746,3.1573336,4.2994876,5.1659493,5.0576415,3.1540515,2.612513,2.487795,3.4888208,4.9887185,5.0182567,4.1222568,6.0160003,8.576,9.682052,7.243488,5.668103,7.325539,9.258667,9.45559,6.8562055,7.6931286,8.034462,7.282872,6.426257,8.044309,7.3780518,6.298257,7.062975,7.860513,2.8192823,5.674667,7.722667,9.498257,11.418258,13.804309,12.527591,8.795898,4.6933336,1.8970258,1.6738462,1.7394873,1.6213335,1.5983591,1.8806155,2.6223593,2.1070771,2.2416413,2.9144619,3.6496413,3.620103,4.844308,7.1122055,6.1013336,2.3466668,1.2504616,0.47589746,0.17394873,0.0951795,0.07876924,0.06564103,0.06564103,0.07548718,0.07876924,0.08533334,0.10502565,0.128,0.13784617,0.14441027,0.14769232,0.12143591,0.128,0.15097436,0.20020515,0.25928208,0.28225642,0.19692309,0.16738462,0.16082053,0.15425642,0.15425642,0.16410258,0.17066668,0.17394873,0.17723078,0.18707694,0.18707694,0.20020515,0.2231795,0.24287182,0.256,0.29210258,0.318359,0.33805132,0.34789747,0.34789747,0.34789747,0.3511795,0.35774362,0.36758977,0.39056414,0.5349744,0.90256417,1.2668719,1.401436,1.0699488,0.5940513,0.44307697,0.5152821,0.92553854,2.0217438,2.937436,3.9286156,4.821334,5.5597954,6.186667,7.3386674,8.736821,9.757539,9.813334,8.369231,6.928411,6.1440005,5.481026,4.821334,4.466872,4.266667,3.754667,2.7437952,1.5031796,0.761436,0.57764107,0.5349744,0.5481026,0.56451285,0.56451285,0.61374366,0.6629744,0.69907695,0.72861546,0.77456415,0.8533334,0.9616411,1.1158975,1.3489232,1.7033848,1.9035898,1.7723079,1.4112822,1.014154,0.86646163,0.0,0.0,0.0,0.0,0.0,0.0,0.049230773,0.14441027,0.23630771,0.2855385,0.25928208,0.18707694,0.068923086,0.0,0.0032820515,0.016410258,0.052512825,0.14441027,0.14441027,0.049230773,0.0,0.0,0.0,0.036102567,0.08205129,0.04594872,0.36430773,1.8609232,2.6847181,2.477949,2.3794873,2.5764105,2.7437952,2.7569232,2.3466668,1.1126155,0.90584624,1.3029745,1.7624617,2.1530259,2.7766156,2.5206156,1.4867693,0.761436,0.56451285,0.25928208,0.40697438,0.40697438,0.7187693,1.1355898,0.79425645,1.3062565,1.654154,1.5064616,0.99774367,0.7187693,1.2668719,2.1070771,2.4549747,1.9068719,0.44307697,0.35774362,0.15097436,0.01969231,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.101743594,0.36430773,0.6071795,0.4135385,0.58420515,3.6726158,4.1124105,1.9429746,2.8225644,2.6289232,2.7175386,3.0096412,3.4198978,3.8596926,3.895795,3.5478978,3.5380516,3.826872,3.629949,2.556718,2.4615386,2.3696413,1.9167181,1.3423591,1.463795,1.7985642,1.8510771,2.15959,4.273231,4.6276927,2.4910772,0.9353847,0.77456415,0.58092314,0.702359,0.8336411,0.69251287,0.36758977,0.3052308,0.6104616,0.7975385,1.020718,1.3817437,1.9068719,1.3095386,0.47261542,0.016410258,0.036102567,0.12143591,0.072205134,0.02297436,0.0,0.0,0.0,0.0,0.0,0.029538464,0.06564103,0.029538464,0.006564103,0.009846155,0.02297436,0.029538464,0.029538464,0.006564103,0.0,0.0,0.0032820515,0.016410258,0.07548718,0.13784617,0.15425642,0.20676924,0.48902568,0.49887183,0.37415388,0.2100513,0.07548718,0.016410258,0.0032820515,0.0,0.0,0.02297436,0.108307704,0.27897438,0.28225642,0.16082053,0.055794876,0.21333335,0.5546667,0.5481026,0.2986667,0.013128206,0.0,0.0,0.0,0.013128206,0.052512825,0.13784617,0.101743594,0.055794876,0.01969231,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016410258,0.07548718,0.016410258,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06235898,0.029538464,0.0,0.0,0.0,0.0,0.055794876,0.055794876,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07876924,0.15753847,0.0,0.049230773,0.02297436,0.02297436,0.049230773,0.0,0.0,0.055794876,0.108307704,0.118153855,0.04594872,0.0951795,0.07876924,0.036102567,0.013128206,0.06235898,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01969231,0.049230773,0.06235898,0.08533334,0.08205129,0.101743594,0.14441027,0.16738462,0.15425642,0.28882053,0.49230772,0.67938465,0.7778462,0.6071795,0.3446154,0.13784617,0.03938462,0.016410258,0.016410258,0.006564103,0.0,0.0,0.0,0.013128206,0.006564103,0.0,0.0,0.0,0.0,0.0,0.006564103,0.016410258,0.016410258,0.016410258,0.016410258,0.02297436,0.029538464,0.029538464,0.029538464,0.029538464,0.02297436,0.026256412,0.07548718,0.12471796,0.18379489,0.23958977,0.27897438,0.28882053,0.28882053,0.25271797,0.17394873,0.08205129,0.04594872,0.068923086,0.10502565,0.1148718,0.101743594,0.07548718,0.15097436,0.23302566,0.29210258,0.318359,0.3052308,0.26912823,0.18707694,0.11158975,0.072205134,0.06235898,0.072205134,0.07548718,0.101743594,0.14769232,0.18379489,0.318359,0.5349744,0.79097444,1.0601027,1.3259488,1.7296412,2.0217438,2.412308,2.7569232,2.546872,1.9626669,2.156308,2.556718,2.9440002,3.4330258,3.6660516,4.0336413,4.325744,4.6769233,5.5532312,4.5423594,3.3903592,4.092718,5.9602056,5.6320004,5.5696416,4.5029745,3.9351797,4.965744,8.283898,10.164514,9.143796,7.7259493,7.716103,10.194052,9.350565,5.2414365,2.5862565,2.8553848,4.273231,6.38359,9.337437,16.210052,21.871592,12.983796,6.7971287,4.3716927,3.0030773,1.719795,1.2832822,1.4276924,1.5556924,1.7263591,1.913436,1.9987694,2.4516926,4.5423594,6.7577443,7.5881033,5.5236926,5.937231,7.131898,6.5411286,4.4734364,4.1189747,1.5556924,0.45620516,0.15753847,0.15097436,0.09189744,0.09189744,0.09189744,0.09189744,0.09189744,0.09189744,0.06564103,0.07876924,0.1148718,0.15753847,0.18379489,0.15753847,0.15097436,0.15753847,0.17066668,0.18379489,0.19692309,0.19692309,0.18707694,0.16738462,0.16738462,0.16738462,0.18707694,0.19692309,0.19692309,0.19692309,0.19692309,0.19692309,0.20348719,0.21989745,0.24287182,0.28225642,0.33476925,0.37743592,0.39712822,0.39712822,0.39712822,0.4135385,0.446359,0.49887183,0.6104616,1.3292309,2.6190772,3.5413337,3.5249233,2.3663592,1.2537436,0.77456415,0.95835906,1.654154,2.5337439,3.4133337,4.391385,5.3694363,6.2818465,7.125334,8.103385,9.363693,10.5780525,10.820924,8.576,5.8157954,3.442872,1.6902566,0.7450257,0.7318975,0.7089231,0.65641034,0.6268718,0.6268718,0.6268718,0.5874872,0.5973334,0.6170257,0.6268718,0.6268718,0.67282057,0.69579494,0.7089231,0.7253334,0.761436,0.8598975,0.9944616,1.2077949,1.5425643,2.044718,2.2153847,2.1300514,1.910154,1.6738462,1.5261539,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.029538464,0.04594872,0.055794876,0.052512825,0.036102567,0.013128206,0.0032820515,0.016410258,0.026256412,0.026256412,0.032820515,0.029538464,0.013128206,0.02297436,0.06235898,0.118153855,0.23630771,0.4594872,0.81394875,1.6016412,1.5688206,1.5622566,1.6443079,1.086359,1.9462565,3.0851285,3.0391798,2.1136413,2.3827693,3.1803079,2.4451284,1.3161026,0.63343596,0.9353847,1.4769232,1.8609232,1.8707694,1.7526156,2.1891284,2.1891284,2.5107694,2.8717952,2.5173335,0.23302566,0.5973334,0.8960001,0.93866676,0.8598975,1.0962052,1.6344616,1.5097437,1.4211283,1.5097437,1.332513,2.0086155,2.2744617,1.4802053,0.15753847,0.0,0.009846155,0.04266667,0.0951795,0.118153855,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.026256412,0.13456412,0.08533334,0.049230773,0.072205134,0.12143591,0.08205129,0.118153855,0.73517954,0.92553854,0.9616411,2.409026,3.5610259,4.841026,4.4800005,2.8389745,2.409026,3.8498464,5.58277,5.408821,3.4921029,2.349949,2.789744,2.553436,2.2383592,2.100513,2.0742567,1.2800001,1.5130258,2.3269746,3.1409233,3.2722054,2.9604106,2.4746668,2.3729234,2.4943593,1.9462565,1.394872,1.7985642,2.2416413,2.100513,1.024,0.6268718,0.6826667,0.85005134,1.1224617,1.8215386,1.8182565,0.955077,0.24615386,0.03938462,0.036102567,0.016410258,0.0032820515,0.0,0.0032820515,0.013128206,0.013128206,0.013128206,0.02297436,0.036102567,0.01969231,0.013128206,0.049230773,0.07876924,0.068923086,0.029538464,0.016410258,0.0032820515,0.029538464,0.08205129,0.12471796,0.07876924,0.055794876,0.03938462,0.04266667,0.098461546,0.101743594,0.16410258,0.19692309,0.16738462,0.07548718,0.026256412,0.0032820515,0.0,0.118153855,0.5940513,0.6498462,0.38400003,0.13128206,0.16082053,0.6892308,1.2865642,1.0043077,0.5021539,0.15753847,0.08533334,0.318359,0.26256412,0.14112821,0.072205134,0.03938462,0.02297436,0.032820515,0.026256412,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.006564103,0.0,0.0,0.0,0.049230773,0.108307704,0.13456412,0.098461546,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.06235898,0.15753847,0.072205134,0.0,0.0,0.0,0.0,0.029538464,0.029538464,0.013128206,0.06235898,0.013128206,0.0,0.016410258,0.059076928,0.13456412,0.06564103,0.01969231,0.029538464,0.068923086,0.049230773,0.009846155,0.009846155,0.02297436,0.03938462,0.0951795,0.07548718,0.036102567,0.006564103,0.0032820515,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.026256412,0.049230773,0.052512825,0.052512825,0.07548718,0.12143591,0.15425642,0.18379489,0.318359,0.446359,0.5415385,0.6695385,0.5546667,0.37415388,0.19692309,0.07548718,0.03938462,0.01969231,0.006564103,0.0,0.0,0.0,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.026256412,0.026256412,0.04266667,0.049230773,0.04266667,0.04266667,0.032820515,0.02297436,0.016410258,0.02297436,0.052512825,0.101743594,0.15753847,0.2100513,0.25271797,0.31507695,0.3446154,0.26912823,0.16738462,0.08861539,0.068923086,0.0951795,0.12143591,0.14769232,0.17066668,0.18707694,0.4266667,0.50543594,0.46276927,0.35774362,0.256,0.2100513,0.17066668,0.14441027,0.128,0.08533334,0.07876924,0.08205129,0.098461546,0.12471796,0.17066668,0.27569234,0.5284103,0.8795898,1.1979488,1.2898463,1.6443079,1.6311796,1.6377437,1.7099489,1.5589745,1.4998976,1.723077,2.097231,2.7208207,3.9220517,5.5893335,5.9569235,5.435077,4.857436,5.4941545,4.529231,3.9975388,5.0084105,7.634052,10.929232,11.2672825,11.346052,9.284924,6.4623594,7.515898,11.185231,12.396309,11.411694,10.082462,11.828514,12.461949,8.484103,4.71959,3.3214362,3.761231,4.5522056,7.200821,11.211488,14.221129,11.98277,8.274052,4.5423594,2.1169233,1.2635899,1.1946667,2.2416413,3.4888208,4.532513,4.9394875,4.2338467,5.651693,7.6603084,7.3616414,4.7491283,2.7175386,2.4976413,2.9669745,3.370667,3.5052311,3.7185643,2.0611284,0.8402052,0.26256412,0.20020515,0.190359,0.14112821,0.34133336,0.40369233,0.25271797,0.1148718,0.09189744,0.08205129,0.07876924,0.08861539,0.12143591,0.128,0.15097436,0.17066668,0.17723078,0.15753847,0.16082053,0.17723078,0.17723078,0.16738462,0.16738462,0.18707694,0.2100513,0.21661541,0.2100513,0.2100513,0.2100513,0.21661541,0.2231795,0.2231795,0.21989745,0.24615386,0.27569234,0.31507695,0.36758977,0.446359,0.64000005,1.1979488,1.5524104,1.7690258,2.5632823,4.2207184,4.197744,3.620103,3.2886157,3.6726158,4.161641,4.821334,5.7731285,6.8988724,7.8539495,7.962257,7.722667,7.456821,7.433847,7.893334,8.421744,7.827693,7.0531287,6.245744,4.7294364,2.5074873,1.6902566,1.4769232,1.4375386,1.5130258,1.4112822,1.522872,1.657436,1.7066668,1.6377437,1.6705642,1.7033848,1.6311796,1.4375386,1.211077,0.9878975,0.81394875,0.8566154,1.1913847,1.8116925,2.1070771,2.172718,2.4451284,2.8258464,2.6912823,2.2482052,1.7591796,1.2800001,0.9124103,0.8041026,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.036102567,0.06564103,0.036102567,0.016410258,0.006564103,0.006564103,0.013128206,0.006564103,0.029538464,0.08533334,0.35774362,1.2012309,3.4921029,5.684513,6.872616,6.6133337,4.926359,4.516103,4.4012313,3.5544617,2.3072822,2.3466668,2.1333334,2.5961027,2.789744,2.3335385,1.4276924,1.585231,1.0994873,0.48246157,0.101743594,0.190359,0.48574364,0.7811283,0.8598975,0.8205129,1.0666667,1.0535386,1.214359,1.3653334,1.1454359,0.036102567,0.16738462,0.28225642,0.318359,0.32820517,0.47589746,0.69907695,0.8598975,0.82379496,0.85005134,1.6213335,3.1606157,3.2754874,2.356513,1.204513,1.0633847,1.1093334,1.2307693,1.394872,1.4441026,1.0994873,0.512,0.3446154,0.49887183,0.6301539,0.14769232,0.0951795,0.1148718,0.08533334,0.01969231,0.06564103,0.04266667,0.013128206,0.0,0.0,0.0,0.072205134,0.14769232,0.27241027,0.5546667,1.1684103,1.7001027,2.550154,3.3509746,4.069744,5.0116925,5.671385,5.3431797,3.7382567,1.7001027,1.214359,1.5786668,1.4900514,1.2373334,1.0338463,1.0043077,0.65969235,0.84348726,1.3653334,1.8707694,1.8510771,2.2514873,2.7011285,3.0490258,3.5610259,4.9329233,2.7044106,2.412308,3.1113849,3.3575387,1.214359,0.69251287,0.8402052,0.90256417,0.8041026,1.1684103,1.2800001,0.77456415,0.26912823,0.03938462,0.016410258,0.055794876,0.098461546,0.07548718,0.013128206,0.032820515,0.013128206,0.006564103,0.009846155,0.013128206,0.016410258,0.06564103,0.21989745,0.23302566,0.098461546,0.02297436,0.098461546,0.14441027,0.15425642,0.12471796,0.07876924,0.049230773,0.06564103,0.08533334,0.08205129,0.04594872,0.02297436,0.07876924,0.15097436,0.18707694,0.14769232,0.06235898,0.02297436,0.006564103,0.13456412,0.67938465,1.204513,1.0404103,0.7056411,0.56451285,0.8369231,1.1881026,1.1749744,1.1454359,1.5458462,2.917744,4.089436,2.3958976,0.65641034,0.029538464,0.006564103,0.0,0.009846155,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02297436,0.049230773,0.08205129,0.09189744,0.0,0.0,0.0,0.0,0.0,0.0,0.029538464,0.036102567,0.02297436,0.013128206,0.06564103,0.08533334,0.036102567,0.0,0.006564103,0.036102567,0.059076928,0.072205134,0.068923086,0.06564103,0.10502565,0.101743594,0.101743594,0.101743594,0.11158975,0.15753847,0.098461546,0.06564103,0.04594872,0.04266667,0.098461546,0.06235898,0.059076928,0.072205134,0.098461546,0.16082053,0.11158975,0.03938462,0.02297436,0.04266667,0.0,0.0,0.026256412,0.026256412,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.032820515,0.06564103,0.07876924,0.072205134,0.08861539,0.14112821,0.19692309,0.24943592,0.36430773,0.49230772,0.62030774,0.7778462,0.7384616,0.58092314,0.41025645,0.27241027,0.15425642,0.049230773,0.009846155,0.0032820515,0.009846155,0.009846155,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.02297436,0.029538464,0.032820515,0.029538464,0.026256412,0.026256412,0.02297436,0.016410258,0.013128206,0.009846155,0.026256412,0.068923086,0.1148718,0.16738462,0.2297436,0.30194873,0.318359,0.24943592,0.16082053,0.08533334,0.059076928,0.098461546,0.17066668,0.23958977,0.28882053,0.31507695,0.4201026,0.45620516,0.4594872,0.40697438,0.19692309,0.13456412,0.13784617,0.15097436,0.13784617,0.072205134,0.09189744,0.108307704,0.1148718,0.118153855,0.15753847,0.27897438,0.5021539,0.7778462,1.0502565,1.2438976,1.5195899,1.4933335,1.2996924,1.1323078,1.2471796,1.3718976,1.5753847,2.2711797,3.3476925,4.1714873,5.789539,5.658257,4.9460516,4.604718,5.3760004,5.3760004,5.5269747,6.5345645,8.815591,12.481642,12.416001,11.946668,9.580308,6.370462,5.914257,7.9425645,9.737847,10.41395,9.93477,9.114257,11.9860525,8.635077,5.546667,4.9920006,5.041231,4.6276927,5.4547696,7.181129,8.92718,9.288206,8.612103,5.0215387,2.172718,1.3193847,1.3226668,2.3204105,3.31159,4.141949,4.4865646,3.8400004,3.5872824,4.017231,3.508513,2.4681027,3.3411283,1.9364104,1.8412309,2.1267693,2.5074873,3.3247182,2.986667,1.6377437,0.67938465,0.49887183,0.4594872,1.7985642,2.5238976,2.15959,1.0371283,0.29538465,0.16082053,0.118153855,0.101743594,0.09189744,0.098461546,0.118153855,0.14441027,0.16410258,0.17066668,0.16082053,0.14769232,0.14112821,0.128,0.118153855,0.13128206,0.12471796,0.15425642,0.21661541,0.28225642,0.29538465,0.23630771,0.2100513,0.21333335,0.2297436,0.23958977,0.25928208,0.3249231,0.36758977,0.4004103,0.512,0.5513847,0.92553854,1.204513,1.3718976,1.8248206,2.92759,3.367385,3.623385,4.1714873,5.4908724,6.701949,6.665847,6.5247183,7.056411,8.65477,9.537642,9.547488,8.914052,8.01477,7.39118,7.273026,6.616616,5.7665644,4.8836927,3.9778464,2.4549747,2.15959,2.2219489,2.1924105,2.0578463,1.972513,2.0906668,2.2055387,2.2350771,2.2219489,2.2646155,2.4484105,2.7142565,2.9604106,3.062154,2.8849232,2.2613335,1.7165129,1.5556924,1.8642052,2.2055387,2.048,1.975795,2.0775387,1.9462565,1.5392822,1.1585642,0.8041026,0.53825647,0.46933338,0.0,0.0,0.0,0.0032820515,0.006564103,0.006564103,0.016410258,0.009846155,0.013128206,0.036102567,0.06564103,0.036102567,0.07876924,0.101743594,0.072205134,0.013128206,0.02297436,0.27897438,1.3193847,2.4746668,1.8806155,3.8728209,6.0192823,7.0465646,6.4557953,4.529231,3.754667,3.8038976,3.0490258,1.7526156,2.0545642,1.4211283,1.332513,1.5524104,1.5195899,0.35446155,0.108307704,0.055794876,0.04266667,0.009846155,0.006564103,0.0,0.0,0.0,0.006564103,0.029538464,0.068923086,0.052512825,0.02297436,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.01969231,0.108307704,0.64000005,0.79425645,0.7318975,1.5885129,2.4385643,2.284308,1.9462565,1.8412309,1.9823592,2.0086155,1.8707694,1.7099489,1.5688206,1.3784616,1.1782565,1.5097437,1.9528207,1.9561027,0.82379496,0.5284103,0.34133336,0.20676924,0.118153855,0.12143591,0.32164106,0.30851284,0.20348719,0.101743594,0.09189744,0.67610264,0.9419488,0.9353847,0.78769237,0.69251287,0.6695385,0.81394875,1.6968206,3.2361028,4.6769233,5.218462,4.20759,2.3433847,0.7089231,0.8041026,0.86317956,0.78769237,0.5940513,0.37415388,0.28882053,0.29210258,0.42338464,0.5907693,0.7450257,0.8730257,1.591795,2.1103592,2.2514873,2.553436,4.263385,2.8882053,3.1540515,4.0434875,4.309334,2.477949,3.5610259,2.7766156,1.8346668,1.4408206,1.2964103,1.3292309,0.9517949,0.54482055,0.3314872,0.37415388,0.3249231,0.26256412,0.19692309,0.13784617,0.0951795,0.029538464,0.009846155,0.009846155,0.016410258,0.032820515,0.07876924,0.25271797,0.34789747,0.2986667,0.18707694,0.21333335,0.22646156,0.19692309,0.128,0.06235898,0.18707694,0.27241027,0.24943592,0.15425642,0.108307704,0.1148718,0.190359,0.2297436,0.21661541,0.23302566,0.24287182,0.15425642,0.06564103,0.10502565,0.44964105,1.214359,1.1881026,0.8763078,0.6235898,0.6235898,0.8992821,1.3193847,1.7624617,2.409026,3.748103,4.2896414,2.356513,0.5874872,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.029538464,0.14112821,0.029538464,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02297436,0.04266667,0.0,0.0,0.0,0.0,0.0,0.0,0.029538464,0.052512825,0.036102567,0.006564103,0.036102567,0.006564103,0.0,0.0,0.006564103,0.036102567,0.059076928,0.118153855,0.16082053,0.18051283,0.21989745,0.21661541,0.19692309,0.190359,0.17723078,0.09189744,0.068923086,0.059076928,0.032820515,0.013128206,0.072205134,0.059076928,0.10502565,0.14112821,0.15097436,0.17394873,0.09189744,0.029538464,0.02297436,0.04266667,0.0,0.04266667,0.068923086,0.04594872,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.006564103,0.013128206,0.029538464,0.049230773,0.07548718,0.08533334,0.08205129,0.101743594,0.17066668,0.30194873,0.4201026,0.5874872,0.7187693,0.79425645,0.8566154,0.7975385,0.67610264,0.5677949,0.47261542,0.30194873,0.15425642,0.07876924,0.04266667,0.026256412,0.02297436,0.026256412,0.026256412,0.01969231,0.009846155,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.026256412,0.026256412,0.016410258,0.009846155,0.016410258,0.016410258,0.016410258,0.013128206,0.006564103,0.016410258,0.04266667,0.068923086,0.1148718,0.17723078,0.24615386,0.26256412,0.2231795,0.15425642,0.08861539,0.059076928,0.09189744,0.16738462,0.256,0.318359,0.31507695,0.28225642,0.28225642,0.318359,0.31507695,0.12471796,0.07548718,0.0951795,0.118153855,0.108307704,0.055794876,0.07548718,0.10502565,0.12143591,0.13456412,0.17723078,0.31507695,0.5316923,0.77128214,1.020718,1.2931283,1.5064616,1.4473847,1.2012309,0.9878975,1.1749744,1.3029745,1.4998976,2.2416413,3.2229745,3.367385,4.7524104,4.716308,4.2240005,4.20759,5.586052,6.409847,6.8496413,7.1548724,8.36595,12.291283,11.474052,11.362462,10.66995,9.284924,8.277334,7.318975,9.403078,12.35036,13.604104,10.233437,10.568206,9.009232,7.0465646,5.602462,5.041231,5.10359,4.7491283,4.8082056,5.4580517,6.1997952,7.1089234,5.2447186,3.2164104,2.1070771,1.4572309,2.169436,2.3926156,2.556718,2.678154,2.3433847,1.595077,1.4244103,1.4178462,1.8937438,3.895795,3.767795,3.6890259,3.4133337,3.4100516,4.8607183,4.886975,3.259077,1.975795,1.8970258,2.7798977,3.948308,3.9023592,2.861949,1.3883078,0.39384618,0.23958977,0.18051283,0.15425642,0.13456412,0.128,0.13456412,0.14441027,0.15753847,0.16410258,0.16738462,0.14769232,0.14112821,0.13456412,0.12471796,0.108307704,0.07876924,0.09189744,0.15097436,0.22646156,0.26584616,0.23630771,0.18707694,0.17394873,0.2231795,0.31507695,0.32164106,0.35774362,0.36758977,0.36758977,0.446359,0.4004103,0.5907693,1.0502565,1.5031796,1.3718976,1.7132308,2.409026,3.1409233,3.9351797,5.159385,6.9743595,6.9677954,6.370462,6.3277955,7.9228725,9.340718,9.350565,8.349539,6.9349747,5.933949,5.609026,5.3202057,4.8771286,4.269949,3.6857438,2.8225644,2.553436,2.477949,2.3794873,2.2219489,2.3893335,2.553436,2.6518977,2.7011285,2.7700515,2.9407182,3.2000003,3.6102567,4.066462,4.312616,4.0500517,3.0030773,2.0020514,1.4703591,1.4244103,1.6049232,1.4408206,1.2635899,1.1946667,1.1585642,0.9878975,0.8205129,0.6301539,0.45620516,0.39712822,0.0,0.0,0.0,0.0032820515,0.013128206,0.013128206,0.032820515,0.02297436,0.006564103,0.0,0.0,0.0,0.13128206,0.20676924,0.15753847,0.029538464,0.049230773,0.508718,2.4681027,4.240411,1.3784616,0.82379496,0.78769237,0.57764107,0.128,0.013128206,0.0032820515,0.0,0.03938462,0.08861539,0.036102567,0.013128206,0.049230773,0.06235898,0.03938462,0.032820515,0.08861539,0.14441027,0.128,0.052512825,0.02297436,0.0032820515,0.0,0.0,0.013128206,0.06235898,0.13784617,0.108307704,0.04266667,0.0,0.0,0.0,0.013128206,0.02297436,0.029538464,0.04594872,0.3249231,0.97805136,1.4145643,1.5327181,1.7001027,1.1126155,1.1290257,1.7033848,2.3696413,2.2416413,2.3794873,1.8674873,1.083077,0.48246157,0.6235898,1.3620514,2.353231,2.9571285,2.7634873,1.6016412,1.5688206,1.5261539,1.4769232,1.4998976,1.7558975,2.4484105,2.3138463,1.591795,0.827077,0.85005134,1.7788719,2.0906668,1.7755898,1.1651284,0.9616411,1.1552821,1.1126155,0.86317956,0.6826667,1.0994873,2.3663592,2.8356924,2.1136413,0.88287187,0.9189744,0.9714873,0.7581539,0.6071795,0.5677949,0.4135385,0.36102566,0.5218462,0.65312827,0.6859488,0.7187693,1.0371283,1.1290257,0.9616411,0.761436,1.0043077,2.162872,3.6496413,4.46359,4.381539,3.948308,6.8463597,4.9952826,3.2820516,3.2951798,3.318154,2.8160002,2.0775387,1.3981539,1.014154,1.0994873,0.8730257,0.6268718,0.48246157,0.40369233,0.18379489,0.08205129,0.04594872,0.03938462,0.03938462,0.059076928,0.049230773,0.16082053,0.3511795,0.49230772,0.37415388,0.26584616,0.18051283,0.12143591,0.09189744,0.08533334,0.34133336,0.44964105,0.36102566,0.19364104,0.19364104,0.23958977,0.4201026,0.58092314,0.58092314,0.28225642,0.4397949,0.3314872,0.17066668,0.08533334,0.118153855,0.6235898,0.65641034,0.512,0.38728207,0.380718,0.7515898,1.3226668,1.7952822,1.9790771,1.7952822,0.75487185,0.19692309,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.036102567,0.04266667,0.0,0.0,0.006564103,0.032820515,0.059076928,0.055794876,0.2100513,0.21661541,0.118153855,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.01969231,0.0032820515,0.032820515,0.032820515,0.0,0.0,0.06235898,0.04594872,0.026256412,0.08533334,0.34789747,0.08533334,0.01969231,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.029538464,0.036102567,0.013128206,0.0,0.0,0.03938462,0.08861539,0.1148718,0.09189744,0.10502565,0.2100513,0.29538465,0.33805132,0.39712822,0.3249231,0.24943592,0.21661541,0.18707694,0.029538464,0.049230773,0.04594872,0.04594872,0.04594872,0.026256412,0.006564103,0.08861539,0.13784617,0.118153855,0.108307704,0.02297436,0.0,0.0,0.0,0.0,0.08861539,0.08205129,0.036102567,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.013128206,0.032820515,0.04594872,0.055794876,0.06564103,0.07548718,0.07876924,0.101743594,0.17394873,0.36430773,0.5546667,0.81394875,0.92225647,0.8533334,0.75487185,0.6498462,0.6235898,0.64000005,0.6170257,0.41682056,0.26912823,0.16082053,0.09189744,0.049230773,0.03938462,0.049230773,0.059076928,0.049230773,0.026256412,0.0032820515,0.0032820515,0.0032820515,0.0032820515,0.0032820515,0.0032820515,0.01969231,0.026256412,0.016410258,0.0032820515,0.013128206,0.013128206,0.016410258,0.01969231,0.016410258,0.016410258,0.026256412,0.03938462,0.068923086,0.1148718,0.17066668,0.20348719,0.190359,0.15097436,0.10502565,0.07876924,0.08533334,0.12471796,0.19692309,0.256,0.18707694,0.12471796,0.118153855,0.128,0.118153855,0.06235898,0.049230773,0.052512825,0.06564103,0.06564103,0.04266667,0.04266667,0.06564103,0.10502565,0.15753847,0.2297436,0.37415388,0.5907693,0.88615394,1.2209232,1.5064616,1.5425643,1.3489232,1.1651284,1.0994873,1.0994873,1.1323078,1.3817437,1.8609232,2.28759,2.0676925,3.4002054,4.056616,4.010667,4.027077,5.687795,6.452513,6.6428723,6.1374364,6.4295387,10.604308,9.921641,10.840616,12.507898,13.892924,13.778052,11.756309,13.590976,16.787693,18.274464,14.411489,9.609847,9.350565,8.474257,5.979898,5.031385,5.9930263,5.2348723,4.276513,3.9122055,4.2272825,4.7327185,5.0543594,4.7458467,3.7809234,2.546872,2.7667694,2.1300514,1.5786668,1.401436,1.2504616,1.5721027,2.0184617,2.3072822,2.5337439,3.1638978,5.431795,5.8880005,5.467898,5.5007186,7.6964107,6.9809237,5.408821,4.0402055,3.7874875,5.425231,5.149539,3.7021542,2.1366155,1.0075898,0.3446154,0.2986667,0.29538465,0.26256412,0.20676924,0.2231795,0.21661541,0.18379489,0.15425642,0.15097436,0.17066668,0.17066668,0.20348719,0.2297436,0.21333335,0.118153855,0.07876924,0.07876924,0.0951795,0.12471796,0.18051283,0.21333335,0.16082053,0.13128206,0.18379489,0.3511795,0.41025645,0.380718,0.32820517,0.28882053,0.29538465,0.3314872,0.5316923,1.3981539,2.4451284,2.2186668,1.9659488,2.0512822,2.1891284,2.3663592,2.8488207,4.8771286,6.235898,6.7314878,6.7840004,7.433847,8.172308,7.4797955,6.0849237,4.7294364,4.1813335,4.089436,3.9581542,3.7284105,3.3805132,2.934154,2.5337439,2.2022567,2.041436,2.0611284,2.1464617,2.7667694,3.1048207,3.2918978,3.4231799,3.570872,3.8301542,4.0041027,4.204308,4.394667,4.4077954,3.69559,2.4910772,1.5195899,1.0633847,0.9419488,0.90256417,0.94523084,0.96492314,0.9321026,0.88615394,0.86974365,0.80738467,0.6662565,0.49230772,0.4135385,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.026256412,0.06564103,0.07876924,0.029538464,0.029538464,0.029538464,0.01969231,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.128,0.26912823,0.06235898,0.049230773,0.2100513,0.24615386,0.13128206,0.108307704,0.18051283,0.23630771,0.2231795,0.14769232,0.06235898,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06564103,0.068923086,0.02297436,0.04594872,0.62030774,1.6508719,2.6880002,3.2000003,2.5796926,3.114667,4.348718,5.21518,4.7327185,1.9987694,2.878359,2.7503593,1.7723079,0.5874872,0.3052308,0.14769232,0.108307704,0.21661541,0.5513847,1.2373334,3.5183592,5.3792825,6.173539,6.370462,7.568411,9.019077,8.467693,5.940513,3.121231,3.3411283,2.8521028,2.5107694,1.7066668,0.6432821,0.3511795,0.88943595,1.4342566,1.4539489,0.9878975,0.67282057,1.0010257,1.1552821,1.0108719,0.6859488,0.56451285,0.636718,0.508718,0.65641034,0.85005134,0.16738462,0.54482055,1.0338463,1.2307693,1.1552821,1.2668719,1.595077,1.6705642,1.8346668,2.1891284,2.5796926,2.7142565,2.681436,2.481231,2.2514873,2.28759,3.0096412,3.0162053,3.876103,5.8912826,8.103385,5.796103,4.312616,3.0358977,1.9889232,1.8313848,1.6246156,1.4703591,1.1946667,0.7581539,0.24287182,0.18379489,0.15097436,0.108307704,0.059076928,0.04594872,0.059076928,0.21661541,0.25928208,0.15425642,0.108307704,0.0951795,0.06564103,0.03938462,0.02297436,0.0,0.013128206,0.04266667,0.128,0.25271797,0.3511795,0.28882053,0.5316923,1.3193847,1.8313848,0.18379489,0.29210258,0.3117949,0.26256412,0.16738462,0.04594872,0.032820515,0.14112821,0.34789747,0.60061544,0.80738467,0.761436,0.6826667,0.5973334,0.47589746,0.24287182,0.17066668,0.06235898,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.072205134,0.17723078,0.20676924,0.0,0.0,0.036102567,0.15753847,0.2986667,0.27569234,1.0436924,1.079795,0.5907693,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01969231,0.09189744,0.01969231,0.16410258,0.16410258,0.0,0.0,0.3052308,0.23630771,0.12471796,0.15097436,0.33476925,0.15097436,0.098461546,0.055794876,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.036102567,0.072205134,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.029538464,0.06235898,0.0,0.0,0.20020515,0.4397949,0.5677949,0.45620516,0.51856416,0.4594872,0.42994875,0.46933338,0.51856416,0.39712822,0.26584616,0.18051283,0.15097436,0.15097436,0.23958977,0.2231795,0.2231795,0.23630771,0.13784617,0.026256412,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.02297436,0.02297436,0.01969231,0.029538464,0.1148718,0.118153855,0.101743594,0.108307704,0.16738462,0.30194873,0.49887183,0.5874872,0.5218462,0.4135385,0.47261542,0.63343596,0.76800007,0.74830776,0.44307697,0.23630771,0.09189744,0.049230773,0.07548718,0.07548718,0.07548718,0.07548718,0.059076928,0.026256412,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.0032820515,0.009846155,0.016410258,0.013128206,0.0,0.013128206,0.02297436,0.029538464,0.026256412,0.016410258,0.016410258,0.032820515,0.059076928,0.08533334,0.12143591,0.14769232,0.15097436,0.14112821,0.1148718,0.09189744,0.07876924,0.14112821,0.21989745,0.23630771,0.07548718,0.016410258,0.0,0.02297436,0.06235898,0.06235898,0.049230773,0.04594872,0.052512825,0.055794876,0.029538464,0.029538464,0.029538464,0.055794876,0.13128206,0.28882053,0.42338464,0.5677949,0.92225647,1.4572309,1.9232821,1.3718976,1.0535386,1.0469744,1.1716924,0.97805136,0.8041026,1.1946667,1.6935385,2.0578463,2.228513,3.0687182,3.9581542,4.453744,4.5029745,4.457026,3.8334363,3.373949,3.5478978,4.46359,5.904411,8.247795,7.8014364,9.160206,12.983796,15.977027,19.24595,18.471386,15.232001,11.956513,11.933539,9.271795,5.8420515,6.3606157,10.049642,10.633847,8.792616,6.5739493,5.2414365,5.0215387,5.080616,4.092718,4.716308,5.717334,6.416411,6.698667,5.540103,3.9680004,2.8192823,2.3138463,2.044718,1.9954873,2.2678976,2.3696413,2.2383592,2.2121027,2.3105643,3.249231,4.1583595,5.412103,8.635077,7.1581545,7.072821,6.0849237,4.069744,3.0818465,3.6562054,3.121231,1.7558975,0.35774362,0.25928208,0.32164106,0.5284103,0.508718,0.30851284,0.380718,0.44307697,0.30194873,0.16738462,0.13456412,0.18379489,0.23302566,0.3249231,0.36430773,0.30194873,0.16738462,0.118153855,0.15097436,0.23958977,0.3249231,0.3511795,0.2297436,0.15097436,0.1148718,0.118153855,0.16738462,0.4594872,0.54482055,0.46276927,0.3314872,0.32164106,0.3446154,0.39712822,1.2077949,2.5862565,3.4034874,2.1956925,1.4605129,1.1946667,1.2832822,1.5425643,2.1136413,4.7950773,7.2960005,8.362667,7.752206,6.409847,5.139693,4.1682053,3.5478978,3.1442053,3.0687182,2.986667,2.8488207,2.665026,2.5173335,2.284308,2.0808206,1.972513,2.0118976,2.2416413,3.2918978,3.9318976,4.3027697,4.5456414,4.7917953,4.6211286,4.578462,4.522667,4.3716927,4.089436,2.5862565,1.6443079,1.1618463,0.9682052,0.80738467,0.8467693,0.8992821,0.9321026,0.92225647,0.88615394,0.8598975,0.7450257,0.574359,0.4004103,0.28882053,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.013128206,0.016410258,0.006564103,0.016410258,0.01969231,0.009846155,0.0,0.0,0.0,0.013128206,0.02297436,0.026256412,0.036102567,0.04594872,0.032820515,0.03938462,0.052512825,0.013128206,0.029538464,0.118153855,0.17723078,0.16410258,0.068923086,0.12471796,0.16738462,0.18379489,0.16082053,0.08533334,0.036102567,0.009846155,0.0,0.0,0.0,0.0,0.0,0.02297436,0.08861539,0.19692309,0.049230773,0.10502565,0.17394873,1.3554872,6.038975,4.775385,2.733949,1.332513,0.892718,0.6498462,0.8566154,1.1552821,1.3292309,1.2603078,0.9485129,1.3292309,1.2012309,1.0469744,1.7099489,4.4077954,3.1048207,1.6213335,0.7515898,0.571077,0.44307697,2.8127182,3.7809234,3.945026,3.9975388,4.7228723,4.352,3.0129232,1.6049232,0.7318975,0.7187693,0.6498462,0.6104616,0.77456415,0.86974365,0.16738462,1.0666667,1.2635899,1.3883078,1.6082052,1.6246156,1.8248206,1.6213335,1.214359,0.90256417,1.0666667,1.5491283,1.7263591,1.6902566,1.5688206,1.5589745,1.6935385,1.8937438,1.4539489,0.8336411,1.657436,2.9636924,3.2065644,3.314872,3.5544617,3.5544617,2.2350771,1.5622566,2.1136413,3.6430771,5.097026,4.850872,3.817026,2.5961027,1.8937438,2.5107694,3.114667,3.9614363,5.5236926,6.8660517,5.651693,4.9460516,4.457026,3.9614363,3.1507695,1.6114873,1.2373334,1.595077,1.6410258,1.1158975,0.55794877,0.3446154,0.20020515,0.12143591,0.08533334,0.04594872,0.072205134,0.036102567,0.006564103,0.0032820515,0.0,0.072205134,0.2986667,0.40369233,0.2986667,0.0951795,0.13128206,0.3314872,0.74830776,1.1191796,0.86646163,0.90912825,2.0086155,2.281026,1.3850257,0.508718,0.3314872,0.190359,0.14112821,1.529436,7.0104623,7.8112826,5.293949,3.006359,2.4155898,2.917744,1.3981539,0.5481026,0.48246157,0.69907695,0.072205134,0.013128206,0.0,0.0,0.0,0.0,0.01969231,0.016410258,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.0,0.0,0.013128206,0.036102567,0.049230773,0.036102567,0.2231795,0.61374366,0.8533334,0.764718,0.36102566,0.27897438,0.2297436,0.12471796,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.059076928,0.059076928,0.0032820515,0.01969231,0.0032820515,0.032820515,0.14441027,0.2986667,0.37743592,0.24287182,0.19692309,0.17723078,0.20020515,0.3249231,0.38400003,0.37743592,0.2855385,0.13784617,0.0,0.0,0.0,0.02297436,0.049230773,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.04266667,0.08205129,0.0,0.0,0.0,0.0,0.0,0.0,0.18707694,0.45292312,0.60061544,0.56123084,0.40369233,0.24615386,0.2986667,0.41025645,0.47589746,0.446359,0.47589746,0.3446154,0.3052308,0.37743592,0.34789747,0.24615386,0.14769232,0.072205134,0.029538464,0.029538464,0.20348719,0.26912823,0.24615386,0.16738462,0.08861539,0.016410258,0.0,0.0,0.0,0.0,0.0,0.052512825,0.07548718,0.049230773,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.016410258,0.016410258,0.016410258,0.01969231,0.04594872,0.055794876,0.06564103,0.07876924,0.068923086,0.08861539,0.16738462,0.21333335,0.19692309,0.15425642,0.22646156,0.33805132,0.4201026,0.41682056,0.29538465,0.16738462,0.06564103,0.026256412,0.04594872,0.06564103,0.055794876,0.06564103,0.068923086,0.04594872,0.016410258,0.006564103,0.0032820515,0.0032820515,0.0032820515,0.0032820515,0.0,0.0032820515,0.006564103,0.013128206,0.013128206,0.013128206,0.016410258,0.01969231,0.016410258,0.016410258,0.026256412,0.029538464,0.049230773,0.08205129,0.098461546,0.11158975,0.12471796,0.12471796,0.12471796,0.128,0.13456412,0.15097436,0.15753847,0.14112821,0.08861539,0.036102567,0.032820515,0.04594872,0.059076928,0.049230773,0.055794876,0.04266667,0.036102567,0.036102567,0.029538464,0.029538464,0.016410258,0.029538464,0.10502565,0.25271797,0.45620516,0.6465641,0.8533334,1.0962052,1.3850257,1.3718976,1.0929232,1.0043077,1.0535386,0.6826667,0.7975385,1.1749744,1.394872,1.5655385,2.3138463,4.6112823,6.301539,6.5411286,5.408821,3.892513,3.2918978,2.8816411,2.6880002,2.9636924,4.20759,8.477539,7.755488,7.5913854,11.073642,18.819284,19.88595,17.174976,14.27036,13.144616,14.155488,11.697231,7.8736415,5.4908724,5.080616,4.886975,3.882667,4.5456414,8.461129,12.560411,9.133949,8.185436,7.2270775,6.948103,7.762052,9.800206,9.186462,7.9491286,6.616616,5.6385646,5.3891287,6.6002054,7.5585647,7.4010262,6.5247183,6.6067696,11.204924,13.548308,12.189539,10.131693,14.8480015,13.059283,12.704822,11.477334,10.121847,12.445539,13.203693,11.030975,7.1220517,2.9702566,0.380718,0.31507695,0.4397949,0.51856416,0.5677949,0.8566154,1.1520001,1.0338463,0.69579494,0.38728207,0.4135385,0.65969235,1.0896411,1.2898463,1.2077949,1.1323078,0.8402052,0.47589746,0.32164106,0.46933338,0.827077,0.8795898,0.6071795,0.49230772,0.574359,0.44964105,0.3511795,0.48246157,0.5940513,0.57764107,0.47917953,0.4660513,0.46276927,0.6301539,0.9911796,1.4375386,1.332513,1.5261539,2.1103592,2.789744,2.9210258,2.7044106,3.3903592,3.7448208,3.442872,3.0752823,3.0818465,2.9407182,2.6978464,2.5107694,2.6551797,2.7766156,2.8160002,2.789744,2.7044106,2.5665643,2.294154,2.0512822,1.8543591,1.7985642,2.0611284,2.9046156,3.6660516,4.3552823,4.8771286,5.024821,5.1265645,4.9099493,4.699898,4.493129,3.9680004,2.5238976,1.4933335,0.99774367,0.9189744,0.90584624,0.9419488,1.086359,1.204513,1.3292309,1.654154,1.6771283,1.5163078,1.1552821,0.7187693,0.47261542,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.0032820515,0.0,0.0,0.0,0.006564103,0.013128206,0.013128206,0.01969231,0.02297436,0.016410258,0.006564103,0.0,0.0,0.009846155,0.059076928,0.108307704,0.12143591,0.068923086,0.068923086,0.08861539,0.13784617,0.17723078,0.118153855,0.03938462,0.009846155,0.0032820515,0.009846155,0.009846155,0.0032820515,0.0,0.013128206,0.049230773,0.1148718,0.32164106,0.60061544,0.65969235,1.0502565,3.170462,2.3663592,1.2438976,0.47589746,0.20676924,0.07548718,0.118153855,0.14769232,0.14769232,0.15753847,0.27569234,0.37743592,0.3249231,0.3446154,0.7975385,2.172718,1.6705642,1.6016412,1.8838975,2.484513,3.4297438,4.466872,4.0402055,3.817026,4.1517954,4.059898,3.4034874,2.297436,1.2635899,0.571077,0.22646156,0.2855385,0.36430773,0.48902568,0.508718,0.12143591,0.4594872,0.49230772,0.6170257,0.9353847,1.2668719,2.7470772,2.9078977,2.0742567,1.024,0.9714873,1.211077,1.276718,1.339077,1.4342566,1.4769232,1.6607181,2.300718,1.7690258,0.65312827,1.7263591,2.2744617,2.0020514,2.5764105,4.017231,4.6966157,3.3641028,2.4582565,2.3926156,3.0096412,3.5905645,3.2361028,2.409026,1.3095386,0.41682056,0.48246157,1.079795,1.9429746,3.0194874,3.8367183,3.5052311,4.6080003,4.8640003,4.7425647,4.2929235,3.1343591,3.9844105,4.460308,4.210872,3.508513,3.2328207,3.4231799,3.367385,2.0742567,0.23958977,0.23302566,0.12143591,0.16410258,0.36102566,0.5973334,0.6498462,0.764718,0.94523084,0.9353847,0.7253334,0.571077,0.45620516,0.34789747,0.65312827,1.4998976,2.7306669,3.2984617,4.6605134,5.1889234,4.7556925,4.716308,8.034462,6.8004107,4.571898,3.6529233,5.0904617,4.8672824,3.5183592,2.6190772,2.6354873,2.9538465,1.6672822,0.827077,0.4660513,0.37415388,0.09189744,0.01969231,0.0,0.0,0.0,0.0,0.009846155,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.013128206,0.06564103,0.18707694,0.21989745,0.13128206,0.0,0.0,0.02297436,0.03938462,0.029538464,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.059076928,0.101743594,0.2100513,0.30194873,0.13784617,0.3117949,0.27897438,0.24615386,0.35774362,0.69579494,0.9124103,1.0108719,0.9156924,0.6432821,0.28225642,0.068923086,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.072205134,0.2297436,0.19364104,0.0,0.0,0.072205134,0.036102567,0.12471796,0.32820517,0.39056414,0.22646156,0.17723078,0.13128206,0.08533334,0.128,0.17723078,0.17723078,0.13784617,0.068923086,0.0,0.0,0.0,0.013128206,0.02297436,0.0,0.06564103,0.032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016410258,0.032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.09189744,0.22646156,0.29538465,0.318359,0.4201026,0.16738462,0.28882053,0.37743592,0.33476925,0.3511795,0.4266667,0.28882053,0.21333335,0.24943592,0.2231795,0.17723078,0.118153855,0.06564103,0.029538464,0.0,0.07876924,0.11158975,0.13784617,0.14441027,0.0951795,0.07876924,0.029538464,0.0,0.013128206,0.072205134,0.013128206,0.026256412,0.03938462,0.02297436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.006564103,0.006564103,0.016410258,0.01969231,0.026256412,0.04266667,0.06564103,0.06564103,0.052512825,0.108307704,0.190359,0.22646156,0.128,0.13456412,0.14769232,0.18707694,0.21661541,0.15097436,0.07548718,0.032820515,0.016410258,0.029538464,0.068923086,0.059076928,0.052512825,0.04594872,0.036102567,0.006564103,0.009846155,0.009846155,0.009846155,0.009846155,0.009846155,0.0032820515,0.0,0.0032820515,0.006564103,0.016410258,0.006564103,0.006564103,0.013128206,0.02297436,0.016410258,0.01969231,0.02297436,0.03938462,0.07548718,0.101743594,0.11158975,0.108307704,0.10502565,0.108307704,0.128,0.12471796,0.108307704,0.108307704,0.12471796,0.13784617,0.11158975,0.08533334,0.055794876,0.029538464,0.01969231,0.029538464,0.026256412,0.016410258,0.013128206,0.02297436,0.036102567,0.026256412,0.04266667,0.118153855,0.27241027,0.5940513,0.95835906,1.1684103,1.2274873,1.3259488,1.3161026,1.1257436,1.020718,0.9714873,0.6662565,0.7384616,0.9485129,1.3259488,1.8215386,2.3171284,6.0324106,6.5345645,5.5532312,4.266667,3.2853336,3.2229745,3.8596926,4.604718,4.9394875,4.453744,5.970052,7.8441033,9.120821,10.541949,14.532925,12.950975,12.754052,12.09436,11.414975,13.446565,14.211283,9.961026,5.182359,2.3794873,2.048,2.156308,3.876103,7.584821,11.293539,10.650257,12.714667,12.507898,10.725744,8.946873,9.622975,11.759591,9.718155,6.7216415,4.6900516,4.210872,4.7917953,5.835488,6.2687182,6.0619493,6.2227697,8.923898,11.10318,11.825232,11.749744,13.13477,12.343796,13.2562065,11.736616,8.953437,11.398565,11.434668,10.203898,9.005949,7.4830775,3.6332312,1.0305642,0.38728207,0.39056414,0.52512825,1.0962052,1.6410258,1.5753847,1.1191796,0.6235898,0.574359,0.7187693,1.086359,1.7558975,2.6420515,3.498667,2.5435898,1.2898463,0.5874872,0.6629744,1.1388719,1.2800001,1.0272821,0.955077,1.079795,0.8566154,0.69251287,0.6268718,0.60061544,0.55794877,0.46276927,0.571077,0.60389745,0.5907693,0.5907693,0.7187693,0.955077,1.3522053,1.9626669,2.6551797,3.117949,3.1638978,3.9417439,4.1682053,3.820308,4.132103,5.907693,6.7150774,6.5280004,5.684513,4.893539,4.1583595,3.6758976,3.436308,3.3312824,3.1737437,2.8849232,2.537026,2.1431797,1.7755898,1.585231,2.5600002,3.5971284,4.4373336,4.955898,5.172513,5.3005133,5.142975,4.6867695,3.9384618,2.9571285,1.8576412,1.211077,0.9419488,0.9156924,0.93866676,1.014154,1.2373334,1.5130258,1.8412309,2.3236926,2.0578463,1.8642052,1.591795,1.1979488,0.74830776,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.009846155,0.006564103,0.0032820515,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.02297436,0.0032820515,0.0032820515,0.0032820515,0.0,0.0,0.0,0.026256412,0.055794876,0.072205134,0.06564103,0.036102567,0.04266667,0.08861539,0.14769232,0.14441027,0.07548718,0.059076928,0.052512825,0.036102567,0.02297436,0.013128206,0.009846155,0.016410258,0.06564103,0.20020515,0.40697438,0.60061544,0.5940513,0.38400003,0.15425642,0.03938462,0.04266667,0.08205129,0.08861539,0.016410258,0.0032820515,0.006564103,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.13128206,0.8008206,1.529436,2.2547693,3.3312824,3.446154,2.8882053,2.9669745,3.5905645,3.2295387,3.945026,3.9318976,2.7700515,1.020718,0.22646156,0.36758977,0.47261542,0.40697438,0.2100513,0.08533334,0.02297436,0.006564103,0.068923086,0.23302566,0.5415385,2.0217438,2.5206156,2.281026,1.7755898,1.7099489,1.3883078,1.0108719,1.0699488,1.4769232,1.5688206,1.9265642,2.546872,1.9692309,0.8369231,1.9167181,1.9593848,1.1848207,1.5458462,3.1245131,4.128821,3.5446157,3.0391798,2.5304618,1.9987694,1.467077,1.1618463,0.81394875,0.40697438,0.059076928,0.036102567,0.128,0.46933338,0.73517954,1.0436924,1.9298463,3.3509746,3.623385,3.446154,3.1113849,2.5009232,3.639795,4.128821,3.889231,3.2984617,3.1967182,3.495385,3.4231799,2.1103592,0.2986667,0.33476925,0.30851284,0.39712822,0.5415385,0.6695385,0.69251287,0.8041026,0.94523084,1.020718,1.0075898,0.97805136,1.9692309,1.9364104,1.7427694,2.1825643,3.9811285,4.3552823,5.6287184,5.904411,5.0904617,4.9132314,8.129642,7.0465646,4.9526157,3.4658465,2.5271797,1.847795,1.4342566,1.3653334,1.5425643,1.7099489,1.204513,0.65641034,0.23302566,0.026256412,0.06235898,0.013128206,0.0,0.0,0.0,0.006564103,0.009846155,0.06235898,0.08205129,0.04594872,0.013128206,0.10502565,0.28225642,0.45620516,0.5677949,0.60061544,1.0272821,1.8412309,1.723077,0.96492314,1.4572309,2.2580514,2.737231,2.4681027,1.7362052,1.5392822,1.4408206,0.9189744,0.3511795,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.0,0.0032820515,0.0032820515,0.06235898,0.318359,0.2986667,0.16082053,0.068923086,0.10502565,0.2855385,0.892718,1.6508719,2.9210258,3.8071797,2.1333334,1.3850257,0.88287187,0.69579494,0.83035904,1.2438976,1.3751796,1.2307693,0.9517949,0.6465641,0.37743592,0.16738462,0.08205129,0.049230773,0.02297436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.02297436,0.11158975,0.26256412,0.2100513,0.029538464,0.15097436,0.26912823,0.20676924,0.18707694,0.23958977,0.20020515,0.13456412,0.101743594,0.055794876,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08533334,0.15425642,0.16410258,0.108307704,0.14769232,0.06235898,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.04266667,0.21989745,0.072205134,0.20676924,0.28225642,0.23630771,0.28225642,0.38728207,0.3511795,0.28882053,0.23630771,0.15425642,0.12471796,0.11158975,0.118153855,0.13784617,0.17066668,0.12143591,0.04266667,0.036102567,0.09189744,0.101743594,0.11158975,0.04594872,0.013128206,0.049230773,0.1148718,0.02297436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.016410258,0.01969231,0.02297436,0.032820515,0.052512825,0.06564103,0.052512825,0.101743594,0.19364104,0.25271797,0.15753847,0.118153855,0.07548718,0.08861539,0.13456412,0.118153855,0.06564103,0.036102567,0.02297436,0.02297436,0.04594872,0.04266667,0.04594872,0.036102567,0.013128206,0.0,0.006564103,0.013128206,0.016410258,0.013128206,0.009846155,0.0032820515,0.0,0.0,0.0032820515,0.009846155,0.0032820515,0.0,0.013128206,0.029538464,0.02297436,0.02297436,0.013128206,0.026256412,0.055794876,0.08205129,0.098461546,0.09189744,0.08533334,0.08861539,0.098461546,0.09189744,0.068923086,0.08205129,0.17066668,0.35774362,0.38728207,0.24615386,0.0951795,0.016410258,0.0,0.006564103,0.009846155,0.006564103,0.0032820515,0.016410258,0.029538464,0.029538464,0.059076928,0.15425642,0.33805132,0.67610264,0.99774367,1.211077,1.3259488,1.4276924,1.1749744,1.0043077,0.892718,0.7975385,0.65312827,0.67282057,0.77128214,1.1946667,1.8445129,2.2908719,4.841026,4.4373336,3.31159,2.6880002,2.7733335,3.4724104,4.2371287,5.0904617,5.536821,4.5817437,4.6112823,6.8594875,8.100103,7.939283,8.802463,6.810257,7.968821,9.744411,11.467488,14.342566,13.650052,9.363693,5.113436,2.6715899,1.9495386,2.6683078,4.57518,7.643898,10.857026,12.182976,14.293334,14.480412,12.521027,9.4457445,7.5520005,10.308924,8.78277,6.488616,4.9362054,3.6693337,3.9844105,4.276513,4.4832826,4.6178465,4.7392826,5.1298466,6.4557953,8.369231,9.819899,9.045334,8.585847,9.800206,9.288206,7.6996927,9.718155,10.860309,12.212514,12.780309,11.618463,7.834257,2.6978464,0.7778462,0.3249231,0.37743592,0.7844103,1.270154,1.3226668,1.0896411,0.8205129,0.8598975,0.8763078,1.1355898,1.9790771,3.2951798,4.5423594,3.6102567,2.048,0.95835906,0.77456415,1.2668719,1.8051283,1.972513,2.3794873,2.612513,1.2537436,0.9189744,0.65641034,0.5218462,0.48246157,0.43323082,0.574359,0.6498462,0.6695385,0.6498462,0.6301539,0.79097444,1.0010257,1.2964103,1.7066668,2.284308,3.1934361,4.6802053,5.6451287,5.930667,6.3245134,8.228104,9.137232,8.933744,7.893334,6.665847,5.5565133,4.7917953,4.342154,4.092718,3.8465643,3.5413337,3.1606157,2.7109745,2.3105643,2.176,2.9472823,4.0533338,4.923077,5.3234878,5.356308,5.0149746,4.6178465,3.9089234,2.9013336,1.8773335,1.270154,1.0305642,0.97805136,1.0010257,1.0502565,1.1224617,1.3817437,1.7657437,2.2613335,2.9078977,2.6880002,2.409026,2.103795,1.7460514,1.273436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.013128206,0.009846155,0.0,0.0,0.006564103,0.009846155,0.0032820515,0.0032820515,0.0,0.016410258,0.016410258,0.0,0.0,0.0,0.0,0.013128206,0.036102567,0.052512825,0.009846155,0.006564103,0.006564103,0.0,0.0,0.0032820515,0.009846155,0.026256412,0.03938462,0.03938462,0.026256412,0.02297436,0.04266667,0.08533334,0.15425642,0.15753847,0.17394873,0.15425642,0.108307704,0.08861539,0.11158975,0.1148718,0.118153855,0.17066668,0.3708718,0.21989745,0.0951795,0.032820515,0.02297436,0.02297436,0.013128206,0.0032820515,0.0032820515,0.013128206,0.013128206,0.0032820515,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.068923086,0.4004103,1.0108719,1.5983591,1.5491283,3.629949,4.59159,3.442872,1.0305642,0.052512825,0.24615386,0.3314872,0.2855385,0.14769232,0.02297436,0.013128206,0.0032820515,0.0,0.006564103,0.036102567,0.17394873,0.62030774,1.4309745,2.2744617,2.428718,1.7755898,1.0929232,1.017436,1.4867693,1.7165129,2.1267693,2.1924105,1.6082052,0.9714873,1.782154,2.0184617,1.3423591,1.2537436,1.9790771,2.4713848,2.2350771,2.2219489,1.8970258,1.1716924,0.39056414,0.098461546,0.02297436,0.013128206,0.0,0.0,0.049230773,0.14769232,0.34789747,0.8763078,2.1398976,2.1136413,1.6869745,1.1323078,0.63343596,0.29210258,0.63343596,1.3029745,1.6640002,1.5819489,1.4309745,1.214359,0.8041026,0.56123084,0.574359,0.67610264,0.82379496,0.7089231,0.42994875,0.14769232,0.098461546,0.19692309,0.32820517,0.57764107,0.9747693,1.4802053,3.8137438,4.073026,3.2689233,2.7667694,4.276513,4.1911798,5.139693,5.139693,3.7907696,2.2449234,1.2471796,0.97805136,0.955077,1.0962052,1.7394873,1.6475899,1.0075898,0.38728207,0.13784617,0.380718,0.43651286,0.20348719,0.029538464,0.016410258,0.013128206,0.0032820515,0.009846155,0.016410258,0.016410258,0.016410258,0.02297436,0.13128206,0.21333335,0.24615386,0.2986667,0.636718,1.1454359,1.6049232,1.8838975,1.9331284,2.5862565,3.636513,3.2689233,2.284308,4.1156926,6.0061545,6.8594875,5.8486156,3.8334363,3.3280003,3.0982566,1.9626669,0.74830776,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.032820515,0.16738462,0.16738462,0.17723078,0.15753847,0.27897438,0.9353847,1.1454359,0.92225647,0.65312827,0.6695385,1.270154,3.511795,5.85518,7.755488,7.936001,4.388103,2.3729234,1.4145643,1.142154,1.2438976,1.463795,1.4802053,1.3620514,1.1782565,0.955077,0.6662565,0.33476925,0.17394873,0.101743594,0.055794876,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02297436,0.055794876,0.10502565,0.19364104,0.2100513,0.22646156,0.16082053,0.10502565,0.32164106,0.39712822,0.34133336,0.23302566,0.118153855,0.0,0.0,0.0,0.0,0.006564103,0.029538464,0.029538464,0.03938462,0.04594872,0.049230773,0.036102567,0.026256412,0.19364104,0.33805132,0.35446155,0.23630771,0.17723078,0.07876924,0.02297436,0.026256412,0.029538464,0.02297436,0.009846155,0.016410258,0.049230773,0.068923086,0.059076928,0.04266667,0.026256412,0.016410258,0.0,0.07548718,0.049230773,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.059076928,0.0951795,0.13784617,0.190359,0.21989745,0.33805132,0.46276927,0.45292312,0.3052308,0.14441027,0.068923086,0.10502565,0.17066668,0.256,0.42994875,0.3511795,0.18379489,0.072205134,0.06235898,0.08861539,0.08533334,0.049230773,0.052512825,0.098461546,0.12143591,0.02297436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.016410258,0.016410258,0.026256412,0.029538464,0.032820515,0.036102567,0.04594872,0.036102567,0.06235898,0.108307704,0.15753847,0.16082053,0.13456412,0.098461546,0.098461546,0.14769232,0.19692309,0.15097436,0.0951795,0.04594872,0.016410258,0.0032820515,0.009846155,0.04266667,0.03938462,0.0,0.0032820515,0.006564103,0.009846155,0.013128206,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.026256412,0.026256412,0.026256412,0.013128206,0.013128206,0.029538464,0.03938462,0.06235898,0.06564103,0.068923086,0.068923086,0.06235898,0.06235898,0.059076928,0.08533334,0.22646156,0.62030774,0.7581539,0.51856416,0.21989745,0.04266667,0.0032820515,0.0,0.0032820515,0.0032820515,0.0032820515,0.013128206,0.013128206,0.013128206,0.06564103,0.20020515,0.42338464,0.6268718,0.67282057,0.81066674,1.0765129,1.3062565,0.88287187,0.7056411,0.62030774,0.56451285,0.5874872,0.6465641,0.77128214,1.0108719,1.4408206,2.1464617,1.975795,1.7263591,1.6180514,1.7887181,2.294154,3.3017437,3.4100516,3.82359,4.6834874,5.074052,5.674667,5.431795,4.4996924,3.7218463,4.630975,4.4701543,4.886975,8.4053335,14.083283,17.513027,12.1238985,7.9524107,5.691077,4.775385,3.3903592,4.1124105,5.579488,8.759795,12.612924,14.096412,12.763899,12.498053,11.805539,9.829744,6.3606157,6.744616,6.87918,7.5913854,8.234667,6.688821,7.0465646,6.413129,5.737026,5.481026,5.61559,4.663795,4.7491283,5.681231,6.7938466,6.925129,6.498462,6.885744,7.765334,9.009232,10.673231,13.735386,17.447386,18.5239,16.216616,12.35036,4.97559,1.5491283,0.4201026,0.29538465,0.22646156,0.38728207,0.56451285,0.7811283,1.024,1.2340513,1.2077949,1.7394873,2.5928206,3.4166157,3.7415388,3.511795,2.5337439,1.5688206,1.0962052,1.3226668,2.5829747,3.245949,4.1813335,4.6211286,2.1366155,1.3489232,0.80738467,0.5513847,0.5021539,0.46933338,0.51856416,0.5874872,0.65641034,0.7089231,0.69579494,0.7089231,0.67938465,0.67282057,0.80738467,1.2570257,2.930872,4.772103,6.311385,7.1483083,6.9645133,7.253334,7.394462,7.2631803,6.8266673,6.166975,5.805949,5.3891287,4.9985647,4.663795,4.3684106,4.056616,3.7185643,3.4067695,3.2820516,3.626667,3.7809234,4.6539493,5.47118,5.7665644,5.3760004,4.348718,3.4560003,2.6683078,1.9626669,1.3259488,1.142154,1.1126155,1.148718,1.2176411,1.3292309,1.404718,1.9626669,2.733949,3.4822567,4.020513,3.9351797,3.4166157,2.7766156,2.2219489,1.8871796,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.016410258,0.016410258,0.0032820515,0.04594872,0.04594872,0.0,0.0,0.0,0.0,0.013128206,0.026256412,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.013128206,0.016410258,0.016410258,0.016410258,0.016410258,0.0032820515,0.0,0.013128206,0.059076928,0.16738462,0.27897438,0.3052308,0.2855385,0.27241027,0.32164106,0.42994875,0.4955898,0.43323082,0.24943592,0.029538464,0.006564103,0.0,0.0,0.02297436,0.108307704,0.068923086,0.02297436,0.0,0.0,0.0,0.0,0.009846155,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.068923086,0.12471796,0.016410258,0.0032820515,0.04594872,0.059076928,0.02297436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.009846155,0.0,0.0,0.0,0.0,0.0,0.006564103,0.029538464,0.029538464,0.029538464,0.01969231,0.0,0.0,0.013128206,0.508718,1.847795,3.2525132,2.8389745,0.92225647,0.19692309,0.01969231,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.026256412,0.02297436,0.009846155,0.0,0.0,0.63343596,1.9823592,3.442872,4.5062566,4.775385,3.6890259,2.6683078,2.0808206,2.0086155,2.228513,1.9823592,1.0994873,0.33476925,0.02297436,0.06235898,0.26912823,0.18379489,0.14112821,0.80738467,3.190154,3.5807183,3.367385,3.0358977,3.2262566,4.716308,6.1538467,6.294975,7.430565,8.838565,6.774154,3.6857438,1.6508719,0.62030774,0.2855385,0.09189744,0.1148718,0.07548718,0.032820515,0.016410258,0.016410258,0.0032820515,0.036102567,0.072205134,0.072205134,0.0,0.013128206,0.052512825,0.08205129,0.07548718,0.016410258,0.0032820515,0.01969231,0.26256412,0.761436,1.3718976,2.1300514,2.9046156,3.4724104,3.8498464,4.3027697,4.535795,1.9659488,0.41682056,1.7723079,5.9963083,7.680001,7.2861543,4.857436,1.8740515,1.2504616,1.0929232,0.64000005,0.22646156,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.15425642,0.7778462,0.827077,0.8566154,0.75487185,0.764718,1.5097437,2.7437952,3.006359,2.5796926,2.281026,3.4789746,9.216001,13.781334,11.61518,4.585026,1.9823592,1.1290257,1.024,1.2340513,1.4769232,1.6475899,1.6738462,1.5786668,1.4244103,1.2012309,0.82379496,0.34789747,0.09189744,0.01969231,0.036102567,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.118153855,0.28225642,0.47261542,0.71548724,0.65641034,0.5218462,0.3708718,0.2231795,0.07548718,0.016410258,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.029538464,0.15097436,0.15097436,0.190359,0.23302566,0.24287182,0.18379489,0.13456412,0.13128206,0.14441027,0.13784617,0.07548718,0.07548718,0.0951795,0.11158975,0.128,0.15097436,0.1148718,0.04266667,0.08533334,0.23958977,0.3511795,0.30194873,0.20676924,0.13456412,0.08533334,0.0,0.37743592,0.24287182,0.055794876,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.049230773,0.098461546,0.0,0.20676924,0.43323082,0.43323082,0.23958977,0.16738462,0.032820515,0.09189744,0.15097436,0.2100513,0.44307697,0.5284103,0.47589746,0.36758977,0.23630771,0.07548718,0.016410258,0.08205129,0.14441027,0.15753847,0.18379489,0.036102567,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.016410258,0.016410258,0.016410258,0.02297436,0.036102567,0.04594872,0.04594872,0.04594872,0.036102567,0.036102567,0.06564103,0.13784617,0.19692309,0.16738462,0.15425642,0.19692309,0.25928208,0.27241027,0.19364104,0.101743594,0.03938462,0.016410258,0.0032820515,0.009846155,0.009846155,0.0032820515,0.016410258,0.026256412,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.026256412,0.029538464,0.036102567,0.049230773,0.06235898,0.072205134,0.0951795,0.12471796,0.2297436,0.5349744,0.8402052,0.81394875,0.5021539,0.11158975,0.016410258,0.0032820515,0.009846155,0.016410258,0.013128206,0.0,0.0,0.009846155,0.07548718,0.2297436,0.47261542,0.4594872,0.32820517,0.28225642,0.36758977,0.48902568,0.318359,0.32820517,0.38400003,0.45620516,0.6268718,0.7220513,0.95835906,1.0929232,1.1946667,1.6311796,1.8149745,2.0709746,2.2547693,2.172718,1.5885129,1.3915899,2.2416413,4.352,7.0892315,8.956718,7.857231,6.055385,3.9056413,2.2383592,2.3335385,3.5905645,4.8672824,9.396514,16.134565,19.761232,17.024002,12.232206,8.073847,5.586052,4.135385,4.818052,4.7622566,6.12759,9.639385,14.572309,11.191795,11.332924,12.06154,11.766154,10.194052,7.8736415,7.962257,10.056206,12.816411,13.974976,12.291283,12.1468725,11.920411,11.460924,12.084514,7.532308,5.723898,6.189949,8.021334,9.90195,11.9171295,12.547283,11.999181,11.0375395,11.001437,12.051693,15.123693,21.008411,25.242258,18.110361,6.9776416,2.162872,0.67282057,0.446359,0.33476925,0.3117949,0.47917953,0.88287187,1.3292309,1.404718,1.4276924,3.1015387,4.6572313,4.8147697,2.7766156,2.802872,2.8914874,2.7733335,2.3236926,1.5425643,3.5052311,3.895795,4.33559,5.0051284,4.637539,3.186872,1.8806155,1.0371283,0.6892308,0.58092314,0.58092314,0.56123084,0.5546667,0.56123084,0.5481026,0.7089231,0.72861546,0.69907695,0.8533334,1.5885129,2.9669745,4.31918,5.3727183,5.8157954,5.280821,4.082872,3.2262566,2.92759,3.0293336,3.006359,4.2272825,4.6966157,4.818052,4.8311796,4.8049235,4.525949,4.1813335,4.027077,4.089436,4.1517954,3.8071797,4.2994876,4.9952826,5.3169236,4.7294364,3.5938463,2.5862565,2.1366155,2.0808206,1.6771283,1.5425643,1.5556924,1.5753847,1.6114873,1.8313848,2.0512822,3.817026,6.0324106,7.4896417,6.8660517,5.8420515,4.7983594,3.564308,2.422154,2.1070771,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0,0.009846155,0.009846155,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.0032820515,0.0,0.0,0.0032820515,0.013128206,0.013128206,0.0032820515,0.009846155,0.01969231,0.026256412,0.016410258,0.013128206,0.0032820515,0.0032820515,0.02297436,0.0951795,0.34133336,0.5284103,0.69579494,0.86974365,1.0633847,1.1946667,1.0732309,0.77128214,0.41682056,0.17723078,0.12471796,0.04266667,0.0,0.016410258,0.08205129,0.026256412,0.0032820515,0.0,0.0,0.0,0.03938462,0.04266667,0.02297436,0.0032820515,0.013128206,0.013128206,0.0032820515,0.0,0.0,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.026256412,0.0032820515,0.0,0.009846155,0.036102567,0.055794876,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.006564103,0.006564103,0.0032820515,0.0,0.0,0.0032820515,0.101743594,0.3708718,0.6498462,0.5677949,0.18379489,0.03938462,0.0032820515,0.0,0.0,0.0,0.006564103,0.013128206,0.009846155,0.0,0.0,0.013128206,0.052512825,0.15753847,0.39384618,0.7089231,1.1585642,2.3335385,3.6824617,3.515077,1.8937438,3.9089234,5.910975,5.933949,3.7021542,2.284308,1.3095386,0.72861546,0.57764107,0.98133343,1.5195899,1.5031796,1.0765129,0.54482055,0.36758977,0.27241027,0.50543594,1.211077,2.5928206,4.9362054,3.255795,3.5413337,5.4843082,8.03118,9.412924,7.4174366,4.5587697,2.868513,2.5698464,2.0873847,1.4408206,0.75487185,0.318359,0.16082053,0.055794876,0.03938462,0.01969231,0.006564103,0.0032820515,0.0032820515,0.0,0.006564103,0.013128206,0.013128206,0.0,0.013128206,0.04594872,0.049230773,0.036102567,0.06564103,0.11158975,1.6213335,2.284308,2.1858463,3.8038976,5.477744,5.142975,3.6890259,2.1070771,1.4834872,1.1979488,0.49230772,0.101743594,0.37743592,1.2603078,1.6082052,1.5589745,1.0732309,0.44307697,0.2986667,0.23958977,0.13456412,0.04594872,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.055794876,0.27897438,0.24943592,0.2297436,0.2231795,0.36430773,0.9124103,1.6180514,1.6475899,1.214359,0.7384616,0.84348726,1.9987694,3.121231,2.6420515,0.96492314,0.43323082,0.58420515,0.9747693,1.3620514,1.6804104,2.0250258,2.03159,1.6016412,0.9911796,0.446359,0.21333335,0.07876924,0.06235898,0.049230773,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.06235898,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02297436,0.08205129,0.15753847,0.45292312,0.761436,0.86646163,0.7515898,0.5940513,0.80738467,1.079795,0.892718,0.318359,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.08205129,0.14769232,0.14441027,0.029538464,0.098461546,0.17394873,0.22646156,0.30194873,0.52512825,0.4660513,0.27897438,0.15425642,0.14112821,0.15097436,0.12143591,0.12471796,0.15097436,0.17066668,0.1148718,0.07876924,0.029538464,0.016410258,0.049230773,0.08205129,0.06235898,0.04266667,0.026256412,0.016410258,0.0,0.13456412,0.2231795,0.23958977,0.18707694,0.098461546,0.01969231,0.0,0.0,0.0,0.0,0.0,0.0,0.032820515,0.08861539,0.098461546,0.19692309,0.26584616,0.19692309,0.06235898,0.108307704,0.098461546,0.101743594,0.10502565,0.12143591,0.19692309,0.29210258,0.30194873,0.3249231,0.37415388,0.380718,0.19364104,0.19364104,0.20348719,0.17066668,0.14769232,0.029538464,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.016410258,0.016410258,0.009846155,0.013128206,0.02297436,0.02297436,0.02297436,0.026256412,0.026256412,0.02297436,0.026256412,0.03938462,0.032820515,0.049230773,0.07876924,0.052512825,0.15097436,0.17394873,0.118153855,0.036102567,0.052512825,0.07876924,0.06564103,0.03938462,0.032820515,0.06564103,0.04594872,0.016410258,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.013128206,0.006564103,0.0032820515,0.0032820515,0.0032820515,0.0032820515,0.0032820515,0.0032820515,0.006564103,0.016410258,0.016410258,0.01969231,0.013128206,0.013128206,0.036102567,0.049230773,0.055794876,0.101743594,0.21333335,0.4135385,0.571077,0.6498462,0.5677949,0.34789747,0.11158975,0.032820515,0.013128206,0.016410258,0.013128206,0.013128206,0.0032820515,0.0032820515,0.055794876,0.17066668,0.3249231,0.29538465,0.2100513,0.15753847,0.15753847,0.18379489,0.17723078,0.2231795,0.28882053,0.3708718,0.49230772,0.6170257,0.90584624,1.1552821,1.2603078,1.1946667,1.6410258,2.2777438,2.9636924,3.3247182,2.7602053,2.231795,2.858667,4.529231,6.5969234,7.8703594,6.87918,6.186667,4.775385,3.5807183,5.4843082,6.564103,8.625232,11.697231,14.585437,14.841437,12.2617445,10.157949,8.467693,7.2336416,6.6002054,7.0990777,5.156103,4.8738465,7.972103,13.804309,11.096616,12.563693,13.003489,11.208206,9.984001,10.722463,10.518975,10.180923,10.522257,12.36677,15.31077,16.065641,13.797745,10.253129,9.754257,7.181129,5.4383593,6.4754877,10.226872,14.628103,14.785643,12.711386,10.322052,8.845129,8.828718,9.38995,13.111795,18.737232,21.031385,10.774975,6.948103,3.1671798,1.0371283,0.6465641,0.5546667,0.5415385,0.7187693,1.0272821,1.3259488,1.3784616,1.3259488,2.6912823,4.201026,4.8738465,4.0467696,4.9887185,4.8738465,4.1058464,3.0424619,2.0184617,3.2689233,3.5052311,4.128821,5.428513,6.567385,5.85518,4.384821,2.9078977,1.7427694,0.761436,0.55794877,0.45292312,0.40697438,0.4004103,0.4266667,0.63343596,0.7844103,0.8369231,0.85005134,0.97805136,2.2383592,3.2984617,3.7809234,3.6562054,3.2164104,2.605949,2.0939488,1.9495386,2.172718,2.481231,3.1638978,3.367385,3.7185643,4.3290257,4.781949,4.8049235,4.33559,3.817026,3.3936412,2.917744,2.3302567,2.3729234,2.8160002,3.3542566,3.6069746,3.0982566,2.2153847,1.7558975,1.7920002,1.7033848,1.9889232,2.0906668,2.1202054,2.1267693,2.1103592,2.4976413,4.709744,7.709539,9.7903595,8.549745,7.1056414,6.8562055,6.2063594,4.8607183,3.8400004,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.009846155,0.006564103,0.0,0.0,0.0,0.0032820515,0.006564103,0.006564103,0.0,0.0032820515,0.009846155,0.009846155,0.006564103,0.006564103,0.0032820515,0.0,0.009846155,0.049230773,0.24943592,0.571077,0.8795898,1.0535386,0.97805136,1.273436,1.4342566,1.2373334,0.75487185,0.37743592,0.21333335,0.098461546,0.03938462,0.036102567,0.06564103,0.029538464,0.029538464,0.049230773,0.052512825,0.0,0.01969231,0.01969231,0.009846155,0.0,0.006564103,0.01969231,0.052512825,0.08861539,0.101743594,0.06564103,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.026256412,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.026256412,0.04594872,0.055794876,0.06564103,0.072205134,0.08205129,0.08861539,0.2100513,0.67282057,1.2373334,1.7296412,2.4910772,3.242667,3.0949745,2.6584618,3.0884104,3.7185643,3.7218463,2.0873847,1.7591796,1.1454359,0.81066674,1.0075898,1.6869745,2.5600002,3.3050258,3.5544617,3.131077,2.0709746,2.1497438,2.4943593,2.8750772,3.318154,4.089436,4.1189747,4.522667,5.5302567,6.6625648,6.744616,6.518154,5.7534366,4.204308,2.2022567,0.6695385,0.6235898,0.58092314,0.4660513,0.3117949,0.256,0.055794876,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.01969231,0.101743594,0.32164106,0.7220513,0.7122052,0.43323082,0.12471796,0.13128206,0.20676924,1.3522053,2.6322052,3.4330258,3.4494362,3.1573336,2.4451284,1.529436,0.69907695,0.32164106,0.14769232,0.049230773,0.009846155,0.009846155,0.029538464,0.036102567,0.052512825,0.055794876,0.04266667,0.02297436,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01969231,0.098461546,0.108307704,0.101743594,0.098461546,0.15097436,0.36102566,0.71548724,0.81066674,0.574359,0.190359,0.09189744,0.10502565,0.19692309,0.38728207,0.6071795,0.7056411,1.6278975,3.6529233,4.5489235,3.5478978,1.3620514,0.9517949,0.6432821,0.35446155,0.101743594,0.02297436,0.0032820515,0.108307704,0.15425642,0.08861539,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.029538464,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.12471796,0.20348719,0.24943592,0.2855385,0.35446155,0.64000005,0.7581539,0.7318975,0.56123084,0.22646156,0.33805132,0.5152821,0.43651286,0.13784617,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03938462,0.07548718,0.068923086,0.0,0.032820515,0.13456412,0.20676924,0.25271797,0.35446155,0.40369233,0.3708718,0.32820517,0.2986667,0.24943592,0.16082053,0.16082053,0.20348719,0.2100513,0.068923086,0.23958977,0.3052308,0.26584616,0.14769232,0.006564103,0.029538464,0.16410258,0.24287182,0.21661541,0.13784617,0.20348719,0.16082053,0.18379489,0.3249231,0.5152821,0.30194873,0.21333335,0.16410258,0.0951795,0.0,0.0,0.0,0.04594872,0.13456412,0.2231795,0.25271797,0.2297436,0.20676924,0.2297436,0.34789747,0.22646156,0.15425642,0.128,0.14112821,0.19364104,0.26912823,0.28225642,0.34133336,0.4397949,0.4660513,0.32820517,0.29538465,0.25928208,0.18707694,0.13784617,0.026256412,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.009846155,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.006564103,0.006564103,0.016410258,0.026256412,0.032820515,0.032820515,0.052512825,0.055794876,0.03938462,0.026256412,0.006564103,0.0,0.009846155,0.02297436,0.009846155,0.059076928,0.08861539,0.072205134,0.032820515,0.04266667,0.055794876,0.04594872,0.032820515,0.032820515,0.03938462,0.029538464,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.006564103,0.0032820515,0.0,0.0,0.0,0.0,0.006564103,0.006564103,0.0,0.006564103,0.006564103,0.013128206,0.016410258,0.02297436,0.03938462,0.04594872,0.052512825,0.08861539,0.17723078,0.3249231,0.56451285,0.6432821,0.6859488,0.6301539,0.2297436,0.059076928,0.016410258,0.013128206,0.006564103,0.006564103,0.009846155,0.013128206,0.059076928,0.14441027,0.22646156,0.2100513,0.16082053,0.108307704,0.07876924,0.07876924,0.13128206,0.190359,0.25271797,0.32164106,0.39384618,0.46933338,0.67610264,0.98461545,1.3128207,1.5491283,1.5786668,1.8412309,2.2088206,2.3893335,1.9167181,1.6738462,3.442872,5.477744,6.695385,6.6822567,6.5312824,7.1122055,7.00718,6.045539,5.284103,6.055385,7.240206,8.73354,10.843898,14.280207,11.608616,11.408411,11.0145645,9.360411,6.9710774,6.0160003,4.3060517,3.6791797,5.1659493,8.979693,9.705027,11.552821,12.685129,12.324103,10.758565,10.04636,9.242257,8.582564,8.395488,9.107693,13.170873,16.036104,15.448617,12.018872,9.216001,7.3091288,5.8945646,5.8847184,7.394462,9.7214365,9.189744,7.276308,5.47118,4.5489235,4.588308,7.076103,11.953232,17.293129,20.22072,16.94195,13.387488,7.857231,3.2918978,1.020718,0.764718,0.8795898,1.0994873,1.4408206,2.1103592,3.5052311,2.540308,2.3663592,3.2853336,5.175795,7.4765134,9.511385,9.613129,8.060719,5.7435904,4.1517954,5.100308,5.044513,5.041231,5.612308,6.7282057,7.13518,6.557539,5.920821,5.3792825,4.315898,2.294154,1.0272821,0.49230772,0.47261542,0.56123084,0.6629744,0.7417436,0.83035904,0.8960001,0.84348726,1.3357949,2.2514873,2.8980515,2.9768207,2.5895386,2.5009232,2.7602053,3.0162053,3.1671798,3.367385,3.7382567,3.7710772,3.9581542,4.4045134,4.8311796,4.854154,4.263385,3.4592824,2.7076926,2.1333334,1.8609232,1.8871796,2.1858463,2.6880002,3.2886157,3.0752823,2.28759,1.8806155,2.038154,2.1956925,2.6518977,2.9801028,3.1671798,3.2361028,3.242667,4.204308,6.8004107,9.668923,11.296822,10.016821,8.684308,8.004924,7.6996927,7.1515903,5.398975,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.009846155,0.009846155,0.006564103,0.006564103,0.006564103,0.013128206,0.026256412,0.029538464,0.009846155,0.0032820515,0.0,0.0,0.006564103,0.0,0.009846155,0.013128206,0.009846155,0.01969231,0.12471796,0.39056414,0.69251287,0.8992821,0.8730257,1.0404103,1.2635899,1.2307693,0.92553854,0.6301539,0.48902568,0.40369233,0.318359,0.22646156,0.17066668,0.15097436,0.17723078,0.2231795,0.23302566,0.108307704,0.026256412,0.006564103,0.009846155,0.009846155,0.0,0.059076928,0.118153855,0.14441027,0.12471796,0.068923086,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02297436,0.03938462,0.049230773,0.06564103,0.072205134,0.07548718,0.072205134,0.14441027,0.48902568,0.9419488,1.3883078,1.7788719,2.0644104,2.2088206,2.9768207,2.4549747,2.284308,2.5731285,1.8871796,2.1825643,1.9265642,1.913436,2.4418464,3.318154,3.3641028,3.4756925,3.620103,3.501949,2.5862565,2.556718,2.8422565,3.0260515,3.0490258,3.2295387,3.6627696,3.69559,3.5446157,3.2754874,2.789744,3.6627696,4.312616,3.7087183,1.9856411,0.43651286,0.35774362,0.43323082,0.44307697,0.34133336,0.256,0.052512825,0.0,0.0,0.0,0.0,0.0,0.0,0.01969231,0.128,0.45620516,1.3817437,2.1267693,2.1464617,1.4998976,0.85005134,1.7755898,1.8313848,2.1398976,2.5632823,1.6836925,0.6301539,0.16410258,0.029538464,0.029538464,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.036102567,0.072205134,0.08205129,0.08533334,0.09189744,0.128,0.26584616,0.35446155,0.2855385,0.17066668,0.3117949,0.34789747,0.43323082,0.83035904,1.4572309,1.8707694,3.18359,4.640821,4.6276927,2.8816411,0.512,0.101743594,0.02297436,0.04266667,0.04266667,0.0,0.0,0.08861539,0.13128206,0.0951795,0.029538464,0.006564103,0.0,0.013128206,0.02297436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.029538464,0.049230773,0.032820515,0.0,0.0,0.12471796,0.318359,0.38728207,0.33476925,0.35446155,0.42994875,0.38728207,0.3249231,0.23302566,0.0,0.0,0.026256412,0.026256412,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06564103,0.15097436,0.23302566,0.3052308,0.446359,0.50543594,0.6104616,0.69907695,0.4955898,0.3446154,0.27897438,0.27241027,0.2855385,0.25928208,0.41682056,0.47261542,0.4135385,0.26912823,0.12143591,0.19692309,0.3446154,0.4135385,0.36102566,0.24615386,0.3314872,0.14112821,0.098461546,0.318359,0.60061544,0.5284103,0.44964105,0.34789747,0.2231795,0.108307704,0.02297436,0.0,0.04266667,0.12143591,0.17394873,0.17394873,0.14112821,0.20676924,0.3446154,0.38400003,0.3511795,0.3249231,0.2855385,0.25928208,0.30194873,0.37415388,0.43323082,0.48574364,0.5316923,0.5513847,0.5677949,0.49230772,0.34133336,0.17394873,0.08205129,0.016410258,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.013128206,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.013128206,0.02297436,0.032820515,0.032820515,0.052512825,0.06235898,0.055794876,0.052512825,0.026256412,0.009846155,0.0032820515,0.0032820515,0.016410258,0.016410258,0.026256412,0.029538464,0.026256412,0.029538464,0.029538464,0.016410258,0.013128206,0.016410258,0.016410258,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.009846155,0.0,0.0,0.0032820515,0.006564103,0.016410258,0.026256412,0.026256412,0.032820515,0.03938462,0.06564103,0.13128206,0.23958977,0.48902568,0.5874872,0.6629744,0.636718,0.23630771,0.06564103,0.013128206,0.006564103,0.0,0.0,0.006564103,0.026256412,0.068923086,0.12471796,0.15097436,0.15753847,0.13784617,0.098461546,0.06564103,0.06235898,0.14112821,0.19692309,0.23630771,0.26584616,0.29538465,0.3314872,0.44964105,0.8369231,1.4605129,2.0644104,1.9495386,1.9593848,1.8674873,1.5589745,1.0010257,1.1191796,3.6430771,6.226052,7.3321033,6.232616,6.4656415,8.116513,9.252103,8.625232,5.674667,4.9099493,4.886975,5.5269747,7.499488,12.228924,10.801231,11.894155,11.58236,8.736821,5.028103,3.751385,4.2371287,5.6418467,6.8988724,6.7314878,8.874667,12.251899,15.02195,15.622565,12.777026,13.203693,10.955488,8.960001,8.237949,7.8802056,9.957745,12.829539,13.538463,11.825232,10.125129,8.15918,7.1548724,5.979898,5.5532312,8.822155,6.8594875,6.7282057,6.488616,5.8978467,6.409847,9.081436,10.660104,13.423591,17.316103,19.948309,14.585437,9.094564,4.706462,2.1070771,1.4441026,1.3029745,2.041436,2.7273848,3.2262566,4.2272825,3.4789746,2.9210258,3.5905645,5.9995904,10.138257,11.08677,10.689642,9.554052,7.8014364,5.0904617,4.965744,5.546667,5.920821,5.835488,5.7042055,6.5837955,7.3714876,8.188719,8.73354,8.28718,4.7622566,2.2219489,0.9616411,0.7417436,0.8041026,0.761436,0.7253334,0.76800007,0.8533334,0.8533334,0.86317956,1.5163078,2.3663592,2.9669745,2.865231,3.0916924,3.639795,3.9253337,3.8596926,3.8531284,3.9680004,3.9089234,3.882667,3.9876926,4.1911798,3.9942567,3.3903592,2.7175386,2.1792822,1.8576412,1.9068719,1.9954873,2.231795,2.6190772,3.0523078,2.8717952,2.3269746,2.0841026,2.3040001,2.6453335,3.0523078,3.3903592,3.820308,4.352,4.8672824,6.117744,8.674462,10.978462,11.992617,11.188514,10.341744,9.632821,9.517949,9.435898,7.834257,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.016410258,0.0032820515,0.013128206,0.01969231,0.026256412,0.03938462,0.055794876,0.06564103,0.026256412,0.009846155,0.0032820515,0.006564103,0.02297436,0.006564103,0.026256412,0.029538464,0.009846155,0.0,0.04266667,0.12471796,0.33476925,0.6662565,1.0043077,0.8172308,0.7515898,0.77456415,0.8172308,0.79425645,0.7975385,0.764718,0.69251287,0.571077,0.38400003,0.318359,0.3314872,0.37743592,0.38400003,0.23302566,0.06235898,0.016410258,0.016410258,0.01969231,0.0,0.08861539,0.13128206,0.11158975,0.052512825,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.013128206,0.016410258,0.006564103,0.009846155,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0032820515,0.016410258,0.14769232,0.21333335,0.16738462,0.13456412,0.39384618,0.7581539,1.2340513,1.8149745,2.4648206,3.170462,3.05559,3.1671798,3.5610259,3.2853336,3.3378465,3.2984617,3.2754874,3.5511796,4.588308,3.3641028,2.2580514,1.8018463,1.913436,1.8904617,1.529436,1.4145643,1.529436,1.8937438,2.5764105,1.6311796,1.2274873,0.9189744,0.61374366,0.56123084,0.48574364,0.4266667,0.39712822,0.36758977,0.26912823,0.17066668,0.12471796,0.14441027,0.16410258,0.036102567,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.052512825,0.26912823,1.3850257,3.0030773,3.6726158,3.0030773,1.6672822,3.3280003,2.5993848,1.2471796,0.29210258,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.01969231,0.04266667,0.08861539,0.15097436,0.18051283,0.13456412,0.128,0.2855385,0.7450257,0.9156924,1.086359,1.3817437,1.8412309,2.4155898,3.5052311,2.7798977,1.3029745,0.072205134,0.0,0.0,0.04266667,0.108307704,0.128,0.0,0.0,0.009846155,0.032820515,0.06564103,0.108307704,0.049230773,0.029538464,0.03938462,0.049230773,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.059076928,0.0951795,0.06564103,0.0,0.0,0.0,0.22646156,0.2986667,0.17723078,0.15753847,0.032820515,0.0,0.0,0.009846155,0.052512825,0.026256412,0.006564103,0.013128206,0.03938462,0.059076928,0.21989745,0.10502565,0.009846155,0.032820515,0.07548718,0.04266667,0.013128206,0.0,0.0,0.0,0.0,0.006564103,0.07548718,0.2231795,0.4397949,0.6104616,0.574359,0.7384616,1.0043077,0.7778462,0.6071795,0.39384618,0.31507695,0.4135385,0.5874872,0.52512825,0.49887183,0.46276927,0.40697438,0.3708718,0.46933338,0.44964105,0.38728207,0.32820517,0.28225642,0.39712822,0.17066668,0.08533334,0.24287182,0.3511795,0.5349744,0.51856416,0.39384618,0.26256412,0.23958977,0.049230773,0.026256412,0.068923086,0.08205129,0.0,0.0,0.013128206,0.13784617,0.29210258,0.20020515,0.4135385,0.512,0.4955898,0.43323082,0.4660513,0.5546667,0.67282057,0.7220513,0.69907695,0.67938465,0.77128214,0.6301539,0.36758977,0.108307704,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.006564103,0.02297436,0.016410258,0.01969231,0.032820515,0.049230773,0.06235898,0.04594872,0.026256412,0.009846155,0.0032820515,0.016410258,0.01969231,0.02297436,0.029538464,0.03938462,0.04594872,0.036102567,0.016410258,0.0032820515,0.0032820515,0.013128206,0.006564103,0.006564103,0.0032820515,0.0032820515,0.0,0.0,0.009846155,0.013128206,0.009846155,0.0,0.0032820515,0.0032820515,0.0032820515,0.0,0.0,0.0,0.006564103,0.006564103,0.0,0.0,0.009846155,0.0032820515,0.006564103,0.013128206,0.006564103,0.009846155,0.013128206,0.036102567,0.08861539,0.15753847,0.30851284,0.47589746,0.5546667,0.47589746,0.20676924,0.08205129,0.02297436,0.006564103,0.0032820515,0.0,0.0,0.02297436,0.059076928,0.09189744,0.101743594,0.118153855,0.12471796,0.11158975,0.08533334,0.072205134,0.16738462,0.21661541,0.2297436,0.21661541,0.2100513,0.23630771,0.318359,0.82379496,1.719795,2.5764105,2.8455386,3.0687182,2.737231,1.8346668,0.83035904,1.0994873,3.4888208,6.2129235,7.5979495,6.0750775,6.196513,8.375795,10.269539,10.325335,7.8014364,5.5565133,4.634257,4.7458467,5.8256416,8.021334,8.789334,10.400822,9.590155,6.1341543,2.865231,2.5140514,4.7950773,8.914052,12.1468725,9.8363085,10.240001,14.723283,18.20554,18.034874,13.984821,17.34236,14.907078,11.687386,9.82318,8.602257,8.303591,9.301334,9.373539,8.766359,10.187488,8.251078,7.6964107,6.619898,6.5969234,12.681848,10.223591,12.465232,13.328411,11.759591,11.703795,11.920411,8.507077,8.339693,12.245335,15.02195,9.396514,6.449231,4.8147697,3.6332312,2.5271797,2.1070771,3.4330258,4.44718,4.31918,3.4756925,4.5029745,4.903385,5.6943593,7.5881033,10.985026,9.517949,8.041026,8.077128,8.41518,5.1331286,4.210872,5.979898,7.2336416,6.6494365,4.7622566,5.408821,7.709539,9.481847,10.404103,12.012309,7.0498466,3.3903592,1.463795,0.98133343,0.93866676,0.81394875,0.73517954,0.7122052,0.74830776,0.8598975,0.9124103,1.1749744,1.9200002,2.8521028,3.1113849,3.446154,3.761231,3.817026,3.6430771,3.5282054,3.3969233,3.2918978,3.1737437,3.0752823,3.1113849,2.7306669,2.228513,1.9429746,1.9495386,2.0644104,2.1530259,2.231795,2.477949,2.7864618,2.7864618,2.5895386,2.3893335,2.3860514,2.665026,3.1967182,3.4789746,3.5872824,4.164923,5.2676926,6.3507695,7.2894363,9.304616,11.053949,11.910565,11.926975,11.736616,11.680821,11.654565,11.477334,10.883283,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.07876924,0.07876924,0.013128206,0.0,0.036102567,0.06564103,0.059076928,0.026256412,0.016410258,0.026256412,0.02297436,0.016410258,0.02297436,0.04594872,0.02297436,0.02297436,0.01969231,0.0,0.0,0.02297436,0.0951795,0.36430773,0.77128214,1.0535386,0.8467693,0.60061544,0.49230772,0.53825647,0.6104616,0.6235898,0.54482055,0.67282057,0.8730257,0.58092314,0.2986667,0.19364104,0.13784617,0.08533334,0.06235898,0.049230773,0.01969231,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.032820515,0.06564103,0.07548718,0.026256412,0.04266667,0.036102567,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.009846155,0.0032820515,0.016410258,0.07548718,0.7056411,0.9747693,0.7187693,0.5481026,1.404718,1.4342566,1.6475899,2.4418464,3.6004105,3.8564105,4.0303593,4.06318,4.141949,4.716308,4.7261543,4.8049235,3.7776413,2.5271797,3.9680004,3.1606157,3.170462,3.31159,3.1573336,2.546872,2.5107694,1.2406155,0.24287182,0.013128206,0.0,0.013128206,0.052512825,0.052512825,0.013128206,0.0,0.06235898,0.059076928,0.026256412,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.256,0.67610264,1.0502565,1.1651284,0.82379496,0.39712822,0.13456412,0.01969231,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.026256412,0.02297436,0.032820515,0.20676924,0.79425645,1.3554872,1.2570257,0.8795898,0.48574364,0.2297436,0.16738462,0.18051283,0.17394873,0.108307704,0.0,0.0,0.0,0.10502565,0.20676924,0.0,0.0,0.055794876,0.16410258,0.26912823,0.24287182,0.18379489,0.14112821,0.072205134,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.049230773,0.02297436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.052512825,0.25928208,0.12471796,0.036102567,0.06564103,0.19364104,0.28882053,1.0962052,0.51856416,0.04266667,0.16082053,0.380718,0.2100513,0.06564103,0.0,0.0,0.0,0.0,0.026256412,0.026256412,0.049230773,0.24287182,0.4135385,0.28225642,0.24615386,0.44964105,0.7778462,0.7056411,0.27569234,0.22646156,0.57764107,0.6268718,0.5513847,0.7089231,0.8369231,0.81066674,0.64000005,0.6892308,0.446359,0.23302566,0.19692309,0.32164106,0.39384618,0.16410258,0.14112821,0.36430773,0.4135385,0.30194873,0.21989745,0.108307704,0.01969231,0.09189744,0.01969231,0.13784617,0.24615386,0.21989745,0.0,0.0,0.06564103,0.15425642,0.23958977,0.27569234,0.36102566,0.46276927,0.52512825,0.56451285,0.6859488,0.7844103,0.80738467,0.88943595,0.9485129,0.7187693,0.48574364,0.30851284,0.13784617,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.016410258,0.02297436,0.04594872,0.02297436,0.006564103,0.01969231,0.049230773,0.06235898,0.036102567,0.02297436,0.009846155,0.0032820515,0.016410258,0.03938462,0.055794876,0.08533334,0.118153855,0.108307704,0.059076928,0.026256412,0.009846155,0.0,0.0,0.02297436,0.029538464,0.02297436,0.013128206,0.0,0.0,0.009846155,0.009846155,0.0,0.0,0.013128206,0.016410258,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.01969231,0.029538464,0.006564103,0.009846155,0.026256412,0.06235898,0.12143591,0.28225642,0.4955898,0.67282057,0.69579494,0.4266667,0.19692309,0.072205134,0.029538464,0.02297436,0.0,0.0,0.0,0.013128206,0.03938462,0.07548718,0.11158975,0.14112821,0.14769232,0.13456412,0.12143591,0.15753847,0.2231795,0.25271797,0.23630771,0.19692309,0.18707694,0.30194873,0.8992821,2.0250258,3.4166157,4.125539,4.8344617,4.522667,3.0391798,1.0994873,1.270154,3.4002054,5.287385,5.720616,4.5029745,5.100308,6.961231,8.950154,10.180923,10.010257,10.020103,8.43159,6.698667,5.786257,6.163693,7.716103,8.569437,8.001641,6.3212314,4.8672824,4.525949,3.6168208,6.705231,13.167591,17.194668,15.218873,15.136822,14.70359,12.908309,9.980719,9.380103,12.757335,13.768207,10.896411,7.430565,9.409642,10.423796,8.930462,5.9634876,5.159385,4.3651285,4.394667,5.943795,8.264206,9.156924,12.389745,16.777847,16.833643,12.09436,7.125334,4.637539,5.074052,7.722667,10.371283,9.3078985,7.269744,6.2194877,5.425231,4.5029745,3.4166157,3.9056413,4.630975,5.1265645,5.149539,4.6834874,7.9195905,8.598975,9.088,10.131693,10.86359,9.728001,7.962257,7.712821,8.598975,7.719385,9.563898,11.260718,11.090053,8.851693,5.874872,6.4590774,10.341744,11.227899,10.473026,17.089642,8.349539,3.2984617,1.1552821,0.7811283,0.67282057,0.63343596,0.6432821,0.6859488,0.761436,0.88615394,1.0436924,1.0568206,1.3620514,1.8806155,2.0151796,2.3696413,2.7602053,3.1606157,3.442872,3.3575387,3.0884104,2.9669745,2.8324106,2.7208207,2.868513,2.7602053,2.3466668,2.0644104,2.1530259,2.6387694,2.4451284,2.5337439,2.8488207,3.1540515,3.006359,3.1048207,3.0654361,3.2361028,3.7710772,4.637539,4.969026,4.903385,5.284103,6.1538467,6.7905645,6.8988724,8.054154,9.659078,11.155693,12.025436,12.452104,12.612924,12.626052,12.665437,12.970668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.016410258,0.0032820515,0.0,0.006564103,0.013128206,0.013128206,0.006564103,0.016410258,0.04594872,0.059076928,0.049230773,0.02297436,0.009846155,0.0032820515,0.0032820515,0.009846155,0.013128206,0.02297436,0.068923086,0.15097436,0.3446154,0.6498462,0.97805136,0.77128214,0.47589746,0.3117949,0.3314872,0.4135385,0.43651286,0.4201026,0.44964105,0.50543594,0.45620516,0.71548724,0.49887183,0.24943592,0.13128206,0.049230773,0.026256412,0.016410258,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.04266667,0.09189744,0.11158975,0.14112821,0.41025645,0.6695385,0.67282057,0.18379489,0.04594872,0.0032820515,0.0,0.0032820515,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.009846155,0.006564103,0.02297436,0.098461546,0.29538465,0.80738467,1.4900514,1.4309745,0.69907695,0.35446155,0.94523084,0.74830776,0.6235898,0.9682052,1.7099489,3.4691284,5.835488,7.7325134,8.39877,7.4010262,7.637334,5.097026,2.678154,1.654154,1.6607181,1.148718,1.0108719,0.9616411,0.8336411,0.58420515,0.5284103,0.25928208,0.06235898,0.013128206,0.0,0.0032820515,0.009846155,0.009846155,0.0032820515,0.0,0.013128206,0.013128206,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06235898,0.14112821,0.2100513,0.23302566,0.16410258,0.07876924,0.026256412,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.0032820515,0.006564103,0.04266667,0.15753847,0.27241027,0.28882053,0.3052308,0.35446155,0.4135385,0.30194873,0.13456412,0.036102567,0.02297436,0.0,0.0,0.06564103,0.23958977,0.3446154,0.0,0.26256412,0.36102566,0.3511795,0.27897438,0.19692309,0.25271797,0.3117949,0.24943592,0.08861539,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.06235898,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.052512825,0.026256412,0.006564103,0.013128206,0.03938462,0.059076928,0.21989745,0.10502565,0.009846155,0.032820515,0.07548718,0.04266667,0.013128206,0.0,0.013128206,0.072205134,0.16082053,0.07876924,0.006564103,0.009846155,0.049230773,0.08205129,0.055794876,0.068923086,0.14769232,0.25271797,0.21989745,0.08533334,0.19692309,0.67610264,1.4178462,0.8369231,1.211077,1.2504616,0.7253334,0.45620516,0.42994875,0.43651286,0.39384618,0.26584616,0.06564103,0.22646156,0.21661541,0.23958977,0.3314872,0.3511795,0.54482055,0.45620516,0.21989745,0.052512825,0.26256412,0.26584616,0.13456412,0.049230773,0.04266667,0.0,0.15753847,0.17723078,0.2231795,0.3511795,0.5546667,0.5349744,0.5152821,0.61374366,0.8205129,0.9911796,1.020718,1.0568206,1.0699488,0.97805136,0.6695385,0.48574364,0.26912823,0.118153855,0.055794876,0.036102567,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.006564103,0.02297436,0.026256412,0.01969231,0.029538464,0.06235898,0.08533334,0.072205134,0.04266667,0.026256412,0.029538464,0.052512825,0.07548718,0.098461546,0.12471796,0.13456412,0.0951795,0.04594872,0.029538464,0.02297436,0.013128206,0.02297436,0.029538464,0.02297436,0.016410258,0.013128206,0.013128206,0.072205134,0.059076928,0.032820515,0.02297436,0.013128206,0.013128206,0.016410258,0.013128206,0.013128206,0.013128206,0.0032820515,0.006564103,0.006564103,0.0,0.0,0.009846155,0.013128206,0.013128206,0.013128206,0.006564103,0.0,0.009846155,0.016410258,0.032820515,0.08533334,0.16738462,0.26584616,0.50543594,0.7450257,0.574359,0.27241027,0.128,0.068923086,0.04594872,0.013128206,0.0032820515,0.0,0.0032820515,0.013128206,0.03938462,0.06564103,0.1148718,0.16738462,0.21989745,0.256,0.20348719,0.20348719,0.21989745,0.22646156,0.19692309,0.19692309,0.48902568,1.2603078,2.349949,3.2722054,3.6168208,3.9876926,3.1540515,1.4703591,0.86646163,1.3489232,3.5807183,5.402257,5.8814363,5.293949,6.3901544,7.8408213,8.723693,9.16677,10.364718,12.22236,11.592206,9.360411,7.240206,7.77518,12.041847,13.633642,12.104206,8.4972315,5.356308,6.0685134,5.6352825,5.3366156,7.64718,16.256,12.422565,14.7331295,15.126975,11.444513,7.4404106,5.290667,6.3212314,7.680001,7.79159,6.3442054,7.532308,7.6110773,7.6570263,8.444718,10.443488,8.809027,9.977437,10.7158985,10.41395,11.07036,11.884309,11.155693,9.3078985,7.24677,6.370462,9.875693,16.57436,18.714258,14.821745,9.6984625,8.050873,8.241231,8.136206,7.2205133,6.5903597,6.3474874,6.892308,7.4240007,6.885744,3.95159,4.6572313,5.0642056,6.6133337,8.490667,7.640616,7.250052,7.0498466,9.019077,12.058257,12.028719,10.269539,8.802463,7.2894363,6.0291286,5.9602056,8.041026,10.656821,10.925949,9.147078,8.802463,6.1440005,3.9909747,2.6256413,1.8740515,1.1093334,0.69251287,0.6662565,0.761436,0.8402052,0.88615394,1.1323078,1.2406155,1.2800001,1.2898463,1.2570257,1.2800001,1.339077,1.6147693,2.1333334,2.7700515,3.1967182,3.2918978,3.190154,3.0326157,2.9538465,2.7963078,2.6584618,2.4484105,2.2547693,2.3236926,2.4385643,2.5698464,2.7109745,2.8389745,2.8947694,3.4527183,4.2305646,5.4482055,6.87918,7.8736415,6.7577443,6.38359,6.616616,7.0334363,6.925129,6.5280004,7.1581545,8.661334,10.5780525,12.156719,12.908309,13.193847,13.088821,12.800001,12.665437,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.029538464,0.036102567,0.029538464,0.036102567,0.128,0.055794876,0.04266667,0.06564103,0.0951795,0.08533334,0.14112821,0.256,0.40697438,0.56451285,0.6859488,0.6104616,0.36758977,0.2231795,0.256,0.35774362,0.29210258,0.256,0.23958977,0.24287182,0.2986667,0.571077,0.5152821,0.36430773,0.2297436,0.108307704,0.032820515,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.009846155,0.006564103,0.0,0.0,0.0,0.04266667,0.068923086,0.06235898,0.049230773,0.098461546,0.29210258,0.7975385,1.4244103,1.6475899,0.53825647,0.10502565,0.0,0.0,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.016410258,0.052512825,0.072205134,0.006564103,0.0,0.0,0.006564103,0.029538464,0.072205134,0.04266667,0.013128206,0.009846155,0.049230773,0.14769232,0.39712822,0.6892308,0.67938465,0.36758977,0.12143591,0.36758977,0.512,0.92553854,1.4145643,1.2438976,1.7099489,2.7634873,3.820308,4.3684106,3.9876926,3.820308,2.2908719,1.0272821,0.58092314,0.43323082,0.26584616,0.190359,0.15097436,0.108307704,0.036102567,0.013128206,0.006564103,0.006564103,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01969231,0.068923086,0.14112821,0.20020515,0.26256412,0.30851284,0.27897438,0.16082053,0.0,0.0,0.2855385,0.47261542,0.42994875,0.29210258,0.48246157,0.32164106,0.15753847,0.19692309,0.5021539,0.3314872,0.24287182,0.2297436,0.20348719,0.0,0.0,0.0,0.029538464,0.118153855,0.29210258,0.24943592,0.13456412,0.03938462,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016410258,0.055794876,0.098461546,0.08205129,0.016410258,0.27897438,0.27897438,0.006564103,0.029538464,0.108307704,0.052512825,0.0,0.006564103,0.036102567,0.04266667,0.03938462,0.036102567,0.036102567,0.036102567,0.006564103,0.0,0.0,0.0,0.0,0.0,0.009846155,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.108307704,0.14441027,0.08861539,0.108307704,0.29210258,0.318359,0.28882053,0.24943592,0.19364104,0.12471796,0.072205134,0.036102567,0.04266667,0.12143591,0.052512825,0.013128206,0.07548718,0.28225642,0.6465641,0.36430773,0.57764107,0.6104616,0.33476925,0.16410258,0.14441027,0.17394873,0.17394873,0.11158975,0.0,0.101743594,0.3052308,0.3708718,0.31507695,0.4004103,0.5940513,0.508718,0.37415388,0.3708718,0.65312827,0.5316923,0.46933338,0.318359,0.118153855,0.118153855,0.2855385,0.37743592,0.45292312,0.56123084,0.75487185,0.77128214,0.78769237,0.90256417,1.079795,1.1585642,1.0994873,1.0371283,0.9156924,0.7122052,0.46276927,0.3446154,0.19692309,0.08205129,0.029538464,0.01969231,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.016410258,0.016410258,0.01969231,0.029538464,0.04594872,0.06564103,0.08205129,0.06235898,0.052512825,0.059076928,0.07876924,0.08861539,0.09189744,0.108307704,0.1148718,0.0951795,0.04594872,0.01969231,0.016410258,0.02297436,0.026256412,0.029538464,0.02297436,0.016410258,0.016410258,0.016410258,0.016410258,0.04594872,0.036102567,0.026256412,0.01969231,0.016410258,0.02297436,0.02297436,0.01969231,0.016410258,0.016410258,0.009846155,0.013128206,0.009846155,0.0032820515,0.009846155,0.013128206,0.016410258,0.016410258,0.013128206,0.0,0.0,0.009846155,0.01969231,0.029538464,0.049230773,0.08861539,0.256,0.5546667,0.74830776,0.380718,0.26256412,0.13784617,0.06564103,0.04594872,0.016410258,0.0032820515,0.0,0.0,0.0032820515,0.013128206,0.029538464,0.06235898,0.12143591,0.20020515,0.26256412,0.23958977,0.19692309,0.18707694,0.20676924,0.190359,0.20348719,0.4594872,0.92553854,1.4408206,1.7066668,1.7132308,1.8248206,1.3653334,0.5481026,0.46933338,1.148718,3.5314875,5.1298466,5.2020516,4.7622566,5.5269747,6.0258465,6.170257,6.436103,7.8802056,8.5891285,7.9261546,8.093539,9.921641,12.875488,13.863386,14.168616,12.544001,9.350565,6.547693,8.608821,8.726975,6.6133337,5.618872,12.698257,13.075693,11.585642,9.885539,8.602257,7.3452315,6.058667,5.970052,6.2490263,6.301539,5.7698464,7.1909747,8.3134365,8.917334,9.209436,9.842873,10.919386,13.692719,13.912617,11.59877,11.011283,8.67118,5.970052,4.073026,3.6857438,5.0543594,9.156924,13.699283,15.228719,13.666463,12.294565,9.449026,9.521232,10.886565,11.83836,10.571488,8.854975,7.9491286,7.6209235,7.325539,6.2030773,6.2129235,7.141744,8.086975,8.274052,7.066257,6.616616,6.554257,7.6012316,9.334154,10.167795,12.465232,12.3766165,9.380103,5.6385646,5.979898,8.631796,14.319591,18.231796,17.040411,8.881231,8.395488,8.362667,7.1647186,4.647385,2.100513,1.4112822,1.2537436,1.1979488,1.083077,1.014154,1.2832822,1.4998976,1.5327181,1.3981539,1.2964103,1.1913847,1.1355898,1.2209232,1.4736412,1.8379488,2.281026,2.7109745,2.986667,3.0785644,3.0752823,3.0358977,3.0720003,3.131077,3.1048207,2.809436,2.6978464,2.930872,3.2918978,3.6562054,3.9942567,5.0116925,6.1997952,7.837539,9.544206,10.276103,8.621949,7.5454364,7.197539,7.2369237,6.820103,6.741334,7.6307697,9.170052,10.95877,12.504617,13.751796,14.601848,14.418053,13.53518,13.24636,0.0,0.0,0.0032820515,0.006564103,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.009846155,0.006564103,0.026256412,0.128,0.055794876,0.04266667,0.07548718,0.12143591,0.14112821,0.24615386,0.4004103,0.54482055,0.6235898,0.61374366,0.5874872,0.39712822,0.2297436,0.18379489,0.25271797,0.18379489,0.14769232,0.13128206,0.13784617,0.18379489,0.33476925,0.4266667,0.446359,0.39712822,0.318359,0.19364104,0.10502565,0.055794876,0.032820515,0.01969231,0.049230773,0.032820515,0.013128206,0.006564103,0.006564103,0.02297436,0.029538464,0.026256412,0.01969231,0.029538464,0.08533334,0.2231795,0.256,0.15425642,0.072205134,0.059076928,0.12143591,0.50543594,1.1454359,1.6410258,0.7450257,0.44307697,0.3708718,0.32164106,0.23958977,0.08533334,0.0951795,0.08533334,0.03938462,0.12143591,0.25271797,0.2100513,0.098461546,0.009846155,0.0,0.0,0.0,0.0,0.0,0.006564103,0.0,0.0,0.0,0.0,0.0,0.009846155,0.08861539,0.17066668,0.18379489,0.02297436,0.0032820515,0.0,0.006564103,0.029538464,0.072205134,0.036102567,0.009846155,0.0,0.0,0.0,0.0,0.016410258,0.059076928,0.08861539,0.0,0.16410258,1.142154,1.8412309,1.7460514,0.93866676,0.42994875,0.26584616,0.36102566,0.58420515,0.761436,0.47589746,0.2231795,0.06564103,0.006564103,0.0,0.006564103,0.0032820515,0.0032820515,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.01969231,0.13784617,0.27897438,0.29210258,0.16082053,0.0,0.0,0.25271797,0.4004103,0.446359,0.7384616,0.8992821,0.6859488,0.4660513,0.43651286,0.6268718,0.3117949,0.18051283,0.21989745,0.29538465,0.15753847,0.3249231,0.3511795,0.34789747,0.4201026,0.6826667,0.5907693,0.3446154,0.16410258,0.10502565,0.06564103,0.052512825,0.059076928,0.03938462,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.02297436,0.029538464,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03938462,0.0951795,0.07548718,0.0,0.0,0.0,0.016410258,0.055794876,0.11158975,0.16082053,0.032820515,0.27897438,0.318359,0.07876924,0.0,0.101743594,0.052512825,0.04594872,0.128,0.17066668,0.108307704,0.059076928,0.07876924,0.15425642,0.20676924,0.04266667,0.009846155,0.009846155,0.006564103,0.036102567,0.16738462,0.190359,0.128,0.03938462,0.029538464,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.036102567,0.032820515,0.13784617,0.15753847,0.08205129,0.072205134,0.24615386,0.3314872,0.33476925,0.27897438,0.19364104,0.18051283,0.23302566,0.24943592,0.21661541,0.23302566,0.29210258,0.27241027,0.20020515,0.1148718,0.055794876,0.009846155,0.07548718,0.101743594,0.052512825,0.0,0.07876924,0.07548718,0.06235898,0.072205134,0.1148718,0.190359,0.36758977,0.38400003,0.25928208,0.31507695,0.36430773,0.3052308,0.3446154,0.49230772,0.56123084,0.47917953,0.5316923,0.46276927,0.3052308,0.38728207,0.58420515,0.7515898,0.8763078,0.9747693,1.1191796,1.0404103,1.024,1.086359,1.1684103,1.148718,1.0338463,0.88287187,0.65641034,0.39056414,0.20020515,0.15097436,0.09189744,0.03938462,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.0032820515,0.0,0.0,0.0,0.013128206,0.026256412,0.01969231,0.006564103,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.016410258,0.009846155,0.013128206,0.02297436,0.036102567,0.052512825,0.06564103,0.049230773,0.06564103,0.098461546,0.128,0.11158975,0.11158975,0.118153855,0.098461546,0.055794876,0.02297436,0.009846155,0.013128206,0.01969231,0.026256412,0.029538464,0.01969231,0.02297436,0.026256412,0.02297436,0.026256412,0.016410258,0.013128206,0.009846155,0.009846155,0.016410258,0.026256412,0.026256412,0.01969231,0.016410258,0.02297436,0.02297436,0.016410258,0.013128206,0.013128206,0.032820515,0.03938462,0.032820515,0.026256412,0.01969231,0.013128206,0.006564103,0.016410258,0.026256412,0.032820515,0.036102567,0.04594872,0.190359,0.4955898,0.73517954,0.4135385,0.30194873,0.16410258,0.072205134,0.03938462,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.006564103,0.02297436,0.07548718,0.15097436,0.22646156,0.23958977,0.190359,0.16738462,0.18051283,0.190359,0.21989745,0.3446154,0.5152821,0.64000005,0.60061544,0.446359,0.39056414,0.28225642,0.15097436,0.20020515,0.7975385,2.809436,4.135385,4.086154,3.373949,3.6102567,3.7382567,4.128821,4.9887185,6.3606157,6.23918,5.7829747,7.5552826,11.831796,16.62359,14.234258,12.491488,11.835078,12.051693,12.291283,11.145847,9.458873,6.560821,4.673641,8.92718,11.661129,7.9983597,5.802667,7.2664623,8.89436,8.004924,7.509334,7.0334363,6.514872,6.229334,7.3649235,8.674462,9.38995,9.616411,10.328616,12.1698475,15.297642,14.592001,10.673231,9.898667,7.778462,5.586052,3.9351797,3.2722054,3.8990772,6.3212314,9.042052,11.0605135,11.690667,10.594462,9.924924,9.281642,10.305642,12.1698475,11.565949,9.69518,8.073847,6.8627696,6.2818465,6.6002054,8.444718,10.607591,11.116308,9.957745,9.07159,8.960001,7.834257,7.5585647,8.241231,8.251078,10.758565,11.795693,10.223591,7.430565,7.312411,9.77395,18.418873,23.03672,19.715284,10.820924,9.90195,10.272821,8.730257,5.1200004,2.3204105,1.7427694,1.5097437,1.339077,1.1388719,1.014154,1.2176411,1.4900514,1.7066668,1.782154,1.6705642,1.5064616,1.3784616,1.332513,1.3751796,1.463795,1.719795,2.228513,2.8127182,3.2065644,3.0818465,3.2000003,3.4034874,3.6168208,3.6824617,3.3772311,3.3542566,3.7448208,4.2994876,4.9296412,5.720616,7.200821,8.267488,9.524513,10.843898,11.385437,10.279386,8.982975,8.018052,7.466667,6.954667,7.463385,8.809027,10.299078,11.595488,12.71795,14.185027,16.072206,16.78113,16.022976,14.805334,0.0,0.0,0.006564103,0.013128206,0.009846155,0.0,0.0032820515,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0,0.01969231,0.068923086,0.14112821,0.2855385,0.46933338,0.6432821,0.761436,0.7844103,0.7318975,0.55794877,0.318359,0.1148718,0.101743594,0.1148718,0.118153855,0.12471796,0.13128206,0.1148718,0.20020515,0.3249231,0.4594872,0.5513847,0.54482055,0.40369233,0.25271797,0.15097436,0.101743594,0.068923086,0.118153855,0.07548718,0.036102567,0.026256412,0.02297436,0.04594872,0.059076928,0.059076928,0.059076928,0.08205129,0.20348719,0.4135385,0.446359,0.27897438,0.15425642,0.06235898,0.07548718,0.14441027,0.21989745,0.27569234,0.6498462,1.0272821,1.1749744,1.0338463,0.7253334,0.5284103,0.702359,0.6892308,0.5513847,0.955077,0.9714873,0.6629744,0.29210258,0.055794876,0.098461546,0.27241027,0.3052308,0.2297436,0.108307704,0.04266667,0.04594872,0.01969231,0.0032820515,0.013128206,0.029538464,0.12143591,0.46276927,0.6235898,0.44307697,0.06235898,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.25271797,1.7263591,2.1464617,1.1749744,0.39056414,0.13784617,0.03938462,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.029538464,0.029538464,0.0,0.0,0.0032820515,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01969231,0.03938462,0.029538464,0.0,0.0,0.0,0.0,0.07876924,0.3446154,0.9419488,1.1520001,1.1027694,0.9353847,0.72861546,0.52512825,0.25271797,0.22646156,0.3052308,0.38728207,0.43651286,0.82379496,0.86646163,0.78769237,0.79425645,1.0535386,0.9682052,0.7089231,0.50543594,0.4135385,0.27897438,0.23958977,0.21333335,0.14769232,0.06564103,0.07876924,0.07548718,0.06235898,0.04594872,0.032820515,0.032820515,0.036102567,0.04266667,0.04594872,0.049230773,0.07876924,0.07876924,0.032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.0032820515,0.0,0.0,0.0,0.08861539,0.19692309,0.15425642,0.0,0.0,0.013128206,0.006564103,0.0,0.04266667,0.20676924,0.072205134,0.013128206,0.08533334,0.18051283,0.03938462,0.049230773,0.055794876,0.128,0.25271797,0.34133336,0.16738462,0.049230773,0.128,0.35774362,0.508718,0.21333335,0.108307704,0.0951795,0.118153855,0.19364104,0.43323082,0.43651286,0.28882053,0.11158975,0.06235898,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01969231,0.10502565,0.0951795,0.06564103,0.04266667,0.032820515,0.03938462,0.098461546,0.11158975,0.108307704,0.08861539,0.016410258,0.18379489,0.44964105,0.5973334,0.5677949,0.4660513,0.6859488,0.65312827,0.4955898,0.3314872,0.23630771,0.08861539,0.101743594,0.09189744,0.026256412,0.026256412,0.18707694,0.18707694,0.15753847,0.18051283,0.27569234,0.4004103,0.37415388,0.26584616,0.14769232,0.098461546,0.01969231,0.032820515,0.17066668,0.29210258,0.098461546,0.23302566,0.3511795,0.46933338,0.6170257,0.8467693,1.1454359,1.3423591,1.467077,1.5392822,1.5753847,1.2471796,1.0896411,1.0305642,1.0010257,0.9156924,0.8041026,0.6104616,0.37415388,0.14769232,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.006564103,0.0032820515,0.0,0.0032820515,0.032820515,0.059076928,0.052512825,0.02297436,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.006564103,0.006564103,0.009846155,0.0032820515,0.013128206,0.032820515,0.04266667,0.03938462,0.07548718,0.12471796,0.15425642,0.118153855,0.13128206,0.13456412,0.108307704,0.055794876,0.032820515,0.02297436,0.01969231,0.01969231,0.01969231,0.029538464,0.01969231,0.029538464,0.036102567,0.029538464,0.036102567,0.01969231,0.006564103,0.006564103,0.009846155,0.01969231,0.029538464,0.026256412,0.02297436,0.026256412,0.03938462,0.03938462,0.026256412,0.01969231,0.029538464,0.059076928,0.068923086,0.055794876,0.03938462,0.032820515,0.026256412,0.016410258,0.02297436,0.029538464,0.032820515,0.04594872,0.036102567,0.04266667,0.27241027,0.6071795,0.6104616,0.39712822,0.23630771,0.12471796,0.04594872,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.04266667,0.108307704,0.18051283,0.19364104,0.17723078,0.15753847,0.15753847,0.19692309,0.23958977,0.26584616,0.3249231,0.40369233,0.43323082,0.3052308,0.18707694,0.108307704,0.08861539,0.128,0.4201026,1.5195899,2.4582565,2.6190772,1.7493335,1.7099489,2.1398976,3.3509746,5.034667,6.2555904,6.442667,6.5247183,8.018052,11.474052,16.456207,14.139078,11.126155,11.37559,14.851283,17.513027,11.828514,8.257642,5.612308,4.20759,5.835488,7.138462,5.2676926,4.903385,7.213949,9.862565,8.792616,8.356103,7.939283,7.4404106,7.250052,7.4863596,7.7292314,8.077128,8.950154,11.057232,11.546257,14.194873,13.4170265,9.626257,9.216001,9.360411,8.372514,6.7971287,5.077334,3.5446157,4.8049235,8.736821,11.74318,11.227899,5.605744,8.635077,7.6274877,7.269744,8.690872,9.452309,8.946873,7.939283,6.452513,5.1364107,5.287385,9.065026,11.831796,12.438975,11.490462,11.37559,11.670976,10.397539,10.262975,10.906258,8.914052,6.4623594,7.13518,9.078155,10.640411,10.345026,11.552821,18.773335,19.882668,13.850258,10.706052,8.946873,8.470975,6.5739493,3.3805132,1.8379488,1.5753847,1.3620514,1.1815386,1.0404103,0.9485129,1.017436,1.2438976,1.6443079,2.028308,1.9889232,1.8215386,1.6311796,1.5425643,1.5983591,1.7427694,1.8773335,2.1891284,2.7569232,3.242667,2.9144619,3.1770258,3.501949,3.6857438,3.7316926,3.8367183,4.2568207,4.70318,5.32677,6.2227697,7.4141545,9.160206,9.931488,10.466462,11.053949,11.542975,11.569232,10.735591,9.416205,8.136206,7.571693,8.592411,10.082462,11.286975,12.009027,12.62277,14.034052,16.75159,18.665028,18.576412,16.200207,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.016410258,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.006564103,0.006564103,0.01969231,0.029538464,0.06564103,0.23302566,0.4955898,0.74830776,0.80738467,0.892718,0.7318975,0.45620516,0.19692309,0.07548718,0.101743594,0.14441027,0.12471796,0.055794876,0.029538464,0.10502565,0.21333335,0.36758977,0.4955898,0.45620516,0.34789747,0.256,0.20020515,0.18051283,0.16738462,0.108307704,0.055794876,0.049230773,0.068923086,0.04594872,0.068923086,0.07548718,0.08205129,0.0951795,0.108307704,0.16738462,0.21989745,0.18379489,0.08205129,0.04594872,0.02297436,0.08861539,0.30194873,0.54482055,0.51856416,0.98133343,1.7493335,2.162872,1.9593848,1.2504616,1.7755898,2.546872,2.609231,2.359795,3.5544617,2.3236926,1.2176411,0.45620516,0.18379489,0.48902568,1.3554872,1.5261539,1.148718,0.5316923,0.15097436,0.21333335,0.09189744,0.01969231,0.06564103,0.15097436,0.50543594,1.6114873,1.8904617,1.0502565,0.06235898,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.08861539,0.17066668,0.06235898,0.02297436,0.016410258,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.006564103,0.0,0.0,0.0,0.013128206,0.016410258,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.052512825,0.25928208,0.27241027,0.108307704,0.0,0.13456412,0.67282057,0.37743592,0.34133336,0.45620516,0.5940513,0.5940513,0.8763078,0.80738467,0.764718,0.9419488,1.3587693,1.4309745,1.4112822,1.2603078,0.99774367,0.7187693,0.6695385,0.47261542,0.33805132,0.33476925,0.39712822,0.38400003,0.30851284,0.2231795,0.16738462,0.16738462,0.18051283,0.2100513,0.2231795,0.20020515,0.15097436,0.10502565,0.036102567,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.049230773,0.02297436,0.0,0.0,0.0,0.049230773,0.02297436,0.0,0.0,0.0,0.072205134,0.036102567,0.0,0.049230773,0.24287182,0.19692309,0.072205134,0.04266667,0.12471796,0.19692309,0.24615386,0.27897438,0.17394873,0.072205134,0.36758977,0.17066668,0.049230773,0.22646156,0.62030774,0.8402052,0.71548724,0.4397949,0.36758977,0.5218462,0.5940513,0.48574364,0.39384618,0.28882053,0.15753847,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.029538464,0.15097436,0.16410258,0.06564103,0.06235898,0.16082053,0.19692309,0.15097436,0.055794876,0.06564103,0.15097436,0.07548718,0.380718,0.6235898,0.76800007,0.80738467,0.74830776,0.67282057,0.53825647,0.46933338,0.5152821,0.6268718,0.3314872,0.18707694,0.13784617,0.13784617,0.13784617,0.15097436,0.17066668,0.18379489,0.190359,0.21333335,0.39712822,0.31507695,0.13784617,0.0,0.0,0.0,0.16410258,0.16410258,0.036102567,0.18379489,0.36758977,0.5874872,0.8795898,1.2242053,1.5425643,1.9692309,2.1398976,2.1530259,2.0250258,1.7099489,1.2438976,0.96492314,0.7515898,0.56123084,0.4266667,0.35446155,0.13456412,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.026256412,0.029538464,0.01969231,0.0032820515,0.016410258,0.016410258,0.032820515,0.052512825,0.052512825,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.02297436,0.029538464,0.029538464,0.006564103,0.0,0.013128206,0.029538464,0.029538464,0.01969231,0.04266667,0.09189744,0.13128206,0.108307704,0.118153855,0.16738462,0.16738462,0.108307704,0.04594872,0.032820515,0.029538464,0.029538464,0.029538464,0.029538464,0.01969231,0.016410258,0.016410258,0.013128206,0.0,0.013128206,0.016410258,0.026256412,0.04266667,0.029538464,0.029538464,0.03938462,0.04594872,0.052512825,0.07548718,0.07548718,0.049230773,0.036102567,0.04594872,0.04594872,0.04594872,0.04594872,0.04594872,0.03938462,0.016410258,0.016410258,0.02297436,0.029538464,0.032820515,0.04594872,0.04594872,0.055794876,0.07876924,0.14769232,0.3052308,0.40369233,0.3446154,0.21661541,0.08861539,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.032820515,0.108307704,0.13128206,0.13784617,0.13784617,0.14769232,0.18379489,0.256,0.3117949,0.33476925,0.3249231,0.27569234,0.22646156,0.17723078,0.128,0.09189744,0.09189744,0.14112821,0.33476925,0.50543594,0.5907693,0.6268718,0.86974365,1.332513,2.481231,3.9745643,4.670359,4.634257,4.532513,5.3858466,7.824411,12.084514,14.5263605,12.803283,11.460924,11.07036,8.224821,7.968821,9.386667,8.648206,5.408821,2.809436,2.930872,3.692308,4.4077954,5.113436,6.5936418,7.4469748,7.5421543,7.243488,7.00718,7.384616,7.4469748,7.4174366,6.311385,4.4274874,3.3411283,5.5532312,9.426052,12.675283,13.574565,10.985026,8.677744,6.6822567,5.671385,5.366154,4.5456414,7.6734366,12.435693,14.546052,12.160001,5.874872,5.435077,5.5532312,6.921847,8.546462,7.765334,8.51036,8.625232,7.817847,6.8266673,7.4010262,7.6209235,7.7948723,7.9163084,8.274052,9.4457445,8.395488,11.867898,14.358975,13.748514,11.306667,7.5946674,8.726975,11.595488,13.971693,14.496821,12.629334,9.9282055,7.968821,7.250052,7.200821,7.2861543,6.5870776,5.2381544,3.570872,2.1070771,1.7263591,1.5491283,1.3850257,1.2176411,1.204513,1.1093334,1.1749744,1.4244103,1.7591796,1.9528207,1.9396925,1.782154,1.6902566,1.7558975,1.9364104,2.1202054,2.284308,2.409026,2.5009232,2.609231,3.0490258,3.239385,3.4067695,3.761231,4.532513,4.9821544,5.077334,5.8781543,7.3419495,8.329846,9.734565,10.883283,11.474052,11.628308,11.871181,12.445539,12.278154,11.073642,9.403078,8.681026,10.023385,10.8996935,11.500309,11.926975,12.20595,13.745232,15.694771,16.866463,16.662975,15.074463,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.01969231,0.013128206,0.006564103,0.032820515,0.108307704,0.21989745,0.32164106,0.3314872,0.43651286,0.54482055,0.49887183,0.30851284,0.13784617,0.12143591,0.12471796,0.11158975,0.07548718,0.04266667,0.08533334,0.13784617,0.19364104,0.26256412,0.3708718,0.3511795,0.318359,0.3249231,0.3708718,0.38728207,0.30851284,0.18379489,0.098461546,0.06564103,0.02297436,0.026256412,0.026256412,0.029538464,0.03938462,0.08205129,0.12471796,0.13456412,0.11158975,0.068923086,0.032820515,0.03938462,0.08205129,0.21333335,0.3314872,0.190359,0.23302566,0.380718,0.51856416,0.56451285,0.48246157,0.65641034,0.9747693,1.2012309,1.2898463,1.3817437,0.86317956,0.75487185,0.9156924,1.0043077,0.48902568,4.1878977,6.245744,6.560821,5.408821,3.4494362,3.1573336,3.387077,2.2482052,0.20348719,0.055794876,0.29210258,0.42338464,0.46276927,0.38400003,0.098461546,0.01969231,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.032820515,0.013128206,0.0032820515,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.013128206,0.01969231,0.049230773,0.098461546,0.10502565,0.08533334,0.052512825,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01969231,0.059076928,0.101743594,0.07548718,0.026256412,0.108307704,0.36758977,0.7581539,0.30851284,0.44307697,0.7253334,0.955077,1.1815386,1.3357949,1.083077,0.85005134,0.7975385,0.8205129,0.86646163,0.9124103,1.2274873,1.6311796,1.4867693,0.95835906,0.75487185,0.90256417,1.204513,1.2274873,0.8041026,0.44307697,0.25928208,0.23630771,0.21661541,0.25928208,0.26584616,0.256,0.21661541,0.128,0.03938462,0.006564103,0.0,0.016410258,0.08533334,0.08533334,0.08533334,0.072205134,0.03938462,0.0,0.009846155,0.0032820515,0.0,0.0,0.0,0.009846155,0.0032820515,0.02297436,0.049230773,0.0,0.013128206,0.006564103,0.0,0.009846155,0.049230773,0.03938462,0.013128206,0.029538464,0.08533334,0.15097436,0.20676924,0.12471796,0.2297436,0.5481026,0.79425645,0.36430773,0.256,0.2855385,0.32820517,0.31507695,0.318359,0.23302566,0.14769232,0.10502565,0.118153855,0.098461546,0.07876924,0.12471796,0.20348719,0.17066668,0.032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.059076928,0.029538464,0.0,0.006564103,0.029538464,0.032820515,0.013128206,0.055794876,0.12143591,0.03938462,0.098461546,0.08861539,0.15097436,0.28225642,0.3446154,0.37743592,0.380718,0.3511795,0.34133336,0.4660513,0.4135385,0.39056414,0.48574364,0.5973334,0.44307697,0.571077,0.5349744,0.41682056,0.30851284,0.30851284,0.26256412,0.26256412,0.25271797,0.2297436,0.21333335,0.2297436,0.3052308,0.28882053,0.17723078,0.108307704,0.13784617,0.18707694,0.23958977,0.35774362,0.67282057,1.1191796,1.3686155,1.6902566,2.103795,2.3696413,2.5337439,2.4352822,2.228513,1.9495386,1.5130258,0.892718,0.6170257,0.48246157,0.39384618,0.36758977,0.128,0.026256412,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.009846155,0.009846155,0.013128206,0.016410258,0.006564103,0.006564103,0.009846155,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.01969231,0.01969231,0.013128206,0.026256412,0.04266667,0.049230773,0.029538464,0.03938462,0.07548718,0.10502565,0.118153855,0.13128206,0.14441027,0.17066668,0.17394873,0.14441027,0.0951795,0.072205134,0.04594872,0.026256412,0.016410258,0.006564103,0.0032820515,0.009846155,0.016410258,0.013128206,0.0,0.013128206,0.02297436,0.03938462,0.055794876,0.055794876,0.04594872,0.04594872,0.049230773,0.059076928,0.06564103,0.06564103,0.06564103,0.068923086,0.072205134,0.08205129,0.072205134,0.068923086,0.068923086,0.06564103,0.03938462,0.029538464,0.029538464,0.026256412,0.02297436,0.032820515,0.052512825,0.08205129,0.1148718,0.15753847,0.21989745,0.318359,0.318359,0.21333335,0.072205134,0.026256412,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.02297436,0.059076928,0.09189744,0.12143591,0.13128206,0.13456412,0.17066668,0.25271797,0.28225642,0.27241027,0.24287182,0.21333335,0.19364104,0.16082053,0.13128206,0.11158975,0.09189744,0.09189744,0.15097436,0.2297436,0.30851284,0.39384618,0.5513847,0.77128214,1.1224617,1.529436,1.7755898,2.3926156,4.4274874,4.9362054,5.2315903,10.889847,12.521027,12.219078,11.900719,11.631591,9.6295395,8.306872,8.096821,8.228104,8.362667,8.605539,5.7403083,4.0402055,3.3444104,4.201026,7.88677,11.592206,12.1928215,11.762873,11.871181,13.59754,11.139283,10.57477,9.32759,8.129642,11.008,11.011283,10.840616,10.732308,10.404103,9.058462,7.90318,6.7807183,6.813539,8.349539,10.9686165,11.789129,14.240822,14.339283,11.378873,7.9130263,6.9842057,4.6966157,3.8137438,4.644103,5.044513,4.0303593,4.4734364,5.2348723,5.9470773,7.0104623,6.741334,6.62318,7.6209235,9.238976,9.544206,9.6754875,12.652308,15.396104,16.466053,16.055796,10.939077,9.734565,11.053949,12.918155,12.750771,11.34277,10.243283,10.259693,10.722463,9.472001,8.152616,7.017026,6.186667,5.32677,3.6693337,3.4264617,3.5478978,2.868513,1.591795,1.2668719,1.1585642,1.1290257,1.1881026,1.3587693,1.6738462,1.8740515,1.9462565,1.8674873,1.7558975,1.8412309,2.2777438,2.5993848,2.7273848,2.7273848,2.8291285,3.006359,2.993231,3.0391798,3.3608208,4.128821,4.6966157,5.5696416,6.7282057,7.834257,8.208411,8.979693,10.121847,11.090053,11.59877,11.628308,11.733335,11.644719,11.119591,10.361437,10.013539,11.024411,11.575796,11.992617,12.245335,11.949949,12.337232,13.1872835,13.699283,13.522053,12.744206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.01969231,0.016410258,0.026256412,0.052512825,0.07548718,0.11158975,0.15097436,0.15097436,0.17723078,0.32820517,0.45292312,0.47261542,0.35446155,0.20348719,0.190359,0.17723078,0.12143591,0.06564103,0.055794876,0.08205129,0.12471796,0.17723078,0.25928208,0.3117949,0.26584616,0.27569234,0.35774362,0.39712822,0.3117949,0.19692309,0.10502565,0.055794876,0.04266667,0.049230773,0.02297436,0.006564103,0.009846155,0.029538464,0.052512825,0.055794876,0.055794876,0.059076928,0.059076928,0.09189744,0.108307704,0.12143591,0.11158975,0.04266667,0.026256412,0.068923086,0.12143591,0.16410258,0.21661541,0.6235898,2.162872,3.7054362,4.529231,4.31918,4.7589746,5.687795,4.785231,2.28759,0.9747693,4.7294364,5.277539,4.417641,3.5774362,3.8071797,3.9023592,3.498667,2.3433847,0.9321026,0.49887183,0.30851284,0.20348719,0.36102566,0.56451285,0.19692309,0.04594872,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016410258,0.08205129,0.016410258,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.01969231,0.055794876,0.1148718,0.07548718,0.055794876,0.04594872,0.032820515,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.09189744,0.20676924,0.26256412,0.190359,0.04266667,0.036102567,0.13128206,0.3117949,0.5874872,0.84348726,1.3062565,1.8904617,2.665026,3.817026,3.2131286,1.8182565,0.75487185,0.41025645,0.40369233,0.6892308,0.9419488,1.3062565,1.7952822,2.300718,1.785436,1.2832822,1.0305642,1.017436,0.98461545,0.6432821,0.33805132,0.20348719,0.2100513,0.15425642,0.20348719,0.21989745,0.21333335,0.20020515,0.17723078,0.18051283,0.17066668,0.18379489,0.21661541,0.24287182,0.30194873,0.3117949,0.2855385,0.24615386,0.21989745,0.22646156,0.20676924,0.18051283,0.16410258,0.16410258,0.15753847,0.14441027,0.15097436,0.16410258,0.15425642,0.029538464,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.08861539,0.33805132,0.13456412,0.29210258,0.43651286,0.4594872,0.5152821,0.3511795,0.256,0.18051283,0.108307704,0.072205134,0.08861539,0.072205134,0.06235898,0.052512825,0.0,0.0,0.026256412,0.06235898,0.098461546,0.15097436,0.072205134,0.02297436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.029538464,0.052512825,0.052512825,0.029538464,0.0,0.029538464,0.013128206,0.0,0.0,0.0,0.0,0.15425642,0.17723078,0.04266667,0.0,0.032820515,0.03938462,0.068923086,0.13784617,0.21989745,0.23302566,0.22646156,0.19692309,0.17394873,0.21333335,0.19364104,0.3052308,0.51856416,0.67610264,0.5152821,0.40369233,0.4266667,0.4397949,0.4135385,0.45292312,0.45620516,0.47261542,0.42994875,0.3314872,0.23958977,0.33476925,0.4201026,0.35774362,0.19692309,0.19364104,0.25928208,0.38400003,0.6268718,1.0043077,1.4998976,1.910154,2.15959,2.359795,2.5140514,2.550154,2.5238976,2.28759,1.9364104,1.5327181,1.0994873,0.61374366,0.44964105,0.30851284,0.14112821,0.14112821,0.029538464,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0032820515,0.006564103,0.006564103,0.0,0.0,0.0032820515,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.0032820515,0.0032820515,0.006564103,0.016410258,0.016410258,0.032820515,0.055794876,0.06564103,0.049230773,0.04594872,0.055794876,0.072205134,0.098461546,0.13784617,0.16410258,0.15097436,0.13456412,0.13128206,0.12471796,0.13128206,0.098461546,0.06235898,0.036102567,0.009846155,0.0032820515,0.009846155,0.016410258,0.013128206,0.0,0.01969231,0.032820515,0.04594872,0.052512825,0.052512825,0.06235898,0.07548718,0.08861539,0.098461546,0.098461546,0.07548718,0.09189744,0.10502565,0.101743594,0.101743594,0.0951795,0.098461546,0.11158975,0.118153855,0.101743594,0.052512825,0.029538464,0.016410258,0.013128206,0.049230773,0.052512825,0.068923086,0.108307704,0.16738462,0.22646156,0.3446154,0.36758977,0.256,0.08861539,0.02297436,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.036102567,0.059076928,0.08533334,0.10502565,0.12143591,0.15097436,0.22646156,0.25271797,0.25271797,0.23958977,0.20676924,0.17394873,0.14769232,0.12143591,0.0951795,0.09189744,0.12471796,0.19692309,0.30194873,0.4004103,0.41025645,0.4201026,0.48902568,0.5973334,0.7253334,0.85005134,1.2504616,2.3827693,2.8291285,3.8400004,9.317744,10.322052,10.679795,10.686359,10.305642,9.199591,8.553026,8.582564,9.140513,9.908514,10.374565,6.951385,5.3891287,4.630975,5.2578464,9.508103,12.596514,14.001232,14.171899,13.804309,13.860104,11.556104,8.402052,6.2523084,6.8299494,11.733335,13.272616,12.435693,11.021129,9.655796,7.8080006,6.449231,6.665847,8.083693,9.954462,11.116308,16.502155,14.569027,10.597744,7.9524107,8.103385,8.4283085,7.7948723,6.921847,5.930667,4.3290257,3.3575387,3.3214362,4.013949,5.21518,6.6822567,7.017026,5.9536414,6.5280004,8.851693,10.108719,9.245539,10.105436,12.73436,16.111591,18.15631,12.242052,9.563898,9.95118,11.920411,12.672001,11.536411,11.067078,10.755282,10.466462,10.423796,11.841642,10.994873,8.6580515,5.910975,4.1222568,3.7316926,3.9023592,3.3641028,2.103795,1.3653334,1.1881026,1.1454359,1.1946667,1.3357949,1.6213335,1.9068719,2.0906668,2.044718,1.8346668,1.7427694,2.03159,2.3958976,2.7142565,2.917744,2.9833848,2.9046156,2.9735386,2.9636924,2.9636924,3.387077,4.1025643,5.5269747,6.892308,7.748924,7.968821,8.438154,9.31118,10.151385,10.6469755,10.587898,10.47959,10.71918,10.79795,10.59118,10.33518,11.021129,11.513436,11.772718,11.733335,11.300103,11.296822,11.510155,11.523283,11.204924,10.696206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.029538464,0.02297436,0.009846155,0.006564103,0.013128206,0.02297436,0.04594872,0.04594872,0.04594872,0.055794876,0.068923086,0.06564103,0.055794876,0.13784617,0.27241027,0.39056414,0.38400003,0.28882053,0.26912823,0.21989745,0.13128206,0.08205129,0.03938462,0.04594872,0.08205129,0.12471796,0.15425642,0.2231795,0.19364104,0.20020515,0.26584616,0.3052308,0.32820517,0.24615386,0.14112821,0.06564103,0.049230773,0.052512825,0.01969231,0.0,0.0,0.0,0.006564103,0.009846155,0.016410258,0.029538464,0.04594872,0.07548718,0.08205129,0.049230773,0.0,0.006564103,0.02297436,0.08205129,0.12143591,0.15425642,0.26584616,0.8402052,2.2219489,3.5610259,4.3060517,4.1911798,4.890257,5.907693,5.0510774,2.7109745,1.8773335,3.6496413,4.1846156,4.2863593,4.5817437,5.5138464,4.6802053,3.495385,2.409026,1.529436,0.6268718,0.32164106,0.27569234,0.40369233,0.48902568,0.18051283,0.04266667,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016410258,0.08205129,0.016410258,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.049230773,0.098461546,0.032820515,0.006564103,0.0032820515,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.026256412,0.01969231,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.026256412,0.013128206,0.0,0.0,0.0,0.0,0.09189744,0.19692309,0.23958977,0.17723078,0.036102567,0.052512825,0.18051283,0.4660513,1.0436924,2.7766156,4.161641,4.650667,4.420923,4.391385,3.2754874,1.7033848,0.5907693,0.20676924,0.16410258,0.5481026,0.69579494,0.85005134,1.2077949,1.9396925,1.8642052,1.5524104,1.214359,0.9485129,0.7122052,0.48574364,0.2986667,0.23630771,0.27241027,0.25928208,0.29210258,0.3117949,0.318359,0.33805132,0.39056414,0.5218462,0.6301539,0.73517954,0.8008206,0.71548724,0.8008206,0.7384616,0.6498462,0.6071795,0.60389745,0.5874872,0.51856416,0.44307697,0.39712822,0.39712822,0.41025645,0.37743592,0.32164106,0.26256412,0.24615386,0.13784617,0.1148718,0.10502565,0.07876924,0.049230773,0.04266667,0.016410258,0.0,0.06564103,0.32164106,0.108307704,0.48574364,0.7187693,0.65312827,0.72861546,0.65641034,0.36102566,0.128,0.052512825,0.029538464,0.006564103,0.0,0.04266667,0.098461546,0.06235898,0.06564103,0.055794876,0.026256412,0.029538464,0.15097436,0.07548718,0.02297436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.029538464,0.052512825,0.052512825,0.029538464,0.0,0.0,0.0,0.0,0.0,0.0,0.03938462,0.27241027,0.31507695,0.128,0.0,0.0,0.036102567,0.036102567,0.026256412,0.13456412,0.15753847,0.15097436,0.16738462,0.2100513,0.24287182,0.24943592,0.31507695,0.51856416,0.7220513,0.571077,0.26912823,0.26912823,0.34133336,0.39056414,0.446359,0.46933338,0.49887183,0.47261542,0.39712822,0.3314872,0.49230772,0.5546667,0.512,0.45292312,0.54482055,0.7089231,0.9682052,1.3489232,1.8412309,2.4024618,2.7831798,2.917744,2.7437952,2.4024618,2.228513,2.0775387,1.9035898,1.6016412,1.1815386,0.7581539,0.4201026,0.29538465,0.16082053,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.0032820515,0.0,0.0032820515,0.016410258,0.01969231,0.032820515,0.055794876,0.08533334,0.10502565,0.12143591,0.108307704,0.098461546,0.10502565,0.12471796,0.13128206,0.108307704,0.09189744,0.11158975,0.16082053,0.23630771,0.21661541,0.15097436,0.08205129,0.03938462,0.016410258,0.013128206,0.016410258,0.013128206,0.006564103,0.029538464,0.04594872,0.055794876,0.06564103,0.06564103,0.08861539,0.108307704,0.12143591,0.128,0.12143591,0.09189744,0.108307704,0.14112821,0.15097436,0.12471796,0.13128206,0.12143591,0.12471796,0.13128206,0.118153855,0.06564103,0.029538464,0.013128206,0.016410258,0.055794876,0.055794876,0.06564103,0.108307704,0.17066668,0.21333335,0.2986667,0.318359,0.23302566,0.09189744,0.02297436,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.02297436,0.04266667,0.059076928,0.07876924,0.101743594,0.13784617,0.23630771,0.26912823,0.29210258,0.3117949,0.3052308,0.21661541,0.15753847,0.1148718,0.0951795,0.1148718,0.17066668,0.25271797,0.33476925,0.39056414,0.36102566,0.35446155,0.380718,0.42994875,0.512,0.6498462,0.80738467,0.9485129,1.2832822,2.550154,6.0291286,7.9819493,10.610872,10.709334,8.3823595,7.026872,7.955693,8.835282,9.321027,9.380103,9.271795,7.8802056,7.8145647,7.5388722,7.197539,8.605539,13.098668,15.681643,15.133539,12.199386,9.5835905,8.690872,5.7501545,3.9680004,5.077334,9.334154,12.27159,11.82195,10.121847,8.28718,6.419693,5.5138464,6.4754877,8.448001,10.102155,9.609847,13.912617,12.619488,9.330873,7.0826674,8.3593855,8.621949,8.635077,8.402052,7.581539,5.4941545,4.027077,3.1671798,3.6102567,5.3037953,7.456821,8.260923,6.62318,6.3967185,8.283898,9.833026,8.730257,8.608821,10.384411,13.380924,15.343591,11.195078,8.592411,8.930462,11.362462,12.780309,12.140308,12.425847,12.196103,11.575796,12.25518,14.427898,13.37436,10.039796,6.1472826,4.1911798,4.141949,5.2447186,5.346462,3.9647183,2.2678976,1.6508719,1.4998976,1.591795,1.7723079,1.9364104,1.9561027,2.0611284,2.169436,2.1956925,2.048,2.048,2.3302567,2.678154,2.92759,2.9735386,2.9636924,3.114667,3.0982566,3.006359,3.3641028,4.132103,5.35959,6.485334,7.250052,7.6931286,8.096821,8.585847,9.002667,9.209436,9.104411,9.068309,9.43918,9.842873,10.06277,10.029949,10.47959,10.860309,10.981745,10.811078,10.476309,10.476309,10.476309,10.276103,9.750975,8.851693,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.026256412,0.06235898,0.049230773,0.01969231,0.0032820515,0.0032820515,0.016410258,0.036102567,0.006564103,0.0,0.0032820515,0.009846155,0.0,0.009846155,0.01969231,0.052512825,0.11158975,0.19364104,0.30851284,0.318359,0.23630771,0.128,0.101743594,0.055794876,0.049230773,0.068923086,0.098461546,0.098461546,0.118153855,0.128,0.14112821,0.16410258,0.18707694,0.36430773,0.36758977,0.26256412,0.12471796,0.049230773,0.01969231,0.009846155,0.006564103,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.009846155,0.009846155,0.01969231,0.03938462,0.09189744,0.18707694,0.3314872,0.54482055,0.90584624,0.96492314,0.8041026,0.5874872,0.57764107,1.1520001,1.467077,1.7690258,2.169436,2.6584618,2.409026,4.5456414,6.875898,7.962257,7.1023593,4.95918,3.626667,2.553436,1.4441026,0.28225642,0.21333335,0.24615386,0.17394873,0.01969231,0.049230773,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0032820515,0.04266667,0.07876924,0.068923086,0.02297436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.036102567,0.06564103,0.009846155,0.0032820515,0.0,0.0,0.0,0.0032820515,0.009846155,0.016410258,0.013128206,0.009846155,0.016410258,0.08533334,0.08861539,0.06235898,0.036102567,0.01969231,0.009846155,0.0032820515,0.0,0.009846155,0.036102567,0.006564103,0.04266667,0.27897438,1.0010257,2.6551797,5.362872,7.0104623,6.6494365,4.585026,2.3827693,1.4375386,0.8598975,0.52512825,0.3249231,0.18707694,0.49230772,0.3511795,0.27569234,0.46933338,0.85005134,1.3029745,1.5983591,1.6607181,1.5195899,1.2996924,1.079795,0.88943595,0.7778462,0.74830776,0.72861546,0.6892308,0.6695385,0.6695385,0.7056411,0.8041026,1.020718,1.2996924,1.4900514,1.4998976,1.3193847,1.3522053,1.1979488,1.0568206,1.0043077,0.99774367,0.9189744,0.79097444,0.67282057,0.5973334,0.5874872,0.64000005,0.60061544,0.48902568,0.36102566,0.29210258,0.380718,0.43323082,0.4201026,0.35446155,0.27897438,0.14769232,0.04594872,0.0,0.013128206,0.072205134,0.101743594,0.45292312,0.7581539,0.9419488,1.2438976,1.0633847,0.508718,0.17066668,0.14769232,0.06235898,0.02297436,0.006564103,0.032820515,0.09189744,0.12143591,0.13128206,0.052512825,0.0032820515,0.04594872,0.17394873,0.036102567,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.032820515,0.036102567,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.101743594,0.26584616,0.3446154,0.26256412,0.0032820515,0.029538464,0.08861539,0.08205129,0.052512825,0.190359,0.20020515,0.20020515,0.25271797,0.36102566,0.46933338,0.44964105,0.4201026,0.571077,0.77456415,0.571077,0.30851284,0.2231795,0.26256412,0.35774362,0.45292312,0.380718,0.4004103,0.446359,0.49230772,0.54482055,0.6892308,0.7581539,0.86646163,1.0436924,1.2274873,1.5163078,1.8642052,2.2383592,2.6157951,2.9768207,3.2984617,3.2295387,2.7437952,2.0742567,1.7362052,1.4506668,1.3850257,1.2242053,0.88287187,0.48902568,0.25271797,0.1148718,0.036102567,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.013128206,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0,0.006564103,0.016410258,0.026256412,0.029538464,0.049230773,0.09189744,0.14441027,0.19364104,0.18051283,0.14769232,0.118153855,0.108307704,0.07548718,0.06235898,0.072205134,0.108307704,0.17723078,0.30194873,0.30194873,0.2231795,0.12471796,0.07876924,0.04266667,0.026256412,0.01969231,0.01969231,0.02297436,0.049230773,0.068923086,0.08861539,0.10502565,0.101743594,0.118153855,0.13456412,0.14112821,0.13456412,0.1148718,0.0951795,0.12471796,0.17066668,0.19692309,0.14769232,0.15753847,0.13128206,0.11158975,0.108307704,0.0951795,0.068923086,0.036102567,0.016410258,0.016410258,0.036102567,0.06564103,0.08533334,0.12471796,0.17723078,0.19692309,0.21333335,0.22646156,0.17394873,0.07876924,0.026256412,0.026256412,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.036102567,0.052512825,0.068923086,0.0951795,0.14112821,0.25928208,0.30851284,0.35446155,0.41025645,0.446359,0.31507695,0.2100513,0.14769232,0.13784617,0.15753847,0.19692309,0.23630771,0.24615386,0.2297436,0.22646156,0.3052308,0.34133336,0.34133336,0.35774362,0.4955898,0.6826667,0.80738467,0.9616411,1.4473847,2.7700515,6.8430777,11.690667,11.316514,6.521436,4.893539,7.4765134,8.845129,8.740103,7.77518,7.4371285,8.897642,10.151385,10.049642,8.592411,6.9349747,13.866668,17.263592,14.792206,8.3593855,4.089436,4.7524104,4.7622566,4.663795,5.2447186,7.53559,9.869129,9.531077,8.096821,6.5280004,5.156103,5.349744,6.2916927,7.9228725,9.42277,9.229129,6.7774363,9.298052,10.246565,8.763078,9.6754875,8.169026,7.017026,7.4141545,8.549745,7.5881033,4.5128207,3.2361028,4.059898,6.409847,8.835282,9.639385,8.39877,7.4929237,7.8047185,8.704,8.602257,8.805744,9.321027,9.8363085,9.731283,8.956718,7.837539,8.251078,10.161232,11.648001,11.779283,12.832822,13.53518,13.538463,13.403898,13.699283,12.747488,10.28595,7.0826674,4.923077,5.284103,7.325539,7.965539,6.311385,3.6529233,2.428718,2.15959,2.3105643,2.4943593,2.4943593,2.0217438,1.9003079,2.162872,2.5796926,2.6584618,2.5337439,2.5632823,2.6518977,2.737231,2.793026,3.045744,3.2196925,3.2656412,3.387077,4.0402055,4.906667,5.4449234,5.970052,6.616616,7.3419495,7.834257,8.027898,7.9819493,7.788308,7.574975,7.6603084,7.962257,8.43159,8.914052,9.156924,9.426052,9.6065645,9.6754875,9.626257,9.468719,9.544206,9.540924,9.399796,8.845129,7.4108725,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.016410258,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.032820515,0.04594872,0.19364104,0.30194873,0.30851284,0.2231795,0.13784617,0.11158975,0.1148718,0.17723078,0.23302566,0.12143591,0.072205134,0.052512825,0.052512825,0.06564103,0.07548718,0.23630771,0.512,0.51856416,0.256,0.12143591,0.02297436,0.026256412,0.03938462,0.02297436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.029538464,0.029538464,0.04266667,0.17394873,0.49230772,0.88943595,1.083077,0.8763078,1.913436,2.0611284,1.1126155,0.80738467,2.4549747,2.5665643,2.0709746,1.7657437,2.3040001,3.255795,3.9351797,4.027077,3.245949,1.3292309,1.4506668,1.3161026,0.86974365,0.29210258,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.009846155,0.0032820515,0.016410258,0.06564103,0.13128206,0.16082053,0.12143591,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.026256412,0.18707694,0.3249231,0.04594872,0.009846155,0.0,0.0,0.0032820515,0.016410258,0.052512825,0.07876924,0.072205134,0.03938462,0.016410258,0.17394873,0.31507695,0.30851284,0.17723078,0.09189744,0.04266667,0.013128206,0.006564103,0.02297436,0.06235898,0.013128206,0.026256412,0.3511795,1.7624617,5.586052,6.3277955,4.601436,2.5042052,1.1881026,0.86974365,0.77128214,0.8467693,0.8041026,0.6268718,0.56451285,0.9682052,1.0502565,1.0568206,1.0962052,1.1454359,1.595077,1.9922053,2.2613335,2.605949,3.508513,3.3378465,2.937436,2.4943593,2.0841026,1.6935385,1.4375386,1.2898463,1.2471796,1.2898463,1.3883078,1.595077,1.9396925,1.9331284,1.5983591,1.463795,1.3423591,1.3029745,1.2800001,1.2307693,1.1454359,0.99774367,0.8598975,0.7450257,0.6629744,0.6268718,0.6859488,0.65641034,0.62030774,0.5973334,0.5481026,0.84348726,1.0338463,1.0699488,0.98461545,0.8992821,0.30194873,0.06235898,0.0,0.0,0.0,0.0,0.0,0.0,0.098461546,0.48902568,0.5973334,0.24943592,0.14112821,0.28225642,0.0,0.06235898,0.029538464,0.0,0.0,0.0,0.0,0.0,0.02297436,0.052512825,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.072205134,0.16410258,0.18379489,0.0,0.0,0.0,0.0,0.013128206,0.06235898,0.12143591,0.13784617,0.101743594,0.03938462,0.016410258,0.15097436,0.072205134,0.036102567,0.10502565,0.15097436,0.26256412,0.45620516,0.571077,0.5546667,0.45620516,0.2986667,0.58092314,0.88615394,0.9616411,0.7187693,0.37415388,0.20676924,0.3249231,0.6465641,0.9156924,0.6104616,0.6071795,0.7187693,0.8369231,0.94523084,1.0929232,1.2570257,1.4834872,1.7624617,2.044718,2.3630772,2.6880002,2.934154,2.9768207,2.6715899,2.5238976,2.3302567,2.28759,2.225231,1.6016412,1.0043077,0.73517954,0.49887183,0.20676924,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.016410258,0.016410258,0.016410258,0.006564103,0.0,0.0,0.0,0.013128206,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.016410258,0.006564103,0.006564103,0.016410258,0.016410258,0.016410258,0.02297436,0.029538464,0.032820515,0.04594872,0.04594872,0.036102567,0.036102567,0.059076928,0.108307704,0.0951795,0.06564103,0.06564103,0.09189744,0.09189744,0.128,0.13784617,0.13128206,0.1148718,0.09189744,0.055794876,0.04594872,0.03938462,0.032820515,0.04594872,0.08205129,0.118153855,0.15097436,0.16082053,0.13784617,0.12471796,0.15097436,0.15425642,0.128,0.09189744,0.09189744,0.14769232,0.18379489,0.17066668,0.12143591,0.13456412,0.13784617,0.13128206,0.118153855,0.108307704,0.068923086,0.04266667,0.01969231,0.0,0.0,0.049230773,0.08861539,0.13784617,0.20676924,0.3052308,0.35446155,0.35774362,0.24615386,0.07548718,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.026256412,0.049230773,0.07876924,0.1148718,0.15097436,0.21333335,0.29210258,0.36758977,0.4201026,0.45620516,0.39712822,0.33476925,0.27569234,0.21989745,0.18379489,0.18379489,0.21989745,0.26256412,0.2855385,0.27569234,0.27569234,0.256,0.23302566,0.22646156,0.27569234,0.5316923,0.76800007,0.98133343,1.782154,4.394667,9.521232,10.866873,8.2904625,4.7491283,6.2851286,9.764103,10.597744,9.412924,7.7423596,8.011488,9.452309,10.013539,8.848411,7.6898465,10.86359,13.794462,16.101746,12.786873,5.5171285,2.6256413,4.1878977,4.850872,5.799385,7.5454364,9.964309,9.865847,9.035488,8.516924,7.90318,5.3398976,5.280821,6.1440005,7.578257,9.265231,10.925949,8.533334,7.240206,6.75118,7.7981544,12.130463,9.432616,8.759795,10.161232,11.58236,8.835282,4.2436924,4.0041027,5.9995904,8.224821,8.772923,9.665642,9.970873,8.602257,6.774154,7.9950776,8.165744,7.604513,7.4896417,7.899898,7.827693,8.146052,8.956718,7.765334,5.7764106,7.890052,8.792616,9.275078,9.93477,10.243283,8.546462,9.193027,11.441232,11.936821,10.013539,7.706257,6.925129,7.030154,7.0367184,6.2162056,4.1058464,2.809436,2.7995899,3.062154,3.0916924,2.8849232,2.1891284,1.847795,1.8937438,2.2908719,2.9768207,3.2328207,2.7569232,2.3893335,2.4155898,2.546872,2.6453335,2.9636924,3.190154,3.4560003,4.332308,5.737026,6.114462,6.12759,6.242462,6.744616,7.4404106,7.640616,7.4404106,6.9776416,6.439385,6.183385,6.6494365,7.1876926,7.460103,7.460103,7.4732313,7.6143594,7.8408213,8.041026,8.041026,7.9819493,7.817847,7.8539495,7.8112826,6.8365135,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0032820515,0.0,0.0,0.02297436,0.02297436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.059076928,0.059076928,0.12471796,0.17066668,0.15753847,0.101743594,0.10502565,0.13128206,0.17066668,0.24615386,0.39056414,0.4004103,0.3117949,0.21661541,0.16082053,0.16082053,0.25271797,0.3511795,0.3249231,0.190359,0.13456412,0.06564103,0.03938462,0.02297436,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.02297436,0.01969231,0.01969231,0.009846155,0.24615386,0.88615394,1.7099489,2.1070771,1.7066668,1.8609232,1.9922053,1.7066668,0.7975385,3.7349746,4.086154,3.3509746,2.8225644,3.5872824,4.969026,4.9985647,4.1124105,2.9965131,2.5862565,1.595077,1.0994873,0.7089231,0.318359,0.12143591,0.2100513,0.20348719,0.108307704,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0032820515,0.016410258,0.016410258,0.026256412,0.032820515,0.02297436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01969231,0.08205129,0.21989745,0.49230772,0.3117949,0.098461546,0.01969231,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.14112821,0.26912823,0.04594872,0.009846155,0.0,0.0,0.006564103,0.03938462,0.06564103,0.07548718,0.052512825,0.006564103,0.0032820515,0.04594872,0.11158975,0.13456412,0.098461546,0.04266667,0.032820515,0.1148718,0.21661541,0.2297436,0.013128206,0.0032820515,0.006564103,0.068923086,0.35774362,1.142154,1.3193847,0.9682052,0.5284103,0.256,0.2100513,0.2100513,0.23958977,0.30194873,0.3511795,0.25928208,0.446359,0.79097444,1.2307693,1.6672822,1.9495386,2.5009232,3.18359,3.9351797,4.4964104,4.414359,4.378257,3.9975388,3.8301542,3.8432825,3.4133337,2.8455386,2.5928206,2.3204105,1.9561027,1.6804104,1.4998976,1.4834872,1.4473847,1.3850257,1.463795,1.5885129,1.7329233,1.8445129,1.7920002,1.3653334,1.1093334,0.9321026,0.8041026,0.7220513,0.67282057,0.7056411,0.7253334,0.6859488,0.56451285,0.37743592,0.37743592,0.39384618,0.35446155,0.256,0.18051283,0.059076928,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.01969231,0.098461546,0.27569234,0.24615386,0.14441027,0.072205134,0.072205134,0.12471796,0.055794876,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.0032820515,0.059076928,0.029538464,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.101743594,0.17066668,0.15753847,0.12143591,0.14112821,0.059076928,0.0,0.0032820515,0.02297436,0.026256412,0.14441027,0.3708718,0.5481026,0.35774362,0.21661541,0.072205134,0.006564103,0.08533334,0.34789747,0.3708718,0.4660513,0.446359,0.32164106,0.3117949,0.32820517,0.39056414,0.45620516,0.48902568,0.44964105,0.4594872,0.6629744,0.52512825,0.24943592,0.7811283,0.74830776,0.7844103,0.86646163,0.9714873,1.0929232,1.2964103,1.5721027,1.9265642,2.2777438,2.4713848,2.809436,2.7667694,2.556718,2.2580514,1.8149745,1.4933335,1.214359,1.0929232,1.0896411,1.0043077,0.62030774,0.45620516,0.26912823,0.04266667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.016410258,0.016410258,0.006564103,0.0,0.0,0.0,0.0,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0,0.006564103,0.016410258,0.016410258,0.016410258,0.009846155,0.009846155,0.01969231,0.02297436,0.03938462,0.029538464,0.02297436,0.04266667,0.08205129,0.07876924,0.059076928,0.059076928,0.08533334,0.1148718,0.1148718,0.11158975,0.12471796,0.15097436,0.16410258,0.22646156,0.26256412,0.21333335,0.11158975,0.0951795,0.11158975,0.13456412,0.13784617,0.118153855,0.11158975,0.11158975,0.1148718,0.11158975,0.0951795,0.06564103,0.08533334,0.118153855,0.14769232,0.16738462,0.15753847,0.16082053,0.16082053,0.15097436,0.13128206,0.118153855,0.072205134,0.04266667,0.02297436,0.013128206,0.013128206,0.032820515,0.04266667,0.06564103,0.13128206,0.26912823,0.42338464,0.46933338,0.36430773,0.16410258,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.036102567,0.06235898,0.07548718,0.098461546,0.16410258,0.18707694,0.26256412,0.3511795,0.4135385,0.4201026,0.4004103,0.39056414,0.3708718,0.32164106,0.256,0.20676924,0.24615386,0.3511795,0.45620516,0.43323082,0.40369233,0.35774362,0.30194873,0.26256412,0.26256412,0.4201026,0.7515898,1.1027694,1.6049232,2.6847181,8.818872,11.483898,9.317744,4.4307694,2.4057438,4.2338467,5.467898,4.97559,4.397949,8.132924,10.157949,9.314463,8.077128,8.641642,12.937847,12.041847,11.539693,10.571488,8.100103,2.8914874,3.7710772,2.678154,2.4451284,4.535795,9.025641,8.749949,8.044309,8.247795,9.284924,9.649232,8.67118,8.03118,8.214975,9.051898,9.718155,6.2785645,5.6320004,5.7632823,5.8157954,6.088206,4.972308,5.1856413,6.8562055,8.228104,5.6352825,3.1277952,2.989949,4.5456414,6.918565,9.028924,10.341744,11.526565,9.964309,6.5772314,5.835488,7.781744,9.42277,10.020103,9.298052,7.4371285,6.4656415,5.7042055,5.32677,5.6385646,7.059693,7.318975,7.6307697,8.372514,9.314463,9.619693,10.850462,11.782565,11.047385,8.690872,6.180103,6.1997952,6.9743595,7.6635904,7.584821,6.2030773,5.1167183,3.945026,2.9735386,2.3762052,2.2383592,2.225231,2.1366155,2.044718,2.0217438,2.156308,2.3072822,2.3827693,2.412308,2.4320002,2.5009232,2.605949,2.7208207,2.7963078,3.0391798,3.9187696,5.6451287,6.380308,6.4722056,6.416411,6.87918,7.3583593,7.463385,7.0367184,6.2720003,5.6943593,5.3398976,5.586052,6.0685134,6.482052,6.5706673,6.669129,6.5772314,6.6494365,6.9054365,7.003898,7.069539,6.882462,6.8332314,6.8693337,6.4689236,0.0,0.006564103,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.026256412,0.02297436,0.0,0.0,0.0,0.0,0.009846155,0.03938462,0.09189744,0.068923086,0.04266667,0.036102567,0.055794876,0.08861539,0.052512825,0.068923086,0.09189744,0.09189744,0.072205134,0.07876924,0.09189744,0.12471796,0.20676924,0.39384618,0.5874872,0.6826667,0.6432821,0.4955898,0.34789747,0.3249231,0.33476925,0.3249231,0.28225642,0.23958977,0.17723078,0.13784617,0.08861539,0.032820515,0.01969231,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.01969231,0.036102567,0.036102567,0.006564103,0.0,0.10502565,0.39712822,0.7778462,0.9747693,0.79425645,0.77128214,0.82379496,0.764718,0.32820517,1.6607181,2.0250258,2.03159,1.9954873,1.9200002,2.5009232,2.8192823,2.9965131,3.0523078,2.8914874,2.103795,2.806154,2.4549747,1.083077,1.3161026,2.2678976,1.6738462,0.73517954,0.14441027,0.06564103,0.036102567,0.026256412,0.016410258,0.0032820515,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.009846155,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.032820515,0.04266667,0.04266667,0.029538464,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.04266667,0.118153855,0.24943592,0.15753847,0.049230773,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.052512825,0.101743594,0.01969231,0.0032820515,0.0,0.0,0.0032820515,0.01969231,0.029538464,0.029538464,0.01969231,0.0,0.0,0.0032820515,0.02297436,0.04266667,0.052512825,0.03938462,0.068923086,0.13784617,0.16082053,0.11158975,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.026256412,0.06564103,0.11158975,0.12143591,0.036102567,0.06235898,0.055794876,0.07876924,0.13456412,0.15425642,0.318359,0.636718,1.2373334,2.0775387,2.9472823,3.508513,4.023795,4.388103,4.6572313,5.0609236,4.604718,4.1485133,4.0992823,4.3684106,4.3684106,4.3651285,4.4865646,3.5511796,1.9462565,1.6082052,1.394872,1.3259488,1.3029745,1.3226668,1.463795,1.7788719,1.9561027,2.0053334,1.910154,1.6016412,1.394872,1.2504616,1.1191796,0.9878975,0.88943595,0.8467693,0.8369231,0.764718,0.57764107,0.26256412,0.19692309,0.16410258,0.108307704,0.029538464,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.07876924,0.098461546,0.059076928,0.006564103,0.036102567,0.055794876,0.06235898,0.049230773,0.029538464,0.04594872,0.009846155,0.0,0.0,0.0,0.0,0.059076928,0.055794876,0.04266667,0.029538464,0.0,0.0,0.03938462,0.03938462,0.0,0.0,0.0,0.04266667,0.068923086,0.06235898,0.06235898,0.101743594,0.049230773,0.009846155,0.009846155,0.006564103,0.04594872,0.20020515,0.41025645,0.5546667,0.4594872,0.37743592,0.25928208,0.24943592,0.35446155,0.42338464,0.50543594,0.4266667,0.32820517,0.27569234,0.26584616,0.318359,0.4266667,0.5940513,0.8795898,1.3883078,0.8336411,0.69579494,0.5940513,0.49230772,0.7122052,0.7122052,0.8533334,1.0502565,1.214359,1.2471796,1.4539489,1.7394873,2.0217438,2.1858463,2.0939488,2.2383592,2.0939488,1.7624617,1.339077,0.9156924,0.67282057,0.6071795,0.6301539,0.6268718,0.44307697,0.2297436,0.15425642,0.08533334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.032820515,0.04266667,0.01969231,0.006564103,0.0,0.0,0.0032820515,0.009846155,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.013128206,0.006564103,0.01969231,0.01969231,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.02297436,0.032820515,0.049230773,0.072205134,0.06235898,0.072205134,0.098461546,0.11158975,0.09189744,0.0951795,0.1148718,0.15097436,0.18379489,0.28225642,0.42994875,0.38728207,0.18051283,0.098461546,0.0951795,0.101743594,0.108307704,0.108307704,0.108307704,0.098461546,0.08533334,0.068923086,0.055794876,0.052512825,0.068923086,0.08533334,0.108307704,0.13456412,0.14112821,0.13456412,0.14769232,0.16082053,0.15753847,0.13128206,0.098461546,0.07548718,0.055794876,0.03938462,0.032820515,0.029538464,0.029538464,0.04266667,0.08205129,0.18707694,0.26584616,0.36102566,0.33476925,0.18379489,0.032820515,0.006564103,0.006564103,0.009846155,0.013128206,0.026256412,0.006564103,0.0,0.0,0.0032820515,0.016410258,0.03938462,0.059076928,0.06564103,0.072205134,0.0951795,0.128,0.21661541,0.3708718,0.5021539,0.4201026,0.3511795,0.34133336,0.3511795,0.35446155,0.33805132,0.30851284,0.31507695,0.3511795,0.380718,0.3708718,0.36430773,0.3446154,0.3249231,0.3052308,0.2855385,0.33476925,0.5284103,0.8172308,1.2438976,1.9462565,6.0258465,13.689437,14.713437,8.2904625,3.0358977,4.06318,5.366154,5.4383593,5.5926156,9.977437,12.002462,7.8145647,5.474462,7.8736415,12.754052,10.650257,9.222565,8.3134365,6.944821,3.3280003,2.5993848,1.6705642,1.6738462,3.4330258,7.4797955,7.4765134,7.138462,7.056411,7.4469748,8.162462,7.768616,6.6461544,6.2687182,6.547693,5.8256416,4.640821,3.8859491,3.6529233,3.6332312,3.121231,2.5042052,2.9210258,4.44718,5.986462,5.2578464,3.05559,2.4188719,3.2196925,4.9460516,6.685539,7.456821,8.484103,7.830975,5.9634876,5.733744,7.0793853,8.333129,9.481847,10.118565,9.4457445,8.218257,6.7249236,6.173539,6.665847,7.207385,6.2884107,6.3540516,9.521232,13.512206,11.680821,11.641437,11.864616,11.224616,9.347282,6.633026,6.806975,8.454565,10.269539,11.204924,10.463181,9.193027,7.197539,5.3760004,3.9712822,2.550154,2.2547693,2.2613335,2.2416413,2.0808206,1.8609232,1.8871796,2.1431797,2.3860514,2.5074873,2.5337439,2.6289232,2.678154,2.6945643,2.8324106,3.373949,4.71959,5.8781543,6.242462,6.0619493,6.426257,6.6625648,6.685539,6.3376417,5.7468724,5.3169236,5.2381544,5.431795,5.5630774,5.5302567,5.4514875,5.6451287,5.792821,5.933949,6.1046157,6.314667,6.514872,6.629744,6.7610264,6.7872825,6.370462,0.0,0.006564103,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.013128206,0.009846155,0.0,0.0,0.0,0.0,0.009846155,0.04266667,0.098461546,0.17394873,0.13128206,0.1148718,0.15753847,0.16738462,0.08861539,0.055794876,0.04594872,0.04266667,0.04266667,0.049230773,0.072205134,0.11158975,0.17394873,0.26584616,0.48902568,0.6826667,0.7318975,0.63343596,0.50543594,0.40697438,0.4201026,0.4266667,0.37743592,0.2986667,0.25271797,0.24615386,0.2297436,0.18051283,0.128,0.04594872,0.009846155,0.0,0.0,0.0,0.0,0.009846155,0.026256412,0.029538464,0.0,0.0,0.0,0.0032820515,0.013128206,0.026256412,0.032820515,0.06564103,0.08533334,0.08205129,0.08205129,0.11158975,0.27241027,0.5677949,0.761436,0.35774362,0.34789747,0.71548724,1.3653334,2.0250258,2.2186668,2.5271797,3.9745643,3.95159,2.4516926,2.0709746,2.6518977,2.1858463,1.6180514,1.3751796,1.3653334,1.7362052,1.5589745,0.9189744,0.24615386,0.3249231,0.06564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.006564103,0.029538464,0.0951795,0.059076928,0.029538464,0.013128206,0.01969231,0.02297436,0.01969231,0.013128206,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.029538464,0.04266667,0.04266667,0.029538464,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.02297436,0.03938462,0.08205129,0.101743594,0.06235898,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.07876924,0.19692309,0.27241027,0.15097436,1.086359,0.90912825,0.4594872,0.22646156,0.36430773,0.6235898,0.8172308,1.2504616,2.0939488,3.370667,3.639795,3.9680004,3.9614363,3.9712822,5.0674877,4.4406157,3.8596926,3.7120004,4.013949,4.391385,4.9952826,5.4547696,4.4242053,2.3893335,1.6738462,1.4933335,1.4309745,1.3620514,1.3029745,1.4145643,1.7362052,1.8149745,1.7755898,1.6738462,1.4933335,1.3784616,1.2931283,1.2012309,1.086359,0.9616411,0.90584624,0.8566154,0.77128214,0.60389745,0.32820517,0.26256412,0.23302566,0.190359,0.13784617,0.13456412,0.10502565,0.068923086,0.04266667,0.029538464,0.02297436,0.0032820515,0.0,0.016410258,0.04594872,0.06235898,0.098461546,0.12143591,0.13128206,0.13456412,0.14112821,0.12471796,0.15753847,0.17723078,0.17066668,0.16082053,0.1148718,0.098461546,0.08205129,0.052512825,0.02297436,0.032820515,0.068923086,0.068923086,0.032820515,0.0,0.02297436,0.049230773,0.03938462,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.049230773,0.029538464,0.009846155,0.006564103,0.0,0.101743594,0.25271797,0.4266667,0.5481026,0.48574364,0.38400003,0.29538465,0.318359,0.40369233,0.37415388,0.53825647,0.4135385,0.26912823,0.23630771,0.32164106,0.702359,0.74830776,0.8008206,1.0305642,1.4506668,0.81394875,0.5481026,0.53825647,0.6235898,0.60061544,0.6498462,0.8566154,1.1355898,1.3915899,1.522872,1.6640002,1.8346668,1.9265642,1.8510771,1.5392822,1.3653334,1.1618463,0.9156924,0.62030774,0.27569234,0.2231795,0.3249231,0.42994875,0.41025645,0.13784617,0.026256412,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.052512825,0.055794876,0.013128206,0.0,0.0,0.0,0.0032820515,0.009846155,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.006564103,0.01969231,0.01969231,0.016410258,0.016410258,0.016410258,0.0032820515,0.006564103,0.016410258,0.026256412,0.029538464,0.052512825,0.055794876,0.072205134,0.101743594,0.11158975,0.09189744,0.10502565,0.13784617,0.17066668,0.190359,0.24943592,0.39712822,0.380718,0.20348719,0.108307704,0.068923086,0.059076928,0.068923086,0.08205129,0.08205129,0.059076928,0.049230773,0.03938462,0.036102567,0.052512825,0.06564103,0.07548718,0.098461546,0.128,0.14112821,0.118153855,0.128,0.15425642,0.17394873,0.15425642,0.14112821,0.12471796,0.098461546,0.068923086,0.04594872,0.032820515,0.032820515,0.04266667,0.06235898,0.101743594,0.11158975,0.20348719,0.2297436,0.16082053,0.04594872,0.013128206,0.006564103,0.009846155,0.013128206,0.026256412,0.006564103,0.0,0.0032820515,0.006564103,0.009846155,0.029538464,0.03938462,0.04594872,0.04594872,0.03938462,0.07876924,0.14112821,0.26912823,0.39384618,0.34789747,0.29538465,0.2855385,0.29210258,0.30851284,0.3249231,0.32820517,0.3249231,0.30194873,0.27241027,0.256,0.27241027,0.29538465,0.30851284,0.29538465,0.26256412,0.256,0.3446154,0.54482055,0.88615394,1.4211283,3.1409233,9.711591,11.54954,7.1154876,2.9210258,3.9975388,5.546667,5.9995904,5.927385,8.054154,9.485129,5.2480006,3.3214362,6.629744,13.02318,9.921641,7.466667,5.677949,4.309334,2.8192823,1.7460514,1.5360001,2.0512822,3.4855387,6.3868723,7.8834877,8.861539,8.198565,6.416411,5.677949,5.536821,4.4832826,4.073026,4.5095387,4.6605134,5.175795,4.378257,3.2918978,2.425436,1.7723079,1.5031796,1.8806155,3.314872,5.5105643,7.4436927,4.07959,4.20759,5.681231,6.951385,7.069539,7.2369237,7.936001,8.024616,7.4436927,7.204103,7.1844106,7.1056414,7.463385,8.339693,9.403078,9.147078,7.6570263,7.0925136,7.890052,8.740103,7.1844106,6.738052,9.813334,13.617231,10.151385,10.016821,10.95877,11.332924,10.473026,8.717129,9.498257,11.641437,13.830565,15.015386,14.41477,13.515489,11.844924,9.829744,7.394462,3.9614363,2.4484105,2.1202054,2.1169233,2.0020514,1.7624617,1.7033848,1.9331284,2.2055387,2.3860514,2.4418464,2.550154,2.6880002,2.7470772,2.7733335,2.9735386,3.7382567,4.906667,5.4875903,5.408821,5.504,5.4843082,5.5565133,5.612308,5.602462,5.543385,5.4941545,5.4613338,5.228308,4.841026,4.6080003,4.7392826,4.965744,5.149539,5.297231,5.546667,5.8486156,6.2785645,6.626462,6.7085133,6.373744,0.016410258,0.013128206,0.006564103,0.0032820515,0.0,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.01969231,0.21661541,0.18051283,0.17066668,0.23630771,0.24287182,0.13784617,0.072205134,0.032820515,0.013128206,0.016410258,0.026256412,0.068923086,0.1148718,0.13784617,0.13128206,0.23958977,0.37743592,0.49230772,0.56123084,0.60061544,0.48246157,0.5513847,0.5546667,0.42338464,0.27569234,0.27569234,0.3249231,0.37415388,0.380718,0.29210258,0.128,0.03938462,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.06235898,0.101743594,0.118153855,0.15097436,0.15097436,0.06564103,0.006564103,0.0,0.0032820515,0.013128206,0.029538464,0.072205134,0.29538465,0.97805136,2.1497438,3.1967182,3.6135387,3.1606157,1.8642052,1.214359,1.5786668,2.2711797,2.7700515,2.7109745,3.442872,3.1081028,1.8576412,0.5284103,0.6432821,0.128,0.0,0.0,0.0,0.0,0.02297436,0.04266667,0.098461546,0.16738462,0.190359,0.10502565,0.032820515,0.0032820515,0.04266667,0.17066668,0.10502565,0.068923086,0.0951795,0.16082053,0.16738462,0.098461546,0.052512825,0.01969231,0.006564103,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.04266667,0.0951795,0.06564103,0.02297436,0.0,0.0,0.0,0.009846155,0.013128206,0.009846155,0.006564103,0.026256412,0.098461546,0.2297436,0.34133336,0.28225642,2.1366155,1.8674873,1.0043077,0.48574364,0.64000005,0.9682052,1.0404103,1.148718,1.6147693,2.7864618,2.7995899,3.1277952,3.0949745,3.0030773,4.1452312,3.9187696,3.4625645,3.2656412,3.43959,3.7152824,4.2305646,4.647385,4.1714873,2.9013336,1.8543591,1.7460514,1.7001027,1.6082052,1.4998976,1.5753847,1.6311796,1.5491283,1.4244103,1.2898463,1.0929232,1.0371283,0.99774367,0.9682052,0.9353847,0.86646163,0.8730257,0.8566154,0.79097444,0.69579494,0.6170257,0.5284103,0.48574364,0.45292312,0.4201026,0.40369233,0.33476925,0.24615386,0.18051283,0.14112821,0.11158975,0.06235898,0.052512825,0.098461546,0.17723078,0.23302566,0.33805132,0.4004103,0.43323082,0.44307697,0.44964105,0.42338464,0.39056414,0.39056414,0.40697438,0.35774362,0.3249231,0.3052308,0.25271797,0.16410258,0.0951795,0.049230773,0.07876924,0.1148718,0.1148718,0.06235898,0.07548718,0.03938462,0.006564103,0.0,0.0,0.0032820515,0.0032820515,0.02297436,0.04266667,0.02297436,0.06235898,0.04266667,0.013128206,0.0,0.0,0.17394873,0.2855385,0.4397949,0.574359,0.45620516,0.256,0.18051283,0.18051283,0.21989745,0.2855385,0.44307697,0.4201026,0.3052308,0.24287182,0.4266667,1.1684103,1.0765129,0.86974365,0.78769237,0.5973334,0.48246157,0.4660513,0.48246157,0.49887183,0.49230772,0.65641034,0.88287187,1.1618463,1.4736412,1.785436,1.8051283,1.7723079,1.6311796,1.3718976,1.014154,0.62030774,0.39712822,0.2986667,0.2231795,0.0,0.10502565,0.20020515,0.256,0.22646156,0.072205134,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02297436,0.03938462,0.029538464,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.013128206,0.02297436,0.02297436,0.013128206,0.006564103,0.016410258,0.01969231,0.009846155,0.0032820515,0.006564103,0.016410258,0.02297436,0.026256412,0.036102567,0.059076928,0.098461546,0.13128206,0.118153855,0.14112821,0.18379489,0.21661541,0.19692309,0.17723078,0.23302566,0.24615386,0.190359,0.14112821,0.059076928,0.032820515,0.036102567,0.04266667,0.049230773,0.026256412,0.02297436,0.02297436,0.032820515,0.055794876,0.068923086,0.08533334,0.1148718,0.15753847,0.17394873,0.12143591,0.108307704,0.12471796,0.15097436,0.16410258,0.17723078,0.17066668,0.13784617,0.0951795,0.059076928,0.04266667,0.04266667,0.049230773,0.052512825,0.03938462,0.055794876,0.09189744,0.128,0.12471796,0.04594872,0.02297436,0.006564103,0.0,0.0032820515,0.0,0.0032820515,0.0032820515,0.006564103,0.013128206,0.0,0.009846155,0.013128206,0.01969231,0.029538464,0.036102567,0.055794876,0.068923086,0.09189744,0.14441027,0.22646156,0.25928208,0.256,0.23958977,0.2231795,0.2297436,0.24615386,0.24943592,0.23302566,0.20348719,0.17723078,0.21333335,0.27569234,0.29538465,0.256,0.20020515,0.19692309,0.2855385,0.45292312,0.67610264,0.92225647,1.3292309,1.6016412,1.6278975,1.4408206,1.2307693,2.809436,4.9329233,5.4908724,4.2863593,3.0162053,3.5380516,2.4418464,2.3236926,5.1265645,12.166565,8.802463,6.1472826,3.9089234,2.228513,1.657436,1.4441026,1.6968206,2.5173335,4.007385,6.242462,9.570462,11.792411,10.630565,6.8332314,4.1452312,3.4560003,2.8455386,2.8258464,3.7448208,5.7764106,6.340924,6.157129,4.6933336,2.5665643,1.522872,1.4834872,1.6508719,2.9144619,5.5302567,9.107693,5.412103,7.5421543,10.55836,11.713642,10.469745,10.125129,10.781539,11.1064625,10.509129,9.120821,8.569437,7.5388722,6.189949,5.428513,6.8988724,7.9819493,6.99077,6.957949,8.67118,10.673231,9.478565,8.562873,8.94359,9.593436,7.4404106,9.061745,10.660104,11.779283,12.182976,11.864616,13.587693,16.246155,17.96595,18.110361,17.243898,16.764719,16.384,14.9628725,11.9171295,7.210667,3.9286156,2.5337439,2.044718,1.8543591,1.7329233,1.6311796,1.785436,2.03159,2.2514873,2.3762052,2.5238976,2.7437952,2.8160002,2.7536411,2.802872,3.2229745,4.092718,4.7524104,4.9132314,4.6211286,4.378257,4.6211286,5.21518,5.904411,6.301539,6.058667,5.7009234,5.2545643,4.778667,4.3684106,4.263385,4.3027697,4.46359,4.709744,4.9493337,5.277539,5.796103,6.2227697,6.3967185,6.2851286,0.07548718,0.06564103,0.032820515,0.009846155,0.0032820515,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.01969231,0.029538464,0.04266667,0.026256412,0.03938462,0.098461546,0.18379489,0.23302566,0.17066668,0.072205134,0.0032820515,0.016410258,0.016410258,0.006564103,0.013128206,0.04594872,0.108307704,0.25271797,0.380718,0.5415385,0.6859488,0.6859488,0.57764107,0.64000005,0.63343596,0.46933338,0.21333335,0.3249231,0.3708718,0.4004103,0.4135385,0.36758977,0.21989745,0.101743594,0.026256412,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.016410258,0.006564103,0.0,0.0032820515,0.016410258,0.016410258,0.1148718,0.1148718,0.013128206,0.0,0.0,0.11158975,0.41682056,0.8402052,1.1454359,1.1552821,1.7460514,1.9889232,1.5261539,0.5481026,0.20676924,0.20348719,0.25271797,0.20348719,0.04594872,0.009846155,0.0,0.0,0.0,0.0,0.108307704,0.21989745,0.48902568,0.8369231,0.94523084,0.46933338,0.14112821,0.0,0.0,0.0,0.013128206,0.098461546,0.33476925,0.6071795,0.5940513,0.30194873,0.108307704,0.029538464,0.032820515,0.04594872,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01969231,0.09189744,0.21333335,0.13456412,0.036102567,0.0,0.0,0.0,0.04594872,0.06564103,0.04266667,0.029538464,0.07876924,0.13784617,0.15425642,0.12471796,0.07548718,0.16082053,0.42994875,0.5152821,0.39712822,0.39712822,0.51856416,0.4955898,0.5021539,0.67610264,1.1126155,1.7624617,2.281026,2.3040001,2.0086155,2.1070771,2.678154,3.170462,3.5314875,3.56759,2.9440002,2.0676925,1.8937438,1.7952822,1.5983591,1.5885129,1.8182565,1.9790771,2.166154,2.3794873,2.5009232,2.0020514,1.7952822,1.4998976,1.0929232,0.88615394,0.8008206,0.761436,0.7417436,0.7581539,0.8533334,0.93866676,1.079795,1.079795,0.98133343,1.0666667,0.92225647,0.81066674,0.7450257,0.7089231,0.67282057,0.6235898,0.5546667,0.48902568,0.41682056,0.32164106,0.25928208,0.26256412,0.3249231,0.4266667,0.5481026,0.6826667,0.8008206,0.8598975,0.86317956,0.8402052,0.86317956,0.76800007,0.67282057,0.6268718,0.6268718,0.56451285,0.5316923,0.43323082,0.28882053,0.2297436,0.20348719,0.13456412,0.2855385,0.52512825,0.3052308,0.13456412,0.072205134,0.036102567,0.0,0.0,0.013128206,0.016410258,0.108307704,0.21989745,0.12143591,0.12143591,0.12143591,0.072205134,0.0,0.0,0.28225642,0.3314872,0.27897438,0.22646156,0.27569234,0.2986667,0.24943592,0.24287182,0.2986667,0.33476925,0.2855385,0.36758977,0.48246157,0.5481026,0.48902568,0.67282057,0.80738467,0.8992821,0.9288206,0.8533334,0.7089231,0.69907695,0.67282057,0.60061544,0.56451285,0.761436,1.0371283,1.3292309,1.5655385,1.6640002,1.5163078,1.3259488,0.9944616,0.5874872,0.3052308,0.14769232,0.13456412,0.09189744,0.0,0.0,0.08533334,0.08861539,0.08861539,0.08533334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.006564103,0.006564103,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.026256412,0.049230773,0.06235898,0.06235898,0.032820515,0.016410258,0.01969231,0.029538464,0.029538464,0.02297436,0.016410258,0.013128206,0.0,0.013128206,0.016410258,0.04594872,0.108307704,0.16738462,0.15425642,0.17066668,0.21333335,0.24287182,0.18379489,0.14769232,0.21989745,0.256,0.21333335,0.15097436,0.09189744,0.049230773,0.029538464,0.036102567,0.06235898,0.098461546,0.068923086,0.032820515,0.01969231,0.029538464,0.055794876,0.07876924,0.1148718,0.16082053,0.19692309,0.08861539,0.06235898,0.06235898,0.06564103,0.09189744,0.15097436,0.18707694,0.18051283,0.14441027,0.108307704,0.08205129,0.059076928,0.03938462,0.026256412,0.016410258,0.03938462,0.072205134,0.098461546,0.0951795,0.04594872,0.02297436,0.006564103,0.006564103,0.013128206,0.0,0.013128206,0.016410258,0.016410258,0.013128206,0.0,0.0,0.0,0.006564103,0.02297436,0.06235898,0.06235898,0.06235898,0.08533334,0.14112821,0.21333335,0.23958977,0.22646156,0.20020515,0.18051283,0.16738462,0.15425642,0.15097436,0.14769232,0.14112821,0.15097436,0.23958977,0.34133336,0.36758977,0.2986667,0.21333335,0.190359,0.27569234,0.47589746,0.71548724,0.82379496,0.90912825,1.2340513,1.4834872,1.5589745,1.5721027,3.318154,6.1341543,6.3901544,3.8465643,1.6475899,1.5261539,1.339077,1.5885129,2.5600002,4.31918,4.8804107,6.705231,5.802667,2.5107694,1.5097437,1.083077,1.2865642,2.3991797,4.4012313,6.987488,9.905231,10.545232,8.992821,5.940513,2.6551797,1.5064616,1.8445129,2.605949,3.0785644,2.8849232,3.4592824,4.9362054,5.0215387,3.6102567,2.793026,2.0118976,1.4867693,1.7558975,2.8553848,4.332308,5.4449234,8.871386,11.441232,12.143591,12.130463,10.801231,11.713642,12.36677,11.625027,9.7214365,11.063796,10.44677,8.516924,6.373744,5.5696416,6.436103,6.0947695,6.7117953,8.681026,10.633847,10.624001,10.098872,9.852718,10.601027,12.970668,16.498873,14.880821,14.506668,16.210052,15.258258,16.94195,21.494156,22.951385,20.772104,19.820309,17.808413,18.49436,18.474669,16.538258,13.656616,8.772923,5.218462,3.1376412,2.2449234,1.8313848,1.7099489,1.8904617,2.284308,2.7076926,2.8521028,2.9997952,2.9636924,2.793026,2.6420515,2.7766156,3.4724104,4.378257,5.080616,5.2545643,4.670359,4.338872,4.706462,5.579488,6.5936418,7.2172313,7.2172313,6.9054365,6.4590774,5.85518,4.8672824,4.4996924,4.5029745,4.7589746,5.1331286,5.4613338,5.681231,5.910975,6.1374364,6.2096415,5.8453336,0.15097436,0.128,0.07876924,0.03938462,0.02297436,0.016410258,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.01969231,0.029538464,0.036102567,0.036102567,0.032820515,0.049230773,0.059076928,0.07548718,0.06564103,0.036102567,0.026256412,0.026256412,0.01969231,0.009846155,0.016410258,0.059076928,0.108307704,0.256,0.47589746,0.7089231,0.8467693,0.67610264,0.58092314,0.574359,0.60061544,0.5316923,0.41682056,0.44307697,0.49230772,0.49887183,0.45292312,0.33476925,0.2231795,0.12471796,0.052512825,0.02297436,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.02297436,0.01969231,0.006564103,0.0,0.0032820515,0.0032820515,0.02297436,0.02297436,0.0032820515,0.0,0.0,0.059076928,0.21661541,0.43323082,0.58420515,0.7220513,1.2471796,1.5392822,1.3423591,0.7581539,1.782154,1.204513,0.4397949,0.098461546,0.009846155,0.0032820515,0.0,0.0,0.013128206,0.06235898,0.6892308,1.0371283,1.017436,0.73517954,0.48246157,0.33805132,0.26584616,0.25928208,0.256,0.15753847,0.11158975,0.27897438,0.60389745,0.92553854,0.9616411,0.5513847,0.22646156,0.1148718,0.16410258,0.15425642,0.059076928,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.06564103,0.20020515,0.28225642,0.24287182,0.1148718,0.036102567,0.04594872,0.059076928,0.052512825,0.06564103,0.190359,0.5513847,0.5481026,0.3314872,0.101743594,0.101743594,0.28225642,0.37743592,0.33805132,0.20676924,0.128,0.190359,0.36430773,0.47261542,0.5349744,0.761436,1.017436,1.7460514,2.1366155,1.9232821,1.3850257,1.1782565,1.0043077,1.0535386,1.3423591,1.7362052,1.4736412,1.2537436,1.1290257,1.148718,1.3915899,1.9167181,2.3302567,2.6190772,2.6420515,2.1497438,2.0086155,1.9200002,1.7690258,1.4966155,1.0929232,1.0371283,0.9517949,0.83035904,0.7318975,0.7811283,0.8467693,0.80738467,0.76800007,0.7778462,0.82379496,0.8041026,0.7844103,0.76800007,0.7515898,0.7450257,0.7253334,0.8566154,0.93866676,0.9156924,0.8566154,0.8566154,0.8205129,0.82379496,0.88615394,0.9878975,1.0732309,1.142154,1.1684103,1.1388719,1.0469744,1.0896411,0.96492314,0.8533334,0.80738467,0.761436,0.6498462,0.5152821,0.4004103,0.3117949,0.23958977,0.18707694,0.16082053,0.22646156,0.33476925,0.32820517,0.2855385,0.26256412,0.20348719,0.128,0.14769232,0.17723078,0.2297436,0.32164106,0.42338464,0.46276927,0.5021539,0.2986667,0.14769232,0.17394873,0.32820517,0.512,0.48246157,0.42338464,0.4135385,0.43323082,0.380718,0.39056414,0.571077,0.8205129,0.8467693,0.54482055,0.4004103,0.40369233,0.5415385,0.79425645,0.8402052,0.9517949,1.0305642,1.0929232,1.2340513,1.0962052,1.1323078,1.1093334,1.0108719,1.0535386,1.1323078,1.1946667,1.273436,1.3554872,1.394872,1.0338463,0.6695385,0.4201026,0.26256412,0.06235898,0.029538464,0.04266667,0.072205134,0.07876924,0.0,0.07548718,0.04594872,0.016410258,0.016410258,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.016410258,0.02297436,0.013128206,0.0032820515,0.0,0.0,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.016410258,0.01969231,0.013128206,0.02297436,0.01969231,0.009846155,0.0032820515,0.006564103,0.016410258,0.009846155,0.0032820515,0.0032820515,0.0,0.0032820515,0.009846155,0.029538464,0.068923086,0.118153855,0.118153855,0.13456412,0.17723078,0.22646156,0.24287182,0.24615386,0.24943592,0.24287182,0.24287182,0.2986667,0.2297436,0.12471796,0.049230773,0.02297436,0.036102567,0.052512825,0.04266667,0.026256412,0.016410258,0.01969231,0.052512825,0.07876924,0.09189744,0.09189744,0.101743594,0.059076928,0.04266667,0.04266667,0.055794876,0.07876924,0.13128206,0.15425642,0.15753847,0.14441027,0.118153855,0.08533334,0.059076928,0.036102567,0.01969231,0.026256412,0.04266667,0.059076928,0.068923086,0.06564103,0.04594872,0.029538464,0.01969231,0.009846155,0.0032820515,0.0,0.0032820515,0.016410258,0.026256412,0.02297436,0.013128206,0.013128206,0.01969231,0.04594872,0.072205134,0.06235898,0.052512825,0.072205134,0.1148718,0.16410258,0.190359,0.18379489,0.17066668,0.15753847,0.14441027,0.14441027,0.15097436,0.16738462,0.18707694,0.20020515,0.20020515,0.23958977,0.256,0.29210258,0.3446154,0.38400003,0.3314872,0.38728207,0.55794877,0.79097444,0.95835906,0.8205129,0.9485129,1.1158975,1.2307693,1.3522053,2.356513,4.1583595,4.890257,3.8564105,1.5491283,1.2635899,0.93866676,0.9124103,1.3161026,2.097231,2.6683078,2.8324106,2.5632823,2.2121027,2.5107694,1.6049232,1.3620514,1.8412309,3.0785644,5.07077,6.4065647,6.124308,4.8738465,3.242667,1.7263591,1.6738462,2.1070771,2.3138463,2.097231,1.785436,2.038154,2.4320002,2.4418464,2.2153847,2.609231,2.4320002,1.7460514,1.4769232,1.8642052,2.4418464,4.381539,8.113232,11.749744,13.489232,11.592206,9.705027,9.3078985,9.078155,8.208411,6.413129,7.2270775,8.572719,9.31118,9.176616,8.792616,8.214975,6.7938466,6.49518,8.395488,12.675283,14.027489,14.841437,14.191591,13.095386,14.496821,16.978052,18.153027,17.8839,16.659693,15.599591,18.048002,17.322668,16.17395,15.921232,16.466053,16.177233,16.390566,16.968206,17.522873,17.414566,13.627078,9.892103,6.9645133,4.9394875,3.2361028,2.7700515,2.7995899,3.2656412,3.9417439,4.4406157,4.1682053,3.892513,3.511795,3.1343591,3.0949745,3.4002054,4.1058464,4.827898,5.182359,4.7917953,4.345436,4.578462,5.3792825,6.449231,7.315693,7.6964107,7.9852314,7.936001,7.4765134,6.7117953,6.226052,6.058667,6.2063594,6.5772314,6.9776416,6.747898,6.482052,6.226052,5.9995904,5.8190775,0.14112821,0.18051283,0.118153855,0.049230773,0.01969231,0.006564103,0.006564103,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.009846155,0.03938462,0.04594872,0.029538464,0.006564103,0.006564103,0.01969231,0.026256412,0.016410258,0.013128206,0.013128206,0.013128206,0.013128206,0.009846155,0.01969231,0.029538464,0.10502565,0.23958977,0.42338464,0.636718,0.5513847,0.41025645,0.3249231,0.32820517,0.35446155,0.380718,0.46933338,0.48574364,0.45292312,0.5284103,0.36102566,0.26256412,0.18707694,0.1148718,0.049230773,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01969231,0.06564103,0.13456412,0.17723078,0.28225642,0.50543594,0.7384616,1.0075898,1.4867693,1.5261539,0.8730257,0.27569234,0.036102567,0.0,0.0,0.0,0.0,0.01969231,0.10502565,0.62030774,1.1815386,1.2865642,0.9911796,0.8960001,0.7778462,0.574359,0.45292312,0.51856416,0.8205129,0.71548724,0.69251287,0.7056411,0.702359,0.64000005,0.36102566,0.18379489,0.15753847,0.2231795,0.21989745,0.08861539,0.02297436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.016410258,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.032820515,0.0951795,0.23302566,0.3117949,0.28225642,0.19364104,0.118153855,0.059076928,0.03938462,0.08205129,0.2100513,0.446359,0.7450257,0.82379496,0.67282057,0.53825647,0.8336411,0.8336411,0.62030774,0.35774362,0.3249231,0.49887183,0.57764107,0.5940513,0.6465641,0.88287187,1.3981539,2.1267693,2.297436,1.6836925,0.60061544,0.41025645,0.2297436,0.20676924,0.38728207,0.7187693,0.7778462,0.72861546,0.7515898,0.892718,1.0601027,1.1454359,1.2274873,1.3259488,1.4441026,1.5655385,1.9856411,2.0545642,1.8084104,1.4145643,1.1913847,1.339077,1.3095386,1.1355898,0.9517949,1.0108719,0.955077,0.9616411,0.97805136,0.9911796,1.0272821,1.0338463,0.90912825,0.82379496,0.90256417,1.2012309,1.2274873,1.3161026,1.4802053,1.6738462,1.8051283,1.6935385,1.591795,1.467077,1.3620514,1.4112822,1.4408206,1.4572309,1.4408206,1.3817437,1.2635899,1.1946667,1.0601027,0.9419488,0.86646163,0.7844103,0.69907695,0.5940513,0.48246157,0.37743592,0.28882053,0.28882053,0.33476925,0.42338464,0.48902568,0.4266667,0.43651286,0.39712822,0.3314872,0.31507695,0.48574364,0.7253334,0.8467693,0.85005134,0.827077,0.9419488,1.0075898,0.69251287,0.46933338,0.52512825,0.7417436,0.79097444,0.6498462,0.56451285,0.6170257,0.74830776,0.5349744,0.6498462,0.90256417,1.1355898,1.1946667,0.81394875,0.51856416,0.38728207,0.44964105,0.67610264,0.85005134,1.0043077,1.1848207,1.3751796,1.5195899,1.5819489,1.467077,1.2570257,1.0502565,0.9747693,1.1027694,1.0469744,1.0108719,1.024,0.9517949,0.44964105,0.20348719,0.108307704,0.08205129,0.04594872,0.052512825,0.11158975,0.15753847,0.16082053,0.128,0.15753847,0.06564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.02297436,0.026256412,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.0032820515,0.0,0.0032820515,0.006564103,0.0032820515,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0032820515,0.01969231,0.04266667,0.06235898,0.052512825,0.059076928,0.07548718,0.10502565,0.15097436,0.17723078,0.18707694,0.18379489,0.18707694,0.24287182,0.23630771,0.17394873,0.09189744,0.029538464,0.02297436,0.026256412,0.01969231,0.016410258,0.026256412,0.032820515,0.055794876,0.07548718,0.08205129,0.08861539,0.0951795,0.108307704,0.07876924,0.049230773,0.03938462,0.049230773,0.08205129,0.10502565,0.1148718,0.118153855,0.12143591,0.07876924,0.059076928,0.04594872,0.032820515,0.029538464,0.036102567,0.03938462,0.04594872,0.052512825,0.055794876,0.055794876,0.03938462,0.01969231,0.009846155,0.009846155,0.02297436,0.029538464,0.029538464,0.026256412,0.006564103,0.006564103,0.01969231,0.052512825,0.08861539,0.1148718,0.15425642,0.22646156,0.30194873,0.35446155,0.33805132,0.28882053,0.23630771,0.20020515,0.20348719,0.256,0.3052308,0.3249231,0.318359,0.30194873,0.29538465,0.34133336,0.3511795,0.4004103,0.49887183,0.574359,0.5284103,0.5316923,0.60061544,0.7384616,0.9353847,0.79425645,0.764718,0.77128214,0.81394875,0.97805136,1.463795,2.3236926,2.8521028,2.540308,1.0601027,0.83035904,0.6268718,0.5316923,0.61374366,0.8992821,1.270154,1.2307693,1.2307693,1.4276924,1.7001027,1.4211283,1.1848207,1.211077,1.6836925,2.733949,3.0523078,2.7536411,2.2055387,1.657436,1.2570257,1.5195899,1.8182565,1.7952822,1.4998976,1.401436,1.2209232,1.2832822,1.4933335,1.8642052,2.5435898,2.3663592,2.484513,2.169436,1.6672822,2.1956925,3.9581542,7.709539,10.66995,10.971898,7.650462,5.8092313,7.00718,8.136206,7.643898,5.5204105,4.8114877,5.4613338,6.445949,7.322257,8.234667,8.766359,8.342975,9.238976,12.028719,15.589745,14.628103,12.891898,11.556104,11.1294365,11.45436,12.6063595,15.602873,18.402462,19.797335,19.419899,18.330257,15.832617,14.204719,14.582155,16.971489,19.242668,18.914463,17.578669,16.554668,16.89272,13.184001,9.603283,7.384616,6.4754877,5.5171285,4.3585644,3.754667,3.7120004,4.161641,4.9362054,4.5522056,4.013949,3.4888208,3.1409233,3.1376412,3.3608208,3.6890259,4.1780515,4.6769233,4.850872,4.3290257,4.525949,5.0609236,5.7534366,6.6067696,7.1122055,7.640616,7.9130263,7.8080006,7.3649235,6.9382567,6.99077,7.2303596,7.496206,7.75877,7.4371285,6.875898,6.311385,5.8781543,5.5762057,0.128,0.18051283,0.15097436,0.08205129,0.01969231,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.026256412,0.03938462,0.026256412,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.013128206,0.01969231,0.016410258,0.02297436,0.013128206,0.02297436,0.055794876,0.14112821,0.29538465,0.30194873,0.20348719,0.108307704,0.072205134,0.108307704,0.2100513,0.29210258,0.3117949,0.318359,0.4594872,0.33476925,0.256,0.190359,0.12143591,0.06235898,0.02297436,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.026256412,0.02297436,0.0,0.0,0.0,0.0,0.0,0.0,0.036102567,0.055794876,0.16738462,0.48902568,1.1618463,0.65641034,0.28882053,0.08205129,0.006564103,0.0,0.0,0.0,0.0,0.013128206,0.072205134,0.29538465,0.7220513,0.90912825,0.88615394,1.1585642,0.93866676,0.5973334,0.37743592,0.4201026,0.74830776,0.7220513,0.7811283,0.7778462,0.6465641,0.4201026,0.256,0.15753847,0.13784617,0.16410258,0.16410258,0.06235898,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.009846155,0.01969231,0.026256412,0.049230773,0.15753847,0.256,0.29538465,0.25271797,0.15425642,0.055794876,0.01969231,0.052512825,0.118153855,0.17723078,0.48246157,0.67282057,0.65312827,0.5973334,0.8402052,0.8041026,0.574359,0.32820517,0.31507695,0.47917953,0.4660513,0.42338464,0.45620516,0.62030774,1.0929232,1.5130258,1.4802053,0.92553854,0.118153855,0.08861539,0.068923086,0.14769232,0.32164106,0.512,0.5874872,0.5316923,0.512,0.56451285,0.6071795,0.43323082,0.33805132,0.318359,0.43651286,0.827077,1.276718,1.3784616,1.1815386,0.88615394,0.8730257,1.2307693,1.7788719,1.8871796,1.6311796,1.7920002,1.5983591,1.5163078,1.4506668,1.3686155,1.273436,1.2077949,1.2340513,1.4802053,1.7788719,1.6607181,1.463795,1.6607181,2.0086155,2.2186668,1.9528207,1.8707694,1.782154,1.6508719,1.522872,1.5425643,1.5622566,1.5622566,1.5327181,1.463795,1.3423591,1.1815386,1.0765129,0.9944616,0.9124103,0.8205129,0.764718,0.7318975,0.702359,0.6498462,0.55794877,0.39384618,0.37743592,0.5152821,0.6892308,0.6465641,0.54482055,0.42994875,0.37415388,0.4660513,0.8041026,1.3522053,1.585231,1.4276924,1.0371283,0.8336411,0.88287187,0.77128214,0.78769237,0.9878975,1.1979488,1.014154,0.88287187,0.97805136,1.2406155,1.3751796,1.017436,1.0075898,1.1355898,1.2406155,1.1848207,0.78769237,0.56451285,0.42338464,0.37743592,0.53825647,0.78769237,0.95835906,1.2209232,1.5491283,1.719795,1.6935385,1.4211283,1.0962052,0.8730257,0.86974365,0.8336411,0.72861546,0.65641034,0.6104616,0.48246157,0.15425642,0.029538464,0.0,0.009846155,0.04594872,0.052512825,0.13128206,0.19364104,0.21661541,0.21989745,0.14769232,0.052512825,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.013128206,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.006564103,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.01969231,0.01969231,0.009846155,0.009846155,0.009846155,0.016410258,0.04594872,0.07876924,0.12471796,0.14769232,0.14441027,0.17723078,0.190359,0.16410258,0.11158975,0.055794876,0.016410258,0.016410258,0.009846155,0.016410258,0.032820515,0.03938462,0.052512825,0.072205134,0.08533334,0.09189744,0.08861539,0.11158975,0.08205129,0.04594872,0.029538464,0.02297436,0.03938462,0.055794876,0.068923086,0.07876924,0.098461546,0.072205134,0.06235898,0.055794876,0.049230773,0.029538464,0.029538464,0.029538464,0.032820515,0.03938462,0.04266667,0.06564103,0.068923086,0.055794876,0.03938462,0.032820515,0.06235898,0.052512825,0.032820515,0.016410258,0.013128206,0.032820515,0.032820515,0.055794876,0.11158975,0.17723078,0.29538465,0.47589746,0.64000005,0.7187693,0.6432821,0.5316923,0.446359,0.36758977,0.30851284,0.318359,0.3511795,0.380718,0.39712822,0.40697438,0.44964105,0.5874872,0.6104616,0.60389745,0.6235898,0.69579494,0.67282057,0.6235898,0.5874872,0.6170257,0.77128214,0.75487185,0.63343596,0.508718,0.47261542,0.60389745,0.79097444,1.0371283,1.2438976,1.2176411,0.67282057,0.48574364,0.40697438,0.36430773,0.3446154,0.38728207,0.508718,0.57764107,0.65969235,0.77128214,0.892718,1.1782565,1.2209232,1.1684103,1.2438976,1.7329233,1.4834872,1.1946667,0.9616411,0.8369231,0.84348726,1.014154,1.1093334,1.0371283,0.8960001,0.9616411,0.73517954,0.8369231,1.204513,1.7788719,2.5074873,2.7536411,3.3608208,2.9735386,1.8970258,2.1070771,3.308308,6.5772314,8.418462,7.4929237,4.6112823,3.7185643,4.923077,6.3376417,6.5870776,4.788513,3.8301542,3.6824617,4.0303593,4.775385,6.0291286,7.3583593,8.04759,9.6525135,12.20595,14.230975,12.166565,10.072617,9.540924,10.210463,9.7673855,8.864821,10.249847,12.796719,15.159796,15.780104,14.04718,13.13477,12.724514,13.08554,15.074463,17.257027,17.001026,15.868719,15.300924,16.630156,11.264001,7.653744,6.2916927,6.5870776,6.87918,5.7009234,4.450462,3.636513,3.7120004,5.0543594,4.906667,3.8465643,2.92759,2.6157951,2.7700515,3.190154,3.515077,3.8695388,4.348718,5.031385,4.4865646,4.4045134,4.5522056,4.886975,5.5565133,6.0783596,6.6461544,7.1023593,7.318975,7.204103,7.1548724,7.3714876,7.6143594,7.8112826,8.067283,7.906462,7.3321033,6.626462,5.9963083,5.605744,0.13128206,0.18379489,0.19364104,0.13128206,0.04266667,0.026256412,0.006564103,0.0032820515,0.0032820515,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016410258,0.029538464,0.032820515,0.01969231,0.016410258,0.006564103,0.0032820515,0.0,0.0032820515,0.0032820515,0.016410258,0.02297436,0.01969231,0.049230773,0.036102567,0.016410258,0.0032820515,0.0032820515,0.02297436,0.06235898,0.049230773,0.01969231,0.0032820515,0.0032820515,0.009846155,0.01969231,0.06235898,0.14769232,0.24943592,0.24943592,0.19692309,0.128,0.072205134,0.049230773,0.032820515,0.013128206,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.029538464,0.055794876,0.052512825,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.026256412,0.098461546,0.21989745,0.4397949,0.86317956,0.65969235,0.36102566,0.16738462,0.1148718,0.059076928,0.14769232,0.45292312,0.7253334,0.81066674,0.63343596,0.5874872,0.38728207,0.20020515,0.101743594,0.06564103,0.01969231,0.009846155,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.02297436,0.036102567,0.049230773,0.04594872,0.072205134,0.10502565,0.128,0.13784617,0.15753847,0.118153855,0.04266667,0.0,0.0,0.0,0.0,0.0,0.0,0.04266667,0.20676924,0.26584616,0.2297436,0.14769232,0.06235898,0.02297436,0.04266667,0.04266667,0.036102567,0.02297436,0.013128206,0.052512825,0.068923086,0.04594872,0.009846155,0.02297436,0.18379489,0.26912823,0.40697438,0.62030774,0.83035904,0.78769237,0.5874872,0.35446155,0.190359,0.18707694,0.14769232,0.18051283,0.20348719,0.20676924,0.2231795,0.22646156,0.24615386,0.25928208,0.27569234,0.3314872,0.7122052,1.7985642,2.2744617,2.0676925,2.3302567,2.156308,1.975795,1.8051283,1.6344616,1.4408206,1.2931283,1.5556924,2.1989746,2.6584618,1.8215386,1.3423591,1.7066668,2.2022567,2.2416413,1.3620514,1.4572309,1.4506668,1.4145643,1.394872,1.4145643,1.4572309,1.4703591,1.4506668,1.3915899,1.2800001,1.1158975,1.0568206,1.020718,0.9616411,0.88615394,0.8402052,0.8533334,0.8992821,0.92553854,0.8467693,0.49887183,0.35774362,0.46933338,0.7056411,0.761436,0.5513847,0.4135385,0.40697438,0.5940513,1.014154,1.8379488,2.1366155,1.7755898,0.9714873,0.27569234,0.31507695,0.571077,0.9156924,1.2471796,1.4933335,1.1881026,1.1224617,1.4375386,1.9265642,2.0217438,1.6738462,1.404718,1.2898463,1.2537436,1.0502565,0.6826667,0.60389745,0.53825647,0.46276927,0.6268718,0.7844103,0.86317956,1.0765129,1.4309745,1.7296412,1.3193847,0.97805136,0.69579494,0.55794877,0.75487185,0.44307697,0.36102566,0.3117949,0.22646156,0.15097436,0.14769232,0.059076928,0.0,0.0,0.0,0.0,0.052512825,0.13456412,0.20348719,0.18379489,0.036102567,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0032820515,0.013128206,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01969231,0.09189744,0.15097436,0.17394873,0.20020515,0.17066668,0.13456412,0.11158975,0.08861539,0.02297436,0.013128206,0.013128206,0.01969231,0.026256412,0.02297436,0.04266667,0.072205134,0.09189744,0.08205129,0.06564103,0.059076928,0.04266667,0.029538464,0.02297436,0.016410258,0.013128206,0.02297436,0.032820515,0.04266667,0.055794876,0.06564103,0.06235898,0.059076928,0.052512825,0.026256412,0.029538464,0.029538464,0.029538464,0.029538464,0.02297436,0.052512825,0.09189744,0.098461546,0.072205134,0.06564103,0.09189744,0.068923086,0.032820515,0.006564103,0.02297436,0.072205134,0.06235898,0.08205129,0.15097436,0.2100513,0.3446154,0.60061544,0.84348726,0.9616411,0.8566154,0.7089231,0.62030774,0.5021539,0.35446155,0.25271797,0.23302566,0.27241027,0.34133336,0.42338464,0.5284103,0.7417436,0.7811283,0.702359,0.6170257,0.71548724,0.71548724,0.6465641,0.56123084,0.51856416,0.574359,0.7318975,0.65969235,0.47589746,0.3249231,0.36430773,0.41025645,0.42994875,0.47589746,0.54482055,0.5677949,0.36430773,0.31507695,0.3314872,0.33805132,0.28225642,0.21989745,0.2297436,0.2986667,0.4397949,0.6662565,0.9714873,1.2340513,1.3292309,1.3751796,1.723077,1.3653334,0.99774367,0.702359,0.5284103,0.48246157,0.47917953,0.44307697,0.39712822,0.39384618,0.48574364,0.55794877,0.71548724,1.0305642,1.5458462,2.2678976,3.2131286,3.6890259,3.2164104,2.162872,1.7394873,2.2777438,4.388103,5.3858466,4.7261543,4.010667,4.4800005,3.7316926,3.7874875,4.5456414,3.767795,4.0434875,3.889231,3.7284105,3.8301542,4.315898,4.97559,5.7403083,6.925129,8.434873,9.764103,8.55959,8.700719,9.856001,11.021129,10.532104,8.083693,6.2490263,5.58277,6.0816417,7.194257,8.139488,9.619693,10.548513,10.640411,10.404103,10.236719,10.748719,12.3076935,14.752822,17.38831,10.295795,6.6461544,5.605744,6.2129235,7.394462,6.9152827,5.2480006,3.7973337,3.8006158,6.3179493,5.865026,4.017231,2.5665643,2.1924105,2.4713848,3.1015387,3.761231,4.2240005,4.6276927,5.467898,5.1200004,4.6211286,4.2994876,4.315898,4.670359,5.156103,5.6976414,6.2227697,6.619898,6.7216415,7.1515903,7.394462,7.5585647,7.752206,8.090257,8.109949,7.7325134,7.0465646,6.370462,6.23918,0.108307704,0.37415388,0.26912823,0.13456412,0.101743594,0.07548718,0.016410258,0.009846155,0.016410258,0.016410258,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.04594872,0.0951795,0.1148718,0.09189744,0.029538464,0.016410258,0.009846155,0.0032820515,0.016410258,0.016410258,0.016410258,0.009846155,0.0,0.0,0.036102567,0.026256412,0.009846155,0.0,0.0,0.0,0.01969231,0.02297436,0.016410258,0.016410258,0.0032820515,0.0,0.0,0.006564103,0.029538464,0.029538464,0.02297436,0.016410258,0.013128206,0.0,0.013128206,0.016410258,0.016410258,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.016410258,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.03938462,0.118153855,0.28225642,0.4135385,0.2297436,0.48574364,0.39384618,0.28225642,0.26584616,0.2297436,0.14441027,0.10502565,0.22646156,0.574359,1.1585642,1.5622566,1.1520001,0.6301539,0.3249231,0.15097436,0.055794876,0.049230773,0.036102567,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02297436,0.059076928,0.068923086,0.059076928,0.04594872,0.032820515,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.016410258,0.013128206,0.0,0.013128206,0.032820515,0.03938462,0.049230773,0.12143591,0.9156924,1.0962052,0.90584624,0.6104616,0.48902568,0.56123084,0.5152821,0.3249231,0.101743594,0.07548718,0.07548718,0.10502565,0.18379489,0.27241027,0.25928208,0.18707694,0.17723078,0.21989745,0.27241027,0.25928208,0.25928208,0.29538465,0.43651286,0.6465641,0.79425645,1.0371283,1.3718976,1.5195899,1.5130258,1.7099489,1.6114873,1.394872,1.3456411,1.467077,1.4802053,1.3226668,1.3653334,1.5031796,1.5819489,1.3718976,1.5064616,1.5031796,1.4441026,1.3784616,1.3423591,1.3554872,1.3686155,1.3423591,1.2800001,1.204513,1.1191796,1.0436924,0.98133343,0.9353847,0.88615394,0.8598975,0.8172308,0.7318975,0.6268718,0.56451285,0.6859488,0.7089231,0.58092314,0.3708718,0.27569234,0.39712822,0.49887183,0.6235898,0.8172308,1.1585642,2.0644104,2.15959,1.6311796,0.82379496,0.27569234,0.4201026,0.6695385,0.73517954,0.74830776,1.2373334,1.4178462,1.2274873,1.2209232,1.5458462,1.9364104,1.9495386,1.7329233,1.5064616,1.404718,1.463795,1.2340513,0.9288206,0.78769237,0.86974365,1.0535386,1.017436,0.84348726,0.761436,0.9124103,1.3259488,0.7417436,0.38400003,0.190359,0.108307704,0.108307704,0.02297436,0.04594872,0.04594872,0.026256412,0.13784617,0.026256412,0.0,0.0,0.0,0.0,0.0,0.0,0.02297436,0.049230773,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.016410258,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.04594872,0.16082053,0.2986667,0.33476925,0.27569234,0.20348719,0.16082053,0.13128206,0.04594872,0.009846155,0.0,0.006564103,0.013128206,0.0,0.036102567,0.072205134,0.08533334,0.07548718,0.07548718,0.052512825,0.036102567,0.01969231,0.0032820515,0.016410258,0.0032820515,0.009846155,0.016410258,0.01969231,0.029538464,0.04266667,0.04594872,0.04594872,0.03938462,0.016410258,0.026256412,0.029538464,0.029538464,0.032820515,0.04594872,0.059076928,0.068923086,0.068923086,0.06564103,0.09189744,0.06564103,0.032820515,0.016410258,0.013128206,0.0,0.049230773,0.08861539,0.13784617,0.18707694,0.19692309,0.13784617,0.21333335,0.35446155,0.47917953,0.5021539,0.44307697,0.35446155,0.256,0.16738462,0.108307704,0.108307704,0.108307704,0.15097436,0.2231795,0.25928208,0.29538465,0.36102566,0.39712822,0.446359,0.64000005,0.64000005,0.6301539,0.60061544,0.56123084,0.5481026,0.8533334,1.0962052,0.9124103,0.44964105,0.3511795,0.33805132,0.3446154,0.40697438,0.50543594,0.58092314,0.4955898,0.41025645,0.36102566,0.35446155,0.36758977,0.256,0.20020515,0.19692309,0.23958977,0.33476925,0.36102566,0.29210258,0.256,0.27241027,0.25928208,0.3708718,0.50543594,0.574359,0.5677949,0.58092314,0.6170257,0.6268718,0.60061544,0.6071795,0.7778462,0.8992821,0.8205129,0.8566154,1.1093334,1.4506668,2.0250258,2.422154,2.4057438,2.044718,1.7394873,1.4112822,1.5753847,2.1366155,3.1081028,4.6080003,5.546667,4.667077,3.895795,3.8531284,3.8301542,4.9526157,4.821334,4.7556925,5.097026,5.218462,4.315898,3.7973337,4.7425647,7.1056414,9.705027,7.9228725,7.604513,8.320001,9.409642,9.993847,9.432616,8.891078,9.065026,9.7214365,9.6754875,10.246565,9.970873,9.636104,9.340718,8.500513,7.9491286,9.416205,12.2847185,15.2155905,16.144411,11.346052,8.490667,7.282872,7.50277,9.019077,9.019077,7.1680007,5.7042055,6.498462,11.076924,7.939283,5.2611284,3.6693337,3.2032824,3.3247182,3.692308,4.397949,5.149539,5.7731285,6.226052,6.629744,6.1440005,5.287385,4.571898,4.4865646,4.8771286,5.4153852,6.0192823,6.491898,6.514872,6.941539,7.3714876,7.6767187,7.834257,7.9195905,7.821129,7.568411,7.1220517,6.872616,7.6307697,0.508718,0.6301539,0.6268718,0.60389745,0.5316923,0.23630771,0.10502565,0.03938462,0.009846155,0.0032820515,0.0032820515,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.02297436,0.036102567,0.029538464,0.009846155,0.0032820515,0.0032820515,0.0,0.0032820515,0.0032820515,0.0032820515,0.0032820515,0.0,0.0,0.006564103,0.006564103,0.0032820515,0.0,0.0,0.0,0.0032820515,0.01969231,0.03938462,0.03938462,0.026256412,0.03938462,0.03938462,0.01969231,0.006564103,0.006564103,0.013128206,0.009846155,0.0032820515,0.0,0.013128206,0.006564103,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.016410258,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.036102567,0.08205129,0.1148718,0.1148718,0.059076928,0.14769232,0.13128206,0.09189744,0.06235898,0.04594872,0.029538464,0.029538464,0.07548718,0.21661541,0.5021539,0.72861546,0.5349744,0.2855385,0.13784617,0.055794876,0.016410258,0.009846155,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.016410258,0.02297436,0.036102567,0.04266667,0.02297436,0.01969231,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.15425642,0.24943592,0.19692309,0.049230773,0.06235898,0.068923086,0.059076928,0.08861539,0.26912823,0.60389745,0.64000005,0.49230772,0.29210258,0.15753847,0.15425642,0.12471796,0.098461546,0.08205129,0.07548718,0.28225642,0.36758977,0.39384618,0.41025645,0.4660513,0.5513847,0.48574364,0.46276927,0.4660513,0.24615386,0.24615386,0.27569234,0.32820517,0.42338464,0.6104616,0.81394875,0.9517949,0.9419488,0.8598975,0.9288206,1.2012309,1.1782565,1.1257436,1.1782565,1.3587693,1.276718,1.3554872,1.6180514,1.8313848,1.5064616,1.7591796,1.7920002,1.657436,1.4834872,1.4769232,1.4605129,1.3686155,1.4080001,1.4998976,1.2800001,1.086359,0.94523084,0.85005134,0.7811283,0.71548724,0.65969235,0.764718,0.9485129,1.1224617,1.1979488,0.82379496,0.5874872,0.56123084,0.71548724,0.92225647,1.014154,1.0371283,1.2668719,1.7591796,2.356513,3.05559,2.8882053,2.0742567,1.0305642,0.38400003,0.39384618,0.58420515,0.7844103,0.9321026,1.0765129,1.3587693,1.3423591,1.1684103,1.0043077,1.0699488,1.1815386,1.5163078,1.4309745,1.0108719,1.0633847,0.95835906,0.77128214,0.64000005,0.57764107,0.4660513,0.4201026,0.53825647,0.5907693,0.48574364,0.26584616,0.14769232,0.09189744,0.06235898,0.03938462,0.02297436,0.0032820515,0.009846155,0.009846155,0.006564103,0.026256412,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0032820515,0.013128206,0.013128206,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.006564103,0.0032820515,0.013128206,0.013128206,0.013128206,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.08205129,0.20676924,0.3117949,0.25928208,0.16410258,0.10502565,0.098461546,0.068923086,0.02297436,0.0032820515,0.0,0.0032820515,0.013128206,0.029538464,0.03938462,0.04594872,0.052512825,0.052512825,0.036102567,0.02297436,0.009846155,0.0032820515,0.016410258,0.0032820515,0.0032820515,0.0032820515,0.0032820515,0.006564103,0.009846155,0.02297436,0.032820515,0.036102567,0.03938462,0.032820515,0.029538464,0.036102567,0.049230773,0.068923086,0.06235898,0.03938462,0.029538464,0.03938462,0.055794876,0.049230773,0.029538464,0.016410258,0.01969231,0.036102567,0.055794876,0.101743594,0.14112821,0.14769232,0.101743594,0.08861539,0.13456412,0.19692309,0.24943592,0.28225642,0.26256412,0.22646156,0.17723078,0.128,0.108307704,0.098461546,0.08861539,0.08205129,0.08205129,0.08861539,0.10502565,0.14441027,0.19364104,0.26584616,0.3708718,0.4594872,0.5546667,0.67938465,0.79425645,0.7811283,0.73517954,0.6892308,0.5907693,0.46933338,0.44964105,0.4266667,0.5021539,0.5874872,0.65312827,0.7253334,0.7384616,0.71548724,0.60061544,0.45292312,0.4135385,0.2855385,0.23302566,0.21333335,0.20676924,0.22646156,0.28882053,0.2986667,0.2855385,0.27241027,0.27241027,0.3708718,0.45620516,0.5021539,0.52512825,0.5546667,0.58092314,0.574359,0.54482055,0.5316923,0.5940513,0.7450257,0.8369231,0.9747693,1.214359,1.5360001,1.8149745,2.1431797,2.5304618,2.6945643,2.0578463,1.3554872,1.2307693,1.3587693,1.6180514,2.0939488,2.5271797,2.8947694,3.4625645,4.066462,4.1091285,2.937436,3.3411283,4.57518,6.114462,7.6242056,6.76759,5.208616,4.1091285,4.5554876,7.5552826,10.033232,10.755282,10.627283,10.397539,10.689642,10.791386,11.234463,11.306667,10.988309,10.981745,12.091078,11.221334,9.895386,9.80677,12.832822,13.397334,12.898462,13.072412,13.863386,13.433437,11.585642,10.059488,9.133949,8.89436,9.225847,8.697436,7.3091288,6.803693,7.318975,7.4043083,5.4383593,3.7021542,2.868513,2.9046156,3.0949745,3.6168208,4.345436,5.1364107,5.943795,6.8233852,6.7183595,6.3179493,5.7632823,5.2447186,5.0215387,5.080616,5.425231,5.9470773,6.452513,6.6625648,6.961231,7.24677,7.4863596,7.6570263,7.762052,8.083693,7.650462,6.954667,6.560821,7.0925136,0.7384616,0.73517954,0.8172308,0.95835906,0.9944616,0.6235898,0.39384618,0.20348719,0.08205129,0.02297436,0.009846155,0.006564103,0.0032820515,0.0,0.0,0.0,0.0,0.006564103,0.006564103,0.0032820515,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.006564103,0.009846155,0.013128206,0.013128206,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.01969231,0.01969231,0.029538464,0.03938462,0.032820515,0.01969231,0.009846155,0.0032820515,0.0032820515,0.0032820515,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0,0.006564103,0.0032820515,0.0,0.0,0.0,0.006564103,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.029538464,0.04266667,0.036102567,0.016410258,0.006564103,0.026256412,0.026256412,0.016410258,0.006564103,0.009846155,0.098461546,0.15097436,0.190359,0.27241027,0.46276927,0.6104616,0.39712822,0.16738462,0.059076928,0.02297436,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.036102567,0.108307704,0.21661541,0.24287182,0.16082053,0.04266667,0.04266667,0.07548718,0.08861539,0.06564103,0.04266667,0.01969231,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06564103,0.3446154,0.51856416,0.41682056,0.04266667,0.055794876,0.059076928,0.068923086,0.098461546,0.15753847,0.26256412,0.26912823,0.2100513,0.1148718,0.029538464,0.036102567,0.08533334,0.12471796,0.128,0.08533334,0.2100513,0.36430773,0.48246157,0.51856416,0.446359,0.43651286,0.42338464,0.39056414,0.35446155,0.3708718,0.29210258,0.19364104,0.19692309,0.3117949,0.45620516,0.51856416,0.5546667,0.54482055,0.55794877,0.7417436,0.83035904,0.7318975,0.7089231,0.86646163,1.1454359,0.98133343,0.9419488,1.0962052,1.2832822,1.1191796,1.2176411,1.2635899,1.2471796,1.1946667,1.1716924,1.1191796,1.0732309,1.079795,1.1126155,1.0765129,0.9616411,0.80738467,0.72861546,0.7220513,0.6629744,0.5513847,0.56123084,0.6826667,0.8369231,0.8730257,0.69579494,0.62030774,0.6662565,0.8205129,1.0272821,1.2537436,1.3883078,1.7493335,2.4024618,3.186872,3.5610259,3.186872,2.5009232,1.8674873,1.5458462,1.529436,1.273436,1.142154,1.2274873,1.3751796,1.6508719,1.7033848,1.4342566,1.0371283,0.9747693,0.8960001,0.9189744,0.85005134,0.7122052,0.761436,0.5973334,0.45292312,0.34133336,0.26584616,0.2297436,0.25928208,0.3052308,0.27241027,0.15097436,0.0,0.006564103,0.009846155,0.016410258,0.026256412,0.04594872,0.02297436,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.0032820515,0.0,0.006564103,0.016410258,0.016410258,0.006564103,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.009846155,0.006564103,0.0,0.006564103,0.006564103,0.0032820515,0.0032820515,0.016410258,0.016410258,0.01969231,0.02297436,0.016410258,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.02297436,0.08205129,0.15753847,0.30851284,0.3511795,0.32164106,0.25271797,0.20348719,0.08205129,0.026256412,0.013128206,0.016410258,0.016410258,0.013128206,0.013128206,0.01969231,0.026256412,0.026256412,0.016410258,0.009846155,0.0032820515,0.0032820515,0.016410258,0.009846155,0.013128206,0.01969231,0.01969231,0.026256412,0.006564103,0.006564103,0.01969231,0.032820515,0.036102567,0.032820515,0.026256412,0.026256412,0.03938462,0.059076928,0.052512825,0.029538464,0.02297436,0.032820515,0.036102567,0.036102567,0.02297436,0.01969231,0.032820515,0.06564103,0.09189744,0.0951795,0.098461546,0.108307704,0.11158975,0.128,0.16082053,0.20020515,0.2297436,0.2297436,0.19364104,0.15753847,0.118153855,0.08205129,0.068923086,0.06564103,0.072205134,0.068923086,0.055794876,0.055794876,0.06564103,0.098461546,0.14112821,0.18707694,0.21333335,0.30194873,0.38728207,0.5316923,0.7089231,0.83035904,0.69579494,0.5907693,0.50543594,0.44307697,0.43651286,0.6104616,0.8467693,0.9747693,0.93866676,0.8008206,0.81394875,0.8369231,0.7581539,0.5907693,0.48246157,0.4135385,0.4266667,0.40697438,0.33805132,0.318359,0.37743592,0.4004103,0.4201026,0.44964105,0.4955898,0.5415385,0.56123084,0.5546667,0.5284103,0.47589746,0.44964105,0.46933338,0.5152821,0.571077,0.61374366,0.73517954,0.8730257,1.0502565,1.2209232,1.2832822,1.3718976,1.6902566,2.1398976,2.4057438,1.9364104,1.3620514,1.142154,1.1191796,1.204513,1.3653334,1.4408206,1.7033848,2.681436,4.161641,5.1954875,3.4822567,3.4560003,4.44718,5.874872,7.2631803,6.5969234,5.4843082,4.516103,4.381539,5.85518,7.9327188,8.710565,8.973129,9.170052,9.426052,11.145847,11.867898,12.544001,13.282462,13.348104,13.105232,12.475078,11.467488,10.564924,10.738873,11.090053,10.512411,10.870154,11.9860525,11.648001,10.282667,8.953437,8.464411,8.644924,8.352821,8.257642,7.857231,8.067283,8.395488,6.9349747,4.893539,3.190154,2.3827693,2.428718,2.678154,3.1081028,3.7087183,4.46359,5.5532312,7.3386674,7.312411,6.8299494,6.196513,5.674667,5.504,5.467898,5.6385646,5.943795,6.2884107,6.550975,6.741334,6.921847,7.0793853,7.2664623,7.6012316,7.824411,7.4043083,6.8496413,6.5017443,6.547693,1.4145643,1.1191796,1.4900514,1.7001027,1.5031796,1.2570257,1.0994873,0.80738467,0.52512825,0.30194873,0.108307704,0.029538464,0.0032820515,0.0,0.0,0.0,0.0,0.006564103,0.006564103,0.006564103,0.016410258,0.006564103,0.006564103,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.026256412,0.029538464,0.013128206,0.006564103,0.006564103,0.006564103,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01969231,0.029538464,0.029538464,0.026256412,0.026256412,0.016410258,0.0032820515,0.0,0.0,0.0,0.009846155,0.013128206,0.013128206,0.009846155,0.0,0.006564103,0.006564103,0.009846155,0.016410258,0.006564103,0.01969231,0.016410258,0.013128206,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.02297436,0.016410258,0.006564103,0.0,0.0,0.0,0.0,0.0,0.006564103,0.032820515,0.27897438,0.41025645,0.5152821,0.7318975,1.2570257,1.9561027,1.910154,1.2832822,0.508718,0.28225642,0.15097436,0.068923086,0.02297436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.006564103,0.006564103,0.006564103,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0032820515,0.029538464,0.108307704,0.20348719,0.18379489,0.24615386,0.3052308,0.28225642,0.16738462,0.04266667,0.049230773,0.0951795,0.13128206,0.118153855,0.055794876,0.01969231,0.0032820515,0.0032820515,0.009846155,0.01969231,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.072205134,0.27569234,0.4004103,0.3249231,0.01969231,0.026256412,0.026256412,0.052512825,0.08533334,0.072205134,0.068923086,0.068923086,0.06564103,0.04594872,0.006564103,0.068923086,0.34789747,0.49887183,0.41025645,0.21333335,0.21661541,0.4004103,0.6268718,0.7515898,0.60389745,0.4201026,0.36430773,0.3117949,0.30851284,0.574359,0.512,0.28882053,0.24287182,0.36430773,0.28225642,0.30194873,0.3446154,0.39056414,0.46933338,0.636718,0.5940513,0.571077,0.6432821,0.79425645,0.8992821,0.702359,0.56451285,0.5677949,0.6695385,0.6859488,0.6859488,0.7187693,0.764718,0.827077,0.94523084,0.8467693,0.892718,0.9189744,0.88615394,0.86317956,0.83035904,0.7187693,0.6892308,0.7417436,0.73517954,0.5973334,0.5218462,0.56451285,0.7089231,0.8467693,1.0305642,0.9321026,0.9353847,1.1618463,1.4802053,1.5786668,1.585231,1.7952822,2.294154,2.9407182,2.868513,2.605949,2.3302567,2.2153847,2.4320002,2.3893335,1.9495386,1.6246156,1.5556924,1.5097437,1.6213335,1.7591796,1.5721027,1.1290257,0.92553854,0.6859488,0.44964105,0.3708718,0.42338464,0.4004103,0.36430773,0.23302566,0.1148718,0.06564103,0.101743594,0.15753847,0.13784617,0.068923086,0.0,0.0,0.013128206,0.013128206,0.013128206,0.02297436,0.04594872,0.02297436,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.0032820515,0.0,0.0032820515,0.009846155,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.006564103,0.013128206,0.013128206,0.0,0.013128206,0.013128206,0.009846155,0.006564103,0.009846155,0.009846155,0.01969231,0.032820515,0.04266667,0.03938462,0.013128206,0.0032820515,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.009846155,0.04266667,0.21989745,0.3511795,0.380718,0.32820517,0.26584616,0.13456412,0.08205129,0.07548718,0.072205134,0.02297436,0.0032820515,0.006564103,0.013128206,0.016410258,0.016410258,0.006564103,0.0032820515,0.0032820515,0.016410258,0.03938462,0.06564103,0.04266667,0.02297436,0.026256412,0.032820515,0.013128206,0.009846155,0.01969231,0.029538464,0.029538464,0.026256412,0.016410258,0.016410258,0.026256412,0.03938462,0.03938462,0.026256412,0.01969231,0.02297436,0.02297436,0.01969231,0.013128206,0.016410258,0.032820515,0.068923086,0.101743594,0.0951795,0.09189744,0.118153855,0.18051283,0.190359,0.21661541,0.24615386,0.256,0.2231795,0.17394873,0.128,0.098461546,0.08205129,0.07548718,0.07548718,0.08205129,0.08861539,0.09189744,0.09189744,0.0951795,0.14112821,0.20020515,0.24287182,0.22646156,0.22646156,0.24287182,0.32164106,0.48246157,0.7089231,0.7187693,0.6268718,0.5152821,0.44964105,0.4660513,0.7417436,1.017436,1.1454359,1.0699488,0.8172308,0.7975385,0.9747693,1.024,0.88943595,0.7811283,0.69251287,0.69907695,0.6498462,0.51856416,0.39056414,0.41025645,0.42994875,0.47917953,0.53825647,0.5677949,0.56123084,0.57764107,0.5907693,0.56123084,0.43323082,0.36758977,0.38728207,0.446359,0.51856416,0.5940513,0.7318975,0.8467693,0.93866676,0.9714873,0.88615394,0.90256417,1.1881026,1.5688206,1.8346668,1.7165129,1.4244103,1.2307693,1.2077949,1.3751796,1.7066668,1.5392822,1.3161026,1.9003079,3.4034874,5.1659493,4.3585644,4.5095387,5.5532312,6.8988724,7.4141545,6.1046157,5.2742567,4.772103,4.709744,5.4547696,6.669129,7.13518,7.466667,8.021334,8.87795,11.441232,12.655591,13.771488,14.857847,14.8250265,13.971693,13.929027,13.673027,12.777026,11.428103,10.236719,9.764103,10.637129,12.11077,12.051693,10.794667,9.324308,8.772923,9.065026,8.920616,9.91836,10.555078,10.541949,9.609847,7.5388722,5.333334,3.4067695,2.3269746,2.162872,2.477949,2.8389745,3.2984617,3.8695388,4.781949,6.498462,7.204103,7.460103,6.9382567,6.0028725,5.737026,5.7042055,5.8420515,6.1013336,6.4032826,6.633026,6.554257,6.5969234,6.8627696,7.2172313,7.2960005,7.1614366,6.9054365,6.6494365,6.3967185,6.0258465,2.1234872,1.6869745,2.353231,2.5238976,1.9528207,1.7329233,1.8346668,1.529436,1.1027694,0.69251287,0.2855385,0.12471796,0.052512825,0.026256412,0.016410258,0.0,0.0,0.0,0.006564103,0.016410258,0.016410258,0.016410258,0.016410258,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.026256412,0.036102567,0.02297436,0.02297436,0.013128206,0.013128206,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.02297436,0.032820515,0.04266667,0.03938462,0.026256412,0.009846155,0.0,0.0,0.0,0.032820515,0.03938462,0.032820515,0.01969231,0.0,0.0,0.009846155,0.032820515,0.052512825,0.032820515,0.052512825,0.055794876,0.049230773,0.036102567,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.0,0.013128206,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.0032820515,0.0,0.0,0.0032820515,0.0,0.0,0.0,0.01969231,0.08861539,0.5152821,0.7417436,0.9156924,1.3029745,2.300718,4.0008206,4.6178465,3.6463592,1.8084104,1.083077,0.5349744,0.22646156,0.072205134,0.013128206,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016410258,0.036102567,0.032820515,0.013128206,0.016410258,0.0032820515,0.009846155,0.013128206,0.009846155,0.013128206,0.052512825,0.190359,0.39056414,0.5218462,0.3446154,0.28882053,0.18379489,0.07876924,0.016410258,0.026256412,0.08205129,0.101743594,0.14441027,0.16738462,0.049230773,0.009846155,0.01969231,0.04594872,0.068923086,0.059076928,0.03938462,0.01969231,0.006564103,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.029538464,0.029538464,0.01969231,0.013128206,0.009846155,0.0032820515,0.0,0.0,0.01969231,0.052512825,0.072205134,0.036102567,0.01969231,0.02297436,0.032820515,0.013128206,0.2231795,0.69579494,0.92225647,0.761436,0.4397949,0.32820517,0.4397949,0.67282057,0.8533334,0.7581539,0.508718,0.380718,0.32164106,0.36430773,0.6268718,0.69251287,0.56123084,0.48574364,0.44964105,0.15753847,0.23302566,0.318359,0.41025645,0.49887183,0.55794877,0.64000005,0.80738467,0.90256417,0.8598975,0.7122052,0.58420515,0.4201026,0.32820517,0.35774362,0.47917953,0.57764107,0.702359,0.80738467,0.9419488,1.2603078,1.1388719,1.2012309,1.2635899,1.211077,0.99774367,0.955077,0.8960001,0.92225647,1.0436924,1.1716924,1.0535386,0.8960001,0.8730257,1.0568206,1.4473847,1.8773335,1.6935385,1.6508719,1.9593848,2.2908719,1.9626669,1.7033848,1.6311796,1.8018463,2.1792822,1.6475899,1.7493335,1.8904617,1.9692309,2.3729234,2.409026,2.359795,2.1858463,1.8740515,1.4276924,1.3259488,1.4473847,1.3357949,0.93866676,0.6104616,0.4004103,0.26912823,0.21661541,0.18051283,0.049230773,0.24287182,0.14769232,0.029538464,0.0,0.0,0.009846155,0.032820515,0.04266667,0.036102567,0.029538464,0.049230773,0.055794876,0.03938462,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.0,0.013128206,0.02297436,0.02297436,0.013128206,0.0,0.0,0.009846155,0.029538464,0.055794876,0.06564103,0.029538464,0.009846155,0.009846155,0.009846155,0.0,0.0,0.0,0.0,0.006564103,0.016410258,0.032820515,0.118153855,0.20348719,0.23958977,0.21661541,0.14112821,0.128,0.13456412,0.118153855,0.02297436,0.0032820515,0.013128206,0.01969231,0.016410258,0.016410258,0.013128206,0.009846155,0.029538464,0.06564103,0.08861539,0.12143591,0.059076928,0.016410258,0.016410258,0.01969231,0.016410258,0.01969231,0.02297436,0.026256412,0.026256412,0.016410258,0.006564103,0.006564103,0.016410258,0.026256412,0.026256412,0.01969231,0.013128206,0.013128206,0.013128206,0.0032820515,0.0032820515,0.01969231,0.049230773,0.08205129,0.0951795,0.118153855,0.13784617,0.16082053,0.22646156,0.21333335,0.21661541,0.22646156,0.23302566,0.21989745,0.18707694,0.14769232,0.128,0.13128206,0.14112821,0.15097436,0.15097436,0.15753847,0.17066668,0.17066668,0.16738462,0.23958977,0.33476925,0.40369233,0.38728207,0.26912823,0.19364104,0.190359,0.28882053,0.5152821,0.761436,0.7515898,0.6859488,0.6695385,0.74830776,0.8566154,0.96492314,1.0272821,1.0075898,0.8763078,0.8598975,1.1881026,1.404718,1.3587693,1.1848207,1.0371283,0.9485129,0.84348726,0.67938465,0.44307697,0.39712822,0.39056414,0.4397949,0.49230772,0.4201026,0.37415388,0.42994875,0.5218462,0.55794877,0.43323082,0.37415388,0.4004103,0.43651286,0.47261542,0.56123084,0.69251287,0.73517954,0.6892308,0.6104616,0.58420515,0.574359,0.7384616,1.0075898,1.2865642,1.4703591,1.4506668,1.3784616,1.401436,1.6475899,2.1891284,2.03159,1.7394873,1.6508719,2.1792822,3.7940516,4.332308,5.3431797,7.0531287,8.730257,8.674462,6.308103,4.919795,4.33559,4.5390773,5.677949,6.8233852,6.948103,6.770872,7.069539,8.65477,11.053949,12.872206,14.155488,14.91036,15.100719,14.775796,14.989129,15.425642,15.855591,16.144411,13.39077,12.389745,12.832822,13.75836,13.53518,12.484924,11.227899,10.499283,10.811078,12.458668,13.643488,13.88636,12.402873,9.6754875,7.4765134,5.927385,4.2535386,2.8947694,2.2186668,2.5435898,2.917744,3.2787695,3.5840003,3.9384618,4.6112823,6.042257,7.568411,7.5913854,6.3310776,5.8420515,5.7698464,5.9503593,6.3343596,6.7774363,7.0367184,6.7314878,6.5837955,6.8594875,7.256616,6.8988724,6.5083084,6.3967185,6.3442054,6.1505647,5.6320004,1.404718,1.8051283,2.1530259,2.3302567,2.1234872,1.2209232,1.6246156,1.4309745,1.0338463,0.67610264,0.45620516,0.3249231,0.20676924,0.13456412,0.08533334,0.0,0.0,0.0,0.006564103,0.016410258,0.016410258,0.016410258,0.016410258,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.026256412,0.052512825,0.059076928,0.04594872,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.02297436,0.026256412,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.06235898,0.06564103,0.036102567,0.0,0.0,0.0,0.009846155,0.052512825,0.108307704,0.108307704,0.15425642,0.15097436,0.101743594,0.036102567,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.01969231,0.029538464,0.006564103,0.036102567,0.04266667,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.0032820515,0.0,0.006564103,0.052512825,0.19692309,0.77128214,1.079795,1.1848207,1.3850257,2.228513,4.4734364,6.445949,6.262154,4.194462,2.6715899,1.204513,0.45620516,0.15097436,0.06564103,0.029538464,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.036102567,0.118153855,0.101743594,0.0032820515,0.016410258,0.0032820515,0.01969231,0.036102567,0.049230773,0.06235898,0.20676924,0.6662565,0.86646163,0.6498462,0.25928208,0.07548718,0.013128206,0.0,0.016410258,0.07548718,0.29538465,0.23958977,0.18051283,0.17066668,0.06235898,0.013128206,0.09189744,0.20676924,0.25271797,0.108307704,0.15425642,0.0951795,0.032820515,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.04266667,0.09189744,0.07876924,0.03938462,0.009846155,0.0032820515,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.013128206,0.006564103,0.006564103,0.013128206,0.0,0.56123084,0.7187693,0.7318975,0.7089231,0.6104616,0.24287182,0.12471796,0.13784617,0.17066668,0.12143591,0.14769232,0.22646156,0.27569234,0.24615386,0.13784617,0.28225642,0.78769237,0.7515898,0.23302566,0.24287182,0.28225642,0.318359,0.4135385,0.6071795,0.8992821,1.1552821,1.1552821,0.8992821,0.60061544,0.6859488,0.636718,0.46933338,0.33476925,0.3446154,0.56451285,0.90584624,1.4966155,2.0217438,2.3466668,2.5173335,2.4451284,2.3072822,2.2088206,2.1333334,1.9364104,1.7657437,1.6705642,1.7591796,2.0512822,2.4418464,2.3433847,1.8970258,1.5491283,1.5688206,2.044718,2.5829747,3.1015387,3.3509746,3.1967182,2.609231,1.8904617,1.8838975,1.975795,2.0939488,2.7175386,1.9593848,2.2547693,2.425436,2.03159,1.3718976,1.8871796,2.793026,2.9013336,2.15959,1.6475899,1.5753847,1.1913847,0.702359,0.29210258,0.12143591,0.14769232,0.19692309,0.19692309,0.12143591,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.072205134,0.17723078,0.15097436,0.20020515,0.18707694,0.101743594,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.016410258,0.016410258,0.013128206,0.0,0.0,0.009846155,0.02297436,0.029538464,0.029538464,0.029538464,0.029538464,0.01969231,0.0,0.0,0.0,0.0,0.006564103,0.016410258,0.016410258,0.0032820515,0.009846155,0.03938462,0.0951795,0.16738462,0.08205129,0.052512825,0.03938462,0.02297436,0.0,0.0,0.0,0.006564103,0.016410258,0.016410258,0.0032820515,0.026256412,0.0951795,0.16082053,0.13784617,0.052512825,0.02297436,0.016410258,0.01969231,0.029538464,0.01969231,0.006564103,0.0,0.0032820515,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.006564103,0.0,0.0,0.0,0.0,0.009846155,0.068923086,0.15425642,0.16738462,0.13128206,0.15097436,0.17394873,0.17723078,0.15097436,0.14112821,0.09189744,0.072205134,0.12143591,0.24287182,0.28225642,0.24287182,0.190359,0.16410258,0.21333335,0.27569234,0.2986667,0.3052308,0.3052308,0.3052308,0.34133336,0.4135385,0.50543594,0.58420515,0.5940513,0.43651286,0.27897438,0.23958977,0.3314872,0.44307697,0.73517954,1.0568206,1.276718,1.394872,1.5425643,1.1618463,0.95835906,0.90256417,0.9747693,1.1454359,1.2668719,1.4080001,1.7165129,1.9035898,1.2209232,1.2209232,1.0732309,0.9156924,0.7975385,0.6859488,0.5513847,0.43651286,0.44307697,0.48246157,0.27569234,0.190359,0.21333335,0.2986667,0.38400003,0.39712822,0.39712822,0.56123084,0.7384616,0.83035904,0.79425645,0.67282057,0.5677949,0.54482055,0.5940513,0.65641034,0.508718,0.43651286,0.508718,0.7253334,1.0075898,1.2504616,1.404718,1.4834872,1.5425643,1.6640002,2.103795,2.7700515,2.6289232,1.9987694,2.546872,3.1474874,4.3027697,6.0717955,7.965539,8.940309,6.928411,4.46359,3.3247182,3.7251284,4.348718,4.5062566,4.31918,4.0992823,4.2601027,5.3103595,7.788308,9.186462,11.0605135,13.574565,15.504412,15.002257,14.263796,15.222155,17.450668,18.15631,16.449642,14.345847,13.400617,13.449847,12.619488,10.689642,10.620719,11.024411,12.875488,19.515078,17.135592,13.052719,8.969847,6.1472826,5.402257,5.9995904,5.8486156,4.338872,2.422154,2.5928206,2.8882053,3.1442053,3.3214362,3.43959,3.5872824,4.342154,6.0980515,7.0137444,6.7085133,6.2555904,5.9503593,5.98318,6.363898,6.9776416,7.5979495,7.634052,7.27959,6.705231,6.301539,6.669129,6.5706673,6.2884107,6.052103,5.865026,5.5236926,2.3696413,3.8564105,3.6036925,3.2820516,3.43959,3.501949,3.2032824,2.2121027,1.5458462,1.401436,1.142154,0.7515898,0.49230772,0.3511795,0.28225642,0.20676924,0.052512825,0.01969231,0.016410258,0.006564103,0.016410258,0.006564103,0.0032820515,0.0032820515,0.0,0.0,0.009846155,0.013128206,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.009846155,0.026256412,0.036102567,0.006564103,0.0,0.0,0.0,0.0,0.0,0.006564103,0.009846155,0.013128206,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.006564103,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.032820515,0.052512825,0.04266667,0.013128206,0.013128206,0.02297436,0.032820515,0.055794876,0.11158975,0.2297436,0.25928208,0.24615386,0.18379489,0.09189744,0.02297436,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.0,0.006564103,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.0032820515,0.0,0.0,0.0,0.0032820515,0.0,0.006564103,0.029538464,0.08861539,0.23630771,0.58420515,0.92553854,0.96492314,0.7778462,0.8008206,1.2964103,1.8510771,2.0151796,1.7033848,1.1946667,0.5874872,0.24287182,0.08205129,0.04594872,0.06564103,0.101743594,0.118153855,0.08205129,0.01969231,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.016410258,0.01969231,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.02297436,0.01969231,0.0,0.0032820515,0.009846155,0.03938462,0.13784617,0.29538465,0.4135385,0.190359,0.2100513,0.2231795,0.14112821,0.052512825,0.016410258,0.0032820515,0.0,0.006564103,0.026256412,0.16082053,0.26584616,0.23302566,0.0951795,0.02297436,0.12143591,0.19364104,0.16410258,0.059076928,0.02297436,0.029538464,0.01969231,0.006564103,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02297436,0.08861539,0.17394873,0.21333335,0.17066668,0.12471796,0.059076928,0.0,0.0032820515,0.0,0.0,0.0032820515,0.009846155,0.0,0.0032820515,0.0,0.0,0.0032820515,0.0,0.12143591,0.18707694,0.22646156,0.27241027,0.34133336,0.4135385,0.28225642,0.18707694,0.20348719,0.24287182,0.38728207,0.42994875,0.33476925,0.17394873,0.11158975,0.11158975,0.21333335,0.25928208,0.2231795,0.20676924,0.28225642,0.41025645,0.5415385,0.7318975,1.1323078,1.0962052,1.1257436,1.1520001,1.270154,1.7362052,2.1169233,2.048,2.0086155,2.300718,3.0654361,3.4756925,3.8695388,4.092718,4.073026,3.82359,3.5544617,3.2164104,2.8389745,2.5600002,2.609231,2.556718,2.4057438,2.3860514,2.5829747,2.9538465,3.2656412,3.1803079,2.9046156,2.878359,3.764513,4.263385,3.9876926,3.2722054,2.5731285,2.4746668,2.4582565,2.553436,2.7044106,2.7798977,2.5829747,1.8346668,1.6410258,1.529436,1.3226668,1.142154,1.0666667,1.2504616,1.214359,0.8992821,0.65969235,0.5973334,0.49887183,0.38728207,0.26256412,0.108307704,0.07548718,0.08205129,0.08205129,0.055794876,0.013128206,0.04266667,0.055794876,0.0951795,0.118153855,0.0,0.049230773,0.02297436,0.013128206,0.059076928,0.15097436,0.06564103,0.036102567,0.01969231,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.0032820515,0.0,0.0,0.0,0.0032820515,0.009846155,0.009846155,0.0032820515,0.013128206,0.02297436,0.01969231,0.016410258,0.01969231,0.01969231,0.01969231,0.026256412,0.02297436,0.009846155,0.0,0.0,0.0,0.006564103,0.016410258,0.026256412,0.026256412,0.026256412,0.06235898,0.14441027,0.26584616,0.27897438,0.20676924,0.12143591,0.055794876,0.013128206,0.013128206,0.013128206,0.01969231,0.026256412,0.016410258,0.013128206,0.026256412,0.032820515,0.036102567,0.03938462,0.013128206,0.0032820515,0.013128206,0.029538464,0.029538464,0.009846155,0.0,0.0032820515,0.009846155,0.0032820515,0.0032820515,0.0032820515,0.0032820515,0.0032820515,0.0032820515,0.0032820515,0.0,0.009846155,0.02297436,0.013128206,0.032820515,0.04594872,0.059076928,0.08861539,0.16738462,0.17066668,0.14769232,0.128,0.118153855,0.10502565,0.08205129,0.052512825,0.04266667,0.09189744,0.23302566,0.27897438,0.29538465,0.30851284,0.33805132,0.39712822,0.48574364,0.5481026,0.5874872,0.60389745,0.5874872,0.61374366,0.7056411,0.78769237,0.8205129,0.8041026,0.6629744,0.4660513,0.28882053,0.18051283,0.17394873,0.3511795,0.5316923,0.7253334,0.94523084,1.1979488,1.1520001,1.0765129,1.1126155,1.2406155,1.2537436,1.2012309,1.2077949,1.3161026,1.3489232,0.93866676,0.88287187,0.98461545,1.0601027,1.0338463,0.9419488,0.80738467,0.6498462,0.5513847,0.512,0.4201026,0.42338464,0.446359,0.43651286,0.36102566,0.23958977,0.20020515,0.30851284,0.52512825,0.7089231,0.6235898,0.39384618,0.26256412,0.26256412,0.34789747,0.4004103,0.36102566,0.32820517,0.34789747,0.4201026,0.4955898,0.8763078,1.1881026,1.339077,1.3489232,1.332513,1.4900514,1.7591796,2.9111798,4.388103,4.2830772,3.8629746,4.135385,5.037949,6.3343596,7.6242056,6.547693,5.85518,5.3103595,5.0642056,5.668103,5.4547696,4.565334,3.6726158,3.370667,4.1747694,5.7632823,6.941539,8.188719,9.833026,12.025436,12.967385,12.672001,12.225642,12.885334,16.082052,19.255796,20.352001,20.647387,20.46031,19.160616,17.056822,13.974976,11.812103,11.211488,11.595488,9.849437,8.129642,6.8365135,6.436103,7.4404106,8.408616,6.994052,5.540103,4.9132314,4.4996924,4.1452312,3.5380516,3.121231,3.1081028,3.501949,4.1025643,4.97559,6.294975,7.4404106,6.987488,6.547693,6.3540516,6.442667,6.774154,7.269744,7.5585647,7.5454364,7.1220517,6.491898,6.1538467,5.920821,5.7534366,5.5729237,5.3398976,5.0477953,2.609231,3.8465643,4.4340515,4.1911798,3.623385,3.9351797,3.2918978,2.609231,2.1891284,2.0118976,1.7427694,1.014154,0.827077,0.7318975,0.58092314,0.54482055,0.3052308,0.14441027,0.04594872,0.0,0.006564103,0.009846155,0.009846155,0.006564103,0.0,0.0,0.0032820515,0.013128206,0.013128206,0.016410258,0.04594872,0.009846155,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.026256412,0.01969231,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.009846155,0.013128206,0.013128206,0.006564103,0.0,0.009846155,0.036102567,0.052512825,0.049230773,0.032820515,0.02297436,0.026256412,0.032820515,0.06235898,0.15097436,0.88287187,0.53825647,0.15097436,0.07876924,0.02297436,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.0,0.0,0.0032820515,0.006564103,0.0,0.0,0.009846155,0.02297436,0.049230773,0.1148718,0.24943592,0.48246157,0.574359,0.46933338,0.3249231,0.3117949,0.38728207,0.54482055,0.7253334,0.8041026,0.61374366,0.43323082,0.34133336,0.3117949,0.2231795,0.15425642,0.14112821,0.118153855,0.06564103,0.026256412,0.01969231,0.006564103,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.01969231,0.052512825,0.072205134,0.108307704,0.17066668,0.23958977,0.08861539,0.04266667,0.02297436,0.0032820515,0.0,0.0,0.006564103,0.03938462,0.118153855,0.25271797,0.24615386,0.24287182,0.17066668,0.052512825,0.006564103,0.06564103,0.098461546,0.068923086,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.01969231,0.059076928,0.09189744,0.01969231,0.03938462,0.068923086,0.12471796,0.20348719,0.26256412,0.24287182,0.12471796,0.029538464,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.009846155,0.029538464,0.026256412,0.02297436,0.026256412,0.026256412,0.055794876,0.118153855,0.21333335,0.318359,0.4201026,0.29538465,0.18707694,0.29538465,0.5349744,0.5316923,0.38728207,0.27569234,0.20348719,0.16410258,0.15097436,0.16082053,0.39056414,0.6465641,0.8369231,0.95835906,1.2635899,1.5983591,1.913436,2.166154,2.353231,2.5862565,2.9013336,3.2328207,3.5511796,3.8564105,3.7448208,4.3060517,4.9329233,5.3070774,5.3760004,5.2315903,5.093744,4.844308,4.460308,4.0041027,3.3805132,2.7470772,2.3105643,2.2580514,2.7503593,2.7831798,2.5271797,2.3072822,2.412308,3.1015387,3.0752823,3.117949,3.0654361,3.1638978,4.0500517,4.598154,4.0500517,3.2886157,3.0326157,3.8432825,3.1573336,2.733949,2.4418464,2.1497438,1.7329233,1.3620514,1.3161026,1.0469744,0.5907693,0.5874872,0.47917953,0.56123084,0.61374366,0.5284103,0.32164106,0.29538465,0.25928208,0.23302566,0.20348719,0.108307704,0.07876924,0.04266667,0.02297436,0.029538464,0.068923086,0.032820515,0.029538464,0.0951795,0.17723078,0.108307704,0.098461546,0.04266667,0.009846155,0.01969231,0.06235898,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.013128206,0.016410258,0.009846155,0.006564103,0.0032820515,0.0,0.0032820515,0.009846155,0.0032820515,0.0032820515,0.0032820515,0.0032820515,0.016410258,0.01969231,0.02297436,0.016410258,0.006564103,0.016410258,0.036102567,0.06235898,0.068923086,0.049230773,0.009846155,0.016410258,0.013128206,0.026256412,0.055794876,0.07548718,0.06235898,0.04594872,0.055794876,0.09189744,0.15097436,0.21989745,0.2100513,0.19364104,0.19364104,0.190359,0.101743594,0.04594872,0.026256412,0.026256412,0.006564103,0.013128206,0.02297436,0.02297436,0.009846155,0.016410258,0.009846155,0.009846155,0.013128206,0.02297436,0.02297436,0.0032820515,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.02297436,0.032820515,0.036102567,0.03938462,0.055794876,0.08533334,0.13128206,0.1148718,0.07876924,0.06235898,0.06564103,0.04594872,0.049230773,0.049230773,0.052512825,0.09189744,0.23958977,0.3511795,0.35446155,0.36758977,0.44307697,0.56123084,0.702359,0.82379496,0.892718,0.9156924,0.92225647,0.92553854,0.9714873,1.0108719,1.0043077,0.9353847,0.78769237,0.60389745,0.41025645,0.2297436,0.108307704,0.15097436,0.2100513,0.318359,0.48574364,0.702359,0.86974365,1.0108719,1.204513,1.3850257,1.3456411,1.2471796,1.1126155,1.0601027,1.0535386,0.9156924,0.9517949,1.0469744,1.1126155,1.0962052,0.9517949,1.0075898,1.0272821,0.9747693,0.81394875,0.512,0.43323082,0.48246157,0.51856416,0.48246157,0.380718,0.29538465,0.29210258,0.34789747,0.40369233,0.3511795,0.21333335,0.15425642,0.18051283,0.25271797,0.27241027,0.26584616,0.26912823,0.29210258,0.33476925,0.37415388,0.5415385,0.78769237,0.97805136,1.0633847,1.0601027,1.1158975,1.204513,1.9462565,3.0687182,3.4231799,3.564308,3.8334363,4.0369234,4.4340515,5.72718,5.297231,5.832206,5.61559,4.6080003,4.460308,5.221744,5.041231,4.352,3.751385,3.9909747,5.543385,6.1046157,6.685539,7.716103,9.02236,10.210463,10.791386,11.050668,11.625027,13.505642,16.676104,19.072002,19.951591,18.87836,15.727591,12.727796,10.246565,8.582564,8.070564,9.081436,9.281642,10.161232,10.312206,9.485129,8.582564,8.677744,7.325539,6.3967185,6.265436,5.805949,5.8814363,5.4547696,4.571898,3.6594875,3.5347695,4.0303593,4.529231,5.540103,6.7840004,7.181129,6.99077,6.918565,6.872616,6.8562055,6.9776416,7.351795,7.680001,7.5913854,7.076103,6.4754877,6.1046157,5.9602056,5.7435904,5.4153852,5.1856413,2.5009232,3.6135387,4.5522056,4.3027697,3.367385,3.7776413,3.367385,2.7864618,2.3138463,1.9922053,1.6213335,1.0305642,1.0633847,1.1060513,0.9517949,0.8008206,0.42994875,0.21661541,0.0951795,0.026256412,0.006564103,0.01969231,0.026256412,0.016410258,0.0,0.006564103,0.006564103,0.013128206,0.016410258,0.02297436,0.052512825,0.016410258,0.006564103,0.006564103,0.006564103,0.006564103,0.006564103,0.006564103,0.0032820515,0.0,0.0,0.0032820515,0.006564103,0.009846155,0.013128206,0.016410258,0.052512825,0.068923086,0.059076928,0.029538464,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0,0.006564103,0.01969231,0.01969231,0.013128206,0.006564103,0.0,0.01969231,0.04594872,0.06564103,0.06564103,0.049230773,0.029538464,0.016410258,0.026256412,0.101743594,0.90256417,0.6071795,0.2297436,0.13128206,0.032820515,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.006564103,0.013128206,0.006564103,0.0,0.006564103,0.013128206,0.01969231,0.036102567,0.06564103,0.20676924,0.3446154,0.41025645,0.36758977,0.37743592,0.3314872,0.33476925,0.4594872,0.7515898,0.88615394,0.88287187,0.7581539,0.5415385,0.27241027,0.13128206,0.0951795,0.08205129,0.055794876,0.026256412,0.01969231,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.006564103,0.0032820515,0.01969231,0.052512825,0.06235898,0.049230773,0.029538464,0.04266667,0.016410258,0.029538464,0.07548718,0.1148718,0.08533334,0.036102567,0.016410258,0.03938462,0.1148718,0.24615386,0.19692309,0.13456412,0.072205134,0.026256412,0.02297436,0.036102567,0.02297436,0.009846155,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.01969231,0.06564103,0.1148718,0.09189744,0.098461546,0.098461546,0.11158975,0.14769232,0.17066668,0.16738462,0.06564103,0.0,0.0,0.0,0.0032820515,0.009846155,0.009846155,0.013128206,0.032820515,0.04594872,0.032820515,0.032820515,0.049230773,0.059076928,0.108307704,0.2297436,0.38728207,0.48574364,0.35446155,0.128,0.072205134,0.24287182,0.4955898,0.47589746,0.24943592,0.1148718,0.118153855,0.21661541,0.26256412,0.23958977,0.50543594,0.8205129,1.0994873,1.3915899,2.2580514,2.9078977,3.3608208,3.629949,3.7021542,4.066462,4.4832826,4.965744,5.5105643,6.0783596,6.048821,6.626462,7.1154876,7.138462,6.6461544,6.091488,5.677949,5.3825645,5.028103,4.273231,3.4133337,2.8750772,2.6978464,2.8389745,3.1770258,2.8553848,2.5304618,2.2350771,2.228513,3.0162053,2.678154,2.674872,2.8258464,3.2065644,4.1485133,5.211898,4.7950773,4.0992823,3.895795,4.5390773,3.4921029,2.6453335,1.9396925,1.3357949,0.8041026,0.7515898,0.8566154,0.69579494,0.35446155,0.42338464,0.30851284,0.318359,0.35774362,0.3446154,0.2100513,0.190359,0.17066668,0.17723078,0.19692309,0.18051283,0.14769232,0.08861539,0.032820515,0.013128206,0.06564103,0.026256412,0.013128206,0.06564103,0.13784617,0.108307704,0.072205134,0.029538464,0.009846155,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.016410258,0.02297436,0.009846155,0.006564103,0.0032820515,0.0,0.0032820515,0.009846155,0.0032820515,0.0,0.0,0.0032820515,0.016410258,0.016410258,0.01969231,0.016410258,0.006564103,0.016410258,0.04594872,0.08533334,0.09189744,0.06564103,0.026256412,0.03938462,0.036102567,0.04594872,0.068923086,0.08205129,0.06235898,0.04266667,0.029538464,0.032820515,0.049230773,0.118153855,0.17066668,0.19692309,0.2100513,0.24943592,0.13784617,0.055794876,0.01969231,0.016410258,0.006564103,0.01969231,0.02297436,0.01969231,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.01969231,0.016410258,0.0032820515,0.0,0.0,0.0,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.026256412,0.026256412,0.032820515,0.04266667,0.059076928,0.068923086,0.049230773,0.02297436,0.016410258,0.026256412,0.016410258,0.029538464,0.049230773,0.08205129,0.13128206,0.19692309,0.32820517,0.37743592,0.44964105,0.5874872,0.7450257,0.9288206,1.0929232,1.204513,1.2635899,1.2865642,1.2471796,1.2406155,1.2274873,1.1618463,0.97805136,0.7975385,0.6268718,0.45620516,0.29210258,0.15097436,0.13128206,0.11158975,0.13456412,0.21989745,0.36102566,0.5284103,0.7318975,0.9747693,1.1881026,1.211077,1.1290257,0.9124103,0.79425645,0.8041026,0.8041026,0.9189744,1.0108719,1.0568206,1.020718,0.8598975,1.0108719,1.1881026,1.214359,1.0075898,0.5973334,0.44307697,0.46276927,0.51856416,0.5284103,0.49230772,0.446359,0.4266667,0.39712822,0.34133336,0.27241027,0.20676924,0.18051283,0.2100513,0.26256412,0.24615386,0.23302566,0.24615386,0.27897438,0.318359,0.36430773,0.36758977,0.48574364,0.6301539,0.7515898,0.8336411,0.90912825,1.0305642,1.2931283,1.7263591,2.300718,3.6135387,4.9362054,5.3037953,5.037949,5.72718,6.2129235,6.764308,6.1078978,4.46359,3.5183592,4.076308,4.7622566,5.0674877,4.854154,4.345436,5.2381544,5.5204105,6.0324106,6.8496413,7.282872,7.9327188,9.005949,10.331899,11.54954,12.100924,13.197129,15.442053,17.348925,17.371899,13.883078,10.259693,8.769642,8.346257,8.608821,9.856001,10.86359,11.989334,11.943385,10.433641,8.178872,7.9917955,7.463385,7.4141545,7.8080006,7.748924,8.119796,7.778462,6.4722056,4.7458467,3.9548721,4.240411,4.604718,5.218462,6.0619493,6.925129,7.197539,7.3452315,7.250052,6.9809237,6.8004107,7.204103,7.702975,7.824411,7.463385,6.8430777,6.4754877,6.3442054,6.124308,5.7632823,5.4908724,2.1103592,3.5380516,4.1091285,3.7776413,3.1671798,3.5774362,3.6562054,2.8553848,2.100513,1.6410258,1.0699488,1.2898463,1.5097437,1.522872,1.273436,0.86974365,0.446359,0.26256412,0.15425642,0.06564103,0.016410258,0.03938462,0.052512825,0.036102567,0.006564103,0.013128206,0.013128206,0.013128206,0.016410258,0.016410258,0.01969231,0.01969231,0.01969231,0.016410258,0.013128206,0.013128206,0.013128206,0.013128206,0.009846155,0.0032820515,0.0032820515,0.009846155,0.013128206,0.016410258,0.02297436,0.01969231,0.07548718,0.13128206,0.13456412,0.08205129,0.026256412,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.013128206,0.0,0.0,0.006564103,0.013128206,0.013128206,0.02297436,0.009846155,0.013128206,0.026256412,0.049230773,0.08861539,0.10502565,0.08861539,0.049230773,0.032820515,0.1148718,0.28225642,0.38400003,0.35774362,0.2231795,0.07876924,0.04594872,0.01969231,0.006564103,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.0032820515,0.0032820515,0.013128206,0.01969231,0.0032820515,0.0,0.009846155,0.068923086,0.24287182,0.48246157,0.6892308,0.8008206,0.83035904,0.8566154,1.0765129,0.92225647,0.67610264,0.5677949,0.761436,1.1126155,1.2274873,1.0108719,0.5677949,0.19692309,0.0951795,0.08533334,0.101743594,0.12471796,0.17723078,0.21661541,0.16082053,0.08533334,0.032820515,0.016410258,0.01969231,0.016410258,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.01969231,0.013128206,0.0,0.0,0.009846155,0.013128206,0.006564103,0.0032820515,0.02297436,0.072205134,0.24943592,0.35446155,0.30851284,0.17066668,0.072205134,0.01969231,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.049230773,0.059076928,0.02297436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.055794876,0.15097436,0.118153855,0.08205129,0.06235898,0.052512825,0.013128206,0.0032820515,0.0,0.0,0.0,0.0032820515,0.013128206,0.026256412,0.029538464,0.036102567,0.09189744,0.08533334,0.08205129,0.07876924,0.07876924,0.072205134,0.128,0.27569234,0.4594872,0.50543594,0.12471796,0.055794876,0.06564103,0.1148718,0.16082053,0.16082053,0.15097436,0.12143591,0.15425642,0.24943592,0.3446154,0.29210258,0.42994875,0.7089231,1.0272821,1.2307693,2.5107694,3.4330258,4.0500517,4.4110775,4.5456414,4.519385,4.588308,4.923077,5.664821,6.9120007,7.77518,7.824411,7.5520005,7.2369237,6.957949,6.2851286,6.2227697,6.432821,6.3606157,5.211898,4.266667,3.9942567,4.027077,4.023795,3.6562054,2.917744,2.6420515,2.5665643,2.678154,3.2164104,2.8258464,2.665026,2.8553848,3.43959,4.3749747,6.1013336,6.2687182,5.5696416,4.601436,3.8662567,3.2361028,2.3991797,1.6082052,0.9419488,0.3117949,0.3052308,0.34133336,0.4135385,0.508718,0.5973334,0.4397949,0.30194873,0.19692309,0.13128206,0.13128206,0.08861539,0.101743594,0.14769232,0.20348719,0.24287182,0.19692309,0.16082053,0.09189744,0.016410258,0.02297436,0.052512825,0.03938462,0.036102567,0.03938462,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.013128206,0.0,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.006564103,0.01969231,0.013128206,0.013128206,0.013128206,0.013128206,0.016410258,0.036102567,0.068923086,0.068923086,0.03938462,0.04594872,0.06235898,0.07548718,0.07548718,0.06564103,0.06235898,0.059076928,0.04594872,0.02297436,0.009846155,0.032820515,0.07876924,0.14112821,0.14441027,0.11158975,0.15097436,0.108307704,0.052512825,0.02297436,0.01969231,0.01969231,0.026256412,0.01969231,0.013128206,0.013128206,0.01969231,0.016410258,0.016410258,0.01969231,0.02297436,0.013128206,0.0032820515,0.0,0.0,0.0032820515,0.013128206,0.0032820515,0.0,0.0,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.026256412,0.02297436,0.0032820515,0.013128206,0.013128206,0.0032820515,0.0,0.006564103,0.016410258,0.016410258,0.052512825,0.12471796,0.190359,0.14112821,0.23302566,0.40697438,0.636718,0.8730257,1.0568206,1.2307693,1.3850257,1.5261539,1.6344616,1.6607181,1.5753847,1.522872,1.4572309,1.3128207,1.0108719,0.75487185,0.57764107,0.43651286,0.318359,0.2297436,0.21661541,0.17723078,0.15753847,0.17723078,0.25271797,0.29538465,0.4397949,0.6235898,0.8008206,0.9353847,0.8960001,0.67610264,0.5513847,0.5677949,0.55794877,0.6629744,0.8008206,0.86317956,0.8205129,0.7253334,0.8467693,1.0962052,1.1585642,0.95835906,0.65969235,0.508718,0.46933338,0.47261542,0.47589746,0.4594872,0.48574364,0.571077,0.61374366,0.5677949,0.44307697,0.36430773,0.30194873,0.28882053,0.30851284,0.27897438,0.27897438,0.29210258,0.3052308,0.31507695,0.33476925,0.3446154,0.36758977,0.40369233,0.47261542,0.6235898,0.7581539,0.9878975,1.3357949,1.7657437,2.169436,3.757949,6.0258465,7.315693,7.2927184,6.9021544,8.536616,8.681026,7.387898,5.3037953,3.6758976,3.1573336,3.9220517,5.0642056,5.664821,4.7917953,4.5390773,4.955898,5.8092313,6.6395903,6.75118,6.564103,7.394462,9.035488,10.781539,11.411694,10.8767185,12.396309,15.8654375,18.963694,17.152,13.033027,11.703795,12.120616,12.826258,11.96636,11.723488,10.975181,9.813334,8.425026,7.1023593,7.7325134,8.001641,8.480822,9.258667,9.947898,10.203898,9.465437,7.781744,5.7698464,4.6145644,4.667077,4.962462,5.349744,5.799385,6.416411,7.0826674,7.4075904,7.3386674,6.99077,6.665847,7.0104623,7.5191803,7.7981544,7.650462,7.0826674,6.738052,6.518154,6.2752824,5.9569235,5.61559,1.204513,2.537026,3.508513,3.7054362,3.3214362,3.1737437,3.1245131,2.865231,2.5304618,2.0841026,1.3259488,2.8160002,2.9505644,2.2547693,1.3095386,0.74830776,0.73517954,0.47589746,0.21333335,0.06564103,0.016410258,0.08861539,0.108307704,0.07548718,0.02297436,0.0,0.0,0.009846155,0.016410258,0.01969231,0.029538464,0.04266667,0.036102567,0.01969231,0.0,0.0,0.013128206,0.006564103,0.006564103,0.016410258,0.016410258,0.0032820515,0.0,0.0,0.006564103,0.029538464,0.01969231,0.052512825,0.08861539,0.101743594,0.07548718,0.06564103,0.02297436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01969231,0.02297436,0.013128206,0.0,0.0,0.0,0.0,0.009846155,0.04594872,0.032820515,0.02297436,0.016410258,0.026256412,0.07548718,0.16082053,0.21989745,0.17066668,0.055794876,0.029538464,0.07876924,0.13784617,0.18051283,0.190359,0.15097436,0.128,0.07548718,0.026256412,0.0,0.0,0.0,0.009846155,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.029538464,0.006564103,0.0,0.02297436,0.256,1.0371283,2.0873847,2.678154,2.6551797,2.2482052,2.0906668,2.7011285,2.349949,1.6836925,1.1618463,1.0535386,1.1027694,0.88615394,0.6104616,0.380718,0.19692309,0.2231795,0.30194873,0.42994875,0.6170257,0.88615394,1.079795,0.8008206,0.4201026,0.16082053,0.07548718,0.101743594,0.08861539,0.052512825,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.06235898,0.35446155,0.9944616,1.024,0.40369233,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.026256412,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.016410258,0.032820515,0.04594872,0.07876924,0.21333335,0.27569234,0.318359,0.2855385,0.18379489,0.06235898,0.036102567,0.08533334,0.15097436,0.19692309,0.19692309,0.13784617,0.18707694,0.28882053,0.35774362,0.25928208,0.3446154,0.32164106,0.2100513,0.11158975,0.19692309,0.3708718,0.7318975,1.276718,1.6213335,1.020718,1.4605129,2.349949,3.4658465,4.384821,4.4701543,3.4691284,2.6715899,2.4451284,2.993231,4.348718,5.874872,6.12759,6.2490263,6.7150774,7.325539,6.3474874,7.4043083,8.342975,8.116513,6.774154,5.664821,4.9099493,4.2929235,3.6562054,2.8980515,2.861949,2.806154,3.3805132,4.352,4.6080003,4.1189747,3.751385,3.7021542,3.9253337,4.1189747,5.609026,7.0531287,6.7610264,4.71959,2.609231,2.4385643,2.0020514,1.5130258,1.0666667,0.64000005,0.4201026,0.35774362,0.35774362,0.35446155,0.3052308,0.4397949,0.49887183,0.37743592,0.15425642,0.108307704,0.0951795,0.09189744,0.07876924,0.06235898,0.06235898,0.06235898,0.12471796,0.13128206,0.08205129,0.108307704,0.118153855,0.059076928,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.016410258,0.016410258,0.016410258,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.016410258,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.016410258,0.01969231,0.029538464,0.006564103,0.0,0.0,0.0032820515,0.016410258,0.016410258,0.016410258,0.009846155,0.009846155,0.04594872,0.08205129,0.13784617,0.16082053,0.14769232,0.12143591,0.15753847,0.14112821,0.07876924,0.02297436,0.04594872,0.068923086,0.11158975,0.14441027,0.13784617,0.07548718,0.11158975,0.11158975,0.108307704,0.09189744,0.029538464,0.01969231,0.016410258,0.009846155,0.006564103,0.029538464,0.01969231,0.016410258,0.016410258,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.016410258,0.016410258,0.026256412,0.08533334,0.15753847,0.21333335,0.21333335,0.2855385,0.5874872,0.99774367,1.3981539,1.6771283,1.7263591,1.7755898,1.8740515,1.9889232,2.0151796,1.9298463,1.8346668,1.7001027,1.4998976,1.204513,0.81394875,0.6170257,0.4955898,0.38728207,0.28882053,0.27897438,0.28225642,0.27241027,0.23958977,0.2297436,0.28882053,0.58092314,0.7450257,0.7515898,0.88615394,0.9353847,0.7450257,0.5546667,0.4594872,0.4135385,0.44964105,0.4955898,0.512,0.50543594,0.51856416,0.7253334,1.079795,1.0994873,0.7811283,0.6104616,0.53825647,0.51856416,0.512,0.48574364,0.4135385,0.33805132,0.5021539,0.69251287,0.77128214,0.6859488,0.5874872,0.49230772,0.38728207,0.30194873,0.28882053,0.43651286,0.47261542,0.44307697,0.38400003,0.33476925,0.3249231,0.32164106,0.30851284,0.3052308,0.36758977,0.5021539,0.63343596,1.2635899,2.3269746,3.2196925,2.1333334,2.7044106,4.772103,6.695385,5.3398976,7.6964107,9.275078,8.766359,6.373744,3.7842054,4.466872,3.8695388,3.895795,4.7294364,4.850872,4.71959,5.097026,5.7009234,6.262154,6.5312824,5.737026,5.7140517,6.4590774,7.686565,8.835282,9.334154,10.880001,15.507693,21.02154,20.995283,15.258258,14.043899,14.916924,15.530668,13.627078,10.709334,8.989539,7.5191803,6.5903597,7.7357955,9.468719,9.517949,8.891078,8.753231,10.436924,10.791386,9.53436,7.6307697,5.8847184,4.9427695,5.0543594,5.290667,5.5171285,5.7074876,5.9503593,6.547693,6.9809237,7.072821,6.810257,6.3474874,6.3606157,6.948103,7.762052,8.241231,7.643898,6.9349747,6.2916927,5.786257,5.4580517,5.3103595,2.2908719,2.8816411,3.9745643,5.4449234,6.4557953,5.481026,4.6211286,4.1813335,3.9384618,3.6726158,3.170462,2.9997952,2.6617439,2.156308,1.6147693,1.2964103,1.1979488,1.0043077,0.764718,0.512,0.24615386,0.15425642,0.101743594,0.1148718,0.14769232,0.08533334,0.026256412,0.02297436,0.032820515,0.032820515,0.006564103,0.009846155,0.013128206,0.016410258,0.013128206,0.013128206,0.0032820515,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.006564103,0.0032820515,0.009846155,0.016410258,0.026256412,0.03938462,0.06564103,0.06564103,0.04594872,0.02297436,0.013128206,0.0032820515,0.0,0.0032820515,0.009846155,0.0,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.013128206,0.0032820515,0.0,0.009846155,0.013128206,0.013128206,0.016410258,0.032820515,0.068923086,0.06235898,0.036102567,0.016410258,0.016410258,0.06235898,0.101743594,0.108307704,0.07548718,0.029538464,0.049230773,0.072205134,0.07876924,0.07876924,0.09189744,0.08533334,0.055794876,0.029538464,0.02297436,0.02297436,0.013128206,0.013128206,0.013128206,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.036102567,0.026256412,0.032820515,0.06235898,0.14769232,0.34789747,0.73517954,0.9682052,0.97805136,1.0929232,2.0512822,2.7700515,2.7503593,2.1792822,1.4506668,1.1749744,1.2471796,1.1454359,1.0305642,1.0535386,1.332513,1.4506668,1.0896411,0.5677949,0.256,0.5874872,1.8346668,2.5993848,2.6584618,2.2711797,2.1792822,3.8990772,5.139693,4.4438977,2.3368206,1.332513,0.9189744,0.6432821,0.4201026,0.20676924,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.013128206,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.08205129,0.20348719,0.20348719,0.08205129,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.013128206,0.016410258,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.016410258,0.016410258,0.032820515,0.07548718,0.13128206,0.17723078,0.190359,0.19692309,0.21661541,0.24943592,0.29210258,0.23958977,0.23630771,0.23630771,0.26256412,0.41682056,0.48246157,0.45620516,0.34789747,0.2297436,0.2100513,0.27569234,0.27569234,0.2100513,0.12143591,0.101743594,0.2231795,0.5284103,1.0732309,1.4080001,0.5940513,1.7165129,2.9013336,4.06318,5.1265645,6.0324106,6.117744,5.280821,4.2962055,3.8859491,4.70318,5.2020516,5.3891287,5.9470773,7.020308,8.214975,7.755488,7.3386674,7.7357955,8.4512825,7.716103,5.1987696,3.4034874,2.3236926,1.9659488,2.3630772,2.1497438,2.0578463,2.681436,3.9680004,5.2315903,4.8016415,4.2338467,3.9351797,3.9614363,4.010667,4.824616,5.602462,5.602462,4.5489235,2.6322052,2.0611284,1.6147693,1.2340513,0.92553854,0.761436,0.67938465,0.571077,0.48574364,0.39712822,0.17066668,0.3052308,0.43323082,0.50543594,0.49887183,0.4004103,0.13456412,0.0951795,0.1148718,0.101743594,0.072205134,0.072205134,0.09189744,0.08533334,0.049230773,0.04594872,0.029538464,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0032820515,0.006564103,0.0,0.006564103,0.013128206,0.036102567,0.12471796,0.16410258,0.19692309,0.20020515,0.19364104,0.2297436,0.3249231,0.32164106,0.29538465,0.27241027,0.20676924,0.20348719,0.17066668,0.128,0.10502565,0.118153855,0.0951795,0.14112821,0.17066668,0.15753847,0.12471796,0.12143591,0.11158975,0.101743594,0.0951795,0.09189744,0.07876924,0.06235898,0.03938462,0.01969231,0.006564103,0.0032820515,0.0032820515,0.006564103,0.016410258,0.02297436,0.02297436,0.016410258,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.02297436,0.009846155,0.0,0.006564103,0.026256412,0.029538464,0.055794876,0.09189744,0.128,0.17723078,0.27897438,0.44964105,0.8041026,1.332513,1.8871796,2.1202054,2.1858463,2.162872,2.0906668,1.9790771,1.8838975,1.7788719,1.6377437,1.4605129,1.2668719,1.0601027,0.88615394,0.7515898,0.7187693,0.9124103,0.7450257,0.65969235,0.5874872,0.49230772,0.36430773,0.36430773,0.44964105,0.571077,0.7122052,0.88615394,1.079795,1.083077,0.9156924,0.6662565,0.4594872,0.54482055,0.54482055,0.49887183,0.4660513,0.50543594,0.7056411,0.9616411,1.0436924,0.9124103,0.7318975,0.571077,0.47261542,0.43323082,0.42338464,0.4004103,0.35446155,0.3511795,0.4135385,0.5316923,0.6498462,0.7384616,0.7220513,0.62030774,0.46933338,0.33805132,0.35774362,0.3117949,0.27241027,0.27241027,0.3117949,0.318359,0.33476925,0.36102566,0.4004103,0.45292312,0.41025645,0.4135385,0.56123084,1.0010257,1.9003079,2.1333334,2.0020514,3.058872,4.768821,4.4996924,6.931693,7.817847,6.9120007,5.0051284,3.9318976,3.6758976,2.865231,2.5698464,2.9636924,3.3378465,3.5938463,4.1222568,4.6867695,5.1659493,5.543385,4.699898,4.6112823,5.3136415,6.419693,7.138462,7.50277,10.266257,15.123693,20.81149,25.08472,20.86072,18.084105,16.823795,16.393847,15.346873,12.596514,10.194052,8.316719,7.000616,6.1374364,6.560821,6.245744,6.121026,7.0957956,10.059488,11.497026,10.299078,7.906462,5.533539,4.161641,4.4077954,4.7622566,5.159385,5.5269747,5.792821,6.12759,6.692103,7.02359,6.951385,6.6034875,6.196513,6.298257,6.672411,7.003898,6.925129,6.498462,5.9930263,5.540103,5.2447186,5.175795,2.7109745,3.0162053,4.33559,6.1341543,7.276308,6.012718,4.598154,4.2338467,4.0500517,3.7120004,3.4133337,3.4494362,3.3050258,2.9571285,2.5206156,2.2580514,2.2022567,1.595077,1.079795,0.84348726,0.6432821,0.4594872,0.26584616,0.15097436,0.11158975,0.052512825,0.016410258,0.016410258,0.01969231,0.013128206,0.0,0.0,0.0032820515,0.006564103,0.006564103,0.016410258,0.0032820515,0.0,0.0032820515,0.009846155,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.006564103,0.0032820515,0.0,0.0032820515,0.013128206,0.049230773,0.06235898,0.059076928,0.04266667,0.02297436,0.013128206,0.009846155,0.013128206,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0,0.013128206,0.016410258,0.013128206,0.009846155,0.02297436,0.055794876,0.07876924,0.059076928,0.013128206,0.009846155,0.02297436,0.03938462,0.049230773,0.052512825,0.03938462,0.04594872,0.049230773,0.04266667,0.029538464,0.03938462,0.068923086,0.08205129,0.072205134,0.049230773,0.049230773,0.02297436,0.026256412,0.032820515,0.026256412,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.026256412,0.036102567,0.013128206,0.0,0.0,0.009846155,0.07548718,0.29210258,0.8041026,0.48574364,0.24943592,0.15097436,0.2100513,0.41025645,0.83035904,1.3029745,1.3817437,1.1881026,1.3981539,1.657436,1.5425643,1.1520001,0.7056411,0.52512825,0.43323082,0.36758977,0.36102566,0.47261542,0.8008206,0.9189744,0.72861546,0.52512825,0.67938465,1.6213335,2.8849232,2.6945643,1.9265642,1.2668719,1.2406155,2.166154,2.740513,2.3236926,1.2340513,0.7417436,0.51856416,0.38728207,0.27897438,0.15425642,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.026256412,0.049230773,0.052512825,0.01969231,0.0032820515,0.006564103,0.009846155,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0,0.013128206,0.06564103,0.12143591,0.12143591,0.06564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.006564103,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.01969231,0.052512825,0.12471796,0.32164106,0.2297436,0.14112821,0.14769232,0.15753847,0.15753847,0.16410258,0.19692309,0.25928208,0.31507695,0.2100513,0.24943592,0.3249231,0.39384618,0.46276927,0.44307697,0.36758977,0.23958977,0.13128206,0.15097436,0.20676924,0.23302566,0.24943592,0.2855385,0.36102566,0.39712822,0.6432821,0.9189744,1.0502565,0.8730257,1.5721027,2.3433847,3.4264617,4.916513,6.7544622,7.5618467,7.4765134,7.4896417,7.8802056,8.234667,7.5979495,7.8408213,9.344001,11.1294365,10.84718,8.612103,6.803693,6.1013336,6.229334,5.973334,4.4734364,2.6847181,1.8445129,2.100513,2.5206156,2.169436,1.782154,1.8806155,2.6322052,3.8400004,4.31918,4.0467696,3.820308,3.9122055,4.066462,4.529231,4.9460516,4.7228723,3.764513,2.4746668,1.8248206,1.6804104,1.7362052,1.723077,1.3981539,0.9517949,0.6235898,0.41682056,0.2855385,0.118153855,0.17394873,0.24615386,0.2986667,0.30194873,0.23630771,0.11158975,0.06235898,0.049230773,0.04594872,0.029538464,0.059076928,0.072205134,0.052512825,0.02297436,0.03938462,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.01969231,0.029538464,0.052512825,0.12471796,0.15097436,0.15753847,0.17066668,0.20348719,0.24615386,0.3117949,0.37743592,0.41682056,0.4201026,0.38400003,0.26912823,0.24943592,0.256,0.24615386,0.20020515,0.18707694,0.25928208,0.27241027,0.20676924,0.18379489,0.13456412,0.11158975,0.098461546,0.08205129,0.08861539,0.10502565,0.098461546,0.06564103,0.02297436,0.0,0.013128206,0.02297436,0.029538464,0.029538464,0.013128206,0.01969231,0.016410258,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.016410258,0.01969231,0.013128206,0.006564103,0.006564103,0.029538464,0.052512825,0.07548718,0.11158975,0.17066668,0.26912823,0.2986667,0.3708718,0.6235898,1.083077,1.654154,2.0020514,2.231795,2.3040001,2.2219489,2.03159,1.8904617,1.8379488,1.7624617,1.6147693,1.4375386,1.2570257,1.0896411,0.95835906,0.9156924,1.0305642,0.9616411,0.81394875,0.67282057,0.56123084,0.42338464,0.4135385,0.446359,0.54482055,0.7056411,0.90256417,1.2242053,1.2438976,1.086359,0.86974365,0.7187693,0.76800007,0.6301539,0.50543594,0.5021539,0.6695385,0.88615394,0.9485129,0.8795898,0.7384616,0.5973334,0.5481026,0.54482055,0.5677949,0.58420515,0.5349744,0.42338464,0.33805132,0.31507695,0.3511795,0.4201026,0.52512825,0.5907693,0.57764107,0.48902568,0.3511795,0.3249231,0.24287182,0.17723078,0.16410258,0.19692309,0.25271797,0.32820517,0.42338464,0.50543594,0.51856416,0.4397949,0.39056414,0.36430773,0.4660513,0.892718,1.3095386,1.3259488,1.6935385,2.3729234,2.546872,4.1156926,4.4767184,4.345436,4.2469745,4.516103,4.1156926,3.3772311,2.8160002,2.6880002,2.9965131,3.6791797,4.6802053,5.2447186,5.024821,4.0500517,3.6791797,4.013949,4.7917953,5.4941545,5.35959,5.2414365,7.2205133,11.59877,18.113642,25.951181,23.798155,19.35754,16.49559,16.8599,19.859694,18.021746,14.381949,10.768411,8.323282,7.50277,7.975385,6.705231,5.8945646,6.6560006,9.028924,13.676309,12.58995,8.815591,5.175795,4.269949,4.571898,4.9362054,5.3169236,5.6254363,5.723898,5.979898,6.6002054,7.128616,7.2664623,6.9054365,6.226052,5.9995904,6.0619493,6.226052,6.294975,6.189949,6.0258465,5.8125134,5.5532312,5.2611284,2.3729234,2.8389745,4.0402055,5.346462,5.98318,5.034667,3.9187696,3.698872,3.515077,3.0982566,2.789744,3.757949,3.9811285,3.8071797,3.5511796,3.4921029,3.4297438,2.5009232,1.6508719,1.214359,0.9124103,0.6826667,0.48574364,0.30851284,0.15425642,0.052512825,0.029538464,0.029538464,0.026256412,0.013128206,0.013128206,0.016410258,0.01969231,0.013128206,0.006564103,0.016410258,0.0032820515,0.0,0.006564103,0.013128206,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.006564103,0.0032820515,0.0,0.0,0.0,0.02297436,0.032820515,0.04266667,0.04594872,0.036102567,0.029538464,0.026256412,0.026256412,0.01969231,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.009846155,0.006564103,0.006564103,0.016410258,0.03938462,0.068923086,0.059076928,0.01969231,0.016410258,0.016410258,0.016410258,0.02297436,0.032820515,0.03938462,0.03938462,0.03938462,0.026256412,0.009846155,0.009846155,0.03938462,0.068923086,0.07876924,0.068923086,0.07876924,0.04266667,0.03938462,0.04594872,0.04266667,0.02297436,0.029538464,0.02297436,0.013128206,0.006564103,0.006564103,0.006564103,0.0032820515,0.0,0.0,0.0,0.032820515,0.15097436,0.15753847,0.052512825,0.01969231,0.009846155,0.04266667,0.17066668,0.46933338,1.0502565,0.72861546,0.4660513,0.27241027,0.18707694,0.24943592,0.5021539,0.86974365,0.93866676,0.69251287,0.5021539,0.508718,0.45620516,0.3511795,0.23958977,0.21333335,0.2297436,0.27241027,0.26912823,0.3446154,0.79425645,0.6826667,0.446359,0.39712822,0.77128214,1.7066668,2.4484105,1.719795,0.761436,0.2855385,0.45292312,0.60389745,0.36758977,0.14441027,0.08861539,0.08205129,0.068923086,0.07548718,0.07548718,0.052512825,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02297436,0.04594872,0.052512825,0.01969231,0.0032820515,0.006564103,0.009846155,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016410258,0.07548718,0.15097436,0.13456412,0.06564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.006564103,0.006564103,0.02297436,0.049230773,0.08533334,0.14441027,0.3511795,0.256,0.18707694,0.28225642,0.48246157,0.6104616,0.5284103,0.37415388,0.25271797,0.25928208,0.16082053,0.28882053,0.4660513,0.574359,0.53825647,0.4004103,0.26584616,0.16738462,0.118153855,0.12143591,0.15753847,0.2231795,0.36430773,0.6268718,1.0502565,0.8533334,0.9517949,1.1618463,1.3817437,1.6246156,1.6246156,1.8018463,2.7109745,4.312616,5.9667697,7.381334,8.5202055,9.8592825,11.362462,12.49477,13.548308,11.057232,10.039796,11.247591,11.168821,8.63836,6.166975,4.598154,4.0303593,3.82359,3.242667,2.0709746,1.6147693,1.9889232,2.1300514,1.8576412,1.5195899,1.5195899,2.1136413,3.4133337,4.013949,3.9089234,3.8432825,4.056616,4.2896414,4.457026,4.670359,4.1846156,3.05559,2.1333334,1.6213335,1.723077,1.9659488,1.972513,1.4703591,0.9288206,0.5677949,0.3511795,0.24615386,0.19692309,0.18379489,0.19692309,0.2297436,0.24287182,0.16738462,0.12471796,0.04594872,0.0,0.0,0.0,0.03938462,0.128,0.12471796,0.036102567,0.026256412,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.013128206,0.006564103,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.006564103,0.006564103,0.013128206,0.016410258,0.026256412,0.049230773,0.0951795,0.12143591,0.1148718,0.12143591,0.16082053,0.19692309,0.29210258,0.44964105,0.49887183,0.42994875,0.38400003,0.24615386,0.21333335,0.25271797,0.31507695,0.34789747,0.38728207,0.43651286,0.4135385,0.33476925,0.2986667,0.18051283,0.13128206,0.098461546,0.07548718,0.08861539,0.17066668,0.190359,0.17066668,0.11158975,0.02297436,0.032820515,0.03938462,0.036102567,0.029538464,0.006564103,0.013128206,0.013128206,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.016410258,0.016410258,0.026256412,0.029538464,0.032820515,0.032820515,0.049230773,0.07548718,0.09189744,0.13456412,0.22646156,0.3708718,0.3708718,0.41682056,0.571077,0.8598975,1.2504616,1.6705642,2.0775387,2.3105643,2.3105643,2.1070771,2.03159,2.0808206,2.0906668,1.9889232,1.8084104,1.595077,1.4342566,1.2800001,1.1355898,1.0568206,1.0666667,0.9321026,0.764718,0.63343596,0.56451285,0.51856416,0.53825647,0.5940513,0.6695385,0.77456415,1.0469744,1.1093334,1.142154,1.1946667,1.2077949,0.9878975,0.702359,0.5021539,0.47917953,0.69907695,1.1060513,1.086359,0.88943595,0.65312827,0.4266667,0.380718,0.42338464,0.5021539,0.56451285,0.5415385,0.42994875,0.36758977,0.34133336,0.33805132,0.318359,0.36430773,0.45620516,0.53825647,0.56451285,0.5152821,0.45620516,0.34133336,0.24943592,0.20348719,0.19692309,0.24287182,0.31507695,0.40697438,0.48574364,0.48246157,0.47261542,0.4397949,0.380718,0.3314872,0.35774362,0.6268718,0.9682052,1.204513,1.3062565,1.4145643,2.5271797,2.674872,2.7963078,3.3050258,4.089436,4.0500517,3.8531284,3.7874875,4.0992823,4.9920006,5.940513,6.816821,7.207385,6.701949,4.890257,4.2240005,4.279795,5.146257,5.9667697,4.9362054,4.8344617,6.567385,10.112,15.809642,24.359386,25.698463,21.609028,17.463797,16.833643,21.513847,22.75118,20.246977,15.320617,10.41395,9.104411,10.154668,8.723693,7.128616,6.8299494,8.444718,12.983796,11.575796,7.7390776,4.44718,4.1222568,4.460308,4.821334,5.21518,5.5532312,5.664821,5.8190775,6.370462,6.997334,7.3682055,7.1122055,6.4032826,5.9569235,5.7632823,5.720616,5.654975,5.671385,5.720616,5.7107697,5.546667,5.139693,1.8576412,2.7602053,3.6693337,4.204308,4.204308,3.751385,3.3280003,3.1770258,3.0030773,2.6847181,2.2711797,3.6463592,4.073026,4.2436924,4.466872,4.6802053,4.4832826,3.6758976,2.789744,2.038154,1.2996924,0.9747693,0.81394875,0.6268718,0.36758977,0.14441027,0.07876924,0.059076928,0.04266667,0.026256412,0.02297436,0.036102567,0.03938462,0.029538464,0.016410258,0.016410258,0.006564103,0.0032820515,0.0032820515,0.013128206,0.009846155,0.006564103,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.026256412,0.036102567,0.03938462,0.03938462,0.032820515,0.02297436,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.013128206,0.032820515,0.03938462,0.036102567,0.02297436,0.013128206,0.013128206,0.013128206,0.01969231,0.026256412,0.02297436,0.02297436,0.02297436,0.016410258,0.0032820515,0.0,0.0032820515,0.01969231,0.052512825,0.09189744,0.12143591,0.09189744,0.07548718,0.06235898,0.052512825,0.06235898,0.072205134,0.06564103,0.049230773,0.036102567,0.029538464,0.016410258,0.009846155,0.01969231,0.04266667,0.072205134,0.13128206,0.27241027,0.25271797,0.09189744,0.072205134,0.032820515,0.068923086,0.18707694,0.36430773,0.5349744,0.5546667,0.5349744,0.3708718,0.12143591,0.026256412,0.07876924,0.108307704,0.09189744,0.049230773,0.049230773,0.052512825,0.04594872,0.04594872,0.098461546,0.28225642,0.6695385,1.0108719,1.0502565,0.9353847,1.204513,0.7778462,0.34789747,0.18707694,0.36102566,0.7220513,0.9156924,0.58420515,0.24615386,0.18379489,0.4266667,0.5546667,0.23302566,0.0032820515,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.006564103,0.0032820515,0.006564103,0.026256412,0.055794876,0.02297436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.013128206,0.01969231,0.04594872,0.07548718,0.08205129,0.049230773,0.07548718,0.09189744,0.19692309,0.45292312,0.8992821,1.1848207,0.9878975,0.6104616,0.30194873,0.25271797,0.20348719,0.35446155,0.53825647,0.65312827,0.6465641,0.51856416,0.3708718,0.26584616,0.21333335,0.14441027,0.14441027,0.23302566,0.47261542,0.955077,1.8116925,1.5622566,1.591795,1.9593848,2.4516926,2.5665643,1.9790771,1.7066668,2.3236926,3.5052311,4.0402055,5.658257,7.5979495,9.45559,11.270565,13.522053,17.473642,11.782565,7.02359,6.99077,8.697436,7.565129,5.1331286,3.442872,2.934154,2.4549747,1.9396925,1.4802053,1.2504616,1.2406155,1.2406155,1.2800001,1.2438976,1.7296412,2.92759,4.634257,4.57518,4.3027697,4.1813335,4.352,4.7458467,4.4045134,4.3027697,3.6890259,2.5731285,1.7394873,1.5491283,1.7755898,1.8018463,1.4473847,0.955077,0.7844103,0.6826667,0.5874872,0.49230772,0.44964105,0.42338464,0.36758977,0.36758977,0.380718,0.24287182,0.14769232,0.049230773,0.0,0.0,0.0,0.01969231,0.18707694,0.20348719,0.059076928,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.006564103,0.0032820515,0.0,0.0,0.0,0.009846155,0.016410258,0.013128206,0.013128206,0.013128206,0.0032820515,0.013128206,0.049230773,0.0951795,0.128,0.14112821,0.14112821,0.13456412,0.13784617,0.28882053,0.46276927,0.45620516,0.30194873,0.28882053,0.19692309,0.14769232,0.20020515,0.3511795,0.5316923,0.5940513,0.571077,0.508718,0.4397949,0.38400003,0.2231795,0.14441027,0.0951795,0.068923086,0.108307704,0.23958977,0.30194873,0.3117949,0.25928208,0.0951795,0.059076928,0.03938462,0.02297436,0.013128206,0.013128206,0.013128206,0.006564103,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.013128206,0.016410258,0.02297436,0.04594872,0.06235898,0.07548718,0.08205129,0.08533334,0.098461546,0.10502565,0.15425642,0.25928208,0.42338464,0.43651286,0.508718,0.6104616,0.7417436,0.9321026,1.401436,1.8904617,2.2219489,2.3236926,2.225231,2.349949,2.5074873,2.5862565,2.5304618,2.359795,2.1169233,1.9495386,1.7263591,1.4375386,1.1946667,1.1355898,1.0601027,0.9353847,0.8172308,0.8336411,0.7089231,0.6826667,0.67610264,0.6465641,0.5874872,0.67282057,0.82379496,1.1257436,1.4867693,1.6180514,1.086359,0.72861546,0.4955898,0.4135385,0.571077,1.1060513,1.142154,0.9878975,0.761436,0.37743592,0.18379489,0.15753847,0.22646156,0.318359,0.36430773,0.3446154,0.3708718,0.40697438,0.4201026,0.36430773,0.33476925,0.40369233,0.53825647,0.67938465,0.7318975,0.6465641,0.51856416,0.4135385,0.36430773,0.3511795,0.35774362,0.37415388,0.39056414,0.40369233,0.39384618,0.4594872,0.4955898,0.49230772,0.42994875,0.27569234,0.41025645,0.8402052,1.2996924,1.5819489,1.529436,2.5435898,2.7076926,2.609231,2.6551797,3.0851285,3.373949,3.7776413,4.525949,5.72718,7.397744,8.1755905,8.845129,9.232411,8.966565,7.4699492,5.904411,5.169231,5.927385,7.1614366,6.193231,6.121026,7.7292314,10.236719,14.355694,22.294975,28.901747,27.40513,22.180105,17.900309,19.551182,22.724924,22.665848,18.665028,13.00677,10.981745,11.697231,10.453334,8.438154,7.125334,8.297027,9.531077,7.788308,5.287385,3.5807183,3.56759,3.7054362,3.95159,4.3684106,4.8705645,5.218462,5.3169236,5.730462,6.340924,6.9054365,7.0465646,6.554257,6.0356927,5.687795,5.4974365,5.2414365,5.1167183,5.10359,5.113436,5.031385,4.7294364,2.3958976,3.7251284,4.919795,5.366154,4.9952826,4.2863593,3.446154,3.190154,3.2262566,3.2722054,3.0523078,2.9538465,3.2689233,4.20759,5.290667,5.3398976,4.890257,4.785231,4.6145644,3.9975388,2.5928206,1.9462565,1.4572309,1.0535386,0.67938465,0.28882053,0.118153855,0.049230773,0.02297436,0.013128206,0.0,0.013128206,0.016410258,0.016410258,0.016410258,0.016410258,0.026256412,0.013128206,0.0,0.009846155,0.04594872,0.032820515,0.02297436,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.009846155,0.0,0.0,0.013128206,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.016410258,0.013128206,0.0,0.0,0.009846155,0.016410258,0.013128206,0.0,0.0,0.0,0.013128206,0.02297436,0.0,0.013128206,0.02297436,0.06235898,0.12143591,0.18379489,0.18379489,0.17394873,0.12471796,0.06235898,0.06235898,0.072205134,0.0951795,0.11158975,0.1148718,0.09189744,0.01969231,0.01969231,0.09189744,0.21989745,0.36758977,0.318359,0.13128206,0.026256412,0.072205134,0.18379489,0.08533334,0.02297436,0.006564103,0.02297436,0.04594872,0.19364104,0.37415388,0.3249231,0.08861539,0.016410258,0.026256412,0.03938462,0.026256412,0.0,0.0,0.013128206,0.016410258,0.016410258,0.15753847,0.7318975,1.8445129,2.6420515,2.6715899,1.8510771,0.47261542,0.0951795,0.0,0.0,0.0032820515,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.036102567,0.036102567,0.02297436,0.016410258,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.036102567,0.06564103,0.059076928,0.02297436,0.0,0.036102567,0.09189744,0.19692309,0.36430773,0.5940513,0.7417436,0.61374366,0.5152821,0.508718,0.4135385,0.3511795,0.28225642,0.256,0.34133336,0.6104616,0.7581539,0.74830776,0.60061544,0.38728207,0.2297436,0.18051283,0.21333335,0.38400003,0.85005134,1.8609232,2.5206156,2.9505644,3.3050258,3.5314875,3.370667,2.2383592,1.7690258,1.9232821,2.3433847,2.3794873,3.0030773,3.8367183,4.525949,5.074052,5.8453336,7.7259493,5.933949,4.699898,5.3891287,6.5017443,5.1331286,2.7667694,1.9068719,2.5009232,1.9528207,1.6738462,1.4178462,1.2307693,1.1454359,1.204513,1.6443079,1.3423591,2.2219489,4.342154,5.904411,6.038975,5.4514875,4.6933336,4.453744,5.540103,4.2207184,3.2951798,2.546872,1.9232821,1.5556924,1.9232821,2.3991797,2.0939488,1.1749744,0.86974365,1.1881026,1.4867693,1.4998976,1.2176411,0.8992821,0.92553854,0.6826667,0.38400003,0.14769232,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.016410258,0.009846155,0.0,0.0,0.0,0.009846155,0.016410258,0.013128206,0.0,0.0,0.0,0.02297436,0.08205129,0.16738462,0.14441027,0.19364104,0.2100513,0.16082053,0.07548718,0.101743594,0.13456412,0.14112821,0.20348719,0.5349744,0.36430773,0.36758977,0.45620516,0.5677949,0.64000005,0.5677949,0.5021539,0.40697438,0.2855385,0.21333335,0.14112821,0.07548718,0.052512825,0.068923086,0.108307704,0.18051283,0.27241027,0.3249231,0.31507695,0.2297436,0.108307704,0.049230773,0.01969231,0.0,0.0,0.013128206,0.016410258,0.02297436,0.02297436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.02297436,0.04594872,0.068923086,0.0951795,0.108307704,0.108307704,0.12143591,0.13456412,0.16410258,0.23302566,0.3249231,0.4135385,0.3249231,0.42338464,0.54482055,0.67282057,0.9321026,1.4309745,1.8412309,2.1103592,2.284308,2.5173335,2.8488207,3.058872,3.1507695,3.114667,2.9440002,2.7142565,2.481231,2.169436,1.7952822,1.463795,1.2077949,1.0994873,1.0929232,1.1388719,1.1749744,0.9419488,0.8041026,0.77128214,0.7844103,0.6859488,0.6629744,0.79425645,1.0436924,1.2865642,1.3128207,0.95835906,0.69579494,0.5316923,0.47261542,0.5349744,0.5218462,0.58420515,0.74830776,0.8533334,0.5481026,0.256,0.15425642,0.13784617,0.14441027,0.16738462,0.2297436,0.318359,0.37743592,0.37415388,0.28882053,0.20348719,0.2297436,0.38728207,0.5874872,0.6104616,0.574359,0.49887183,0.45292312,0.4594872,0.5349744,0.62030774,0.6301539,0.60061544,0.5415385,0.44307697,0.42994875,0.56451285,0.77128214,0.8467693,0.45620516,0.34789747,0.47589746,0.8795898,1.4309745,1.847795,1.6377437,1.7329233,2.7273848,4.023795,3.8301542,3.6102567,3.6824617,3.9712822,4.457026,5.1889234,5.028103,7.325539,8.802463,8.4972315,7.752206,6.311385,5.8486156,5.973334,6.669129,8.316719,6.498462,4.7228723,5.907693,11.798975,22.980925,36.480003,38.104618,32.019695,23.332104,18.097233,14.043899,12.691693,13.728822,15.694771,15.977027,13.338258,10.371283,8.12636,7.1515903,7.4929237,7.896616,7.125334,5.284103,3.3969233,3.4330258,2.665026,2.3893335,2.5961027,3.131077,3.692308,4.082872,4.4832826,4.9526157,5.58277,6.485334,6.373744,6.045539,5.8190775,5.7534366,5.6320004,5.21518,4.900103,4.650667,4.450462,4.3027697,1.2242053,1.7920002,2.2022567,2.5928206,2.9472823,3.0785644,2.9997952,3.058872,2.9997952,2.7109745,2.1956925,2.284308,3.1967182,4.4964104,5.5663595,5.5958977,3.9548721,2.9013336,2.6256413,2.8717952,2.9243078,2.7831798,2.5796926,2.4385643,2.1891284,1.3883078,0.67938465,0.2986667,0.15425642,0.13784617,0.14769232,0.098461546,0.0951795,0.072205134,0.032820515,0.052512825,0.055794876,0.04266667,0.026256412,0.013128206,0.009846155,0.016410258,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.013128206,0.0032820515,0.0032820515,0.0032820515,0.0,0.0,0.0032820515,0.009846155,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0032820515,0.0,0.0,0.0032820515,0.0032820515,0.0032820515,0.013128206,0.02297436,0.02297436,0.016410258,0.0032820515,0.0,0.0032820515,0.032820515,0.072205134,0.108307704,0.17066668,0.2100513,0.22646156,0.24943592,0.27241027,0.23302566,0.19692309,0.15425642,0.13128206,0.13128206,0.1148718,0.072205134,0.04266667,0.049230773,0.08205129,0.108307704,0.09189744,0.049230773,0.01969231,0.013128206,0.036102567,0.016410258,0.072205134,0.09189744,0.059076928,0.04594872,0.0951795,0.128,0.13456412,0.11158975,0.07548718,0.059076928,0.049230773,0.04266667,0.032820515,0.013128206,0.0032820515,0.009846155,0.15097436,0.36430773,0.39056414,0.446359,0.58092314,0.571077,0.3708718,0.0951795,0.01969231,0.256,0.42338464,0.3314872,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.32820517,0.32164106,0.15753847,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.01969231,0.029538464,0.026256412,0.013128206,0.03938462,0.18051283,0.318359,0.38400003,0.3511795,0.42994875,0.28225642,0.39056414,0.80738467,1.1684103,0.9321026,0.4594872,0.17066668,0.17723078,0.28225642,0.50543594,0.8369231,1.017436,0.9747693,0.81394875,0.8041026,0.6432821,0.764718,1.1815386,1.4834872,1.8871796,2.6880002,3.7284105,4.630975,4.7622566,4.0467696,3.2984617,4.309334,6.678975,7.8014364,6.9677954,6.7249236,5.6254363,4.1813335,4.893539,6.7610264,6.8430777,6.196513,5.47118,4.900103,3.5741541,2.4320002,1.7723079,1.5031796,1.1585642,1.2209232,1.3817437,1.4178462,1.4145643,1.7657437,2.1169233,2.5862565,3.4756925,4.5390773,4.9887185,4.089436,3.754667,3.8564105,4.010667,3.5741541,3.045744,2.7306669,2.3105643,1.7165129,1.1158975,1.2012309,1.4802053,1.3357949,0.74830776,0.29538465,0.47589746,0.84348726,0.76800007,0.35446155,0.44964105,0.8336411,0.78769237,0.47261542,0.118153855,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0032820515,0.0,0.0,0.029538464,0.03938462,0.052512825,0.16738462,0.20348719,0.20020515,0.17394873,0.13456412,0.08861539,0.17066668,0.21333335,0.23302566,0.3249231,0.65641034,1.0896411,1.142154,0.9124103,0.7515898,1.276718,0.9878975,0.57764107,0.32164106,0.27569234,0.24943592,0.17723078,0.12143591,0.10502565,0.14441027,0.23958977,0.3052308,0.256,0.16738462,0.108307704,0.118153855,0.06564103,0.03938462,0.029538464,0.02297436,0.013128206,0.013128206,0.006564103,0.02297436,0.052512825,0.036102567,0.026256412,0.032820515,0.02297436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.026256412,0.02297436,0.009846155,0.032820515,0.068923086,0.118153855,0.15753847,0.18379489,0.19692309,0.128,0.15425642,0.23630771,0.3446154,0.44964105,0.5284103,0.64000005,0.69251287,0.7220513,0.88287187,1.2471796,1.7526156,2.2711797,2.6847181,2.9078977,3.170462,3.1803079,3.1934361,3.2131286,2.993231,2.7142565,2.5337439,2.3269746,2.0545642,1.7952822,1.6738462,1.5983591,1.4900514,1.3522053,1.2603078,1.3883078,1.4802053,1.394872,1.1881026,1.1027694,0.9616411,0.79097444,0.6695385,0.62030774,0.60389745,0.571077,0.45620516,0.4201026,0.5513847,0.8763078,1.1093334,1.0404103,1.1060513,1.2242053,0.7811283,0.48902568,0.3446154,0.26584616,0.21333335,0.16738462,0.17066668,0.27241027,0.32820517,0.28882053,0.20348719,0.17723078,0.2297436,0.32164106,0.4201026,0.512,0.52512825,0.49887183,0.48574364,0.508718,0.58420515,0.6695385,0.6498462,0.57764107,0.5021539,0.49230772,0.48902568,0.5316923,0.6170257,0.6859488,0.6170257,0.5152821,0.5513847,0.8369231,1.3095386,1.723077,1.6836925,1.5097437,1.4375386,1.7723079,2.9144619,3.0851285,3.4034874,3.8301542,4.1517954,3.9548721,3.9318976,4.9887185,6.3277955,7.4929237,8.349539,7.817847,6.8955903,6.3343596,6.485334,7.3025646,5.717334,4.7524104,5.7403083,9.238976,15.02195,21.376001,28.642464,34.048004,35.840004,33.270157,24.421745,16.764719,13.869949,16.25272,21.395695,21.083899,15.658668,10.203898,7.529026,8.162462,9.45559,8.579283,6.8266673,4.972308,3.2623591,2.4746668,2.3105643,2.4943593,2.8160002,3.1442053,3.318154,3.5905645,3.9154875,4.332308,4.972308,5.3891287,5.586052,5.5762057,5.5269747,5.7764106,5.586052,5.159385,4.772103,4.571898,4.571898,1.1520001,1.1126155,1.214359,1.5195899,1.9035898,2.0644104,1.8051283,1.6771283,1.6344616,1.6147693,1.5261539,1.529436,1.9003079,2.546872,3.3641028,4.2601027,4.348718,3.8990772,3.318154,2.92759,2.9702566,2.6715899,2.737231,2.7470772,2.4418464,1.7362052,1.4145643,1.1913847,0.83035904,0.38728207,0.20020515,0.11158975,0.08205129,0.059076928,0.029538464,0.02297436,0.04594872,0.049230773,0.032820515,0.013128206,0.0,0.0032820515,0.0032820515,0.009846155,0.029538464,0.04594872,0.029538464,0.02297436,0.01969231,0.02297436,0.016410258,0.0032820515,0.006564103,0.009846155,0.006564103,0.0,0.0,0.0032820515,0.0032820515,0.0032820515,0.009846155,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.026256412,0.01969231,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.03938462,0.04266667,0.02297436,0.0,0.0,0.006564103,0.029538464,0.049230773,0.06235898,0.08533334,0.15753847,0.19364104,0.2100513,0.20348719,0.14769232,0.13456412,0.128,0.12143591,0.108307704,0.0951795,0.07876924,0.049230773,0.026256412,0.01969231,0.026256412,0.20676924,0.21661541,0.128,0.02297436,0.009846155,0.0032820515,0.03938462,0.068923086,0.072205134,0.055794876,0.04266667,0.04266667,0.08533334,0.14112821,0.101743594,0.055794876,0.032820515,0.026256412,0.026256412,0.016410258,0.016410258,0.02297436,0.08533334,0.16738462,0.12143591,0.03938462,0.026256412,0.01969231,0.0,0.0,0.0,0.128,0.2100513,0.16738462,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.04594872,0.2297436,0.2100513,0.098461546,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.006564103,0.0,0.0,0.0,0.006564103,0.006564103,0.0032820515,0.01969231,0.068923086,0.190359,0.20348719,0.098461546,0.04266667,0.029538464,0.0951795,0.190359,0.30851284,0.48246157,0.7122052,0.5481026,0.5218462,0.7778462,1.0929232,0.98133343,0.6301539,0.38728207,0.35446155,0.4004103,0.636718,0.827077,0.8960001,0.8960001,1.017436,1.2931283,1.3522053,1.3029745,1.2438976,1.2406155,1.6278975,2.3663592,3.570872,5.0084105,6.0717955,5.346462,4.824616,5.2414365,6.3442054,6.8955903,6.941539,6.298257,5.21518,4.4898467,5.477744,6.701949,6.51159,5.280821,3.8071797,3.3280003,3.255795,2.9144619,2.297436,1.5655385,1.0535386,1.1979488,1.4375386,1.7460514,2.100513,2.484513,2.9965131,3.508513,3.9122055,4.0992823,3.9548721,2.7667694,2.2449234,2.3368206,2.7241027,2.8356924,2.806154,2.3466668,1.8412309,1.595077,1.8674873,1.9298463,1.6968206,1.204513,0.6301539,0.28882053,0.23958977,0.3314872,0.26584616,0.08205129,0.15097436,0.3446154,0.3446154,0.2100513,0.04594872,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.01969231,0.009846155,0.009846155,0.016410258,0.026256412,0.026256412,0.026256412,0.009846155,0.0,0.0,0.0,0.0,0.013128206,0.01969231,0.026256412,0.07548718,0.12471796,0.13128206,0.12143591,0.108307704,0.108307704,0.17723078,0.27897438,0.36102566,0.40369233,0.40369233,0.79097444,0.9747693,0.8763078,0.69579494,0.9124103,0.76800007,0.51856416,0.36102566,0.32164106,0.24943592,0.21333335,0.20020515,0.21333335,0.25271797,0.3117949,0.41025645,0.35446155,0.2297436,0.12143591,0.13784617,0.072205134,0.12143591,0.14441027,0.101743594,0.052512825,0.029538464,0.009846155,0.013128206,0.032820515,0.026256412,0.02297436,0.029538464,0.029538464,0.01969231,0.01969231,0.0032820515,0.0,0.0,0.0032820515,0.009846155,0.013128206,0.016410258,0.01969231,0.01969231,0.029538464,0.06564103,0.098461546,0.13784617,0.17723078,0.20348719,0.14769232,0.17066668,0.23302566,0.33805132,0.512,0.58420515,0.6170257,0.6301539,0.67282057,0.84348726,1.3193847,1.9200002,2.4352822,2.7437952,2.7864618,2.7241027,2.7011285,2.7864618,2.8980515,2.806154,2.6945643,2.6026669,2.477949,2.300718,2.0775387,2.0151796,2.0676925,1.9856411,1.723077,1.4572309,1.4769232,1.463795,1.204513,0.82379496,0.764718,0.955077,0.9419488,0.764718,0.5152821,0.33476925,0.3249231,0.30194873,0.31507695,0.4266667,0.7220513,1.1257436,1.1684103,1.2012309,1.2077949,0.8205129,0.65312827,0.6104616,0.58092314,0.51856416,0.45292312,0.30851284,0.25928208,0.2231795,0.16738462,0.118153855,0.15753847,0.21989745,0.26584616,0.29210258,0.3511795,0.5284103,0.5940513,0.57764107,0.5349744,0.5481026,0.65641034,0.71548724,0.67610264,0.57764107,0.5415385,0.7318975,0.8402052,0.86646163,0.83035904,0.7844103,0.7515898,0.9353847,1.1618463,1.4441026,1.9692309,2.861949,3.1376412,2.4451284,1.5622566,2.412308,3.2722054,4.073026,4.6080003,4.6802053,4.1124105,3.692308,4.0434875,4.70318,5.4941545,6.5411286,6.170257,6.5805135,7.6931286,9.051898,9.82318,8.129642,6.7872825,6.692103,8.113232,10.706052,14.106257,20.207592,26.998156,32.44636,34.49108,29.994669,24.365952,20.634258,19.337847,18.51077,19.02277,15.684924,12.251899,10.735591,11.408411,11.493745,9.67877,7.381334,5.3431797,3.6036925,3.0391798,2.993231,3.0785644,3.1442053,3.2886157,3.4133337,3.7284105,4.125539,4.5489235,5.0149746,5.366154,5.398975,5.35959,5.402257,5.5762057,5.435077,5.097026,4.8016415,4.6605134,4.6769233,1.5885129,1.3620514,1.3620514,1.6410258,2.0217438,2.1103592,1.9232821,2.0020514,2.3236926,2.7569232,3.0391798,2.5961027,2.2711797,2.3827693,3.0490258,4.194462,4.650667,4.8016415,4.325744,3.446154,2.9210258,2.612513,2.7798977,2.9210258,2.7831798,2.3663592,2.166154,1.9167181,1.4309745,0.7975385,0.40369233,0.27241027,0.2231795,0.190359,0.14441027,0.08533334,0.072205134,0.07548718,0.07548718,0.072205134,0.055794876,0.03938462,0.026256412,0.032820515,0.059076928,0.06564103,0.03938462,0.029538464,0.026256412,0.026256412,0.016410258,0.006564103,0.013128206,0.016410258,0.016410258,0.0,0.0032820515,0.0032820515,0.0,0.0032820515,0.009846155,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.026256412,0.01969231,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.029538464,0.029538464,0.01969231,0.006564103,0.006564103,0.009846155,0.01969231,0.026256412,0.029538464,0.029538464,0.08205129,0.118153855,0.12143591,0.08861539,0.036102567,0.049230773,0.08205129,0.101743594,0.09189744,0.07548718,0.06564103,0.04266667,0.01969231,0.0032820515,0.016410258,0.20676924,0.24287182,0.18051283,0.098461546,0.08861539,0.052512825,0.029538464,0.052512825,0.0951795,0.06564103,0.0951795,0.12471796,0.16738462,0.19692309,0.17394873,0.11158975,0.055794876,0.02297436,0.016410258,0.016410258,0.02297436,0.01969231,0.009846155,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.0032820515,0.0,0.0,0.013128206,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.04594872,0.068923086,0.052512825,0.02297436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0,0.006564103,0.006564103,0.013128206,0.013128206,0.006564103,0.013128206,0.026256412,0.036102567,0.029538464,0.026256412,0.06235898,0.17066668,0.3314872,0.33476925,0.18707694,0.1148718,0.068923086,0.052512825,0.08533334,0.2100513,0.46933338,0.77128214,0.7089231,0.6235898,0.6662565,0.8041026,0.92225647,1.0043077,0.9944616,0.92553854,0.92553854,0.98133343,0.9353847,0.8730257,0.8795898,1.0469744,1.719795,2.0250258,2.0512822,1.9889232,2.1333334,2.5632823,3.0687182,3.7185643,4.4373336,5.024821,4.634257,4.594872,4.6080003,4.588308,4.6769233,5.464616,5.0871797,4.4800005,4.315898,5.0084105,5.723898,5.142975,4.0434875,3.1245131,3.0194874,3.4231799,3.1573336,2.5238976,1.9003079,1.7427694,2.1070771,2.477949,3.3050258,4.2929235,4.394667,4.096,4.2830772,4.309334,3.9417439,3.3312824,2.2514873,1.8149745,1.9954873,2.5271797,2.9144619,2.7175386,1.9265642,1.3883078,1.5163078,2.2711797,2.2711797,1.7263591,1.0929232,0.60389745,0.27241027,0.14112821,0.068923086,0.036102567,0.026256412,0.01969231,0.01969231,0.01969231,0.009846155,0.0032820515,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.01969231,0.016410258,0.02297436,0.036102567,0.04266667,0.026256412,0.026256412,0.009846155,0.0,0.0,0.0,0.0032820515,0.006564103,0.006564103,0.013128206,0.02297436,0.06564103,0.1148718,0.15753847,0.19364104,0.23302566,0.23630771,0.30851284,0.39056414,0.41025645,0.26256412,0.5349744,0.78769237,0.90584624,0.8795898,0.8041026,0.6235898,0.49887183,0.42994875,0.38728207,0.29210258,0.33476925,0.33805132,0.3314872,0.33805132,0.36758977,0.48902568,0.4660513,0.3511795,0.21661541,0.16082053,0.13456412,0.23630771,0.26912823,0.20348719,0.17394873,0.09189744,0.036102567,0.01969231,0.026256412,0.026256412,0.016410258,0.01969231,0.026256412,0.029538464,0.01969231,0.0032820515,0.0032820515,0.006564103,0.006564103,0.016410258,0.009846155,0.006564103,0.013128206,0.026256412,0.036102567,0.068923086,0.08533334,0.11158975,0.14769232,0.17394873,0.16082053,0.18707694,0.23302566,0.32164106,0.50543594,0.5973334,0.6301539,0.65312827,0.7253334,0.88615394,1.3751796,1.9429746,2.3762052,2.5764105,2.5600002,2.4484105,2.4943593,2.5928206,2.6880002,2.7602053,2.8291285,2.789744,2.6912823,2.5600002,2.4320002,2.6223593,2.8422565,2.7536411,2.3302567,1.847795,1.7066668,1.6804104,1.4408206,1.0272821,0.8402052,1.214359,1.3620514,1.1815386,0.764718,0.39056414,0.26912823,0.25928208,0.26912823,0.29538465,0.42994875,0.8369231,1.0436924,1.1290257,1.0896411,0.80738467,0.7122052,0.78769237,0.8730257,0.88615394,0.84348726,0.6104616,0.35446155,0.17066668,0.08205129,0.059076928,0.15097436,0.26256412,0.30851284,0.27897438,0.23630771,0.43323082,0.5973334,0.65641034,0.6170257,0.5677949,0.7056411,0.8598975,0.90256417,0.81066674,0.67282057,0.7515898,0.8467693,1.0043077,1.1848207,1.2307693,1.1454359,1.3193847,1.463795,1.657436,2.359795,3.8662567,4.5095387,3.764513,2.4385643,2.6617439,4.092718,5.5171285,6.160411,5.756718,4.5423594,3.817026,3.7940516,3.9548721,4.2502565,5.080616,4.630975,5.930667,8.274052,10.528821,11.136001,9.416205,7.719385,7.207385,8.323282,10.778257,13.121642,16.137848,20.210873,24.832003,28.612925,29.075695,27.72349,26.377848,24.825438,20.83118,19.715284,16.699078,14.345847,13.705847,14.34913,14.267078,11.464206,8.192,5.671385,4.07959,3.5380516,3.3509746,3.3378465,3.4560003,3.7973337,4.138667,4.529231,4.7983594,4.9296412,5.0642056,5.1987696,5.172513,5.1889234,5.297231,5.3694363,5.3103595,5.0871797,4.827898,4.6211286,4.4996924,1.9528207,1.8543591,1.8379488,2.1070771,2.5665643,2.7963078,3.0654361,3.6102567,4.3684106,5.146257,5.6287184,4.8836927,4.4274874,4.637539,5.362872,5.9470773,4.841026,4.886975,4.8804107,4.2568207,3.0916924,2.9144619,2.9636924,3.1770258,3.3575387,3.1934361,2.6518977,2.162872,1.7099489,1.2603078,0.79097444,0.62030774,0.5513847,0.49887183,0.41025645,0.27569234,0.17066668,0.14769232,0.16738462,0.18707694,0.15425642,0.101743594,0.06235898,0.052512825,0.059076928,0.03938462,0.02297436,0.01969231,0.02297436,0.029538464,0.013128206,0.013128206,0.016410258,0.01969231,0.02297436,0.0,0.013128206,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.013128206,0.0032820515,0.009846155,0.02297436,0.029538464,0.029538464,0.029538464,0.04266667,0.04594872,0.032820515,0.0,0.009846155,0.04266667,0.08205129,0.10502565,0.07876924,0.055794876,0.03938462,0.02297436,0.006564103,0.013128206,0.032820515,0.07548718,0.12143591,0.15425642,0.16738462,0.128,0.101743594,0.118153855,0.14769232,0.101743594,0.190359,0.24615386,0.24615386,0.2231795,0.23302566,0.17723078,0.098461546,0.04266667,0.01969231,0.013128206,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.006564103,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.016410258,0.009846155,0.006564103,0.03938462,0.016410258,0.013128206,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.01969231,0.026256412,0.02297436,0.013128206,0.02297436,0.02297436,0.02297436,0.02297436,0.029538464,0.04266667,0.07548718,0.0951795,0.101743594,0.11158975,0.15425642,0.24615386,0.33476925,0.36430773,0.3249231,0.26912823,0.15753847,0.101743594,0.108307704,0.16410258,0.26584616,0.47917953,0.60061544,0.67282057,0.7318975,0.8041026,0.955077,1.3522053,1.5753847,1.5655385,1.6016412,1.4998976,1.3850257,1.3292309,1.3161026,1.2242053,1.9626669,2.281026,2.5435898,2.92759,3.4330258,4.023795,4.3290257,4.135385,3.5052311,2.7503593,2.9669745,3.2131286,3.2951798,3.318154,3.7054362,4.5489235,4.841026,4.578462,4.076308,3.9811285,4.598154,4.2601027,4.1189747,4.338872,4.1091285,3.7940516,3.1606157,2.6289232,2.4648206,2.7503593,3.245949,3.95159,5.4547696,7.128616,7.1483083,5.671385,5.356308,5.2381544,4.70318,3.501949,2.5895386,2.5829747,3.045744,3.4330258,3.0916924,2.294154,1.3981539,1.0535386,1.339077,1.7690258,1.5556924,1.0962052,0.7384616,0.49887183,0.08533334,0.04594872,0.02297436,0.006564103,0.0,0.0,0.006564103,0.006564103,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.026256412,0.036102567,0.029538464,0.0,0.0032820515,0.0,0.0,0.0,0.0,0.013128206,0.013128206,0.006564103,0.0032820515,0.02297436,0.052512825,0.14112821,0.23302566,0.3052308,0.35446155,0.318359,0.30194873,0.33805132,0.38400003,0.33805132,0.636718,0.9189744,1.1290257,1.1979488,1.017436,0.65312827,0.49230772,0.43651286,0.40697438,0.33476925,0.41682056,0.4266667,0.4135385,0.41682056,0.4660513,0.58092314,0.56123084,0.45620516,0.33476925,0.26256412,0.3249231,0.39056414,0.38400003,0.32820517,0.35774362,0.18379489,0.07876924,0.04266667,0.04594872,0.03938462,0.01969231,0.016410258,0.01969231,0.01969231,0.0,0.0,0.009846155,0.016410258,0.01969231,0.01969231,0.0032820515,0.006564103,0.013128206,0.02297436,0.04594872,0.06564103,0.08205129,0.101743594,0.128,0.15097436,0.17066668,0.20348719,0.25271797,0.32820517,0.46276927,0.64000005,0.77456415,0.86974365,0.9485129,1.0535386,1.4441026,1.8871796,2.2350771,2.4188719,2.4582565,2.5796926,2.6683078,2.6847181,2.6945643,2.8553848,2.9702566,2.9801028,2.9243078,2.8750772,2.930872,3.4264617,3.7448208,3.620103,3.05559,2.3466668,2.1792822,2.3696413,2.356513,2.0053334,1.585231,1.8149745,1.9626669,1.7329233,1.1618463,0.6170257,0.37743592,0.31507695,0.29210258,0.256,0.23302566,0.4955898,0.79097444,0.98133343,0.9911796,0.8008206,0.69907695,0.8467693,1.0371283,1.1454359,1.1520001,0.9156924,0.512,0.20020515,0.068923086,0.036102567,0.14769232,0.3314872,0.4201026,0.36102566,0.21333335,0.256,0.45620516,0.6465641,0.7253334,0.67282057,0.79097444,0.9321026,1.083077,1.2274873,1.3095386,0.8598975,0.6465641,0.90256417,1.4506668,1.7033848,1.5261539,1.4802053,1.5195899,1.8051283,2.7109745,4.0008206,4.8049235,4.7392826,4.059898,3.6562054,4.7655387,6.413129,7.1548724,6.419693,4.529231,3.7349746,3.498667,3.5872824,4.027077,5.097026,4.709744,5.7140517,7.712821,9.744411,10.259693,8.969847,7.4765134,7.4830775,9.573745,13.200411,15.136822,16.59077,18.346668,20.558771,22.738052,23.955694,25.071592,27.044106,29.03631,28.406157,25.252104,20.680206,17.293129,16.164104,16.83036,16.981335,13.403898,9.317744,6.373744,4.673641,3.8104618,3.2262566,3.2098465,3.8400004,5.0084105,5.83877,5.9634876,5.612308,5.077334,4.7294364,4.670359,4.7917953,4.972308,5.1265645,5.1987696,5.32677,5.221744,4.9460516,4.588308,4.2568207,1.6475899,1.5491283,1.6278975,1.7362052,1.9167181,2.3794873,2.5993848,2.7109745,3.1540515,4.027077,5.0674877,5.2611284,5.7140517,6.5312824,7.4371285,7.765334,6.2785645,5.6943593,5.8092313,5.7403083,3.9220517,3.190154,2.9604106,3.0162053,3.117949,3.0227695,2.4713848,2.1070771,1.8051283,1.5097437,1.204513,0.98461545,0.88615394,0.84348726,0.761436,0.51856416,0.34789747,0.27897438,0.27897438,0.28882053,0.2297436,0.108307704,0.049230773,0.02297436,0.016410258,0.016410258,0.026256412,0.029538464,0.036102567,0.036102567,0.0,0.013128206,0.016410258,0.016410258,0.013128206,0.0,0.013128206,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01969231,0.029538464,0.029538464,0.029538464,0.029538464,0.02297436,0.016410258,0.013128206,0.0,0.0,0.009846155,0.059076928,0.1148718,0.09189744,0.06564103,0.052512825,0.03938462,0.02297436,0.0,0.0,0.009846155,0.016410258,0.02297436,0.04594872,0.14441027,0.26912823,0.2986667,0.23630771,0.19692309,0.16082053,0.12471796,0.08861539,0.06235898,0.06235898,0.02297436,0.068923086,0.08205129,0.036102567,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.016410258,0.009846155,0.03938462,0.19692309,0.03938462,0.04594872,0.04594872,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.04594872,0.0951795,0.08861539,0.068923086,0.06235898,0.06235898,0.06235898,0.052512825,0.059076928,0.07876924,0.09189744,0.1148718,0.17723078,0.256,0.3249231,0.3511795,0.21661541,0.2297436,0.41682056,0.63343596,0.5481026,0.23302566,0.13456412,0.18379489,0.27897438,0.28882053,0.37415388,0.5973334,0.9156924,1.2438976,1.463795,1.0371283,1.0043077,1.204513,1.5425643,1.9692309,2.284308,2.3926156,2.3926156,2.284308,1.9692309,1.7001027,1.6508719,1.7920002,2.1267693,2.7011285,3.8498464,4.1091285,3.889231,3.629949,3.8006158,3.9581542,3.639795,3.190154,3.1081028,4.059898,5.6943593,6.5444107,6.6395903,6.2785645,5.9963083,6.678975,6.705231,6.678975,6.560821,5.6451287,4.5587697,3.9680004,3.9351797,3.9712822,3.006359,2.7011285,3.8596926,5.802667,7.781744,9.002667,8.4053335,7.4765134,7.072821,6.738052,4.699898,3.698872,3.895795,4.0369234,3.5052311,2.3335385,1.332513,0.8533334,0.761436,0.84348726,0.79425645,0.3052308,0.2100513,0.24615386,0.21989745,0.0,0.0,0.0,0.0,0.0,0.0,0.036102567,0.036102567,0.01969231,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.016410258,0.016410258,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.006564103,0.0,0.0,0.0,0.013128206,0.006564103,0.0,0.0,0.0,0.0,0.072205134,0.14769232,0.18379489,0.18379489,0.24287182,0.3052308,0.38400003,0.43651286,0.3511795,0.6695385,1.1224617,1.2570257,0.955077,0.44307697,0.3314872,0.2855385,0.28225642,0.27569234,0.21333335,0.128,0.23630771,0.4135385,0.57764107,0.6859488,0.77128214,0.69251287,0.56451285,0.51856416,0.702359,0.761436,0.6695385,0.55794877,0.5021539,0.5021539,0.2231795,0.098461546,0.06235898,0.052512825,0.016410258,0.016410258,0.02297436,0.01969231,0.0,0.0,0.0,0.009846155,0.02297436,0.029538464,0.029538464,0.006564103,0.0,0.006564103,0.02297436,0.04594872,0.04594872,0.06564103,0.0951795,0.13784617,0.19692309,0.2100513,0.23958977,0.30851284,0.4135385,0.5481026,0.7450257,0.9944616,1.1782565,1.273436,1.3587693,1.847795,2.2711797,2.5435898,2.6289232,2.5173335,2.6518977,2.5665643,2.5304618,2.612513,2.6847181,2.6617439,2.8192823,3.0391798,3.2820516,3.6004105,3.882667,4.089436,4.0467696,3.6168208,2.7011285,2.6026669,3.1015387,3.2361028,2.806154,2.3794873,2.356513,2.4681027,2.1956925,1.4966155,0.82379496,0.5546667,0.44307697,0.380718,0.318359,0.24287182,0.34133336,0.5940513,0.8205129,0.8960001,0.761436,0.702359,0.8960001,1.079795,1.1520001,1.1749744,0.9321026,0.57764107,0.28225642,0.12143591,0.06235898,0.13456412,0.2986667,0.4266667,0.43323082,0.27569234,0.20020515,0.24615386,0.45620516,0.7187693,0.79425645,0.7581539,0.56451285,0.86974365,1.847795,3.190154,2.0644104,1.0994873,0.8172308,1.1520001,1.4342566,1.4703591,1.2603078,1.2603078,1.7591796,2.868513,3.1737437,4.4767184,6.0258465,6.7085133,5.034667,3.8038976,4.2994876,5.044513,5.041231,3.7842054,2.7963078,2.3926156,2.5698464,3.6069746,6.0717955,6.1472826,6.4590774,7.0859494,8.185436,9.980719,9.869129,9.045334,9.478565,11.369026,13.154463,15.156514,18.530462,21.385847,23.079386,24.214975,20.919796,20.644104,22.18995,24.730259,27.831797,27.257439,25.32759,22.649437,20.614565,21.408823,17.769028,13.400617,9.632821,7.1023593,5.720616,4.342154,3.4034874,3.5807183,5.142975,7.9491286,9.412924,8.352821,6.7117953,5.5007186,4.7917953,4.450462,4.345436,4.516103,4.7950773,4.8049235,5.159385,5.3398976,5.2545643,4.9296412,4.4996924,1.7591796,2.930872,3.5807183,3.1277952,2.041436,1.8313848,1.6804104,1.5885129,1.6278975,1.8806155,2.428718,3.0358977,2.8717952,2.7109745,2.993231,3.8104618,5.0477953,5.907693,5.924103,5.290667,4.84759,3.511795,2.858667,2.5238976,2.2678976,1.9823592,1.8346668,2.0086155,2.1431797,2.0611284,1.7558975,1.4375386,1.1355898,0.85005134,0.67938465,0.8369231,0.508718,0.318359,0.21661541,0.16082053,0.118153855,0.14441027,0.19692309,0.21333335,0.18379489,0.12471796,0.068923086,0.03938462,0.036102567,0.03938462,0.013128206,0.052512825,0.04266667,0.02297436,0.013128206,0.013128206,0.013128206,0.01969231,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.006564103,0.006564103,0.006564103,0.0032820515,0.0032820515,0.0032820515,0.0,0.0,0.0032820515,0.013128206,0.02297436,0.01969231,0.013128206,0.009846155,0.006564103,0.0032820515,0.0,0.009846155,0.006564103,0.0032820515,0.006564103,0.02297436,0.049230773,0.09189744,0.13784617,0.2297436,0.4660513,0.256,0.15097436,0.15425642,0.21333335,0.23302566,0.049230773,0.013128206,0.016410258,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.06235898,0.08205129,0.049230773,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.02297436,0.013128206,0.032820515,0.055794876,0.049230773,0.029538464,0.052512825,0.009846155,0.009846155,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01969231,0.03938462,0.0,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.013128206,0.01969231,0.04594872,0.06564103,0.052512825,0.032820515,0.026256412,0.036102567,0.04594872,0.06235898,0.19364104,0.380718,0.3708718,0.24943592,0.20020515,0.2855385,0.4594872,0.571077,0.318359,0.36758977,0.51856416,0.60389745,0.48902568,0.23958977,0.2100513,0.380718,0.6695385,0.9353847,1.529436,2.0053334,2.228513,2.4549747,3.3214362,2.989949,3.2525132,4.4898467,6.2227697,7.1187696,5.3858466,4.6867695,4.076308,3.515077,3.8596926,3.8367183,3.570872,3.314872,3.121231,2.8356924,3.8367183,4.2338467,3.9712822,3.308308,2.8356924,3.259077,3.6726158,4.3290257,5.431795,7.1483083,9.153642,10.614155,11.0145645,9.800206,6.373744,8.123077,9.452309,9.478565,8.054154,5.792821,4.460308,3.3411283,3.0884104,3.7743592,4.8607183,3.9614363,3.2131286,3.6758976,5.139693,6.1341543,7.4896417,7.532308,7.3485136,7.1548724,6.2851286,4.788513,4.634257,4.2436924,3.2754874,2.6518977,1.9528207,1.339077,0.9189744,0.7122052,0.63343596,0.61374366,0.4397949,0.29538465,0.23958977,0.19692309,0.068923086,0.02297436,0.052512825,0.118153855,0.15753847,0.118153855,0.04594872,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.02297436,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0,0.0,0.0,0.0,0.0032820515,0.0,0.0032820515,0.013128206,0.013128206,0.013128206,0.04266667,0.06564103,0.08861539,0.14769232,0.19692309,0.27897438,0.36758977,0.4135385,0.33805132,1.0568206,1.1585642,0.90584624,0.53825647,0.25928208,0.23630771,0.2855385,0.3446154,0.36102566,0.2986667,0.19364104,0.20676924,0.34133336,0.52512825,0.6268718,0.7515898,0.6235898,0.508718,0.571077,0.8598975,1.086359,0.8960001,0.5940513,0.41025645,0.47917953,0.36430773,0.20676924,0.118153855,0.098461546,0.052512825,0.04266667,0.055794876,0.059076928,0.04266667,0.013128206,0.013128206,0.006564103,0.0032820515,0.016410258,0.055794876,0.059076928,0.032820515,0.009846155,0.0032820515,0.009846155,0.03938462,0.049230773,0.049230773,0.06235898,0.11158975,0.2231795,0.31507695,0.40697438,0.508718,0.63343596,0.9189744,1.2406155,1.522872,1.782154,2.1530259,2.678154,3.0260515,3.1474874,3.114667,3.0916924,3.3050258,2.9538465,2.4746668,2.169436,2.172718,2.3236926,2.540308,2.7700515,3.006359,3.2951798,3.6660516,3.9384618,4.0992823,4.125539,3.9811285,3.945026,4.0533338,3.56759,2.5698464,1.9659488,1.8740515,1.9035898,1.8149745,1.5097437,1.0436924,0.7056411,0.6071795,0.57764107,0.51856416,0.37743592,0.318359,0.47589746,0.6629744,0.75487185,0.6892308,0.5907693,0.65641034,0.8369231,0.9911796,0.9189744,0.8205129,0.6432821,0.45620516,0.30194873,0.18379489,0.21661541,0.48246157,0.702359,0.8008206,0.8960001,0.6465641,0.42338464,0.512,0.9485129,1.4998976,0.95835906,0.6662565,1.5622566,3.6857438,6.193231,5.917539,2.8849232,0.8730257,0.88943595,1.1913847,1.276718,1.0633847,1.1257436,1.7362052,2.8553848,3.7087183,5.2578464,8.093539,11.185231,11.894155,7.5191803,5.654975,4.900103,4.269949,3.1967182,2.3368206,2.537026,3.4494362,4.1091285,2.9243078,3.515077,3.5380516,4.2601027,5.9470773,7.8802056,7.584821,7.680001,7.762052,8.116513,9.724719,11.090053,12.235488,13.820719,16.866463,22.738052,22.675694,20.096,18.428719,19.183592,21.973335,24.22154,25.898668,24.362669,20.919796,20.834463,17.499899,13.078976,9.603283,7.9917955,8.077128,6.23918,4.670359,4.066462,4.637539,6.1078978,8.001641,7.076103,5.989744,5.717334,5.536821,5.3792825,5.1626673,4.896821,4.6244106,4.4045134,4.699898,5.0051284,5.0904617,4.906667,4.588308,2.0873847,2.4352822,2.6289232,2.3335385,1.7394873,1.5753847,1.595077,1.7591796,1.9593848,2.1234872,2.1989746,2.556718,2.8914874,3.3247182,3.6890259,3.5380516,3.1770258,3.3772311,3.764513,4.1878977,4.6966157,3.9318976,3.5938463,3.2984617,2.858667,2.2646155,1.7460514,1.6672822,1.8642052,2.176,2.4516926,2.0939488,1.7001027,1.2996924,0.9714873,0.8598975,0.574359,0.45292312,0.35774362,0.24287182,0.15425642,0.16410258,0.20348719,0.20676924,0.15753847,0.108307704,0.049230773,0.01969231,0.01969231,0.026256412,0.02297436,0.052512825,0.052512825,0.036102567,0.016410258,0.02297436,0.02297436,0.029538464,0.032820515,0.029538464,0.009846155,0.0032820515,0.0,0.0032820515,0.006564103,0.0,0.006564103,0.0032820515,0.0032820515,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.013128206,0.009846155,0.009846155,0.016410258,0.026256412,0.07548718,0.13128206,0.19692309,0.3052308,0.25271797,0.20676924,0.190359,0.190359,0.15425642,0.029538464,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.032820515,0.04266667,0.02297436,0.0,0.006564103,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.01969231,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.02297436,0.016410258,0.006564103,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.006564103,0.03938462,0.059076928,0.049230773,0.01969231,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.01969231,0.0,0.026256412,0.01969231,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.02297436,0.03938462,0.049230773,0.04594872,0.04266667,0.03938462,0.052512825,0.08533334,0.14112821,0.14441027,0.08861539,0.12143591,0.22646156,0.2231795,0.16082053,0.16738462,0.28225642,0.49887183,0.77128214,0.571077,0.5513847,0.61374366,0.6892308,0.7187693,0.7515898,0.6859488,0.7384616,1.0043077,1.4375386,1.8937438,1.9856411,1.8904617,1.9167181,2.5009232,2.4549747,2.9636924,4.007385,5.1659493,5.61559,5.0182567,6.038975,6.685539,6.3573337,5.8453336,5.097026,4.7950773,5.0149746,5.179077,4.0402055,4.1025643,4.3027697,4.381539,4.2436924,3.9318976,3.626667,4.33559,5.228308,5.940513,6.554257,7.1089234,7.755488,9.875693,11.497026,7.282872,7.716103,8.868103,9.468719,8.861539,7.000616,5.4908724,3.9844105,3.501949,4.322462,5.9569235,5.792821,4.378257,3.1113849,2.7995899,3.6594875,4.1025643,4.013949,4.2305646,5.037949,6.170257,6.547693,5.5696416,3.9647183,2.4713848,1.8445129,1.6607181,1.3554872,1.017436,0.8730257,1.3095386,1.1290257,0.6826667,0.3249231,0.17394873,0.108307704,0.108307704,0.07548718,0.068923086,0.101743594,0.13456412,0.0951795,0.032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.016410258,0.02297436,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.0032820515,0.0,0.0032820515,0.009846155,0.01969231,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.009846155,0.009846155,0.0032820515,0.006564103,0.016410258,0.016410258,0.016410258,0.02297436,0.029538464,0.059076928,0.14769232,0.128,0.18051283,0.26256412,0.36430773,0.51856416,0.98461545,0.86974365,0.64000005,0.5284103,0.54482055,0.571077,0.5152821,0.39384618,0.2855385,0.3117949,0.26584616,0.27897438,0.40697438,0.6235898,0.8402052,0.9747693,0.78769237,0.71548724,0.8598975,1.0010257,0.92553854,0.67282057,0.45292312,0.3708718,0.41682056,0.36758977,0.23958977,0.24615386,0.4135385,0.58420515,0.512,0.32164106,0.15425642,0.068923086,0.032820515,0.03938462,0.032820515,0.02297436,0.01969231,0.02297436,0.052512825,0.04266667,0.02297436,0.006564103,0.0,0.02297436,0.049230773,0.049230773,0.04594872,0.108307704,0.2231795,0.3511795,0.51856416,0.6892308,0.764718,0.9682052,1.1913847,1.4112822,1.6771283,2.0939488,2.7273848,3.0260515,3.062154,2.9768207,3.006359,3.1277952,2.8356924,2.412308,2.162872,2.4188719,2.6880002,2.8717952,3.0358977,3.245949,3.5872824,3.9844105,4.312616,4.4865646,4.493129,4.394667,4.2371287,4.0467696,3.5971284,2.9735386,2.5764105,2.3401027,2.169436,1.9790771,1.7001027,1.2898463,0.86317956,0.69251287,0.6465641,0.6104616,0.4955898,0.4266667,0.5546667,0.67938465,0.7122052,0.6629744,0.574359,0.5874872,0.6826667,0.7581539,0.65312827,0.51856416,0.38728207,0.33805132,0.36430773,0.3708718,0.3511795,0.43651286,0.5513847,0.6662565,0.7975385,0.7384616,0.571077,0.571077,0.8730257,1.4408206,1.017436,0.761436,1.7755898,4.1550775,6.987488,7.207385,4.197744,1.6114873,0.827077,0.955077,1.3029745,1.4966155,1.7165129,2.0545642,2.5337439,2.8849232,3.6496413,5.5171285,8.018052,9.527796,7.397744,5.914257,5.1364107,4.713026,3.892513,3.692308,4.535795,5.681231,6.121026,4.598154,4.916513,3.9811285,3.4494362,4.0402055,5.5597954,6.4065647,8.155898,8.789334,8.4283085,9.324308,10.010257,10.463181,11.753027,14.043899,16.57436,17.903591,16.262566,14.539488,14.378668,16.196924,20.762259,26.804514,27.549541,23.102362,20.424206,17.076513,13.321847,10.269539,8.493949,8.044309,6.2752824,5.3431797,5.8256416,7.273026,8.208411,7.7292314,5.85518,4.4438977,4.125539,4.312616,4.598154,4.7228723,4.647385,4.4045134,4.1025643,4.197744,4.460308,4.6966157,4.768821,4.6080003,1.8445129,1.6475899,1.5556924,1.5589745,1.5885129,1.5130258,1.5819489,1.8084104,2.0841026,2.3040001,2.3663592,2.4516926,3.1081028,3.9745643,4.571898,4.263385,3.062154,2.5600002,2.6617439,3.1770258,3.7940516,4.4307694,4.7491283,4.4012313,3.4888208,2.5632823,2.100513,1.9035898,2.0512822,2.487795,3.0227695,2.9210258,2.7241027,2.3269746,1.785436,1.2996924,0.88615394,0.6465641,0.49887183,0.4004103,0.3249231,0.30851284,0.3052308,0.2855385,0.23630771,0.18707694,0.108307704,0.055794876,0.04594872,0.059076928,0.06235898,0.07876924,0.08861539,0.068923086,0.036102567,0.049230773,0.032820515,0.02297436,0.026256412,0.029538464,0.009846155,0.0032820515,0.0032820515,0.013128206,0.01969231,0.006564103,0.009846155,0.0032820515,0.0032820515,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.006564103,0.013128206,0.013128206,0.013128206,0.01969231,0.03938462,0.036102567,0.14769232,0.2297436,0.21661541,0.13456412,0.16738462,0.19692309,0.18707694,0.13456412,0.08205129,0.055794876,0.04594872,0.032820515,0.013128206,0.0,0.0,0.0032820515,0.009846155,0.009846155,0.0,0.0,0.0,0.0,0.0,0.006564103,0.013128206,0.009846155,0.013128206,0.02297436,0.013128206,0.02297436,0.029538464,0.032820515,0.032820515,0.036102567,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.009846155,0.0,0.0,0.0,0.0,0.0,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.02297436,0.016410258,0.006564103,0.0,0.0,0.0032820515,0.02297436,0.02297436,0.009846155,0.029538464,0.052512825,0.04594872,0.026256412,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02297436,0.016410258,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.026256412,0.03938462,0.04266667,0.026256412,0.01969231,0.026256412,0.052512825,0.101743594,0.17066668,0.17723078,0.108307704,0.072205134,0.09189744,0.108307704,0.13128206,0.19692309,0.3117949,0.5415385,1.0108719,0.88287187,0.7450257,0.6826667,0.7450257,0.9288206,1.4900514,1.4736412,1.2898463,1.2438976,1.5031796,1.8248206,1.6114873,1.4309745,1.4900514,1.6410258,1.6804104,2.0512822,2.5337439,2.9111798,2.9833848,3.564308,5.100308,6.157129,6.193231,5.5696416,4.926359,5.2742567,6.229334,6.8562055,5.674667,5.2545643,5.221744,5.1922054,5.0116925,4.7655387,4.2535386,4.7458467,5.2315903,5.333334,5.3103595,5.7140517,5.874872,8.129642,10.79795,8.169026,7.581539,8.077128,9.127385,9.931488,9.416205,7.0892315,4.9821544,4.066462,4.637539,6.311385,7.578257,6.482052,4.391385,2.6289232,2.4615386,2.0873847,2.028308,2.6420515,3.9253337,5.536821,6.3277955,5.07077,3.2525132,1.8313848,1.2340513,1.2307693,1.1651284,1.014154,0.955077,1.3718976,1.0436924,0.63343596,0.318359,0.15097436,0.06564103,0.12471796,0.098461546,0.055794876,0.03938462,0.055794876,0.03938462,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.009846155,0.0,0.0,0.0,0.0032820515,0.006564103,0.0032820515,0.0,0.0032820515,0.0032820515,0.0032820515,0.009846155,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.016410258,0.0032820515,0.0032820515,0.013128206,0.02297436,0.02297436,0.016410258,0.009846155,0.0032820515,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.016410258,0.016410258,0.009846155,0.0032820515,0.0032820515,0.009846155,0.016410258,0.016410258,0.029538464,0.049230773,0.09189744,0.190359,0.21989745,0.27569234,0.3249231,0.42338464,0.6826667,0.8960001,0.8533334,0.827077,0.8598975,0.78769237,0.85005134,0.761436,0.58092314,0.4266667,0.48246157,0.6432821,0.54482055,0.4955898,0.61374366,0.8336411,0.93866676,0.8467693,0.827077,0.90584624,0.85005134,0.5874872,0.38728207,0.32164106,0.37743592,0.4594872,0.40369233,0.33476925,0.41682056,0.64000005,0.81394875,0.67938465,0.40369233,0.20020515,0.13128206,0.0951795,0.068923086,0.04594872,0.026256412,0.016410258,0.006564103,0.04266667,0.049230773,0.036102567,0.01969231,0.013128206,0.02297436,0.06564103,0.07876924,0.08861539,0.19692309,0.25271797,0.35774362,0.51856416,0.6892308,0.77128214,0.8960001,1.0075898,1.1454359,1.3751796,1.8116925,2.5173335,2.8882053,2.9538465,2.8324106,2.7569232,2.7208207,2.5042052,2.2908719,2.284308,2.6880002,3.0293336,3.1671798,3.245949,3.3903592,3.6890259,4.135385,4.571898,4.775385,4.6966157,4.4373336,4.1091285,3.82359,3.6562054,3.4921029,3.0391798,2.5665643,2.1431797,1.8740515,1.7033848,1.4178462,0.9878975,0.7778462,0.761436,0.8205129,0.7450257,0.65312827,0.702359,0.7778462,0.7975385,0.7220513,0.5677949,0.5218462,0.52512825,0.52512825,0.46276927,0.3446154,0.21333335,0.20020515,0.3249231,0.49887183,0.5218462,0.48246157,0.5021539,0.58420515,0.6301539,0.67938465,0.58420515,0.5284103,0.6465641,1.0010257,1.0371283,1.0043077,1.8543591,3.7415388,6.0061545,6.0816417,4.2863593,2.7569232,2.2646155,2.2482052,2.484513,2.6453335,2.92759,3.2984617,3.508513,3.2262566,3.4888208,4.263385,5.3037953,6.1538467,6.3212314,5.874872,5.32677,4.8344617,4.204308,4.1550775,4.9427695,5.76,5.9995904,5.2348723,5.425231,4.919795,4.394667,4.420923,5.4514875,6.5739493,8.306872,9.563898,10.262975,11.329642,12.009027,12.603078,13.298873,13.814155,13.413745,14.539488,14.989129,14.293334,12.895181,12.143591,16.036104,22.846361,25.796925,23.657028,20.755693,18.267899,15.970463,13.5548725,10.965334,8.421744,6.012718,5.474462,6.875898,8.809027,8.392206,8.234667,5.802667,3.623385,2.7864618,2.9636924,3.3411283,3.6627696,3.817026,3.7809234,3.626667,3.5807183,3.7218463,3.9286156,4.1058464,4.1682053,1.5589745,1.6114873,1.6508719,1.7723079,1.8904617,1.7296412,1.6049232,1.6147693,1.6935385,1.8313848,2.1070771,2.1267693,2.5206156,3.1245131,3.7940516,4.388103,4.4077954,4.082872,3.5282054,3.045744,3.114667,4.7360005,5.293949,4.7294364,3.4724104,2.4615386,2.4910772,2.5042052,2.612513,2.8553848,3.1967182,3.5216413,3.6791797,3.4100516,2.7864618,2.2219489,1.5589745,1.0469744,0.73517954,0.60061544,0.5316923,0.50543594,0.49887183,0.50543594,0.48902568,0.4004103,0.25928208,0.15097436,0.108307704,0.108307704,0.098461546,0.1148718,0.12143591,0.098461546,0.068923086,0.07548718,0.04266667,0.02297436,0.016410258,0.016410258,0.016410258,0.009846155,0.013128206,0.01969231,0.02297436,0.013128206,0.0032820515,0.0,0.0,0.0,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.01969231,0.013128206,0.013128206,0.0032820515,0.006564103,0.029538464,0.08205129,0.101743594,0.24287182,0.318359,0.25928208,0.1148718,0.072205134,0.12143591,0.13784617,0.101743594,0.09189744,0.108307704,0.11158975,0.09189744,0.052512825,0.0,0.0,0.009846155,0.02297436,0.029538464,0.013128206,0.009846155,0.0032820515,0.0,0.0032820515,0.013128206,0.016410258,0.026256412,0.052512825,0.07876924,0.068923086,0.08533334,0.09189744,0.09189744,0.09189744,0.08861539,0.02297436,0.0032820515,0.0,0.0,0.0,0.0032820515,0.01969231,0.04266667,0.052512825,0.013128206,0.0032820515,0.0,0.0,0.0032820515,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.049230773,0.052512825,0.026256412,0.06564103,0.06564103,0.026256412,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.013128206,0.006564103,0.0,0.0,0.0,0.006564103,0.02297436,0.049230773,0.09189744,0.13456412,0.14112821,0.13456412,0.14112821,0.16738462,0.23630771,0.3446154,0.446359,0.64000005,1.1355898,1.0666667,0.90584624,0.8205129,0.8763078,1.0371283,2.0053334,2.1956925,1.9462565,1.6016412,1.4998976,1.7558975,1.5064616,1.404718,1.5556924,1.5097437,1.4605129,1.4736412,1.6147693,1.8674873,2.1234872,2.5271797,2.7963078,3.045744,3.318154,3.5741541,3.820308,5.0642056,6.363898,7.017026,6.547693,6.521436,6.567385,5.9963083,4.9952826,4.630975,4.844308,5.1232824,5.1987696,5.139693,5.362872,7.1089234,7.788308,8.592411,9.442462,8.999385,8.36595,8.257642,9.081436,10.384411,10.850462,7.8441033,5.4383593,4.164923,4.2240005,5.504,7.962257,7.837539,6.242462,4.204308,2.6584618,2.5173335,2.8816411,3.6004105,4.378257,4.768821,4.1813335,3.2918978,2.3072822,1.4867693,1.148718,1.014154,0.955077,0.88287187,0.76800007,0.6170257,0.42994875,0.34133336,0.26256412,0.17394873,0.13784617,0.12143591,0.08533334,0.03938462,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.013128206,0.016410258,0.009846155,0.0,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0,0.0,0.0,0.0032820515,0.013128206,0.013128206,0.0032820515,0.006564103,0.01969231,0.026256412,0.016410258,0.013128206,0.013128206,0.006564103,0.0,0.0,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.013128206,0.0032820515,0.0032820515,0.006564103,0.013128206,0.02297436,0.02297436,0.06235898,0.118153855,0.190359,0.27897438,0.41682056,0.47589746,0.49887183,0.5481026,0.71548724,0.8763078,1.0404103,1.1716924,1.1552821,0.79425645,0.90584624,0.9747693,0.9189744,0.7975385,0.80738467,1.1224617,0.9714873,0.761436,0.6695385,0.6268718,0.6695385,0.7187693,0.7318975,0.67938465,0.5349744,0.33476925,0.27569234,0.33805132,0.47589746,0.6235898,0.5677949,0.5415385,0.58092314,0.636718,0.5677949,0.41682056,0.24943592,0.17723078,0.18707694,0.16082053,0.07876924,0.032820515,0.013128206,0.006564103,0.016410258,0.04266667,0.04266667,0.032820515,0.029538464,0.029538464,0.04266667,0.07876924,0.118153855,0.190359,0.3708718,0.36102566,0.380718,0.4266667,0.49887183,0.60389745,0.7056411,0.7778462,0.88287187,1.1257436,1.6443079,2.3466668,2.8258464,2.986667,2.858667,2.605949,2.4976413,2.356513,2.3663592,2.5665643,2.861949,3.0982566,3.1245131,3.1081028,3.1770258,3.4067695,3.9220517,4.450462,4.7360005,4.6867695,4.378257,3.9680004,3.7415388,3.764513,3.748103,3.0129232,2.300718,1.6804104,1.4178462,1.4473847,1.3718976,1.0436924,0.8730257,0.92225647,1.0699488,1.0043077,0.85005134,0.77128214,0.79097444,0.8369231,0.74830776,0.512,0.41025645,0.36758977,0.34789747,0.34789747,0.30851284,0.19692309,0.17394873,0.3052308,0.57764107,0.67282057,0.636718,0.6235898,0.65641034,0.6301539,0.6104616,0.5152821,0.43323082,0.44307697,0.58092314,1.0699488,1.3587693,1.8871796,2.8192823,4.0434875,3.9548721,3.623385,3.7120004,4.141949,4.1222568,3.95159,3.820308,4.4767184,5.7501545,6.564103,6.1374364,6.311385,6.5083084,6.3868723,5.8256416,6.1407185,6.2129235,5.668103,4.6867695,4.027077,3.7382567,3.7940516,3.9680004,4.125539,4.2174363,4.630975,5.5663595,6.3310776,6.7544622,7.200821,7.6767187,8.280616,9.941334,12.396309,14.17518,15.320617,16.636719,16.728617,15.593027,14.592001,14.670771,16.643284,16.90913,14.519796,11.18195,11.559385,15.228719,19.088411,21.490873,22.232616,22.186668,21.556515,19.544617,15.894976,10.889847,7.2237954,6.1472826,7.072821,8.254359,6.7807183,8.349539,6.058667,3.5807183,2.5337439,2.4910772,2.6157951,2.7602053,2.861949,2.9144619,2.9735386,2.8914874,2.878359,2.8980515,2.9833848,3.239385,3.0982566,2.8291285,2.7076926,2.7011285,2.6945643,2.487795,2.3401027,2.3401027,2.2383592,1.9954873,1.8018463,1.7526156,1.8215386,2.0906668,2.605949,3.387077,4.2174363,4.7458467,4.854154,4.6178465,4.2863593,4.325744,3.5741541,3.0129232,2.8291285,2.425436,2.2186668,2.2416413,2.300718,2.3926156,2.6847181,3.1376412,3.370667,3.3378465,3.1507695,3.0523078,2.4648206,1.9790771,1.4572309,0.92225647,0.58092314,0.50543594,0.56123084,0.67610264,0.7417436,0.5940513,0.38728207,0.22646156,0.12143591,0.072205134,0.06235898,0.049230773,0.055794876,0.072205134,0.08861539,0.07548718,0.052512825,0.06564103,0.08205129,0.08861539,0.07548718,0.052512825,0.026256412,0.016410258,0.013128206,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01969231,0.036102567,0.0,0.0,0.0,0.006564103,0.032820515,0.108307704,0.30194873,0.3052308,0.24287182,0.190359,0.15097436,0.128,0.0951795,0.059076928,0.04266667,0.09189744,0.07876924,0.10502565,0.128,0.108307704,0.0,0.0,0.009846155,0.026256412,0.049230773,0.06235898,0.049230773,0.01969231,0.006564103,0.013128206,0.0,0.02297436,0.07548718,0.13128206,0.18051283,0.2297436,0.20348719,0.17066668,0.18379489,0.23630771,0.25928208,0.07548718,0.013128206,0.0,0.0,0.0,0.02297436,0.06564103,0.13456412,0.17066668,0.06235898,0.02297436,0.006564103,0.006564103,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.009846155,0.0,0.0,0.0,0.0,0.006564103,0.01969231,0.029538464,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.01969231,0.029538464,0.190359,0.24615386,0.25271797,0.23958977,0.2297436,0.3249231,0.58092314,0.761436,0.8041026,0.79425645,0.84348726,0.98133343,1.2406155,1.4408206,1.2209232,1.6738462,2.169436,2.487795,2.546872,2.425436,2.1956925,1.8510771,1.394872,0.99774367,1.024,1.1191796,1.2274873,1.591795,2.3072822,3.2951798,2.5271797,2.3335385,2.537026,2.92759,3.2820516,3.3411283,4.31918,4.886975,4.8049235,4.9132314,5.756718,6.560821,5.920821,4.3749747,4.4242053,5.6320004,6.803693,7.5191803,7.6931286,7.584821,9.426052,11.224616,11.976206,11.464206,10.269539,9.255385,8.628513,8.103385,7.506052,6.7610264,5.504,4.46359,3.6594875,3.0720003,2.6715899,4.8672824,5.9569235,5.8486156,4.8311796,3.5872824,3.7185643,4.056616,4.201026,3.9876926,3.4625645,2.865231,2.1956925,1.4933335,0.9517949,0.9156924,0.93866676,0.8467693,0.61374366,0.3117949,0.09189744,0.22646156,0.20348719,0.15097436,0.12471796,0.13784617,0.11158975,0.07876924,0.04266667,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.036102567,0.036102567,0.01969231,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.016410258,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.02297436,0.036102567,0.04594872,0.04594872,0.059076928,0.098461546,0.21333335,0.36430773,0.4135385,0.42338464,0.3708718,0.41025645,0.5316923,0.58092314,0.65312827,0.7089231,0.7318975,0.7187693,0.67282057,0.892718,1.2570257,1.2996924,1.0535386,1.0535386,1.017436,1.3915899,1.6180514,1.4080001,0.74830776,0.7220513,0.6071795,0.5513847,0.58420515,0.5940513,0.38728207,0.4266667,0.5874872,0.7450257,0.79425645,0.86646163,0.8205129,0.67282057,0.46933338,0.27569234,0.20020515,0.16410258,0.14112821,0.12471796,0.13784617,0.06564103,0.026256412,0.02297436,0.026256412,0.016410258,0.0032820515,0.0,0.006564103,0.01969231,0.029538464,0.04266667,0.06564103,0.16082053,0.36102566,0.64000005,0.5907693,0.50543594,0.4135385,0.34789747,0.33476925,0.41025645,0.49887183,0.6662565,0.99774367,1.6311796,2.2547693,2.6486156,2.8192823,2.789744,2.5928206,2.678154,2.9111798,3.1803079,3.387077,3.4494362,3.117949,2.789744,2.612513,2.6978464,3.1113849,3.636513,4.07959,4.33559,4.378257,4.2568207,4.013949,3.761231,3.6430771,3.5249233,2.9768207,2.2547693,1.6443079,1.2603078,1.1290257,1.1913847,1.0075898,0.92553854,0.9321026,0.955077,0.86974365,0.73517954,0.574359,0.46933338,0.44307697,0.44307697,0.39384618,0.33476925,0.29210258,0.26256412,0.21333335,0.1148718,0.101743594,0.24615386,0.5152821,0.74830776,0.69907695,0.5940513,0.5284103,0.5316923,0.58092314,0.5907693,0.5677949,0.48902568,0.43323082,0.58092314,1.1290257,1.5885129,1.6902566,1.6738462,2.2744617,3.4822567,3.9023592,3.5807183,3.0129232,3.1573336,3.0358977,3.5544617,5.8814363,9.383386,11.641437,11.897437,11.349334,10.633847,9.829744,8.438154,7.6701546,7.4863596,6.9743595,5.920821,4.821334,5.175795,4.6244106,4.348718,4.900103,6.196513,6.6592827,7.2336416,7.972103,8.434873,7.6898465,8.65477,10.505847,12.612924,14.395078,15.333745,16.324924,19.11795,20.489847,19.026052,15.107284,14.555899,16.131283,17.046976,16.246155,14.404924,11.218052,11.556104,13.840411,17.923283,25.10113,29.32513,29.298874,26.49272,21.891283,16.006565,11.881026,9.45559,8.103385,7.8670774,9.4916935,6.11118,3.7809234,2.858667,2.9801028,3.0523078,3.186872,2.9440002,2.6453335,2.4582565,2.412308,2.300718,2.1267693,1.9790771,1.9561027,2.1530259,1.7066668,1.9265642,1.9626669,1.8937438,1.9003079,2.281026,2.806154,3.1442053,3.3345644,3.2000003,2.349949,2.4188719,2.5895386,2.858667,3.259077,3.876103,4.3749747,4.519385,4.604718,4.6802053,4.5554876,4.1156926,3.7185643,3.3542566,2.9407182,2.353231,1.9298463,1.8248206,1.9265642,2.038154,1.8937438,2.3729234,2.7798977,3.0884104,3.249231,3.2098465,2.6551797,2.4746668,2.1891284,1.6869745,1.2406155,1.0305642,0.9189744,0.86317956,0.8467693,0.8763078,0.7844103,0.6235898,0.45620516,0.3314872,0.28225642,0.14112821,0.07876924,0.06235898,0.072205134,0.08861539,0.101743594,0.0951795,0.1148718,0.15097436,0.15097436,0.08533334,0.04594872,0.02297436,0.013128206,0.0,0.0,0.0,0.0032820515,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0,0.0,0.0032820515,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.0032820515,0.0032820515,0.006564103,0.0,0.0,0.0,0.0,0.01969231,0.08205129,0.24943592,0.25271797,0.21989745,0.21989745,0.26256412,0.27569234,0.2231795,0.118153855,0.055794876,0.20020515,0.101743594,0.04594872,0.026256412,0.026256412,0.02297436,0.06235898,0.03938462,0.013128206,0.016410258,0.049230773,0.055794876,0.052512825,0.07548718,0.12471796,0.17066668,0.18707694,0.256,0.3314872,0.33476925,0.16738462,0.19364104,0.18707694,0.18707694,0.23630771,0.35774362,0.39712822,0.20020515,0.06235898,0.068923086,0.098461546,0.101743594,0.11158975,0.14769232,0.17723078,0.098461546,0.032820515,0.01969231,0.03938462,0.06235898,0.049230773,0.009846155,0.006564103,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.18707694,0.7975385,2.2121027,2.0545642,0.8533334,0.04594872,0.0,0.0,0.0,0.0,0.01969231,0.059076928,0.09189744,0.01969231,0.108307704,0.13784617,0.06235898,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01969231,0.052512825,0.08861539,0.10502565,0.06564103,0.108307704,0.13128206,0.15097436,0.18379489,0.23958977,0.28882053,0.60389745,0.8992821,1.0633847,1.148718,1.1946667,1.3292309,1.723077,2.4057438,3.2722054,3.1277952,2.6190772,2.0184617,1.6049232,1.6705642,2.8717952,2.6847181,2.1398976,1.785436,1.6804104,1.8281027,2.100513,2.1792822,2.1333334,2.428718,2.0709746,1.7985642,1.7001027,1.8215386,2.1464617,2.1858463,2.6322052,3.0490258,3.3903592,3.9975388,5.622154,6.51159,7.683283,8.592411,7.1483083,6.2752824,7.000616,8.320001,9.235693,8.756514,10.473026,10.866873,10.266257,9.206155,8.438154,9.475283,9.058462,8.27077,7.5913854,6.9054365,5.805949,4.309334,3.058872,2.481231,2.793026,4.2568207,4.7327185,4.210872,3.1507695,2.4615386,2.6847181,3.1442053,3.4330258,3.3017437,2.6584618,1.8051283,1.394872,1.3981539,1.4834872,0.9878975,0.61374366,0.40369233,0.2297436,0.07876924,0.055794876,0.08205129,0.09189744,0.08533334,0.06564103,0.03938462,0.09189744,0.055794876,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.006564103,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.013128206,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.01969231,0.01969231,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.013128206,0.013128206,0.016410258,0.029538464,0.055794876,0.0951795,0.15425642,0.16410258,0.190359,0.25928208,0.3249231,0.35774362,0.38400003,0.42994875,0.46933338,0.4201026,0.50543594,0.58420515,0.61374366,0.65641034,0.892718,0.9944616,1.0436924,1.0043077,0.92225647,0.9321026,0.9321026,1.0338463,1.142154,1.1454359,0.90584624,0.7253334,0.61374366,0.5940513,0.6071795,0.5218462,0.47917953,0.63343596,0.8336411,0.9485129,0.8795898,0.88287187,0.65969235,0.42994875,0.29538465,0.22646156,0.23958977,0.32164106,0.3511795,0.32164106,0.3314872,0.21989745,0.101743594,0.029538464,0.016410258,0.016410258,0.013128206,0.01969231,0.04594872,0.07548718,0.07876924,0.04266667,0.036102567,0.06235898,0.1148718,0.20020515,0.2100513,0.21333335,0.2231795,0.23630771,0.21333335,0.3249231,0.43323082,0.5415385,0.6662565,0.85005134,1.0436924,1.6443079,2.2416413,2.7273848,3.3017437,3.748103,3.879385,4.023795,4.1780515,4.0336413,3.4691284,3.1048207,3.0096412,3.1934361,3.5872824,4.1813335,4.466872,4.391385,4.0467696,3.6726158,3.4756925,3.2656412,2.7241027,1.9659488,1.5360001,1.7033848,1.9889232,2.0053334,1.7132308,1.4211283,1.2865642,1.1881026,1.0535386,0.86646163,0.67282057,0.65641034,0.65641034,0.636718,0.6071795,0.636718,0.6071795,0.5349744,0.4266667,0.3052308,0.17723078,0.108307704,0.108307704,0.24615386,0.5316923,0.9321026,0.86317956,0.7318975,0.64000005,0.6071795,0.5677949,0.6104616,0.6859488,0.67610264,0.6268718,0.761436,1.3915899,1.6902566,1.6836925,1.719795,2.4943593,4.6867695,4.601436,3.6332312,2.7766156,2.6223593,2.5665643,3.373949,5.3694363,8.083693,10.262975,11.398565,11.648001,11.021129,9.616411,7.6077952,7.4043083,8.756514,9.869129,9.964309,9.265231,9.130668,8.769642,8.04759,7.2861543,7.282872,7.5585647,7.1483083,7.0104623,7.250052,7.141744,7.6077952,9.357129,12.025436,14.936617,17.115898,19.02277,19.498669,18.625643,16.538258,13.420309,12.071385,12.596514,14.043899,15.0088215,13.6237955,12.790154,12.882052,13.279181,14.385232,17.618053,23.620924,24.31672,22.626463,20.404514,18.448412,15.386257,14.080001,13.348104,11.943385,8.539898,4.706462,3.1540515,2.793026,2.8849232,3.0260515,3.1507695,3.0752823,2.92759,2.7864618,2.678154,2.550154,2.3926156,2.1891284,1.9987694,1.9692309,2.2186668,2.553436,2.8849232,3.1934361,3.3017437,2.8947694,3.1967182,3.5249233,3.7054362,3.5347695,2.7700515,2.5009232,2.6518977,2.8455386,3.0326157,3.501949,3.7940516,3.570872,3.1409233,2.92759,3.4592824,3.4789746,3.564308,3.6496413,3.6562054,3.5052311,2.789744,2.2055387,1.8740515,1.7493335,1.6377437,1.9003079,2.156308,2.6026669,3.0949745,3.1573336,3.0720003,3.190154,3.1606157,2.865231,2.412308,1.8149745,1.4211283,1.214359,1.1618463,1.211077,1.017436,0.7975385,0.61374366,0.48574364,0.3708718,0.2100513,0.108307704,0.068923086,0.08205129,0.13784617,0.14769232,0.14769232,0.15753847,0.17066668,0.14112821,0.08205129,0.055794876,0.04266667,0.029538464,0.009846155,0.0032820515,0.0,0.006564103,0.013128206,0.0,0.006564103,0.009846155,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.032820515,0.029538464,0.009846155,0.0,0.0,0.0,0.0,0.055794876,0.14441027,0.17723078,0.190359,0.2100513,0.23630771,0.27241027,0.318359,0.23302566,0.13456412,0.055794876,0.036102567,0.118153855,0.16410258,0.16410258,0.12143591,0.06235898,0.013128206,0.032820515,0.01969231,0.0032820515,0.0032820515,0.01969231,0.02297436,0.02297436,0.036102567,0.068923086,0.12143591,0.25271797,0.53825647,0.76800007,0.7844103,0.49230772,0.79097444,0.8369231,0.9124103,1.0043077,0.7844103,0.3314872,0.10502565,0.029538464,0.04266667,0.0951795,0.08861539,0.08533334,0.101743594,0.108307704,0.04266667,0.013128206,0.009846155,0.01969231,0.029538464,0.032820515,0.006564103,0.0032820515,0.02297436,0.04266667,0.036102567,0.02297436,0.02297436,0.036102567,0.03938462,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.02297436,0.026256412,0.01969231,0.0032820515,0.009846155,0.10502565,0.4135385,1.1126155,1.0436924,0.44307697,0.049230773,0.029538464,0.0,0.0,0.055794876,0.118153855,0.14769232,0.08861539,0.016410258,0.06564103,0.09189744,0.055794876,0.02297436,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.01969231,0.029538464,0.055794876,0.08205129,0.08533334,0.059076928,0.068923086,0.08205129,0.11158975,0.16410258,0.25271797,0.37743592,0.73517954,1.0043077,1.1126155,1.2373334,1.6443079,2.3204105,2.930872,3.2754874,3.2886157,3.0391798,2.8291285,2.6551797,2.5600002,2.6256413,2.6847181,2.1333334,1.5622566,1.2537436,1.1782565,1.2406155,1.2800001,1.3784616,1.5753847,1.8642052,1.8806155,1.8248206,1.8182565,1.8904617,1.9889232,1.975795,2.1267693,2.3433847,2.6322052,3.1015387,4.568616,4.2568207,4.384821,5.277539,5.356308,5.605744,6.49518,6.7971287,6.7282057,7.9786673,10.561642,11.795693,11.572514,9.974154,7.256616,8.192,8.165744,7.6635904,7.0104623,6.3376417,5.914257,4.4767184,2.9440002,1.9790771,1.9889232,2.5993848,2.6880002,2.4418464,1.9889232,1.4309745,1.6082052,1.913436,2.1267693,2.1530259,2.0184617,1.7165129,1.276718,1.0371283,0.9944616,0.7778462,0.6235898,0.318359,0.09189744,0.02297436,0.04594872,0.03938462,0.03938462,0.03938462,0.036102567,0.006564103,0.036102567,0.01969231,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.006564103,0.009846155,0.009846155,0.0032820515,0.0,0.0032820515,0.009846155,0.01969231,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.009846155,0.009846155,0.009846155,0.006564103,0.0,0.0032820515,0.009846155,0.009846155,0.006564103,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.006564103,0.013128206,0.026256412,0.04266667,0.098461546,0.27241027,0.46933338,0.45620516,0.318359,0.18379489,0.21333335,0.49230772,0.6465641,0.6268718,0.5513847,0.7187693,0.61374366,0.72861546,0.9616411,1.2438976,1.5491283,1.463795,1.4605129,1.3620514,1.1782565,1.1093334,1.1946667,1.2898463,1.3095386,1.2406155,1.1290257,0.9747693,0.8336411,0.7056411,0.60389745,0.5218462,0.77128214,0.9616411,1.0732309,1.0568206,0.827077,0.60389745,0.46276927,0.34789747,0.3249231,0.5874872,0.58092314,0.508718,0.42994875,0.36102566,0.30851284,0.19364104,0.13784617,0.108307704,0.07876924,0.032820515,0.055794876,0.08205129,0.098461546,0.098461546,0.08205129,0.049230773,0.032820515,0.03938462,0.06235898,0.09189744,0.13128206,0.15753847,0.190359,0.23302566,0.27569234,0.36758977,0.48246157,0.5874872,0.64000005,0.6104616,0.5349744,0.85005134,1.3161026,1.913436,2.865231,3.4166157,3.5511796,3.5610259,3.5774362,3.5577438,3.4560003,3.3969233,3.4297438,3.6036925,3.9647183,4.6539493,4.9854364,4.8640003,4.388103,3.8465643,3.508513,3.1573336,2.4385643,1.5195899,1.1027694,2.0184617,2.6715899,2.7109745,2.169436,1.4539489,1.2570257,1.142154,0.98133343,0.76800007,0.5973334,0.6629744,0.80738467,0.8730257,0.80738467,0.6695385,0.571077,0.53825647,0.5349744,0.48902568,0.3052308,0.17723078,0.13784617,0.20348719,0.380718,0.67610264,0.7778462,0.74830776,0.67610264,0.5973334,0.49230772,0.48902568,0.55794877,0.6104616,0.74830776,1.2570257,1.8313848,2.1464617,2.3729234,2.8225644,3.9384618,5.7009234,4.827898,3.6102567,3.1507695,3.3575387,3.2918978,3.436308,4.066462,5.097026,6.091488,7.680001,8.736821,8.507077,7.0826674,5.4153852,5.7107697,7.282872,8.950154,9.990565,10.148104,9.120821,8.953437,8.553026,7.6077952,6.5837955,6.170257,6.0160003,6.1472826,6.5903597,7.3714876,7.5520005,8.763078,11.0375395,14.053744,17.115898,22.22277,23.27631,21.280823,17.391592,12.937847,11.700514,15.268104,17.988924,17.217642,13.289026,12.225642,12.458668,12.176412,11.713642,13.541744,19.511797,21.044514,20.115694,18.386053,17.217642,16.643284,13.840411,11.648001,10.269539,7.276308,4.342154,3.2886157,3.0260515,2.937436,2.8849232,2.6912823,2.5304618,2.4648206,2.5009232,2.5993848,2.5698464,2.484513,2.3302567,2.1464617,2.03159,2.8291285,3.0523078,3.7021542,4.397949,4.6834874,4.0434875,4.076308,4.397949,4.4406157,3.9811285,3.1507695,2.802872,3.0687182,3.4034874,3.5938463,3.7710772,3.69559,3.1638978,2.428718,1.9364104,2.3138463,2.3302567,2.5238976,2.8127182,3.1442053,3.501949,3.2820516,2.9210258,2.550154,2.2088206,1.8707694,1.7657437,1.7952822,2.1300514,2.6420515,2.9144619,3.3772311,3.7087183,3.8596926,3.7842054,3.4494362,2.6617439,2.097231,1.7165129,1.4834872,1.3686155,1.142154,0.9321026,0.72861546,0.5513847,0.4397949,0.30851284,0.21333335,0.16082053,0.15097436,0.15425642,0.14441027,0.14769232,0.16082053,0.16738462,0.128,0.07548718,0.068923086,0.06564103,0.04594872,0.02297436,0.009846155,0.009846155,0.013128206,0.013128206,0.013128206,0.009846155,0.009846155,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.029538464,0.026256412,0.009846155,0.0,0.0,0.02297436,0.10502565,0.20020515,0.27241027,0.26912823,0.2231795,0.23302566,0.23958977,0.24615386,0.3117949,0.19692309,0.108307704,0.08205129,0.11158975,0.15097436,0.15097436,0.15753847,0.13784617,0.08533334,0.01969231,0.04266667,0.14769232,0.27569234,0.32820517,0.14769232,0.049230773,0.016410258,0.016410258,0.029538464,0.04266667,0.17723078,0.43651286,0.6268718,0.636718,0.43651286,0.7220513,0.77128214,0.8960001,1.0272821,0.7122052,0.15753847,0.006564103,0.0,0.009846155,0.04594872,0.04266667,0.04266667,0.04266667,0.036102567,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.0032820515,0.0,0.02297436,0.055794876,0.04266667,0.029538464,0.032820515,0.04594872,0.04266667,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.0,0.009846155,0.02297436,0.032820515,0.029538464,0.006564103,0.006564103,0.013128206,0.016410258,0.009846155,0.016410258,0.01969231,0.026256412,0.032820515,0.02297436,0.013128206,0.07548718,0.13784617,0.15425642,0.07548718,0.01969231,0.01969231,0.032820515,0.03938462,0.04266667,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0032820515,0.009846155,0.01969231,0.049230773,0.0951795,0.13784617,0.17066668,0.18707694,0.20348719,0.23630771,0.2986667,0.39384618,0.49230772,0.69907695,1.0404103,1.2964103,1.4539489,1.7001027,2.3236926,3.0260515,3.7907696,4.309334,3.9975388,3.7349746,3.6726158,3.515077,3.1967182,2.9046156,2.0841026,1.3456411,0.8467693,0.69579494,0.9517949,0.9714873,0.88943595,0.9616411,1.2865642,1.7985642,2.422154,2.428718,2.2580514,2.1858463,2.3072822,2.356513,2.3729234,2.3827693,2.4648206,2.733949,3.6168208,3.1540515,2.6387694,2.6190772,2.8717952,4.1813335,5.0510774,4.7261543,4.2436924,6.452513,9.921641,12.678565,12.872206,10.361437,6.695385,6.5772314,6.518154,6.232616,5.654975,4.9526157,5.1922054,4.46359,3.2623591,2.1169233,1.5819489,1.7788719,1.972513,2.034872,1.8445129,1.2800001,1.1454359,1.0929232,1.1191796,1.2996924,1.7985642,1.6968206,1.1618463,0.67938465,0.48574364,0.58420515,0.5218462,0.26256412,0.072205134,0.036102567,0.04594872,0.04266667,0.036102567,0.029538464,0.01969231,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.013128206,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.0,0.0,0.0032820515,0.009846155,0.009846155,0.0032820515,0.0,0.0032820515,0.009846155,0.01969231,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.006564103,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.016410258,0.013128206,0.009846155,0.006564103,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.013128206,0.02297436,0.04266667,0.06235898,0.12471796,0.30851284,0.45620516,0.43323082,0.30194873,0.18707694,0.24287182,0.8205129,1.086359,1.0994873,1.0502565,1.2635899,1.142154,1.1618463,1.4506668,1.913436,2.228513,1.9922053,1.8313848,1.5589745,1.2537436,1.2406155,1.339077,1.4506668,1.4309745,1.2931283,1.1946667,1.1093334,1.0404103,0.90912825,0.7581539,0.7417436,1.024,1.1585642,1.142154,1.0010257,0.7975385,0.47917953,0.36758977,0.30194873,0.318359,0.6268718,0.571077,0.446359,0.34133336,0.2855385,0.23958977,0.20020515,0.2100513,0.18379489,0.118153855,0.08861539,0.13128206,0.12471796,0.098461546,0.07548718,0.07548718,0.06235898,0.049230773,0.049230773,0.06564103,0.08533334,0.108307704,0.13456412,0.16082053,0.20020515,0.2855385,0.38400003,0.4955898,0.574359,0.58420515,0.49887183,0.34789747,0.39712822,0.64000005,1.1158975,1.9331284,2.3040001,2.5206156,2.6978464,2.9407182,3.3509746,3.751385,3.9680004,4.066462,4.1517954,4.3684106,4.8377438,5.0543594,4.850872,4.3290257,3.8498464,3.515077,3.170462,2.609231,1.9331284,1.5589745,2.5206156,3.1606157,3.1409233,2.5074873,1.6902566,1.4211283,1.2832822,1.1290257,0.9288206,0.7811283,0.83035904,0.94523084,0.92225647,0.7318975,0.5284103,0.36758977,0.36430773,0.43651286,0.48246157,0.3708718,0.27897438,0.2231795,0.23630771,0.33805132,0.5284103,0.72861546,0.7844103,0.72861546,0.60061544,0.44307697,0.4004103,0.48574364,0.6662565,0.94523084,1.3620514,1.8773335,2.7470772,3.7382567,4.6539493,5.362872,6.373744,5.3169236,4.31918,4.197744,4.457026,4.1714873,3.9680004,3.7316926,3.4658465,3.2886157,4.2305646,5.293949,5.549949,4.8705645,3.9122055,4.082872,4.8836927,5.937231,6.8430777,7.1680007,6.49518,6.875898,7.1089234,6.678975,5.7764106,5.35959,5.4482055,5.5105643,5.7403083,7.026872,7.9852314,9.222565,10.939077,13.285745,16.351181,22.452515,24.95672,24.264208,21.103592,16.52513,14.181745,17.604925,19.925335,18.113642,13.010053,11.040821,10.610872,10.059488,9.708308,11.874462,16.646564,18.773335,18.661745,17.286566,16.17395,16.370872,13.4400015,10.515693,8.5891285,6.518154,4.5390773,3.6069746,3.1934361,2.9472823,2.6880002,2.2711797,2.0020514,1.9265642,1.9987694,2.0873847,2.0611284,2.15959,2.2711797,2.3204105,2.2711797,3.3411283,3.442872,4.325744,5.225026,5.684513,5.58277,5.733744,6.196513,6.163693,5.366154,4.0467696,3.6463592,3.9056413,4.3585644,4.634257,4.44718,4.1091285,3.7054362,3.2525132,2.7766156,2.3204105,1.6836925,1.4605129,1.4900514,1.7066668,2.1530259,2.8455386,3.3017437,3.3805132,3.05559,2.3991797,2.0841026,1.8871796,1.8379488,1.9823592,2.3860514,3.1934361,3.6824617,4.020513,4.20759,4.089436,3.4888208,2.9243078,2.353231,1.8116925,1.4112822,1.211077,1.0568206,0.8467693,0.6268718,0.56451285,0.5021539,0.45620516,0.41682056,0.36758977,0.28225642,0.24615386,0.190359,0.15753847,0.14769232,0.13456412,0.0951795,0.098461546,0.09189744,0.055794876,0.026256412,0.01969231,0.026256412,0.029538464,0.02297436,0.032820515,0.009846155,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0,0.0,0.0,0.0,0.06564103,0.25928208,0.37743592,0.37415388,0.33476925,0.318359,0.27897438,0.21661541,0.18707694,0.3052308,0.24615386,0.19364104,0.18707694,0.23302566,0.29210258,0.108307704,0.052512825,0.052512825,0.06235898,0.036102567,0.08533334,0.29538465,0.5546667,0.7089231,0.56451285,0.5874872,0.5874872,0.512,0.33805132,0.07876924,0.10502565,0.14112821,0.18707694,0.23630771,0.27569234,0.21661541,0.16410258,0.27569234,0.4397949,0.28225642,0.11158975,0.09189744,0.12143591,0.13128206,0.06564103,0.03938462,0.02297436,0.016410258,0.026256412,0.052512825,0.04266667,0.03938462,0.032820515,0.026256412,0.02297436,0.02297436,0.026256412,0.026256412,0.02297436,0.013128206,0.013128206,0.01969231,0.01969231,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.0032820515,0.0,0.0032820515,0.013128206,0.02297436,0.0032820515,0.0,0.0,0.0032820515,0.0,0.0,0.0,0.0,0.009846155,0.049230773,0.032820515,0.04594872,0.068923086,0.08205129,0.06564103,0.052512825,0.059076928,0.06235898,0.06235898,0.072205134,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.01969231,0.052512825,0.032820515,0.013128206,0.013128206,0.036102567,0.12471796,0.2231795,0.318359,0.39056414,0.42994875,0.46276927,0.53825647,0.6629744,0.8041026,0.9124103,1.1618463,1.467077,1.785436,2.1202054,2.5140514,3.0391798,3.1573336,3.764513,4.7491283,4.9887185,4.7261543,4.4832826,3.9417439,3.1048207,2.297436,1.6738462,1.1749744,0.96492314,1.1651284,1.8510771,1.7099489,1.7165129,1.8576412,2.2383592,3.0982566,4.0533338,4.082872,3.826872,3.7120004,3.9680004,4.059898,4.2141542,4.4045134,4.5029745,4.266667,4.4110775,4.850872,4.8738465,4.1780515,2.868513,3.9253337,4.201026,3.882667,3.751385,5.1922054,8.530052,11.930258,11.88759,8.539898,5.677949,4.6572313,4.2863593,4.07959,3.7809234,3.3608208,4.0303593,4.210872,3.7087183,2.7536411,1.9922053,2.1956925,2.6584618,2.7798977,2.422154,1.9364104,1.4966155,1.0962052,0.86974365,1.0010257,1.7263591,1.3686155,0.8566154,0.45292312,0.3052308,0.4266667,0.23302566,0.13456412,0.08205129,0.055794876,0.052512825,0.052512825,0.052512825,0.036102567,0.013128206,0.013128206,0.0032820515,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01969231,0.02297436,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.006564103,0.026256412,0.032820515,0.01969231,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.013128206,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0032820515,0.0032820515,0.009846155,0.01969231,0.026256412,0.04266667,0.055794876,0.1148718,0.20348719,0.26584616,0.19692309,0.16738462,0.21661541,0.3511795,0.54482055,1.2931283,1.6278975,1.782154,1.847795,1.7690258,1.7788719,1.6377437,1.7263591,2.0611284,2.300718,2.0775387,1.7755898,1.3981539,1.1060513,1.2274873,1.2865642,1.332513,1.3128207,1.2471796,1.2274873,1.1913847,1.2242053,1.142154,0.98133343,0.97805136,1.086359,1.1552821,1.0896411,0.94523084,0.9156924,0.6235898,0.40369233,0.26912823,0.2297436,0.28225642,0.23630771,0.21661541,0.2297436,0.27241027,0.3314872,0.3708718,0.35774362,0.24615386,0.11158975,0.13128206,0.18379489,0.118153855,0.049230773,0.032820515,0.06235898,0.06235898,0.052512825,0.049230773,0.052512825,0.06235898,0.052512825,0.068923086,0.08861539,0.12471796,0.23630771,0.36102566,0.44964105,0.47589746,0.44307697,0.39056414,0.28225642,0.27897438,0.41682056,0.69251287,1.0666667,1.1454359,1.4276924,1.9035898,2.5698464,3.43959,4.125539,4.493129,4.630975,4.650667,4.6900516,4.7556925,4.7261543,4.388103,3.82359,3.4264617,3.2754874,3.1606157,2.9833848,2.7208207,2.4352822,2.8127182,3.1540515,3.0490258,2.487795,1.8609232,1.5753847,1.4145643,1.2570257,1.0765129,0.9321026,0.90256417,0.86974365,0.67938465,0.39384618,0.28882053,0.14441027,0.14112821,0.21333335,0.3052308,0.37743592,0.43323082,0.40369233,0.38728207,0.44307697,0.5940513,0.761436,0.8566154,0.827077,0.67938465,0.48246157,0.4201026,0.5513847,0.86974365,1.2077949,1.214359,1.782154,3.190154,4.706462,5.7468724,5.868308,6.485334,6.0750775,5.907693,6.166975,5.976616,4.9887185,4.6834874,4.4734364,3.9844105,3.045744,2.546872,2.9144619,3.511795,3.826872,3.4592824,3.2886157,3.2131286,3.3017437,3.4822567,3.5249233,3.945026,4.604718,5.07077,5.2053337,5.146257,5.435077,5.5893335,5.654975,6.0980515,7.817847,10.230155,11.730052,12.484924,13.233232,15.284514,19.534771,23.017027,25.15036,25.291489,22.724924,18.586258,17.64759,17.54913,16.59077,13.755078,11.953232,10.331899,9.02236,8.779488,10.988309,14.28677,16.81395,17.880617,17.706669,17.414566,16.213335,14.693745,12.245335,9.209436,6.892308,5.1954875,4.141949,3.6332312,3.4691284,3.3378465,2.7634873,2.176,1.7920002,1.6246156,1.4802053,1.3817437,1.6475899,2.0742567,2.4385643,2.5206156,5.172513,5.428513,6.3540516,7.2992826,7.79159,7.522462,8.195283,8.864821,9.048616,8.356103,6.498462,4.890257,4.2305646,4.010667,3.8596926,3.5544617,3.8728209,4.7392826,5.208616,5.0182567,4.578462,3.6496413,2.6945643,2.0709746,1.7887181,1.4966155,1.8740515,2.4615386,2.8160002,2.861949,2.8980515,3.0326157,2.5173335,1.8281027,1.3489232,1.3718976,2.0808206,2.8258464,3.6332312,4.309334,4.457026,4.332308,3.8367183,3.1081028,2.3269746,1.6771283,1.2635899,1.0404103,0.9321026,0.86974365,0.80738467,0.8467693,0.9189744,0.9419488,0.90584624,0.86974365,0.77128214,0.51856416,0.256,0.098461546,0.12143591,0.17066668,0.18379489,0.13456412,0.052512825,0.016410258,0.026256412,0.03938462,0.04594872,0.04594872,0.04594872,0.02297436,0.006564103,0.0,0.0,0.0,0.013128206,0.016410258,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.006564103,0.0,0.0,0.0,0.08533334,0.25271797,0.44307697,0.5546667,0.45620516,0.3249231,0.22646156,0.20676924,0.28225642,0.4266667,0.32820517,0.2231795,0.16738462,0.18379489,0.24287182,0.256,0.19692309,0.10502565,0.02297436,0.0,0.0,0.0,0.0,0.27241027,1.3587693,2.4451284,2.7700515,2.3926156,1.4834872,0.33476925,0.3708718,0.51856416,0.8172308,1.1651284,1.3128207,1.020718,0.7253334,0.79425645,1.017436,0.6268718,0.40697438,0.4594872,0.61374366,0.65312827,0.33476925,0.14112821,0.04594872,0.052512825,0.13784617,0.25928208,0.2100513,0.190359,0.16410258,0.13128206,0.108307704,0.108307704,0.12471796,0.08861539,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.032820515,0.052512825,0.052512825,0.016410258,0.15097436,0.19364104,0.18707694,0.15753847,0.12143591,0.02297436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01969231,0.055794876,0.09189744,0.21333335,0.14441027,0.06564103,0.072205134,0.18379489,0.32820517,0.45620516,0.56123084,0.61374366,0.56451285,0.6268718,0.76800007,0.92225647,1.0601027,1.204513,1.4736412,1.8445129,2.2646155,2.674872,2.989949,3.2722054,3.058872,2.8488207,2.806154,2.7306669,2.7306669,3.0523078,3.5216413,3.6758976,2.7602053,2.225231,2.172718,2.6617439,3.4756925,4.135385,3.2328207,3.2164104,4.132103,5.6976414,7.3091288,7.003898,7.722667,8.756514,9.449026,9.216001,8.897642,9.760821,11.257437,12.028719,9.91836,9.235693,9.275078,9.317744,8.910769,7.8736415,8.129642,7.259898,6.0324106,5.106872,5.0215387,6.1440005,7.716103,7.0793853,4.2863593,2.0742567,1.3292309,1.2077949,1.4703591,2.0184617,2.8849232,3.8498464,4.1091285,3.7218463,3.05559,2.7602053,2.7503593,2.7634873,2.7273848,2.6223593,2.487795,2.425436,2.0250258,1.4769232,1.0305642,1.0075898,0.8730257,0.6301539,0.35446155,0.13456412,0.06235898,0.072205134,0.07548718,0.06564103,0.052512825,0.07548718,0.026256412,0.016410258,0.009846155,0.0,0.0,0.013128206,0.016410258,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.016410258,0.016410258,0.03938462,0.055794876,0.06235898,0.049230773,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.016410258,0.013128206,0.0,0.0,0.0,0.006564103,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.016410258,0.016410258,0.016410258,0.02297436,0.029538464,0.026256412,0.016410258,0.03938462,0.06564103,0.25271797,0.5218462,0.5349744,0.38728207,0.36102566,0.50543594,0.81394875,1.204513,1.8149745,2.1956925,2.4352822,2.428718,1.8904617,1.7460514,1.6443079,1.401436,1.0666667,0.94523084,1.0075898,1.214359,1.2996924,1.2406155,1.2504616,1.3620514,1.2800001,1.2471796,1.3850257,1.6771283,1.7033848,1.5819489,1.276718,0.892718,0.6859488,0.88287187,1.0601027,1.1979488,1.2832822,1.2832822,0.79425645,0.48902568,0.3117949,0.2231795,0.19692309,0.29538465,0.29210258,0.41025645,0.6498462,0.80738467,0.761436,0.5907693,0.33476925,0.0951795,0.04594872,0.108307704,0.06564103,0.01969231,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.032820515,0.052512825,0.11158975,0.32164106,0.40697438,0.46276927,0.46933338,0.4397949,0.4266667,0.32820517,0.3511795,0.45620516,0.60061544,0.74830776,0.80738467,0.92553854,1.1979488,1.719795,2.546872,3.43959,4.020513,4.33559,4.4832826,4.59159,4.6769233,4.6900516,4.4340515,3.8432825,2.9768207,2.9505644,3.1081028,3.2196925,3.1540515,2.8980515,2.7766156,2.5895386,2.1956925,1.6049232,1.0075898,0.8008206,0.62030774,0.47261542,0.3708718,0.32164106,0.27241027,0.23958977,0.19364104,0.13128206,0.108307704,0.108307704,0.12471796,0.19364104,0.32820517,0.5481026,0.7318975,0.7318975,0.6235898,0.508718,0.5349744,0.67938465,0.8730257,0.94523084,0.8467693,0.64000005,0.5316923,0.60389745,0.90912825,1.3718976,1.8018463,2.6322052,3.058872,3.1737437,3.4888208,4.9296412,5.7107697,6.3901544,7.8670774,9.465437,8.940309,6.3540516,4.7917953,4.7491283,5.1954875,3.570872,2.1530259,2.1300514,2.6551797,3.0326157,2.7175386,3.373949,3.767795,4.263385,5.0018463,5.904411,5.5138464,4.565334,3.9253337,3.764513,3.570872,4.1452312,5.1298466,7.5520005,11.175385,14.496821,17.424412,17.762463,15.894976,13.548308,13.794462,16.59077,19.945026,23.289438,25.668924,25.74113,22.33436,18.005335,15.228719,15.205745,17.867489,18.868515,17.26031,13.715693,9.9282055,8.621949,11.283693,14.503386,17.28,19.367386,21.270975,18.743795,16.518566,13.883078,10.981745,8.835282,6.6002054,5.5565133,5.3858466,5.802667,6.560821,5.4383593,3.7120004,2.3302567,1.6738462,1.5425643,1.5425643,1.6771283,2.0151796,2.412308,2.5337439,5.4908724,5.074052,5.0149746,5.152821,5.2053337,4.8016415,5.579488,6.2490263,6.2227697,5.405539,4.204308,4.0303593,3.31159,2.9440002,3.0326157,2.8849232,2.8980515,3.4494362,4.2207184,4.568616,3.501949,3.7284105,3.7185643,3.5380516,3.2689233,3.0326157,2.4155898,2.038154,1.7723079,1.6344616,1.7887181,2.3729234,2.4582565,2.740513,3.0884104,2.556718,2.2022567,2.1956925,2.477949,2.930872,3.3805132,3.9023592,3.895795,3.5282054,3.0391798,2.7634873,1.7920002,1.2471796,0.95835906,0.8205129,0.80738467,0.9124103,0.9878975,1.0338463,1.0469744,1.0404103,0.88287187,0.6170257,0.34789747,0.17723078,0.17066668,0.17066668,0.14112821,0.09189744,0.052512825,0.06564103,0.0951795,0.07548718,0.052512825,0.04594872,0.04594872,0.03938462,0.029538464,0.013128206,0.0,0.0,0.0032820515,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0,0.0,0.0,0.0,0.19364104,0.3511795,0.38728207,0.3446154,0.38400003,0.40697438,0.3117949,0.24287182,0.28225642,0.4397949,0.28225642,0.14769232,0.08205129,0.12143591,0.28225642,0.380718,0.23302566,0.08205129,0.029538464,0.02297436,0.0032820515,0.0,0.0,0.055794876,0.27241027,0.48902568,0.5546667,0.6892308,1.0010257,1.4966155,1.5819489,1.1323078,0.76800007,0.67938465,0.64000005,0.5152821,0.45292312,0.49887183,0.5415385,0.30851284,0.23630771,0.3117949,0.44964105,0.5349744,0.43323082,0.256,0.190359,0.30851284,0.5907693,0.9189744,0.6662565,0.446359,0.31507695,0.25271797,0.18051283,0.12143591,0.14112821,0.13128206,0.07876924,0.036102567,0.016410258,0.013128206,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.01969231,0.029538464,0.029538464,0.0032820515,0.01969231,0.016410258,0.013128206,0.009846155,0.0,0.0,0.006564103,0.009846155,0.0032820515,0.0,0.0,0.006564103,0.02297436,0.032820515,0.013128206,0.013128206,0.01969231,0.032820515,0.052512825,0.06564103,0.09189744,0.07876924,0.06235898,0.072205134,0.12143591,0.02297436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06235898,0.190359,0.3249231,0.45620516,0.4594872,0.47917953,0.5481026,0.5973334,0.5284103,0.5513847,0.6629744,0.78769237,0.80738467,0.93866676,1.2438976,1.591795,1.7788719,1.5360001,1.3161026,1.6443079,2.3269746,2.9538465,2.8816411,2.809436,2.5829747,2.300718,2.048,1.8773335,1.8773335,1.6475899,1.5655385,1.654154,1.5786668,1.7723079,2.034872,2.172718,2.3171284,2.92759,5.0215387,7.1483083,8.979693,10.345026,11.21477,10.978462,11.201642,11.71036,12.373334,13.098668,13.512206,15.504412,16.384,14.608412,9.770667,7.817847,8.887795,11.201642,13.633642,15.711181,15.360002,14.260514,12.662155,10.817642,8.976411,9.337437,9.472001,8.086975,5.3136415,2.733949,2.038154,2.103795,2.3762052,2.6978464,3.31159,3.7874875,3.7120004,3.255795,2.605949,1.9790771,1.7033848,1.7362052,1.8642052,1.8149745,1.2406155,1.5031796,1.4244103,1.0765129,0.6301539,0.36102566,0.3708718,0.34133336,0.27241027,0.17723078,0.072205134,0.036102567,0.01969231,0.016410258,0.01969231,0.016410258,0.006564103,0.009846155,0.01969231,0.026256412,0.036102567,0.03938462,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.02297436,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.013128206,0.013128206,0.006564103,0.0,0.0,0.0,0.006564103,0.006564103,0.0,0.0,0.0,0.0,0.006564103,0.016410258,0.016410258,0.009846155,0.009846155,0.013128206,0.009846155,0.0,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.013128206,0.013128206,0.026256412,0.032820515,0.02297436,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.006564103,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.013128206,0.013128206,0.006564103,0.0,0.0,0.0,0.0032820515,0.0032820515,0.006564103,0.02297436,0.04266667,0.04266667,0.02297436,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.016410258,0.026256412,0.036102567,0.01969231,0.009846155,0.016410258,0.016410258,0.059076928,0.11158975,0.15753847,0.19364104,0.20348719,0.4594872,0.69907695,0.8467693,0.8763078,0.827077,1.6508719,1.8445129,1.7362052,1.5327181,1.3193847,1.1126155,1.276718,1.1782565,0.7811283,0.6301539,0.64000005,0.75487185,0.90584624,1.020718,1.0436924,1.086359,1.2340513,1.3981539,1.4572309,1.2504616,1.2373334,1.4473847,1.5688206,1.5392822,1.5655385,1.3883078,1.3554872,1.4539489,1.6672822,1.9889232,1.5786668,0.90584624,0.43651286,0.29210258,0.25928208,0.26912823,0.27241027,0.40369233,0.65641034,0.892718,0.7581539,0.53825647,0.31507695,0.14769232,0.068923086,0.052512825,0.029538464,0.01969231,0.026256412,0.036102567,0.04594872,0.049230773,0.04266667,0.032820515,0.02297436,0.006564103,0.006564103,0.026256412,0.08205129,0.2100513,0.36430773,0.41682056,0.39384618,0.33805132,0.318359,0.30851284,0.3446154,0.38400003,0.39712822,0.35774362,0.3314872,0.38728207,0.57764107,0.955077,1.5589745,2.4615386,3.1442053,3.5216413,3.6004105,3.5052311,3.698872,4.096,4.1485133,3.6791797,2.8914874,2.5337439,2.5796926,2.9538465,3.2853336,2.9111798,2.172718,1.585231,1.2570257,1.0601027,0.6301539,0.51856416,0.4660513,0.4135385,0.36102566,0.3708718,0.38728207,0.29538465,0.2231795,0.21333335,0.2297436,0.21989745,0.256,0.35774362,0.5874872,1.0633847,1.3226668,1.3062565,1.1716924,1.017436,0.8763078,0.8467693,0.86974365,0.88615394,0.8795898,0.8960001,0.8172308,0.8598975,1.142154,1.5491283,1.7526156,1.7132308,1.7985642,2.103795,2.7602053,3.9286156,4.017231,4.670359,6.626462,9.235693,10.47959,7.315693,5.5138464,5.5105643,6.36718,5.7665644,2.8488207,2.0217438,2.3269746,2.8914874,2.934154,2.6486156,2.6157951,3.2886157,4.9985647,7.9425645,8.530052,8.562873,8.434873,8.809027,10.627283,10.006975,7.7456417,7.634052,11.0375395,16.889437,19.426462,19.974566,18.425438,15.885129,14.674052,15.721026,16.873028,18.753643,21.507284,24.81231,22.99077,20.233849,19.268925,20.601437,22.531284,17.664001,14.043899,11.1294365,9.517949,10.965334,13.361232,14.92677,16.99118,19.334566,20.184616,20.801643,20.63754,17.975796,13.7386675,11.483898,9.3768215,8.395488,7.8145647,7.3091288,6.9645133,4.3749747,2.9046156,2.169436,1.8904617,1.8838975,1.9331284,1.8838975,1.9593848,2.1858463,2.3860514,4.9362054,5.3398976,4.850872,4.4077954,4.273231,4.0369234,4.3027697,4.5817437,4.604718,4.2601027,3.6036925,3.501949,3.2295387,3.2951798,3.7349746,4.1091285,3.9647183,3.9318976,4.0402055,4.0467696,3.4166157,3.623385,3.7874875,4.1124105,4.4373336,4.2338467,3.3575387,3.0326157,2.6354873,2.0742567,1.8051283,2.3663592,3.0293336,3.8695388,4.6276927,4.713026,4.1846156,3.4494362,2.8225644,2.5009232,2.5731285,2.6420515,2.789744,2.8816411,2.8488207,2.6880002,1.9298463,1.3817437,1.0568206,0.9616411,1.1027694,1.1651284,1.148718,1.1158975,1.0568206,0.9189744,0.7778462,0.58420515,0.39712822,0.26256412,0.21989745,0.17066668,0.12143591,0.08533334,0.06564103,0.07548718,0.098461546,0.08861539,0.06564103,0.04266667,0.026256412,0.01969231,0.013128206,0.006564103,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.16738462,0.29538465,0.33805132,0.32820517,0.36758977,0.4135385,0.2986667,0.21333335,0.256,0.40697438,0.40369233,0.26256412,0.17066668,0.19364104,0.28882053,0.49230772,0.5513847,0.3446154,0.036102567,0.059076928,0.1148718,0.118153855,0.08861539,0.052512825,0.04594872,0.009846155,0.0,0.10502565,0.35446155,0.71548724,0.75487185,0.5152821,0.30194873,0.2231795,0.190359,0.15425642,0.15425642,0.17066668,0.17066668,0.09189744,0.07548718,0.108307704,0.16410258,0.20348719,0.18379489,0.12143591,0.10502565,0.16738462,0.29538465,0.43323082,0.3249231,0.27569234,0.25271797,0.21989745,0.13456412,0.068923086,0.06564103,0.068923086,0.055794876,0.026256412,0.016410258,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.01969231,0.016410258,0.013128206,0.01969231,0.02297436,0.009846155,0.098461546,0.16738462,0.17723078,0.1148718,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0032820515,0.01969231,0.036102567,0.032820515,0.049230773,0.06235898,0.09189744,0.13128206,0.14112821,0.08205129,0.03938462,0.016410258,0.01969231,0.049230773,0.009846155,0.009846155,0.013128206,0.009846155,0.009846155,0.009846155,0.0032820515,0.02297436,0.059076928,0.072205134,0.22646156,0.40369233,0.636718,0.82379496,0.7187693,0.5677949,1.3357949,2.0841026,2.2186668,1.4802053,1.2340513,1.4309745,1.8248206,2.1070771,1.8937438,1.9462565,3.1113849,3.5938463,2.8389745,1.5163078,0.8598975,1.1913847,2.2186668,3.0654361,2.284308,2.1792822,1.8838975,1.5589745,1.3456411,1.3718976,1.4080001,1.4441026,1.5655385,1.7526156,1.8937438,2.03159,2.1169233,2.169436,2.5304618,3.8695388,5.1232824,6.1374364,7.351795,8.083693,6.488616,6.2818465,6.114462,6.518154,7.778462,9.931488,9.613129,11.10318,11.365745,9.350565,6.009436,5.1167183,6.49518,8.786052,10.9226675,12.130463,11.513436,10.896411,10.581334,10.322052,9.304616,8.815591,8.362667,7.3419495,5.6352825,3.623385,3.2164104,2.5206156,2.0873847,2.1398976,2.556718,2.7208207,2.349949,1.9593848,1.7690258,1.7132308,1.5327181,1.3784616,1.3981539,1.5031796,1.3981539,1.079795,0.82379496,0.6301539,0.4660513,0.28882053,0.16410258,0.128,0.1148718,0.08205129,0.029538464,0.009846155,0.0032820515,0.0032820515,0.0032820515,0.0,0.0,0.0032820515,0.009846155,0.013128206,0.01969231,0.01969231,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.02297436,0.0032820515,0.0,0.0032820515,0.013128206,0.026256412,0.006564103,0.0,0.0,0.0032820515,0.016410258,0.02297436,0.013128206,0.0032820515,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0,0.006564103,0.0032820515,0.0032820515,0.006564103,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.016410258,0.029538464,0.052512825,0.055794876,0.036102567,0.016410258,0.009846155,0.059076928,0.08861539,0.068923086,0.009846155,0.0032820515,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.006564103,0.006564103,0.0032820515,0.0,0.0,0.013128206,0.013128206,0.009846155,0.009846155,0.013128206,0.029538464,0.02297436,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.02297436,0.03938462,0.06564103,0.055794876,0.026256412,0.006564103,0.006564103,0.016410258,0.04266667,0.07876924,0.12471796,0.19364104,0.31507695,0.55794877,0.90584624,1.1355898,1.1684103,1.0633847,1.3095386,1.394872,1.394872,1.2898463,0.9353847,0.67282057,0.7417436,0.79097444,0.67282057,0.4397949,0.7318975,0.8467693,0.86974365,0.8763078,0.94523084,1.1520001,1.3193847,1.4408206,1.5524104,1.719795,2.0184617,2.0053334,1.8281027,1.6640002,1.719795,1.4605129,1.6672822,2.605949,3.6693337,3.373949,2.8389745,2.1398976,1.5885129,1.2931283,1.1520001,1.0305642,0.7844103,0.63343596,0.65969235,0.81394875,0.82379496,0.6629744,0.44964105,0.25928208,0.13128206,0.101743594,0.12471796,0.15753847,0.16410258,0.108307704,0.09189744,0.0951795,0.108307704,0.12471796,0.11158975,0.04594872,0.009846155,0.009846155,0.059076928,0.18379489,0.37743592,0.38400003,0.32164106,0.26584616,0.26256412,0.3249231,0.4004103,0.4397949,0.4135385,0.31507695,0.28882053,0.31507695,0.39056414,0.5316923,0.7811283,1.529436,2.3072822,2.8750772,3.1442053,3.1803079,3.370667,3.8071797,3.9023592,3.511795,2.934154,2.7798977,2.989949,3.2787695,3.3476925,2.8882053,2.1333334,1.5556924,1.2077949,0.9911796,0.65312827,0.52512825,0.4201026,0.34133336,0.29538465,0.28882053,0.28882053,0.25271797,0.23302566,0.25271797,0.3052308,0.35774362,0.39056414,0.42338464,0.5316923,0.8336411,1.0633847,1.1454359,1.1651284,1.2077949,1.3554872,1.1290257,1.0108719,0.8960001,0.7778462,0.7417436,0.90256417,1.1520001,1.404718,1.5786668,1.6016412,1.522872,1.9396925,3.446154,6.3376417,10.617436,8.385642,6.5739493,7.466667,11.188514,15.717745,12.475078,9.065026,7.506052,7.936001,8.595693,4.647385,2.9013336,2.9735386,3.9876926,4.5390773,4.378257,4.2469745,4.535795,5.290667,6.2096415,6.62318,6.957949,7.4371285,8.710565,11.858052,12.534155,11.579078,10.752001,11.0605135,12.754052,14.683899,14.864411,14.749539,14.805334,14.5263605,14.464001,14.742975,15.655386,17.35877,19.866259,21.083899,21.431797,21.418669,21.074053,19.925335,16.328207,13.161027,11.460924,12.018872,15.386257,17.417847,16.433231,14.523078,13.252924,13.6697445,17.168411,20.096,19.396925,15.199181,10.837335,8.080411,6.5903597,5.5991797,4.778667,4.2436924,2.917744,2.2613335,2.0184617,2.0118976,2.15959,2.3171284,2.2744617,2.3302567,2.4976413,2.5042052,4.5095387,5.0051284,4.417641,3.8662567,3.767795,3.8071797,3.882667,4.240411,4.637539,4.8082056,4.46359,4.1583595,4.2994876,4.8311796,5.536821,6.048821,5.5663595,4.9394875,4.325744,3.95159,4.1452312,4.4865646,4.7261543,4.9427695,5.100308,5.0642056,4.31918,4.092718,3.8006158,3.308308,2.92759,3.1048207,4.1222568,5.1889234,5.901129,6.2555904,6.0160003,4.9526157,3.8006158,2.9243078,2.3236926,1.7263591,1.6410258,1.8379488,2.038154,1.9068719,1.5392822,1.2077949,1.0075898,0.9944616,1.1881026,1.1684103,1.1158975,1.0601027,0.9682052,0.761436,0.58420515,0.43323082,0.31507695,0.23630771,0.21989745,0.2100513,0.20020515,0.20020515,0.19364104,0.118153855,0.08205129,0.068923086,0.059076928,0.03938462,0.016410258,0.006564103,0.0032820515,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.009846155,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.01969231,0.01969231,0.009846155,0.009846155,0.01969231,0.03938462,0.06564103,0.04266667,0.01969231,0.0032820515,0.0,0.0,0.17394873,0.25271797,0.32164106,0.4201026,0.54482055,0.58092314,0.37415388,0.24943592,0.30194873,0.40697438,0.5415385,0.60389745,0.57764107,0.5021539,0.47917953,0.5940513,0.72861546,0.7056411,0.7515898,1.5097437,1.595077,1.1191796,0.5152821,0.09189744,0.04594872,0.009846155,0.0032820515,0.009846155,0.013128206,0.013128206,0.0032820515,0.0,0.0032820515,0.026256412,0.08533334,0.08533334,0.07548718,0.08533334,0.10502565,0.09189744,0.2855385,0.27241027,0.15097436,0.036102567,0.06235898,0.08205129,0.06564103,0.03938462,0.01969231,0.0,0.013128206,0.072205134,0.128,0.13784617,0.06564103,0.01969231,0.013128206,0.02297436,0.032820515,0.02297436,0.02297436,0.016410258,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.049230773,0.032820515,0.009846155,0.0032820515,0.013128206,0.02297436,0.12471796,0.18707694,0.18051283,0.108307704,0.0,0.0,0.0,0.0032820515,0.009846155,0.01969231,0.01969231,0.013128206,0.04266667,0.11158975,0.19692309,0.23302566,0.3511795,0.571077,0.69579494,0.3052308,0.12471796,0.036102567,0.006564103,0.0,0.006564103,0.0,0.032820515,0.08205129,0.118153855,0.11158975,0.14769232,0.4397949,0.53825647,0.44964105,0.63343596,1.1552821,1.7263591,2.2547693,2.3040001,1.086359,0.84348726,1.6804104,2.4943593,2.6486156,1.9561027,2.349949,2.8717952,3.2984617,3.3641028,2.7602053,2.294154,3.2820516,3.495385,2.3762052,1.0338463,0.48574364,0.7253334,1.5655385,2.228513,1.3751796,1.4408206,1.4309745,1.4244103,1.4539489,1.5163078,1.3915899,1.4834872,1.6771283,1.8970258,2.103795,2.2088206,2.169436,2.1891284,2.7995899,4.84759,5.2578464,4.338872,4.0500517,4.2240005,2.5764105,2.546872,2.3729234,2.6617439,3.7152824,5.5302567,6.803693,7.896616,7.817847,6.665847,5.6418467,5.0018463,6.1768208,8.264206,9.96759,9.580308,7.975385,7.955693,8.579283,9.07159,8.828718,7.387898,6.298257,5.789539,5.412103,4.0303593,3.6660516,2.7011285,1.9593848,1.7558975,1.8871796,1.9331284,1.6213335,1.2898463,1.142154,1.2242053,1.2242053,1.1027694,1.2406155,1.5721027,1.5688206,0.88943595,0.4201026,0.23958977,0.25928208,0.2100513,0.06564103,0.02297436,0.01969231,0.02297436,0.02297436,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0032820515,0.009846155,0.0032820515,0.0,0.0032820515,0.013128206,0.026256412,0.006564103,0.0,0.0,0.0032820515,0.009846155,0.026256412,0.016410258,0.0032820515,0.0,0.006564103,0.0,0.0,0.0,0.0,0.006564103,0.01969231,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.009846155,0.02297436,0.026256412,0.04266667,0.055794876,0.059076928,0.032820515,0.01969231,0.06564103,0.0951795,0.07548718,0.026256412,0.01969231,0.013128206,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0,0.006564103,0.03938462,0.068923086,0.059076928,0.016410258,0.0,0.006564103,0.009846155,0.016410258,0.01969231,0.006564103,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0032820515,0.006564103,0.0032820515,0.0,0.009846155,0.0032820515,0.0,0.0,0.0,0.0032820515,0.006564103,0.0032820515,0.0,0.0,0.0032820515,0.016410258,0.029538464,0.03938462,0.055794876,0.03938462,0.01969231,0.013128206,0.026256412,0.052512825,0.03938462,0.03938462,0.14769232,0.35446155,0.5415385,0.6235898,0.76800007,0.892718,0.9682052,1.024,1.024,1.0929232,1.148718,1.0469744,0.56451285,0.56451285,0.5677949,0.6071795,0.6104616,0.41025645,0.7122052,0.92553854,1.017436,1.0568206,1.2012309,1.4441026,1.5327181,1.657436,1.9692309,2.605949,3.2164104,3.117949,2.540308,1.8773335,1.654154,1.4112822,1.9396925,3.2229745,4.4898467,4.2174363,3.9187696,3.5478978,3.0523078,2.4943593,2.0644104,1.7558975,1.2438976,0.7975385,0.574359,0.5940513,0.65969235,0.6071795,0.5546667,0.5349744,0.5284103,0.4397949,0.4201026,0.41682056,0.39384618,0.34133336,0.29538465,0.20348719,0.15097436,0.14769232,0.15097436,0.0951795,0.04266667,0.01969231,0.068923086,0.26256412,0.52512825,0.574359,0.51856416,0.44307697,0.4266667,0.49887183,0.60389745,0.6826667,0.6859488,0.57764107,0.5546667,0.5874872,0.61374366,0.65312827,0.7811283,1.4867693,2.2186668,2.7766156,3.0687182,3.1245131,3.1540515,3.3542566,3.3772311,3.1606157,2.9144619,2.9965131,3.2229745,3.2787695,3.0260515,2.5140514,2.0053334,1.6213335,1.3292309,1.083077,0.8041026,0.51856416,0.3511795,0.2855385,0.28882053,0.30851284,0.37743592,0.57764107,0.636718,0.5973334,0.81066674,0.7253334,0.4955898,0.35774362,0.380718,0.5021539,0.702359,0.9485129,1.1913847,1.4211283,1.6771283,1.3883078,1.1290257,0.8960001,0.7187693,0.65641034,0.8992821,1.2077949,1.4408206,1.522872,1.4178462,1.4506668,2.1891284,4.414359,8.664616,15.232001,12.993642,9.504821,8.470975,11.421539,17.700104,15.366566,11.017847,8.152616,8.14277,10.240001,8.3364105,5.1889234,3.8859491,4.673641,4.9394875,4.8804107,5.0543594,5.290667,5.3169236,4.7524104,4.781949,5.280821,6.377026,8.323282,11.487181,13.082257,13.456411,12.721231,11.319796,10.020103,10.735591,11.040821,11.58236,12.268309,12.245335,12.179693,13.046155,13.942155,14.897232,16.869745,19.111385,20.502975,20.522669,19.072002,16.489027,16.06236,13.922462,12.09436,11.864616,13.781334,14.260514,13.052719,11.063796,9.639385,10.555078,14.03077,17.283283,18.290873,16.482462,12.73436,8.664616,5.228308,3.2295387,2.5632823,2.2121027,1.9528207,1.8018463,1.8051283,1.9823592,2.3302567,2.7798977,3.0391798,3.1277952,3.0129232,2.5862565,4.3618464,4.010667,3.508513,3.186872,3.1606157,3.2951798,3.570872,4.348718,5.1232824,5.533539,5.362872,5.1856413,5.671385,6.3573337,6.921847,7.181129,6.311385,5.3924108,4.634257,4.397949,5.1954875,6.2129235,6.5444107,6.0947695,5.346462,5.353026,4.7458467,4.3716927,4.3290257,4.5489235,4.818052,4.841026,5.789539,6.5805135,6.75118,6.47877,6.380308,5.4416413,4.4406157,3.5807183,2.4681027,1.6508719,1.1913847,1.079795,1.142154,1.0272821,0.96492314,0.90912825,0.8960001,0.94523084,1.0666667,0.9714873,0.92553854,0.8763078,0.78769237,0.6268718,0.4135385,0.29210258,0.21989745,0.190359,0.21989745,0.27241027,0.3052308,0.33805132,0.3314872,0.190359,0.08861539,0.055794876,0.052512825,0.049230773,0.02297436,0.016410258,0.009846155,0.0032820515,0.0032820515,0.0,0.0,0.006564103,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.03938462,0.04266667,0.026256412,0.026256412,0.03938462,0.07548718,0.13456412,0.08533334,0.036102567,0.006564103,0.0,0.0,0.190359,0.30851284,0.38728207,0.49230772,0.7187693,0.83035904,0.63343596,0.48574364,0.48246157,0.44964105,0.56451285,0.86974365,0.98461545,0.84348726,0.7056411,0.7450257,0.92553854,1.2504616,1.8445129,2.930872,2.9702566,2.0151796,0.86646163,0.08861539,0.0,0.0,0.006564103,0.016410258,0.02297436,0.02297436,0.0032820515,0.0,0.009846155,0.055794876,0.17394873,0.17066668,0.14769232,0.16738462,0.21333335,0.18379489,0.60061544,0.5874872,0.3446154,0.108307704,0.14769232,0.16410258,0.108307704,0.049230773,0.016410258,0.009846155,0.01969231,0.02297436,0.04594872,0.07548718,0.03938462,0.02297436,0.02297436,0.036102567,0.049230773,0.055794876,0.055794876,0.055794876,0.04594872,0.029538464,0.013128206,0.009846155,0.009846155,0.009846155,0.009846155,0.009846155,0.013128206,0.016410258,0.016410258,0.009846155,0.009846155,0.009846155,0.006564103,0.0032820515,0.01969231,0.06564103,0.04594872,0.016410258,0.0032820515,0.01969231,0.059076928,0.10502565,0.07548718,0.029538464,0.0,0.0,0.0,0.0,0.013128206,0.03938462,0.06564103,0.055794876,0.04266667,0.11158975,0.27897438,0.47261542,0.58092314,0.827077,1.1881026,1.3259488,0.58092314,0.23630771,0.098461546,0.07548718,0.08205129,0.036102567,0.052512825,0.23302566,0.45292312,0.62030774,0.69579494,0.84348726,1.2077949,1.2996924,1.2438976,1.785436,2.540308,3.2229745,3.7382567,3.4789746,1.3128207,1.2668719,1.3915899,1.4998976,1.5655385,1.7296412,3.2820516,4.010667,4.1124105,3.7710772,3.1507695,2.6453335,2.225231,1.6902566,1.1027694,0.77456415,0.62030774,0.56451285,0.7975385,1.1158975,0.92225647,1.0765129,1.3850257,1.7329233,1.9659488,1.8806155,1.5622566,1.3620514,1.339077,1.5097437,1.8281027,2.03159,2.1530259,2.1924105,2.6354873,4.460308,5.0018463,3.245949,1.9331284,1.9790771,2.4582565,2.6157951,2.6683078,2.7536411,2.8717952,2.9013336,6.7774363,8.129642,8.375795,8.333129,8.2215395,6.9382567,7.9097443,10.200616,12.12718,11.277129,8.470975,8.55959,8.969847,8.664616,8.132924,6.11118,4.585026,4.417641,4.9460516,3.9712822,3.2951798,2.678154,2.1858463,1.8576412,1.723077,1.7690258,1.782154,1.5721027,1.1782565,0.86974365,0.7417436,0.8041026,1.1651284,1.5195899,1.1191796,0.6498462,0.2231795,0.01969231,0.013128206,0.0,0.0,0.0,0.009846155,0.029538464,0.049230773,0.01969231,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.029538464,0.02297436,0.016410258,0.016410258,0.02297436,0.009846155,0.0032820515,0.0032820515,0.0032820515,0.016410258,0.026256412,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.006564103,0.0032820515,0.0,0.0,0.006564103,0.013128206,0.016410258,0.02297436,0.006564103,0.009846155,0.03938462,0.072205134,0.052512825,0.026256412,0.016410258,0.016410258,0.01969231,0.03938462,0.03938462,0.032820515,0.02297436,0.016410258,0.006564103,0.006564103,0.0032820515,0.0032820515,0.0,0.0,0.009846155,0.0032820515,0.0,0.0032820515,0.016410258,0.055794876,0.1148718,0.101743594,0.02297436,0.009846155,0.0032820515,0.013128206,0.032820515,0.04266667,0.013128206,0.0032820515,0.006564103,0.009846155,0.0032820515,0.0,0.0032820515,0.009846155,0.013128206,0.016410258,0.009846155,0.03938462,0.029538464,0.013128206,0.009846155,0.006564103,0.009846155,0.013128206,0.009846155,0.0032820515,0.0,0.013128206,0.013128206,0.013128206,0.009846155,0.0032820515,0.0032820515,0.0,0.016410258,0.052512825,0.098461546,0.098461546,0.13456412,0.3314872,0.6268718,0.79425645,0.67938465,0.47589746,0.36102566,0.4201026,0.636718,0.8369231,0.892718,0.82379496,0.6301539,0.30194873,0.6695385,0.76800007,0.7417436,0.6892308,0.6695385,0.7220513,0.9714873,1.211077,1.4178462,1.7493335,1.9429746,2.0217438,2.2908719,3.0030773,4.3290257,4.8344617,4.59159,3.6168208,2.3663592,1.7526156,1.7165129,2.4451284,3.3345644,3.9942567,4.279795,4.3651285,4.3585644,4.1091285,3.5544617,2.7273848,2.0644104,1.3357949,0.7384616,0.39384618,0.34133336,0.38400003,0.45620516,0.58092314,0.7515898,0.9189744,0.78769237,0.6826667,0.60389745,0.56451285,0.58420515,0.5349744,0.33805132,0.17394873,0.118153855,0.128,0.128,0.08205129,0.04594872,0.118153855,0.4266667,0.8369231,1.0601027,1.086359,0.9714873,0.83035904,0.8533334,0.9419488,1.0404103,1.083077,0.97805136,0.9156924,0.97805136,1.0929232,1.2570257,1.5327181,2.2219489,2.6978464,2.9735386,3.0752823,3.0424619,2.9243078,2.8422565,2.7995899,2.802872,2.865231,2.9669745,2.9801028,2.806154,2.4320002,1.972513,1.7460514,1.5491283,1.3850257,1.2406155,1.0699488,0.6892308,0.5677949,0.57764107,0.6301539,0.69251287,1.0994873,1.7066668,1.8116925,1.4736412,1.5163078,1.079795,0.5284103,0.24943592,0.29538465,0.36758977,0.5316923,0.8730257,1.2537436,1.5556924,1.6869745,1.4802053,1.1651284,0.90256417,0.764718,0.7515898,0.8402052,0.9714873,1.1684103,1.332513,1.2307693,1.2504616,1.9954873,4.066462,8.077128,14.660924,14.102976,10.994873,8.779488,9.731283,14.92677,13.820719,9.93477,7.017026,7.026872,10.128411,11.542975,7.6143594,4.8672824,4.95918,4.673641,4.1911798,4.57518,5.218462,5.651693,5.536821,5.3792825,5.9602056,7.315693,9.206155,11.113027,12.245335,12.665437,12.396309,11.595488,10.548513,10.026668,10.643693,10.794667,10.121847,9.511385,10.095591,11.812103,13.08554,14.027489,16.443079,17.641027,18.290873,18.153027,17.040411,14.808617,15.645539,14.313026,11.913847,9.586872,8.51036,6.514872,6.7183595,8.165744,10.177642,12.340514,14.283488,15.675078,17.063385,17.880617,16.423386,11.313231,5.933949,2.789744,2.1234872,1.8970258,1.6213335,1.463795,1.4900514,1.7362052,2.2088206,2.9801028,3.636513,3.8104618,3.4034874,2.605949,3.8006158,3.4691284,3.1671798,2.8882053,2.612513,2.3204105,2.3204105,2.7602053,3.2164104,3.5052311,3.6758976,4.1156926,5.333334,5.7140517,5.2644105,5.6320004,4.9460516,4.3716927,4.4406157,5.110154,5.7665644,7.453539,7.4075904,6.550975,5.546667,4.7917953,3.9122055,3.564308,3.948308,5.0871797,6.820103,8.004924,8.218257,7.821129,6.954667,5.540103,4.6605134,4.0369234,3.6758976,3.31159,2.3958976,2.2121027,1.8084104,1.3259488,0.9321026,0.80738467,1.0272821,1.0732309,1.1060513,1.1749744,1.2373334,1.1126155,0.9288206,0.71548724,0.5152821,0.380718,0.3446154,0.39056414,0.4266667,0.4135385,0.36758977,0.29210258,0.21989745,0.18379489,0.190359,0.21333335,0.15097436,0.128,0.1148718,0.0951795,0.04594872,0.02297436,0.02297436,0.02297436,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.029538464,0.04266667,0.026256412,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02297436,0.4594872,0.61374366,0.40369233,0.36758977,0.76800007,1.0633847,1.0633847,0.79097444,0.47261542,0.37415388,0.44307697,0.62030774,0.72861546,0.47261542,1.0601027,1.8740515,2.3630772,1.9396925,0.0,0.0,0.055794876,0.07876924,0.049230773,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.13456412,0.19692309,0.20020515,0.17066668,0.12143591,0.06235898,0.036102567,0.029538464,0.032820515,0.04594872,0.0951795,0.108307704,0.08861539,0.06564103,0.07548718,0.08861539,0.08205129,0.068923086,0.07876924,0.15097436,0.16410258,0.15753847,0.13456412,0.098461546,0.06235898,0.049230773,0.04594872,0.04594872,0.04594872,0.04594872,0.059076928,0.08861539,0.08205129,0.04594872,0.04594872,0.04594872,0.026256412,0.02297436,0.029538464,0.029538464,0.01969231,0.006564103,0.01969231,0.068923086,0.16738462,0.15425642,0.098461546,0.036102567,0.0,0.0,0.0,0.0,0.04266667,0.11158975,0.13784617,0.101743594,0.06564103,0.19692309,0.47261542,0.65641034,0.99774367,1.1946667,1.0535386,0.77456415,0.94523084,0.446359,0.32820517,0.38400003,0.39056414,0.12143591,0.24287182,0.9517949,1.6049232,2.0151796,2.4418464,2.8324106,1.6836925,1.3357949,2.3105643,3.31159,3.4198978,2.8816411,2.2153847,1.7033848,1.3718976,1.5327181,1.3423591,1.0568206,0.8992821,1.083077,2.937436,3.3476925,3.0982566,2.9407182,3.6004105,5.674667,3.95159,2.4024618,2.300718,2.228513,1.7394873,1.1060513,1.148718,1.8379488,2.28759,1.9954873,1.585231,1.3456411,1.3193847,1.2832822,1.3062565,1.2570257,1.2931283,1.5097437,1.9364104,1.7427694,2.225231,2.537026,2.3827693,2.028308,1.8215386,1.6771283,1.9298463,2.4451284,2.6387694,2.553436,2.4516926,2.5042052,2.5862565,2.2416413,3.3050258,4.9362054,6.678975,7.512616,5.8289237,5.9634876,7.581539,9.527796,10.935796,11.21477,9.055181,8.139488,7.584821,6.813539,5.5696416,4.2994876,3.9286156,4.263385,4.6900516,4.164923,3.1277952,2.284308,1.7952822,1.6508719,1.6640002,1.6508719,1.7591796,1.972513,2.162872,2.0906668,1.017436,0.8763078,0.7844103,0.44964105,0.16738462,0.068923086,0.072205134,0.06564103,0.02297436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.029538464,0.04266667,0.026256412,0.03938462,0.072205134,0.06235898,0.036102567,0.02297436,0.009846155,0.0032820515,0.016410258,0.016410258,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.032820515,0.03938462,0.02297436,0.0,0.0,0.0,0.006564103,0.013128206,0.0,0.013128206,0.006564103,0.006564103,0.016410258,0.016410258,0.03938462,0.026256412,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.02297436,0.029538464,0.029538464,0.029538464,0.02297436,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.016410258,0.016410258,0.016410258,0.02297436,0.04594872,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.02297436,0.0,0.013128206,0.006564103,0.013128206,0.032820515,0.04594872,0.0951795,0.098461546,0.072205134,0.04266667,0.029538464,0.006564103,0.009846155,0.016410258,0.013128206,0.0,0.013128206,0.006564103,0.0,0.0032820515,0.016410258,0.016410258,0.006564103,0.013128206,0.036102567,0.06235898,0.256,0.571077,0.86317956,1.0732309,1.2209232,0.84348726,0.6104616,0.5316923,0.56451285,0.6268718,0.5874872,0.44307697,0.33805132,0.36430773,0.5349744,0.6071795,0.8533334,1.0633847,1.204513,1.4506668,1.6213335,1.5261539,1.3620514,1.4441026,2.2121027,2.7503593,3.058872,3.5577438,4.9526157,8.224821,7.722667,6.189949,4.381539,2.9243078,2.28759,2.9833848,3.7809234,4.4340515,4.6933336,4.3027697,3.8990772,3.6726158,4.056616,4.4996924,3.4494362,2.03159,1.0272821,0.43651286,0.20676924,0.24287182,0.5481026,0.7187693,0.61374366,0.35774362,0.32164106,0.39384618,0.34789747,0.32820517,0.37415388,0.4135385,0.4135385,0.32820517,0.24943592,0.20020515,0.15097436,0.10502565,0.08205129,0.07548718,0.18379489,0.6104616,1.2931283,1.7755898,1.9593848,1.8051283,1.3423591,1.3062565,1.3161026,1.3259488,1.3095386,1.2373334,1.0666667,1.1585642,1.5130258,2.0086155,2.412308,2.678154,2.6551797,2.5764105,2.6026669,2.8225644,2.9571285,2.9636924,2.9440002,2.9636924,3.0358977,2.9505644,2.7733335,2.4746668,2.1300514,1.9232821,1.9232821,1.7591796,1.6246156,1.6082052,1.6935385,1.6935385,1.8215386,1.8642052,1.7920002,1.7558975,2.9505644,4.06318,4.1025643,2.9702566,1.4802053,0.761436,0.4135385,0.3249231,0.35446155,0.36758977,0.36758977,0.512,0.77456415,1.0896411,1.3587693,1.2471796,1.1552821,1.0338463,0.88615394,0.761436,0.67610264,0.60061544,0.6629744,0.85005134,1.020718,1.020718,1.5425643,3.3017437,6.8233852,12.452104,10.059488,8.700719,8.595693,9.6295395,11.336206,9.957745,7.3419495,5.8223596,6.442667,8.956718,8.749949,7.204103,6.245744,6.514872,7.3682055,6.088206,5.5007186,6.3507695,8.001641,8.454565,8.15918,8.326565,8.930462,9.622975,9.7214365,9.829744,10.975181,11.707078,11.37559,10.131693,9.875693,9.334154,9.383386,10.112,10.817642,11.293539,11.605334,12.087796,12.865642,13.853539,15.307488,17.56554,18.638771,17.408,13.610668,11.451077,11.001437,11.313231,11.831796,12.406155,8.631796,7.27959,7.7292314,9.691898,13.184001,17.51631,19.83672,20.368412,18.855387,14.555899,10.443488,6.87918,3.9778464,2.044718,1.5556924,1.2865642,1.1093334,1.0732309,1.1979488,1.463795,2.1366155,2.806154,3.2787695,3.3509746,2.8389745,6.265436,6.1407185,6.2555904,6.0685134,5.428513,4.578462,4.069744,3.761231,3.495385,3.2623591,3.190154,3.570872,4.2896414,4.7524104,4.716308,4.2994876,3.764513,3.9286156,4.420923,5.0116925,5.622154,7.1023593,7.509334,7.312411,6.7216415,5.681231,4.7556925,3.9417439,3.5577438,3.8334363,4.893539,5.4416413,6.045539,6.951385,7.4929237,6.0750775,4.768821,4.1780515,3.948308,3.7874875,3.4560003,2.3171284,2.0053334,1.8051283,1.463795,1.1749744,1.0043077,0.8795898,0.8467693,0.88615394,0.9189744,0.892718,0.827077,0.67282057,0.48246157,0.41682056,0.508718,0.61374366,0.71548724,0.7844103,0.79425645,0.69251287,0.6235898,0.5973334,0.5874872,0.54482055,0.35446155,0.24943592,0.17066668,0.108307704,0.068923086,0.08533334,0.07548718,0.04594872,0.013128206,0.013128206,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.029538464,0.06235898,0.06564103,0.03938462,0.0,0.0,0.0,0.006564103,0.006564103,0.0032820515,0.02297436,0.059076928,0.20348719,0.30851284,0.38728207,0.63343596,0.8730257,0.86646163,0.81394875,0.7187693,0.4135385,0.24615386,0.20676924,0.32164106,0.58420515,0.9747693,1.2373334,1.0633847,0.77128214,0.48902568,0.15753847,0.108307704,0.17394873,0.18051283,0.14441027,0.28225642,0.5349744,0.5973334,0.44307697,0.18707694,0.098461546,0.07876924,0.06564103,0.036102567,0.0,0.0032820515,0.0,0.036102567,0.072205134,0.072205134,0.013128206,0.068923086,0.101743594,0.108307704,0.098461546,0.098461546,0.15425642,0.2100513,0.21989745,0.17394873,0.108307704,0.07876924,0.049230773,0.026256412,0.02297436,0.06564103,0.055794876,0.04594872,0.032820515,0.029538464,0.055794876,0.055794876,0.08533334,0.12471796,0.14769232,0.108307704,0.068923086,0.06564103,0.068923086,0.072205134,0.08205129,0.0951795,0.059076928,0.029538464,0.02297436,0.02297436,0.02297436,0.026256412,0.01969231,0.006564103,0.006564103,0.0032820515,0.009846155,0.01969231,0.04266667,0.08205129,0.08861539,0.059076928,0.02297436,0.0,0.0,0.0,0.02297436,0.049230773,0.118153855,0.30851284,0.6432821,1.014154,1.1684103,1.1388719,1.2537436,1.4703591,1.522872,1.273436,0.88287187,0.8008206,0.5513847,0.54482055,0.69251287,0.88943595,1.0010257,1.014154,1.8871796,2.3171284,1.8838975,1.0502565,1.0404103,0.702359,0.6892308,1.083077,1.3718976,1.4998976,1.6672822,1.7001027,1.4966155,1.020718,0.8960001,0.76800007,0.6170257,0.47917953,0.44964105,1.0436924,1.1520001,1.3653334,2.0053334,3.1245131,2.484513,1.5458462,1.4080001,1.9790771,1.9823592,0.83035904,0.4266667,0.53825647,0.9156924,1.2865642,1.394872,1.3193847,1.1323078,1.014154,1.2340513,1.8740515,2.1300514,1.9790771,1.7427694,2.1202054,2.8127182,2.3991797,1.595077,0.93866676,0.761436,0.88287187,0.8467693,1.6738462,3.0654361,3.4100516,2.6387694,2.1169233,2.225231,2.678154,2.5107694,2.5862565,2.9013336,3.3050258,3.7382567,4.2305646,4.2863593,4.332308,4.5489235,5.077334,6.0028725,5.737026,5.398975,5.097026,4.818052,4.420923,3.9351797,3.5380516,4.4734364,5.927385,5.031385,3.1442053,2.7109745,2.1497438,1.3161026,1.5031796,2.0086155,2.048,1.6278975,1.0994873,1.1618463,0.5481026,0.29538465,0.17723078,0.09189744,0.04594872,0.06564103,0.07548718,0.059076928,0.02297436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.01969231,0.016410258,0.01969231,0.026256412,0.02297436,0.01969231,0.009846155,0.0032820515,0.0,0.0032820515,0.0032820515,0.0,0.0032820515,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.02297436,0.052512825,0.07876924,0.072205134,0.032820515,0.016410258,0.013128206,0.013128206,0.013128206,0.0032820515,0.0,0.006564103,0.016410258,0.016410258,0.009846155,0.013128206,0.016410258,0.013128206,0.0032820515,0.013128206,0.016410258,0.016410258,0.01969231,0.01969231,0.009846155,0.0032820515,0.006564103,0.013128206,0.013128206,0.013128206,0.0032820515,0.0032820515,0.009846155,0.0032820515,0.013128206,0.016410258,0.01969231,0.029538464,0.032820515,0.016410258,0.013128206,0.02297436,0.032820515,0.02297436,0.06235898,0.072205134,0.055794876,0.026256412,0.013128206,0.02297436,0.032820515,0.032820515,0.029538464,0.02297436,0.029538464,0.02297436,0.01969231,0.01969231,0.01969231,0.04266667,0.049230773,0.04594872,0.032820515,0.0,0.0032820515,0.0,0.0,0.0,0.0032820515,0.013128206,0.013128206,0.01969231,0.04594872,0.108307704,0.42338464,0.62030774,0.63343596,0.5349744,0.52512825,0.48902568,0.51856416,0.5415385,0.5349744,0.5284103,0.47261542,0.42338464,0.40697438,0.39384618,0.30194873,0.36430773,0.508718,0.65312827,0.7811283,0.9353847,0.9321026,1.0338463,1.270154,1.657436,2.2121027,2.7011285,3.1081028,3.4264617,3.636513,3.69559,3.43959,3.6069746,4.1911798,4.9493337,5.3891287,5.3727183,5.8518977,5.973334,5.47118,4.670359,4.1780515,3.7021542,3.5249233,3.4921029,3.0096412,1.7001027,0.96492314,0.6859488,0.6629744,0.6104616,0.52512825,0.56451285,0.571077,0.50543594,0.47917953,0.5415385,0.6268718,0.69579494,0.6629744,0.38728207,0.30851284,0.25928208,0.18051283,0.09189744,0.09189744,0.12143591,0.08205129,0.072205134,0.19364104,0.56123084,1.3817437,1.9922053,2.3236926,2.349949,2.100513,1.6640002,1.3095386,1.1684103,1.204513,1.1979488,1.1848207,1.3193847,1.5097437,1.6738462,1.7165129,1.7493335,1.8642052,2.097231,2.4681027,2.9801028,3.0490258,3.0720003,3.0687182,3.0326157,2.9505644,2.8356924,2.6518977,2.5009232,2.412308,2.3630772,2.1858463,2.028308,2.0053334,2.156308,2.4385643,2.2416413,2.038154,2.8160002,4.453744,5.6976414,5.8880005,5.8125134,4.893539,3.186872,1.394872,0.6826667,0.48902568,0.5349744,0.5940513,0.48902568,0.47917953,0.49230772,0.54482055,0.6465641,0.7975385,0.9616411,0.9944616,0.9747693,0.90584624,0.71548724,0.512,0.4660513,0.5218462,0.64000005,0.8041026,0.90912825,1.1716924,3.0129232,6.314667,9.412924,7.13518,5.7698464,6.5739493,9.048616,10.935796,8.979693,6.5772314,5.684513,6.8988724,9.481847,9.088,7.4830775,6.163693,5.8518977,6.491898,6.419693,6.5247183,7.177847,8.129642,8.503796,8.776206,9.449026,9.941334,10.125129,10.328616,9.4916935,8.651488,7.906462,7.39118,7.240206,7.020308,6.9743595,7.3452315,8.260923,9.731283,11.293539,12.379898,12.895181,12.983796,13.026463,13.568001,14.437745,14.91036,14.546052,13.170873,11.529847,11.529847,12.3306675,13.24636,13.761642,12.107488,10.909539,10.006975,9.734565,10.8996935,14.345847,16.443079,16.987898,15.717745,12.297847,9.757539,7.141744,4.562052,2.3762052,1.214359,1.0043077,0.8795898,0.8467693,0.9321026,1.1716924,1.4244103,1.7493335,2.03159,2.1825643,2.1169233,6.304821,6.121026,5.914257,5.398975,4.7458467,4.5554876,4.7425647,4.5029745,4.0992823,3.7316926,3.5511796,3.9417439,5.579488,6.5706673,6.3540516,5.717334,5.353026,5.1364107,4.97559,5.0051284,5.5762057,6.170257,6.3179493,6.2785645,6.1046157,5.6320004,6.294975,6.012718,5.031385,4.1156926,4.5390773,5.602462,5.910975,6.052103,6.114462,5.723898,6.009436,5.586052,5.405539,5.6352825,5.664821,4.6145644,3.757949,2.8422565,1.9364104,1.4211283,1.1684103,1.020718,0.9878975,0.98461545,0.8402052,0.8041026,0.79097444,0.7384616,0.636718,0.53825647,0.5415385,0.56451285,0.5907693,0.6170257,0.63343596,0.6498462,0.65641034,0.702359,0.74830776,0.63343596,0.3708718,0.19364104,0.108307704,0.08861539,0.06564103,0.06235898,0.059076928,0.049230773,0.029538464,0.016410258,0.02297436,0.026256412,0.02297436,0.01969231,0.01969231,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.029538464,0.03938462,0.0951795,0.108307704,0.059076928,0.0,0.0,0.0032820515,0.0032820515,0.006564103,0.029538464,0.04594872,0.07876924,0.17394873,0.3117949,0.41025645,0.43651286,0.43651286,0.512,0.56123084,0.27897438,0.41025645,0.446359,0.5152821,0.7187693,1.1355898,0.92225647,0.63343596,0.4594872,0.43651286,0.43651286,0.12471796,0.08861539,0.08861539,0.07548718,0.17723078,0.318359,0.3314872,0.23630771,0.101743594,0.049230773,0.04594872,0.049230773,0.03938462,0.036102567,0.06564103,0.026256412,0.47589746,0.8008206,0.6662565,0.006564103,0.01969231,0.036102567,0.04594872,0.052512825,0.06564103,0.10502565,0.16082053,0.16738462,0.13128206,0.11158975,0.108307704,0.108307704,0.08533334,0.059076928,0.07876924,0.06564103,0.049230773,0.026256412,0.009846155,0.029538464,0.04594872,0.0951795,0.14112821,0.13784617,0.049230773,0.052512825,0.13128206,0.190359,0.18379489,0.13784617,0.07548718,0.049230773,0.036102567,0.02297436,0.02297436,0.02297436,0.03938462,0.052512825,0.04594872,0.009846155,0.0032820515,0.049230773,0.1148718,0.15753847,0.1148718,0.08533334,0.049230773,0.026256412,0.016410258,0.009846155,0.0032820515,0.009846155,0.029538464,0.16082053,0.6268718,1.3456411,1.7066668,1.8740515,1.8543591,1.4769232,1.204513,1.1388719,1.2176411,1.211077,0.6892308,0.5349744,0.7417436,0.9517949,1.0765129,1.3226668,1.3751796,1.7427694,1.7755898,1.2898463,0.58420515,0.574359,0.46276927,0.446359,0.5349744,0.5546667,0.5874872,0.7975385,1.1881026,1.4572309,1.0043077,0.7056411,0.65641034,0.65641034,0.5907693,0.41025645,0.44964105,0.41682056,0.6498462,1.273436,2.1924105,1.1716924,0.74830776,0.79097444,1.0075898,0.9419488,0.41682056,0.24943592,0.318359,0.5513847,0.9288206,1.1946667,1.1913847,1.1979488,1.2832822,1.3226668,1.910154,2.2777438,2.100513,1.595077,1.5064616,1.9035898,1.595077,1.1454359,0.9485129,1.2012309,0.955077,1.0404103,1.6935385,2.5993848,2.858667,2.1825643,1.8084104,2.0086155,2.5796926,2.8160002,2.937436,3.1442053,3.6693337,4.585026,5.799385,4.9493337,3.945026,3.7710772,4.46359,5.10359,4.0369234,3.2787695,3.3378465,4.3618464,6.1505647,4.8016415,3.9154875,4.6605134,6.2884107,6.117744,3.0391798,1.9823592,1.4605129,0.9353847,0.82379496,0.93866676,0.9714873,0.7844103,0.48574364,0.446359,0.21661541,0.09189744,0.026256412,0.0,0.006564103,0.049230773,0.059076928,0.03938462,0.009846155,0.0,0.006564103,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.013128206,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.013128206,0.016410258,0.01969231,0.02297436,0.016410258,0.006564103,0.0032820515,0.0,0.0032820515,0.009846155,0.0032820515,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.02297436,0.036102567,0.036102567,0.016410258,0.013128206,0.013128206,0.006564103,0.016410258,0.009846155,0.01969231,0.029538464,0.029538464,0.016410258,0.0032820515,0.0032820515,0.006564103,0.0032820515,0.0,0.013128206,0.016410258,0.016410258,0.016410258,0.016410258,0.0032820515,0.006564103,0.016410258,0.02297436,0.02297436,0.016410258,0.016410258,0.016410258,0.013128206,0.009846155,0.013128206,0.016410258,0.016410258,0.01969231,0.013128206,0.006564103,0.013128206,0.016410258,0.02297436,0.049230773,0.07548718,0.059076928,0.036102567,0.02297436,0.02297436,0.052512825,0.06235898,0.06564103,0.055794876,0.006564103,0.006564103,0.006564103,0.016410258,0.02297436,0.02297436,0.04594872,0.03938462,0.026256412,0.013128206,0.0,0.0,0.006564103,0.009846155,0.013128206,0.026256412,0.04594872,0.06235898,0.06235898,0.08533334,0.23302566,0.5284103,0.6695385,0.6235898,0.47261542,0.42338464,0.39384618,0.4004103,0.4135385,0.41025645,0.38400003,0.3314872,0.4004103,0.4660513,0.446359,0.30851284,0.28882053,0.39712822,0.52512825,0.6301539,0.73517954,0.9714873,1.1290257,1.2537436,1.4309745,1.7920002,2.2678976,2.6157951,2.8225644,2.8488207,2.6190772,2.4516926,2.8750772,3.6562054,4.4800005,4.9394875,4.7950773,4.97559,4.9920006,4.716308,4.3749747,3.7087183,2.917744,2.4451284,2.3171284,2.1300514,1.8084104,1.7755898,1.8149745,1.7887181,1.6344616,1.5392822,1.4900514,1.401436,1.2603078,1.0962052,0.85005134,0.8008206,0.764718,0.5940513,0.190359,0.128,0.101743594,0.072205134,0.04266667,0.03938462,0.052512825,0.03938462,0.055794876,0.14441027,0.33805132,0.86974365,1.4178462,1.9364104,2.294154,2.2514873,1.8674873,1.4441026,1.1716924,1.0929232,1.0896411,1.273436,1.4375386,1.5392822,1.5655385,1.5327181,1.5425643,1.7624617,2.0676925,2.412308,2.8389745,3.0391798,3.1638978,3.170462,3.05559,2.8389745,2.6945643,2.546872,2.3926156,2.2449234,2.1234872,2.0644104,1.9790771,1.9364104,1.9790771,2.1103592,1.8609232,2.162872,3.7218463,6.2916927,8.651488,8.034462,6.675693,4.6933336,2.5238976,0.9353847,0.62030774,0.62030774,0.77456415,0.86974365,0.6465641,0.4955898,0.4135385,0.37415388,0.41025645,0.5907693,0.8763078,1.0469744,1.1290257,1.1060513,0.95835906,0.65969235,0.5284103,0.48574364,0.508718,0.6104616,0.8172308,0.95835906,1.6377437,2.7995899,3.7251284,3.1737437,3.501949,6.3442054,10.962052,14.276924,12.635899,9.110975,6.889026,7.318975,9.895386,8.753231,6.9021544,5.5072823,5.3005133,6.5739493,6.872616,6.961231,6.948103,6.9677954,7.204103,7.77518,8.408616,9.271795,10.377847,11.59877,11.162257,9.593436,7.9195905,6.7905645,6.442667,6.1472826,6.0258465,6.0750775,6.416411,7.3091288,8.283898,9.301334,10.016821,10.236719,9.915077,9.90195,10.994873,12.314258,13.124924,12.822975,11.096616,10.738873,10.548513,10.272821,10.57477,11.136001,11.264001,10.177642,9.3078985,12.327386,13.945437,13.200411,11.575796,9.852718,8.116513,8.218257,6.6592827,4.2469745,1.9954873,1.1552821,0.93866676,0.81066674,0.7384616,0.7384616,0.8598975,0.9616411,1.0699488,1.1684103,1.2504616,1.3062565,5.10359,4.972308,4.6539493,4.453744,4.667077,5.58277,6.5280004,6.514872,6.163693,5.7009234,4.955898,4.388103,5.221744,5.986462,6.3376417,7.066257,6.8594875,6.432821,6.1505647,6.3245134,7.181129,6.764308,6.47877,6.229334,5.917539,5.4547696,6.5083084,6.7840004,6.11118,5.0576415,4.9526157,5.7698464,5.756718,5.1626673,4.601436,5.041231,5.87159,5.3366156,5.097026,5.3792825,4.9985647,4.598154,4.0041027,3.2262566,2.487795,2.2088206,2.1169233,1.7296412,1.3095386,0.97805136,0.73517954,0.74830776,0.7975385,0.79097444,0.69579494,0.54482055,0.47589746,0.446359,0.43651286,0.43651286,0.4397949,0.49887183,0.5284103,0.58420515,0.6235898,0.5316923,0.32164106,0.15753847,0.07876924,0.068923086,0.06235898,0.04594872,0.03938462,0.036102567,0.029538464,0.009846155,0.016410258,0.02297436,0.02297436,0.01969231,0.02297436,0.016410258,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.01969231,0.009846155,0.06564103,0.108307704,0.098461546,0.029538464,0.009846155,0.0032820515,0.0,0.0032820515,0.01969231,0.029538464,0.059076928,0.15425642,0.25271797,0.16410258,0.0951795,0.128,0.24615386,0.3314872,0.18707694,0.56123084,0.7581539,0.8041026,0.77128214,0.78769237,0.45292312,0.34789747,0.37743592,0.42338464,0.3708718,0.17723078,0.30851284,0.3117949,0.12143591,0.06564103,0.055794876,0.032820515,0.013128206,0.006564103,0.0,0.006564103,0.02297436,0.032820515,0.04594872,0.068923086,0.04266667,0.5152821,0.85005134,0.69579494,0.013128206,0.036102567,0.06235898,0.072205134,0.108307704,0.27897438,0.46933338,0.48574364,0.53825647,0.65641034,0.67938465,0.5284103,0.3511795,0.21661541,0.14769232,0.128,0.12143591,0.10502565,0.08205129,0.068923086,0.07876924,0.08533334,0.13456412,0.15425642,0.1148718,0.013128206,0.06235898,0.16410258,0.21333335,0.18379489,0.108307704,0.036102567,0.029538464,0.029538464,0.01969231,0.01969231,0.049230773,0.09189744,0.10502565,0.07548718,0.032820515,0.03938462,0.128,0.23302566,0.26584616,0.10502565,0.055794876,0.032820515,0.026256412,0.026256412,0.009846155,0.006564103,0.07548718,0.20676924,0.48246157,1.0633847,1.6869745,1.5655385,1.4605129,1.4900514,1.1158975,1.0568206,1.4375386,2.0742567,2.2678976,0.8041026,0.5152821,0.77128214,0.9878975,0.9878975,0.9911796,1.0404103,1.0404103,0.955077,0.7844103,0.58420515,0.51856416,0.39384618,0.30851284,0.28225642,0.24287182,0.2855385,0.6826667,1.3883078,1.913436,1.3587693,0.7417436,0.5481026,0.53825647,0.571077,0.58092314,0.42338464,0.38728207,0.6071795,1.0010257,1.2438976,0.69251287,0.5316923,0.46276927,0.36758977,0.30851284,0.3511795,0.39056414,0.6301539,1.0568206,1.4342566,1.2898463,1.1520001,1.3259488,1.6475899,1.5163078,1.5885129,1.7066668,1.6607181,1.4342566,1.214359,1.2964103,1.3357949,1.404718,1.4834872,1.4572309,1.0502565,1.1520001,1.4769232,1.7985642,1.9429746,1.7362052,1.6836925,2.048,2.789744,3.56759,4.1813335,4.663795,5.1364107,5.651693,6.170257,5.0510774,3.9286156,3.639795,4.06318,4.1025643,3.0194874,2.3696413,2.4155898,3.5216413,6.160411,4.565334,3.6529233,3.82359,4.4767184,4.020513,1.7788719,0.8566154,0.56451285,0.44307697,0.24287182,0.1148718,0.13128206,0.17394873,0.16738462,0.098461546,0.06235898,0.03938462,0.016410258,0.0,0.006564103,0.02297436,0.029538464,0.01969231,0.0,0.0,0.006564103,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.013128206,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.026256412,0.032820515,0.013128206,0.009846155,0.013128206,0.016410258,0.009846155,0.0032820515,0.0,0.0,0.0032820515,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.006564103,0.009846155,0.01969231,0.0032820515,0.0,0.0,0.0,0.0,0.0032820515,0.01969231,0.026256412,0.026256412,0.026256412,0.016410258,0.029538464,0.055794876,0.072205134,0.059076928,0.029538464,0.013128206,0.0032820515,0.0,0.0,0.026256412,0.026256412,0.01969231,0.016410258,0.016410258,0.016410258,0.03938462,0.059076928,0.072205134,0.06235898,0.03938462,0.03938462,0.032820515,0.013128206,0.009846155,0.009846155,0.013128206,0.016410258,0.013128206,0.006564103,0.006564103,0.013128206,0.013128206,0.013128206,0.04266667,0.049230773,0.036102567,0.032820515,0.03938462,0.04266667,0.049230773,0.049230773,0.052512825,0.052512825,0.01969231,0.032820515,0.026256412,0.02297436,0.02297436,0.02297436,0.032820515,0.02297436,0.01969231,0.02297436,0.02297436,0.013128206,0.013128206,0.013128206,0.016410258,0.04594872,0.06564103,0.101743594,0.12143591,0.13784617,0.21989745,0.37743592,0.508718,0.52512825,0.43651286,0.3708718,0.34133336,0.27897438,0.23630771,0.23630771,0.24943592,0.26912823,0.38400003,0.47261542,0.46276927,0.3446154,0.29210258,0.380718,0.5218462,0.6826667,0.892718,1.1454359,1.2603078,1.3686155,1.6180514,2.162872,1.8838975,1.9790771,2.2383592,2.5107694,2.7109745,2.540308,2.8225644,3.1573336,3.367385,3.501949,3.4067695,3.255795,3.2295387,3.3542566,3.4789746,2.934154,2.294154,2.0611284,2.3991797,3.1245131,3.3214362,3.7087183,4.0467696,4.0533338,3.4100516,3.1113849,2.740513,2.3171284,1.8740515,1.4572309,1.0535386,0.78769237,0.6662565,0.5677949,0.28225642,0.14769232,0.16738462,0.17394873,0.13128206,0.12471796,0.128,0.12471796,0.14441027,0.16738462,0.15097436,0.3708718,0.6892308,1.0994873,1.4933335,1.6607181,1.5556924,1.2865642,1.0502565,0.9517949,1.0043077,1.2635899,1.529436,1.7329233,1.8346668,1.847795,1.8281027,1.9265642,2.0906668,2.3105643,2.6354873,3.0391798,3.3805132,3.5314875,3.442872,3.1606157,2.9210258,2.6354873,2.2908719,1.9823592,1.9035898,1.8149745,1.8674873,1.910154,1.847795,1.6410258,1.404718,2.0775387,3.446154,5.1922054,6.8627696,6.245744,5.024821,3.373949,1.7165129,0.7253334,0.702359,0.8369231,1.0075898,1.079795,0.92225647,0.69251287,0.512,0.39056414,0.36758977,0.512,0.79097444,0.97805136,1.0732309,1.0929232,1.0633847,0.73517954,0.58420515,0.512,0.48902568,0.5481026,0.7811283,0.83035904,0.7089231,0.52512825,0.49887183,0.93866676,2.1070771,5.5105643,10.765129,15.599591,15.701335,12.370052,8.448001,6.2523084,7.571693,7.50277,7.026872,6.8004107,7.397744,9.301334,11.565949,10.354873,8.234667,6.8332314,6.8463597,7.8834877,8.12636,8.713847,10.000411,11.546257,11.851488,10.834052,9.399796,8.113232,7.210667,6.9120007,6.705231,6.3245134,5.786257,5.398975,5.684513,6.416411,7.509334,8.533334,8.707283,8.874667,9.941334,11.273847,12.2387705,12.189539,10.673231,9.91836,9.074872,8.132924,7.9195905,8.4972315,8.618668,8.096821,8.687591,14.102976,15.248411,13.6237955,11.831796,10.246565,7.02359,6.8529234,5.474462,3.4888208,1.7001027,1.1323078,1.0502565,0.92225647,0.7844103,0.6826667,0.67610264,0.7318975,0.7450257,0.7450257,0.761436,0.8172308,4.3027697,4.3552823,4.3585644,4.923077,6.124308,7.496206,8.503796,8.740103,8.897642,8.999385,8.418462,6.518154,5.142975,4.8082056,5.684513,7.5979495,7.4863596,7.2270775,7.282872,7.8473854,8.835282,8.172308,7.958975,7.6635904,6.9842057,5.8486156,5.720616,6.1078978,6.193231,5.8125134,5.4580517,5.159385,4.9099493,4.2601027,3.5872824,4.0992823,4.2436924,3.639795,3.3772311,3.387077,2.4648206,2.6945643,2.7963078,2.8291285,2.9046156,3.190154,3.318154,2.678154,1.7657437,0.9944616,0.6826667,0.71548724,0.8008206,0.77456415,0.61374366,0.45292312,0.38728207,0.36430773,0.380718,0.41025645,0.4135385,0.40697438,0.39712822,0.38400003,0.37743592,0.39712822,0.32164106,0.23302566,0.15753847,0.10502565,0.08861539,0.07548718,0.049230773,0.029538464,0.016410258,0.0032820515,0.0,0.0032820515,0.0032820515,0.0032820515,0.013128206,0.013128206,0.013128206,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.0,0.0,0.032820515,0.08205129,0.06564103,0.026256412,0.013128206,0.006564103,0.009846155,0.032820515,0.06235898,0.10502565,0.17723078,0.23302566,0.15097436,0.059076928,0.04266667,0.07876924,0.14112821,0.19692309,0.5415385,0.8369231,0.88287187,0.6465641,0.27241027,0.17394873,0.23958977,0.2297436,0.10502565,0.03938462,0.3117949,0.79097444,0.74830776,0.23630771,0.06564103,0.026256412,0.016410258,0.013128206,0.0032820515,0.0,0.0032820515,0.02297436,0.036102567,0.04266667,0.04266667,0.0951795,0.29210258,0.4660513,0.5021539,0.3446154,0.21333335,0.2100513,0.20348719,0.23630771,0.5415385,1.1158975,1.4408206,1.5786668,1.6410258,1.7723079,1.3915899,0.88943595,0.512,0.32164106,0.2100513,0.23630771,0.2855385,0.3249231,0.2986667,0.16738462,0.13784617,0.15425642,0.15097436,0.108307704,0.052512825,0.101743594,0.128,0.11158975,0.06235898,0.013128206,0.0032820515,0.0,0.006564103,0.01969231,0.02297436,0.10502565,0.19692309,0.19364104,0.1148718,0.098461546,0.14769232,0.2297436,0.29210258,0.256,0.029538464,0.009846155,0.013128206,0.032820515,0.049230773,0.052512825,0.14112821,0.508718,0.8041026,0.9682052,1.2242053,1.4112822,0.81066674,0.35774362,0.35774362,0.4955898,1.3522053,2.5993848,3.370667,2.9801028,0.90584624,0.49887183,0.61374366,0.7450257,0.65312827,0.34789747,0.3052308,0.30194873,0.36758977,0.4955898,0.62030774,0.46276927,0.3052308,0.21333335,0.19692309,0.19364104,0.3249231,1.0666667,1.9035898,2.284308,1.6016412,0.7811283,0.41682056,0.30194873,0.36102566,0.6465641,0.55794877,0.6301539,0.8402052,0.97805136,0.6432821,0.512,0.44307697,0.38728207,0.3511795,0.37415388,0.5907693,0.8402052,1.3751796,2.0578463,2.3466668,1.6344616,1.2471796,1.4408206,1.9462565,1.9626669,1.5983591,1.4145643,1.4375386,1.5721027,1.595077,1.785436,2.0118976,2.103795,1.8806155,1.1815386,0.95835906,0.9321026,1.020718,1.1618463,1.3029745,1.5195899,1.6836925,2.162872,3.0687182,4.273231,5.3234878,5.8814363,5.7731285,5.172513,4.57518,4.0041027,3.3444104,2.806154,2.4352822,2.1464617,2.3762052,2.4484105,2.1891284,2.1398976,3.5511796,2.7142565,2.284308,1.9692309,1.3718976,0.0,0.006564103,0.006564103,0.0032820515,0.0032820515,0.013128206,0.032820515,0.013128206,0.009846155,0.029538464,0.052512825,0.04594872,0.036102567,0.029538464,0.026256412,0.026256412,0.006564103,0.006564103,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.026256412,0.049230773,0.049230773,0.009846155,0.0,0.0032820515,0.006564103,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.02297436,0.032820515,0.049230773,0.072205134,0.032820515,0.016410258,0.006564103,0.0032820515,0.0,0.009846155,0.029538464,0.049230773,0.06564103,0.068923086,0.029538464,0.029538464,0.06564103,0.108307704,0.10502565,0.06235898,0.029538464,0.013128206,0.013128206,0.013128206,0.04266667,0.032820515,0.02297436,0.02297436,0.02297436,0.04266667,0.07548718,0.108307704,0.12143591,0.108307704,0.07548718,0.06564103,0.049230773,0.02297436,0.009846155,0.013128206,0.01969231,0.02297436,0.01969231,0.016410258,0.026256412,0.032820515,0.049230773,0.072205134,0.08205129,0.04594872,0.052512825,0.072205134,0.08205129,0.06235898,0.029538464,0.016410258,0.013128206,0.01969231,0.036102567,0.06564103,0.04266667,0.01969231,0.01969231,0.029538464,0.02297436,0.016410258,0.029538464,0.049230773,0.052512825,0.029538464,0.01969231,0.016410258,0.026256412,0.06564103,0.06564103,0.11158975,0.15425642,0.15425642,0.09189744,0.10502565,0.24615386,0.37415388,0.4004103,0.28225642,0.3314872,0.27569234,0.18379489,0.128,0.18379489,0.28882053,0.36102566,0.41025645,0.4135385,0.32820517,0.30194873,0.3708718,0.51856416,0.7515898,1.0929232,1.086359,1.0962052,1.3554872,1.9429746,2.7798977,1.6705642,1.4408206,1.7755898,2.3138463,2.674872,2.4713848,2.665026,2.7175386,2.5271797,2.4385643,2.3401027,1.9561027,1.8543591,2.1202054,2.356513,2.176,1.9954873,2.2153847,3.1015387,4.7950773,4.965744,5.349744,5.789539,5.85518,4.850872,4.2305646,3.5052311,2.7602053,2.0873847,1.5655385,1.2931283,0.9124103,0.7581539,0.83035904,0.78769237,0.6071795,0.69579494,0.69251287,0.54482055,0.5316923,0.48574364,0.4266667,0.36758977,0.28225642,0.09189744,0.16410258,0.21989745,0.28882053,0.42338464,0.702359,0.8566154,0.83035904,0.76800007,0.77456415,0.92553854,1.211077,1.7132308,2.1267693,2.3138463,2.3236926,2.1924105,2.0644104,2.048,2.2055387,2.537026,3.0523078,3.570872,3.882667,3.9023592,3.6562054,3.2918978,2.793026,2.2547693,1.8707694,1.9364104,1.7624617,1.9035898,2.0217438,1.8838975,1.3587693,1.1191796,1.5885129,1.9692309,1.9790771,1.8773335,1.9200002,1.9626669,1.719795,1.2307693,0.86317956,0.88943595,1.0962052,1.2800001,1.3620514,1.3817437,1.1618463,0.86646163,0.60061544,0.4397949,0.43651286,0.6170257,0.7450257,0.8369231,0.90256417,0.97805136,0.7515898,0.64000005,0.574359,0.54482055,0.6104616,0.80738467,0.77128214,0.64000005,0.55794877,0.6465641,0.86317956,1.5130258,3.6529233,7.4141545,11.979488,14.257232,13.111795,9.189744,4.778667,3.8071797,5.677949,7.3583593,8.858257,10.459898,12.704822,16.83036,14.080001,10.098872,8.044309,8.576,10.617436,10.33518,9.898667,10.266257,11.201642,11.378873,10.712616,9.813334,8.907488,7.8539495,7.6143594,7.4174366,6.7807183,5.664821,4.453744,4.6244106,5.1626673,6.498462,8.27077,9.337437,10.466462,11.119591,11.467488,11.533129,11.188514,10.171078,9.370257,8.766359,8.2445135,7.571693,6.948103,7.059693,7.2927184,8.605539,13.51877,15.386257,15.284514,15.27795,14.378668,8.572719,6.226052,4.6966157,3.4198978,2.228513,1.3686155,1.3128207,1.1093334,0.88287187,0.7089231,0.63343596,0.6629744,0.65969235,0.64000005,0.63343596,0.6662565,6.012718,6.0356927,6.2818465,6.6395903,6.885744,6.6527185,6.616616,7.5585647,9.586872,12.498053,15.793232,14.388514,13.167591,11.83836,10.295795,8.635077,8.513641,7.9163084,7.000616,6.11118,5.7829747,6.8562055,8.03118,8.802463,8.717129,7.4010262,6.6067696,6.675693,6.3376417,5.5565133,5.5072823,4.9362054,4.096,3.2164104,2.5731285,2.487795,3.4133337,3.8498464,3.9154875,3.8695388,4.089436,4.2601027,3.314872,2.5928206,2.6026669,3.006359,3.114667,2.9604106,2.484513,1.782154,1.0994873,0.76800007,0.71548724,0.67610264,0.574359,0.48902568,0.40369233,0.3249231,0.30851284,0.35446155,0.4266667,0.39056414,0.3446154,0.3249231,0.3708718,0.51856416,0.48246157,0.4266667,0.36102566,0.28225642,0.19692309,0.12471796,0.07876924,0.049230773,0.026256412,0.016410258,0.0032820515,0.009846155,0.016410258,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.01969231,0.029538464,0.006564103,0.0,0.0,0.0032820515,0.016410258,0.026256412,0.03938462,0.032820515,0.04594872,0.16738462,0.21661541,0.18379489,0.15753847,0.2100513,0.380718,0.12471796,0.02297436,0.055794876,0.17394873,0.32164106,0.3314872,0.46276927,0.54482055,0.5152821,0.44307697,0.44307697,0.5973334,0.4955898,0.16082053,0.07548718,0.5152821,0.90912825,0.6826667,0.052512825,0.016410258,0.06564103,0.08533334,0.06564103,0.02297436,0.0,0.013128206,0.032820515,0.06564103,0.10502565,0.15097436,0.3249231,0.8795898,1.4966155,1.847795,1.6016412,0.69907695,0.48246157,0.4135385,0.28225642,0.19692309,1.2242053,2.92759,3.1343591,2.1398976,2.7011285,2.4549747,1.8642052,1.211077,0.67282057,0.32164106,0.44307697,0.7384616,0.94523084,0.8402052,0.2297436,0.18051283,0.13128206,0.11158975,0.12471796,0.13784617,0.101743594,0.04594872,0.009846155,0.0,0.0,0.0,0.0,0.036102567,0.0951795,0.108307704,0.2297436,0.36102566,0.3708718,0.28225642,0.24287182,0.34133336,0.32164106,0.18707694,0.029538464,0.029538464,0.01969231,0.032820515,0.07548718,0.15097436,0.25928208,0.6629744,1.7887181,2.0250258,1.1520001,0.32164106,0.5284103,0.45292312,0.28225642,0.21333335,0.45620516,1.9232821,3.5971284,2.986667,0.67610264,0.32164106,0.380718,0.37743592,0.26256412,0.1148718,0.15097436,0.029538464,0.036102567,0.08533334,0.15425642,0.28882053,0.5349744,0.40369233,0.318359,0.4135385,0.5349744,0.571077,1.0010257,1.2340513,1.0765129,0.74830776,0.60061544,0.67282057,0.6629744,0.49887183,0.36758977,0.7450257,1.020718,0.88287187,0.5218462,0.65641034,0.6301539,0.5874872,0.56451285,0.55794877,0.5349744,1.1684103,1.7591796,2.2153847,2.481231,2.5173335,2.225231,1.6213335,1.6147693,2.3040001,2.9768207,3.1573336,3.3608208,2.986667,2.2678976,2.2416413,2.6584618,2.8914874,2.5042052,1.7558975,1.5721027,1.2406155,0.9682052,0.827077,0.8992821,1.2668719,1.4244103,1.5392822,1.8248206,2.4549747,3.5413337,4.5522056,4.6605134,4.3716927,4.0369234,3.8301542,3.511795,2.8389745,2.1366155,1.7296412,1.9364104,2.4024618,2.4910772,2.294154,1.8445129,1.0994873,0.574359,0.29538465,0.13128206,0.02297436,0.0,0.036102567,0.036102567,0.01969231,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.026256412,0.10502565,0.14769232,0.12471796,0.07548718,0.016410258,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.026256412,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.026256412,0.059076928,0.108307704,0.15753847,0.18379489,0.13456412,0.07548718,0.032820515,0.013128206,0.0,0.0,0.009846155,0.03938462,0.0951795,0.16738462,0.059076928,0.049230773,0.06235898,0.055794876,0.029538464,0.01969231,0.006564103,0.029538464,0.072205134,0.06235898,0.013128206,0.0,0.01969231,0.049230773,0.06235898,0.049230773,0.055794876,0.06564103,0.08533334,0.12143591,0.098461546,0.08205129,0.068923086,0.059076928,0.04594872,0.059076928,0.06235898,0.055794876,0.03938462,0.016410258,0.07548718,0.101743594,0.18051283,0.30194873,0.3511795,0.16738462,0.12143591,0.12143591,0.108307704,0.06235898,0.049230773,0.055794876,0.04266667,0.013128206,0.0,0.0,0.0,0.006564103,0.029538464,0.09189744,0.055794876,0.026256412,0.009846155,0.0032820515,0.016410258,0.0032820515,0.009846155,0.03938462,0.08861539,0.13784617,0.08861539,0.0951795,0.08861539,0.06564103,0.09189744,0.20020515,0.30194873,0.5349744,0.761436,0.56451285,0.56451285,0.6301539,0.50543594,0.256,0.24287182,0.28225642,0.30851284,0.30851284,0.29210258,0.3052308,0.26912823,0.3052308,0.41025645,0.54482055,0.64000005,0.65312827,0.53825647,0.64000005,0.99774367,1.3292309,1.4506668,1.0962052,1.1454359,1.723077,2.2121027,2.0184617,2.0217438,2.0184617,1.9364104,1.8773335,1.6804104,1.5130258,1.4703591,1.5622566,1.7099489,1.6344616,1.3883078,1.3587693,1.719795,2.425436,3.2328207,3.6069746,3.6332312,3.5347695,3.692308,3.373949,2.8849232,2.4155898,2.1267693,2.1530259,2.1136413,1.8871796,1.6246156,1.4572309,1.4966155,1.7165129,1.8609232,1.7887181,1.5688206,1.4966155,1.1782565,0.92553854,0.67938465,0.4201026,0.15097436,0.22646156,0.20676924,0.18379489,0.20020515,0.27569234,0.41025645,0.5349744,0.55794877,0.54482055,0.7187693,1.3161026,2.1956925,2.6486156,2.5304618,2.2744617,2.0644104,2.0151796,2.1070771,2.3171284,2.609231,2.9997952,3.2820516,3.4264617,3.436308,3.3280003,2.9735386,2.5993848,2.2777438,2.0611284,1.9987694,2.2908719,2.228513,1.9659488,1.5655385,0.9911796,0.6268718,0.44307697,0.380718,0.4135385,0.5349744,0.98461545,1.3357949,1.4408206,1.2668719,0.8992821,0.9747693,1.3029745,1.7427694,2.0906668,2.0906668,1.8215386,1.3981539,0.92225647,0.5218462,0.3511795,0.37415388,0.62030774,0.86974365,1.017436,1.0535386,1.1257436,0.9156924,0.6826667,0.5874872,0.67282057,0.8795898,0.7844103,0.7056411,0.76800007,0.9156924,1.024,1.3456411,2.3171284,3.446154,3.31159,5.717334,7.4174366,7.752206,6.49518,3.8465643,4.210872,5.346462,6.7938466,8.5661545,11.155693,11.178667,9.334154,8.083693,8.930462,12.419283,16.278976,15.593027,14.28677,14.10954,14.631386,12.386462,8.868103,6.439385,5.7042055,5.5072823,5.2020516,4.7622566,4.069744,3.4264617,3.5249233,3.95159,4.3716927,5.156103,6.3245134,7.506052,10.072617,11.506873,11.812103,11.188514,10.039796,8.917334,8.379078,8.228104,8.205129,8.011488,9.242257,14.513232,14.972719,10.259693,8.513641,9.685334,9.82318,9.245539,8.195283,6.8529234,6.449231,6.51159,5.8518977,4.276513,2.5796926,1.7001027,1.1323078,0.7975385,0.63343596,0.6104616,0.65969235,0.6071795,0.5415385,0.4955898,0.45620516,7.893334,7.6734366,8.198565,8.740103,8.868103,8.457847,7.397744,6.7150774,6.6527185,7.2237954,8.224821,8.500513,8.835282,9.77395,11.208206,12.370052,13.010053,13.210258,12.924719,12.166565,11.008,10.256411,9.764103,9.504821,9.321027,8.937026,7.207385,6.0816417,5.349744,4.9296412,4.8607183,4.8738465,4.818052,4.529231,3.9417439,3.0851285,3.495385,4.0041027,4.4373336,4.7425647,4.9788723,4.896821,4.2896414,3.6824617,3.239385,2.7634873,2.930872,3.0687182,2.7044106,1.9265642,1.3784616,1.0305642,0.7450257,0.50543594,0.36758977,0.4266667,0.44964105,0.43651286,0.40697438,0.37743592,0.35446155,0.35774362,0.35774362,0.37743592,0.42994875,0.50543594,0.57764107,0.6235898,0.574359,0.4397949,0.29538465,0.17394873,0.07876924,0.032820515,0.032820515,0.03938462,0.026256412,0.013128206,0.006564103,0.013128206,0.013128206,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.0,0.0,0.0,0.0,0.0032820515,0.07548718,0.09189744,0.08861539,0.08861539,0.14441027,0.12471796,0.08205129,0.04594872,0.04594872,0.101743594,0.128,0.08205129,0.16082053,0.34789747,0.40697438,0.17394873,0.19364104,0.3249231,0.446359,0.44307697,0.38400003,0.34133336,0.26584616,0.190359,0.2231795,0.9156924,1.2931283,1.0568206,0.63343596,1.1618463,1.0732309,0.7975385,0.46276927,0.18707694,0.08533334,0.029538464,0.013128206,0.013128206,0.02297436,0.04266667,0.10502565,0.6498462,1.0699488,1.3062565,1.8346668,2.1234872,1.3981539,1.585231,2.546872,2.0906668,1.3489232,1.020718,0.7187693,0.4397949,0.5513847,0.5021539,0.37743592,0.25271797,0.17723078,0.18707694,0.4266667,0.52512825,0.52512825,0.46933338,0.37415388,0.44307697,0.50543594,0.45292312,0.27897438,0.07548718,0.029538464,0.009846155,0.029538464,0.15753847,0.49887183,0.7844103,0.7811283,0.71548724,0.636718,0.42338464,0.28225642,0.2231795,0.2100513,0.28225642,0.53825647,0.5677949,0.43323082,0.21661541,0.036102567,0.055794876,0.26584616,0.49887183,0.6104616,0.5415385,0.32164106,0.4594872,0.5677949,0.6695385,0.67610264,0.39384618,0.20020515,0.14769232,0.446359,1.0075898,1.4473847,1.3193847,1.214359,0.82379496,0.26256412,0.06564103,0.07548718,0.20020515,0.17723078,0.02297436,0.029538464,0.10502565,0.18707694,0.27241027,0.34133336,0.38728207,0.37743592,0.35774362,0.3511795,0.40697438,0.6071795,1.5819489,1.9298463,1.6705642,1.0699488,0.6629744,0.6826667,0.5907693,0.54482055,0.5349744,0.39056414,0.60389745,1.014154,1.3029745,1.3128207,1.0469744,0.8467693,0.7811283,0.88287187,1.2012309,1.7920002,1.9954873,1.9790771,2.172718,2.9144619,4.4340515,3.2918978,2.7470772,2.6617439,2.8947694,3.2918978,3.9647183,4.20759,3.7907696,3.131077,3.2918978,4.010667,4.0533338,3.4494362,2.5961027,2.2547693,2.041436,1.8576412,1.6902566,1.7362052,2.3762052,1.9692309,1.6246156,1.6246156,2.0151796,2.612513,2.169436,1.9364104,1.7985642,1.6607181,1.4244103,1.0896411,0.892718,0.7515898,0.764718,1.204513,0.9944616,0.75487185,0.55794877,0.41025645,0.23302566,0.118153855,0.07548718,0.04594872,0.013128206,0.0,0.006564103,0.006564103,0.009846155,0.009846155,0.0,0.0,0.006564103,0.006564103,0.0,0.0032820515,0.006564103,0.029538464,0.04594872,0.049230773,0.03938462,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.01969231,0.01969231,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.02297436,0.02297436,0.013128206,0.01969231,0.02297436,0.016410258,0.016410258,0.0032820515,0.0,0.0032820515,0.009846155,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.016410258,0.03938462,0.11158975,0.2231795,0.318359,0.318359,0.256,0.16082053,0.072205134,0.06235898,0.09189744,0.049230773,0.01969231,0.029538464,0.032820515,0.02297436,0.036102567,0.052512825,0.059076928,0.055794876,0.06235898,0.03938462,0.029538464,0.04266667,0.06235898,0.02297436,0.026256412,0.03938462,0.04266667,0.036102567,0.04266667,0.032820515,0.026256412,0.032820515,0.049230773,0.04266667,0.055794876,0.06235898,0.068923086,0.108307704,0.108307704,0.0951795,0.06564103,0.04594872,0.101743594,0.11158975,0.12471796,0.13456412,0.16738462,0.26584616,0.20020515,0.15425642,0.098461546,0.052512825,0.072205134,0.09189744,0.07548718,0.049230773,0.02297436,0.013128206,0.013128206,0.01969231,0.026256412,0.029538464,0.029538464,0.02297436,0.016410258,0.029538464,0.052512825,0.06564103,0.072205134,0.052512825,0.049230773,0.06564103,0.06564103,0.101743594,0.13784617,0.18051283,0.21989745,0.22646156,0.33476925,0.3117949,0.25928208,0.21661541,0.13784617,0.14769232,0.16082053,0.13456412,0.07876924,0.08533334,0.08205129,0.09189744,0.101743594,0.108307704,0.108307704,0.24943592,0.5481026,0.67282057,0.5874872,0.5677949,0.86317956,1.014154,1.0305642,0.9911796,1.0469744,0.98461545,0.8763078,0.88943595,1.0896411,1.4309745,1.273436,1.2537436,1.4145643,1.7099489,1.9987694,1.8215386,1.6311796,1.401436,1.1848207,1.086359,1.1979488,0.88943595,0.764718,0.9878975,1.2668719,1.585231,1.785436,1.7362052,1.5655385,1.6672822,1.5721027,1.5031796,1.522872,1.7526156,2.3827693,2.865231,2.9997952,2.9997952,3.114667,3.620103,3.6036925,3.5840003,3.367385,2.9833848,2.6683078,2.2514873,1.6902566,1.0994873,0.5874872,0.24943592,0.22646156,0.24943592,0.26912823,0.28225642,0.33476925,0.46933338,0.7187693,0.93866676,1.079795,1.1815386,1.6410258,2.176,2.5961027,2.7798977,2.6518977,2.4155898,2.481231,2.737231,3.0687182,3.3411283,3.2820516,3.4067695,3.508513,3.4658465,3.2295387,2.8849232,2.6157951,2.477949,2.3958976,2.156308,2.0611284,1.7165129,1.4998976,1.3817437,0.90584624,0.5021539,0.36102566,0.3314872,0.3314872,0.3249231,0.45620516,0.69579494,0.9288206,1.017436,0.827077,0.764718,0.96492314,1.3259488,1.7132308,1.9692309,1.847795,1.6475899,1.3489232,0.9944616,0.7187693,0.6826667,0.86974365,1.0404103,1.1224617,1.1979488,1.204513,1.0994873,0.90912825,0.69907695,0.6104616,0.61374366,0.6432821,0.69579494,0.78769237,0.96492314,1.4342566,2.7995899,4.5456414,6.1505647,7.069539,8.470975,10.607591,11.490462,10.679795,9.288206,4.8705645,3.249231,3.242667,4.466872,7.3583593,10.47959,12.73436,15.192616,18.22195,21.477745,21.710772,18.326975,13.784616,10.525539,10.971898,11.605334,12.022155,12.455385,12.977232,13.515489,13.062565,11.506873,9.235693,6.6002054,3.9154875,3.8334363,4.125539,4.4701543,4.8836927,5.737026,7.4010262,8.828718,9.616411,9.7903595,9.796924,9.521232,8.165744,6.8693337,6.2588725,6.422975,6.6034875,7.0104623,6.633026,6.3376417,8.868103,13.974976,12.86236,10.266257,8.503796,7.4732313,5.937231,5.1200004,4.3027697,3.259077,2.2383592,1.463795,1.020718,0.77128214,0.6432821,0.5973334,0.5973334,0.56451285,0.5152821,0.46933338,0.43323082,7.207385,7.1844106,7.9130263,8.6580515,9.094564,9.284924,8.628513,7.712821,6.997334,6.6034875,6.340924,6.114462,5.920821,6.2720003,7.4075904,9.29477,10.732308,12.130463,13.128206,13.348104,12.406155,12.347078,11.293539,9.9282055,8.720411,7.9130263,6.7249236,5.717334,5.0215387,4.630975,4.4340515,4.585026,4.844308,4.670359,3.9811285,3.1540515,3.5282054,4.3618464,4.890257,5.031385,5.3760004,4.850872,4.0336413,3.3444104,2.8750772,2.3991797,2.0841026,1.9462565,1.7001027,1.3587693,1.211077,0.8730257,0.6629744,0.53825647,0.47261542,0.4660513,0.58092314,0.60061544,0.5677949,0.512,0.45620516,0.45292312,0.49230772,0.5349744,0.56451285,0.5940513,0.62030774,0.63343596,0.57764107,0.4594872,0.32820517,0.2100513,0.118153855,0.06564103,0.04594872,0.036102567,0.02297436,0.013128206,0.02297436,0.049230773,0.07876924,0.036102567,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.04594872,0.016410258,0.0032820515,0.0,0.0032820515,0.009846155,0.08861539,0.108307704,0.09189744,0.072205134,0.06564103,0.04266667,0.026256412,0.01969231,0.01969231,0.029538464,0.068923086,0.07548718,0.16082053,0.36430773,0.6301539,0.5546667,0.3314872,0.2855385,0.4135385,0.39712822,0.50543594,0.61374366,0.5874872,0.5940513,1.1093334,1.6246156,1.6836925,1.3686155,1.083077,1.5425643,0.8992821,0.571077,0.5316923,0.6662565,0.79425645,0.23630771,0.055794876,0.08205129,0.17066668,0.19692309,0.06564103,0.25271797,0.6235898,1.0075898,1.1782565,1.1355898,0.7089231,0.827077,1.3554872,1.0994873,0.60389745,0.29210258,0.18707694,0.18707694,0.068923086,0.06235898,0.08533334,0.108307704,0.1148718,0.08861539,0.22646156,0.25271797,0.23958977,0.24287182,0.29210258,0.28882053,0.2855385,0.23630771,0.13456412,0.02297436,0.01969231,0.036102567,0.13456412,0.318359,0.52512825,0.6071795,0.5415385,0.47261542,0.42338464,0.30194873,0.20348719,0.15753847,0.17066668,0.28882053,0.62030774,0.5152821,0.3446154,0.23302566,0.3052308,0.7122052,0.9517949,0.9944616,0.8763078,0.65312827,0.39056414,0.3314872,0.3511795,0.5316923,0.80738467,0.9616411,0.8369231,1.2274873,1.8313848,2.2153847,1.8313848,0.90256417,0.48246157,0.41025645,0.49230772,0.5021539,0.7515898,0.9747693,0.6629744,0.059076928,0.14769232,0.23302566,0.30851284,0.36430773,0.3708718,0.28225642,0.3708718,0.3511795,0.31507695,0.37743592,0.6629744,1.9659488,1.8248206,1.4145643,1.394872,1.913436,2.5238976,1.9035898,1.1520001,0.7187693,0.38728207,0.45620516,0.6826667,1.1027694,1.4244103,1.0436924,0.83035904,0.892718,1.1782565,1.5983591,2.041436,2.556718,2.7798977,3.1376412,4.1846156,6.5969234,4.6802053,3.6332312,3.308308,3.5774362,4.325744,5.0084105,4.7556925,4.066462,3.4297438,3.3345644,3.7120004,3.9286156,3.626667,3.2000003,3.7809234,4.1682053,3.4067695,2.4385643,2.0250258,2.7175386,2.8717952,2.7437952,2.4910772,2.172718,1.7394873,1.1027694,0.85005134,0.80738467,0.8041026,0.6695385,0.42994875,0.30851284,0.23958977,0.24943592,0.43651286,0.26912823,0.13128206,0.049230773,0.01969231,0.006564103,0.0,0.006564103,0.013128206,0.013128206,0.009846155,0.0032820515,0.0,0.0032820515,0.006564103,0.009846155,0.009846155,0.006564103,0.0032820515,0.0,0.0,0.0,0.0032820515,0.009846155,0.013128206,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.01969231,0.016410258,0.0032820515,0.0,0.0,0.006564103,0.006564103,0.0032820515,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.01969231,0.01969231,0.01969231,0.02297436,0.029538464,0.02297436,0.029538464,0.04266667,0.04594872,0.03938462,0.02297436,0.013128206,0.009846155,0.026256412,0.049230773,0.036102567,0.029538464,0.02297436,0.013128206,0.009846155,0.016410258,0.006564103,0.013128206,0.052512825,0.118153855,0.17723078,0.23958977,0.36758977,0.40697438,0.31507695,0.14112821,0.14769232,0.15097436,0.12471796,0.06235898,0.0,0.013128206,0.06564103,0.11158975,0.1148718,0.07876924,0.049230773,0.029538464,0.026256412,0.036102567,0.052512825,0.04594872,0.04594872,0.055794876,0.068923086,0.049230773,0.032820515,0.026256412,0.03938462,0.055794876,0.029538464,0.03938462,0.052512825,0.068923086,0.07548718,0.06564103,0.059076928,0.06235898,0.068923086,0.08861539,0.14112821,0.12471796,0.12143591,0.128,0.15097436,0.18051283,0.15097436,0.15097436,0.12471796,0.08205129,0.11158975,0.101743594,0.06564103,0.029538464,0.013128206,0.016410258,0.02297436,0.032820515,0.03938462,0.032820515,0.006564103,0.006564103,0.006564103,0.01969231,0.049230773,0.06564103,0.0951795,0.11158975,0.108307704,0.08533334,0.072205134,0.11158975,0.13456412,0.17394873,0.21989745,0.21333335,0.21989745,0.17723078,0.12471796,0.08533334,0.06564103,0.06564103,0.059076928,0.04266667,0.026256412,0.04594872,0.06235898,0.07548718,0.068923086,0.059076928,0.08861539,0.3446154,0.5907693,0.69907695,0.65312827,0.5677949,0.8533334,1.2176411,1.3259488,1.1158975,0.8041026,0.955077,1.1191796,1.3423591,1.5721027,1.6672822,1.5622566,1.6902566,2.1136413,2.6551797,2.8717952,2.6289232,2.3171284,2.176,2.0939488,1.6344616,1.2668719,1.0010257,1.2603078,1.8543591,1.975795,2.0020514,1.9200002,1.6902566,1.467077,1.5819489,1.5163078,1.5556924,2.0118976,2.8882053,3.889231,3.9844105,4.023795,4.0467696,4.1780515,4.6276927,4.604718,4.2240005,3.636513,2.986667,2.412308,1.9495386,1.4309745,0.9419488,0.571077,0.38400003,0.29210258,0.26912823,0.2986667,0.36758977,0.48902568,0.5874872,0.77456415,1.0305642,1.3357949,1.6902566,2.0578463,2.4943593,2.8816411,3.0851285,2.9571285,2.7634873,2.9604106,3.3444104,3.7218463,3.9187696,3.6890259,3.6168208,3.6594875,3.6069746,3.0654361,2.5862565,2.3269746,2.2055387,2.1398976,2.0512822,2.156308,2.0742567,1.8838975,1.5130258,0.74830776,0.44307697,0.3446154,0.32164106,0.2986667,0.24615386,0.26584616,0.380718,0.51856416,0.6104616,0.58092314,0.60061544,0.71548724,0.97805136,1.3489232,1.6738462,1.8871796,2.041436,1.8937438,1.4703591,1.0469744,0.80738467,0.88615394,1.0666667,1.1881026,1.1716924,0.9485129,0.7975385,0.7056411,0.65641034,0.6301539,0.56123084,0.6498462,0.84348726,1.1290257,1.5261539,2.3794873,3.8859491,5.805949,7.64718,8.631796,9.7214365,12.310975,13.748514,13.147899,11.401847,6.941539,3.9614363,2.7569232,3.436308,5.904411,10.443488,15.527386,20.417643,24.12636,25.4359,22.554258,18.730669,14.306462,10.410667,8.992821,9.938052,11.257437,11.936821,11.529847,10.161232,9.6525135,9.104411,8.2904625,7.0400004,5.2381544,4.7983594,4.086154,3.6004105,3.6758976,4.4898467,6.0685134,7.3550773,8.132924,8.457847,8.65477,8.43159,7.351795,6.0750775,5.3924108,6.229334,9.291488,9.321027,7.2960005,5.3727183,6.87918,12.934566,13.24636,11.280411,9.222565,7.9786673,6.2523084,4.4898467,3.0982566,2.2449234,1.8674873,1.4080001,1.1749744,0.94523084,0.69251287,0.5874872,0.5973334,0.65969235,0.6629744,0.5874872,0.49230772,7.9819493,8.04759,8.293744,8.257642,7.9491286,7.8769236,8.208411,7.8736415,7.53559,7.568411,8.044309,8.021334,7.315693,6.5083084,6.0980515,6.5017443,6.8266673,8.516924,10.328616,11.385437,11.16554,11.585642,11.34277,10.571488,9.508103,8.474257,7.6110773,6.688821,5.6385646,4.8016415,4.9099493,4.535795,4.1517954,3.7251284,3.314872,3.0916924,3.6824617,4.2338467,4.276513,4.027077,4.417641,4.135385,3.5511796,3.0523078,2.7733335,2.5829747,2.2022567,1.6443079,1.211077,1.017436,0.9911796,0.7122052,0.5907693,0.60061544,0.65969235,0.6301539,0.6629744,0.6071795,0.52512825,0.46276927,0.42994875,0.42338464,0.47589746,0.5415385,0.60389745,0.67938465,0.6465641,0.60061544,0.5415385,0.47261542,0.40369233,0.30851284,0.2231795,0.15097436,0.09189744,0.04266667,0.01969231,0.016410258,0.03938462,0.08533334,0.13456412,0.052512825,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.04594872,0.02297436,0.006564103,0.0,0.0032820515,0.016410258,0.059076928,0.07548718,0.06564103,0.04266667,0.02297436,0.01969231,0.016410258,0.01969231,0.029538464,0.04266667,0.06564103,0.108307704,0.16082053,0.3052308,0.702359,0.81066674,0.5973334,0.48246157,0.5316923,0.46933338,0.4955898,0.574359,0.5546667,0.58420515,1.0994873,1.3062565,1.2603078,1.1979488,1.332513,1.8412309,0.78769237,0.4397949,0.512,0.7384616,0.8533334,0.26912823,0.072205134,0.08861539,0.17066668,0.19364104,0.07548718,0.12143591,0.40369233,0.73517954,0.67610264,0.46276927,0.39712822,0.28882053,0.12471796,0.072205134,0.055794876,0.07876924,0.14769232,0.19364104,0.068923086,0.059076928,0.08205129,0.108307704,0.101743594,0.03938462,0.068923086,0.07548718,0.08205129,0.0951795,0.128,0.08533334,0.04594872,0.036102567,0.068923086,0.16410258,0.28225642,0.24615386,0.24615386,0.30851284,0.318359,0.25271797,0.18707694,0.16410258,0.18051283,0.18051283,0.20020515,0.2231795,0.23958977,0.29210258,0.4594872,0.318359,0.19364104,0.17066668,0.33476925,0.7778462,1.017436,1.1782565,1.1552821,0.92225647,0.52512825,0.40369233,0.78769237,1.2865642,1.7329233,2.176,2.3236926,2.231795,2.2416413,2.225231,1.5753847,0.73517954,0.36430773,0.35446155,0.58420515,0.9124103,1.1323078,1.0896411,0.65641034,0.14441027,0.2986667,0.3117949,0.318359,0.33476925,0.36430773,0.40697438,0.48246157,0.39712822,0.34133336,0.4266667,0.67282057,1.5392822,1.3062565,1.2340513,1.847795,2.9440002,3.7218463,3.8137438,3.0851285,1.8412309,0.8336411,0.6465641,0.5415385,0.8336411,1.2898463,1.0994873,0.9517949,1.0010257,1.2537436,1.5622566,1.6278975,2.103795,2.861949,4.2305646,6.052103,7.683283,5.72718,4.3749747,3.7809234,4.020513,5.0674877,5.21518,4.4307694,3.515077,2.9144619,2.7142565,2.6453335,3.43959,4.013949,4.20759,4.7622566,4.781949,4.634257,3.8137438,2.6880002,2.5173335,2.7044106,2.858667,3.0358977,3.058872,2.4910772,1.8576412,1.270154,0.8336411,0.5940513,0.54482055,0.5021539,0.40697438,0.27897438,0.16410258,0.15097436,0.12471796,0.08205129,0.032820515,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.009846155,0.036102567,0.01969231,0.0032820515,0.0032820515,0.009846155,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.006564103,0.006564103,0.0032820515,0.0,0.0,0.006564103,0.009846155,0.006564103,0.0,0.0,0.0,0.006564103,0.006564103,0.0032820515,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.013128206,0.006564103,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0032820515,0.01969231,0.02297436,0.029538464,0.029538464,0.02297436,0.016410258,0.03938462,0.06235898,0.072205134,0.068923086,0.049230773,0.026256412,0.026256412,0.04266667,0.06235898,0.055794876,0.03938462,0.02297436,0.013128206,0.009846155,0.016410258,0.006564103,0.006564103,0.029538464,0.08533334,0.190359,0.27569234,0.380718,0.42338464,0.35446155,0.17066668,0.16738462,0.21333335,0.2297436,0.17723078,0.06235898,0.04266667,0.07548718,0.11158975,0.11158975,0.06235898,0.01969231,0.009846155,0.016410258,0.026256412,0.03938462,0.04266667,0.036102567,0.04594872,0.055794876,0.04266667,0.016410258,0.013128206,0.03938462,0.06235898,0.04266667,0.059076928,0.059076928,0.055794876,0.049230773,0.01969231,0.01969231,0.03938462,0.08205129,0.13128206,0.128,0.12471796,0.13128206,0.15097436,0.16738462,0.16082053,0.108307704,0.118153855,0.118153855,0.09189744,0.08861539,0.06235898,0.032820515,0.009846155,0.0032820515,0.009846155,0.016410258,0.03938462,0.049230773,0.03938462,0.013128206,0.006564103,0.0032820515,0.006564103,0.02297436,0.036102567,0.059076928,0.08861539,0.09189744,0.072205134,0.07876924,0.10502565,0.10502565,0.118153855,0.14441027,0.15097436,0.10502565,0.108307704,0.14112821,0.16410258,0.14112821,0.108307704,0.101743594,0.08533334,0.055794876,0.04594872,0.068923086,0.08861539,0.098461546,0.118153855,0.21661541,0.508718,0.60061544,0.61374366,0.6104616,0.5907693,0.8041026,1.1388719,1.273436,1.1027694,0.7417436,1.0765129,1.4900514,1.910154,2.2186668,2.2580514,2.281026,2.5337439,3.0194874,3.5314875,3.6463592,2.937436,2.4943593,2.3729234,2.3105643,1.7165129,1.463795,2.0644104,3.255795,4.4045134,4.525949,3.3312824,2.6157951,2.1464617,1.9200002,2.172718,2.4155898,2.425436,3.0752823,4.315898,5.1954875,4.919795,4.634257,4.4964104,4.5587697,4.7655387,4.594872,3.9844105,3.239385,2.5435898,1.972513,1.4375386,1.0404103,0.764718,0.574359,0.43323082,0.33476925,0.3511795,0.40697438,0.48574364,0.5907693,0.85005134,1.2340513,1.5327181,1.7165129,1.9396925,2.1891284,2.5796926,2.930872,3.1540515,3.2623591,3.370667,3.639795,3.9351797,4.1747694,4.325744,4.1025643,3.8596926,3.7218463,3.5347695,2.8488207,2.3466668,2.0873847,1.9462565,1.8674873,1.8543591,2.284308,2.422154,2.2219489,1.7066668,0.9747693,0.7318975,0.5021539,0.33805132,0.256,0.2297436,0.24287182,0.26584616,0.29210258,0.318359,0.34789747,0.41025645,0.47589746,0.6235898,0.8795898,1.2077949,1.6672822,2.0578463,2.0644104,1.6771283,1.1881026,0.9288206,0.98133343,1.1815386,1.3653334,1.3718976,1.0305642,0.82379496,0.73517954,0.7122052,0.6695385,0.5481026,0.6859488,1.0633847,1.6311796,2.3204105,3.1113849,4.4406157,6.2818465,8.073847,8.736821,9.186462,12.064821,14.5952835,15.218873,13.590976,10.614155,7.8145647,5.674667,5.0149746,7.0104623,11.208206,16.889437,23.017027,26.857027,23.991796,18.993233,16.282257,14.785643,13.426873,11.122872,9.787078,9.298052,8.612103,7.177847,4.900103,4.338872,4.46359,4.768821,4.8705645,4.532513,4.2962055,3.639795,3.1113849,3.0490258,3.5807183,4.9394875,6.1013336,6.9809237,7.574975,7.958975,7.574975,6.6494365,5.5532312,5.0871797,6.4590774,9.964309,10.443488,8.595693,6.304821,6.633026,10.184206,10.656821,9.429334,7.8637953,7.3353853,6.701949,4.9460516,3.373949,2.6223593,2.6486156,2.4681027,1.9922053,1.394872,0.8598975,0.5907693,0.6170257,0.8763078,0.9616411,0.7778462,0.5513847,10.249847,9.941334,9.206155,7.962257,6.518154,5.5696416,6.36718,6.616616,6.9087186,7.765334,9.6525135,10.758565,10.44677,9.563898,8.418462,6.7807183,5.0018463,5.7435904,7.200821,8.320001,8.802463,8.746667,9.570462,10.30236,10.427077,9.905231,8.805744,7.64718,6.160411,4.9854364,5.677949,4.8344617,3.4592824,2.5665643,2.4910772,2.865231,3.8137438,3.6824617,3.0916924,2.6322052,2.8882053,3.1376412,3.186872,3.2032824,3.255795,3.3280003,3.4921029,3.0260515,2.2449234,1.4703591,1.0699488,0.8008206,0.6498462,0.67282057,0.8041026,0.8730257,0.7253334,0.5316923,0.3708718,0.2855385,0.29538465,0.28225642,0.3052308,0.38728207,0.5316923,0.7187693,0.6826667,0.6235898,0.58092314,0.55794877,0.5349744,0.42994875,0.3249231,0.22646156,0.13456412,0.059076928,0.026256412,0.01969231,0.04594872,0.0951795,0.14112821,0.06235898,0.01969231,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.0032820515,0.009846155,0.02297436,0.032820515,0.02297436,0.02297436,0.036102567,0.059076928,0.101743594,0.1148718,0.055794876,0.016410258,0.02297436,0.059076928,0.13456412,0.19692309,0.18707694,0.20348719,0.5152821,0.69251287,0.7384616,0.7220513,0.6859488,0.6301539,0.39712822,0.23302566,0.18707694,0.26584616,0.4135385,0.38400003,0.41025645,0.69251287,1.2504616,1.9265642,1.024,0.65641034,0.5316923,0.47261542,0.41682056,0.36758977,0.3446154,0.25271797,0.10502565,0.029538464,0.072205134,0.23302566,0.37743592,0.47261542,0.5973334,0.9288206,1.079795,0.6892308,0.036102567,0.006564103,0.02297436,0.026256412,0.026256412,0.02297436,0.013128206,0.0032820515,0.0032820515,0.01969231,0.059076928,0.108307704,0.06564103,0.06564103,0.068923086,0.059076928,0.04594872,0.052512825,0.04266667,0.06235898,0.16082053,0.37415388,0.5874872,0.44964105,0.25928208,0.15097436,0.09189744,0.08205129,0.07876924,0.101743594,0.14112821,0.17723078,0.256,0.31507695,0.31507695,0.25271797,0.18379489,0.12143591,0.14112821,0.21333335,0.30851284,0.38400003,0.6498462,1.1158975,1.401436,1.3128207,0.84348726,0.73517954,1.2570257,1.8937438,2.4320002,2.9472823,3.31159,2.3335385,1.4736412,1.2012309,0.9747693,0.6629744,0.34133336,0.29538465,0.6235898,1.2307693,1.1257436,0.57764107,0.2231795,0.256,0.41682056,0.3511795,0.28225642,0.26584616,0.36430773,0.65641034,0.636718,0.63343596,0.7318975,0.8992821,0.98133343,1.0601027,1.0732309,1.394872,2.1169233,3.0851285,3.764513,5.034667,5.0477953,3.5872824,2.0709746,1.0699488,0.6235898,0.7220513,1.1158975,1.3259488,1.3883078,1.2996924,1.2504616,1.2471796,1.1191796,1.270154,2.4418464,4.9132314,7.3353853,6.7577443,5.5630774,4.6933336,4.269949,4.3618464,4.9920006,4.59159,3.7973337,3.045744,2.5764105,2.428718,2.044718,3.2065644,4.4898467,5.028103,4.525949,3.564308,4.6244106,4.71959,3.259077,2.0611284,1.7755898,2.0644104,2.9604106,4.0500517,4.5062566,3.9909747,2.5993848,1.3161026,0.636718,0.5513847,0.6662565,0.67610264,0.56451285,0.40697438,0.3708718,0.32820517,0.2297436,0.11158975,0.01969231,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.068923086,0.04266667,0.009846155,0.0032820515,0.009846155,0.009846155,0.0032820515,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0032820515,0.0,0.0,0.0032820515,0.016410258,0.01969231,0.013128206,0.02297436,0.016410258,0.016410258,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.02297436,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.009846155,0.009846155,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.009846155,0.0032820515,0.0,0.0,0.0,0.009846155,0.01969231,0.01969231,0.013128206,0.013128206,0.032820515,0.06235898,0.07548718,0.07548718,0.06564103,0.036102567,0.036102567,0.03938462,0.036102567,0.03938462,0.01969231,0.013128206,0.013128206,0.02297436,0.032820515,0.029538464,0.029538464,0.059076928,0.16082053,0.3708718,0.4201026,0.33476925,0.24943592,0.20348719,0.14769232,0.14112821,0.18707694,0.256,0.2855385,0.16410258,0.0951795,0.06235898,0.055794876,0.049230773,0.01969231,0.0032820515,0.0,0.006564103,0.016410258,0.026256412,0.016410258,0.013128206,0.016410258,0.01969231,0.01969231,0.006564103,0.0,0.009846155,0.036102567,0.06564103,0.07548718,0.06564103,0.055794876,0.049230773,0.052512825,0.04266667,0.06564103,0.118153855,0.15097436,0.09189744,0.118153855,0.15097436,0.17394873,0.190359,0.2231795,0.128,0.0951795,0.08205129,0.06235898,0.016410258,0.006564103,0.0,0.0,0.0,0.0,0.0,0.029538464,0.049230773,0.04266667,0.03938462,0.026256412,0.013128206,0.0032820515,0.0032820515,0.0032820515,0.0032820515,0.009846155,0.013128206,0.026256412,0.06235898,0.118153855,0.11158975,0.08533334,0.072205134,0.098461546,0.0951795,0.13456412,0.19364104,0.22646156,0.17723078,0.128,0.14112821,0.13784617,0.10502565,0.068923086,0.08861539,0.118153855,0.15097436,0.21989745,0.3708718,0.6235898,0.6465641,0.57764107,0.5316923,0.5874872,0.7417436,0.88287187,0.9714873,0.99774367,0.98461545,1.3095386,1.8642052,2.3696413,2.7076926,2.9144619,3.1113849,3.3969233,3.69559,3.9253337,4.007385,3.05559,2.5764105,2.3663592,2.2121027,1.8904617,2.409026,4.279795,6.170257,7.24677,7.1876926,4.6178465,3.2098465,2.5304618,2.3335385,2.5731285,3.0818465,3.0654361,3.7021542,4.896821,5.293949,4.9296412,4.3552823,4.017231,4.0041027,4.0336413,3.6332312,3.0851285,2.537026,2.0906668,1.7985642,1.2996924,1.0305642,0.892718,0.76800007,0.5284103,0.41682056,0.508718,0.57764107,0.55794877,0.53825647,1.0043077,1.7591796,2.284308,2.3893335,2.2022567,2.1924105,2.3696413,2.6190772,2.9440002,3.4691284,4.0500517,4.391385,4.519385,4.5423594,4.6572313,4.562052,4.2601027,3.882667,3.446154,2.8324106,2.4582565,2.1825643,1.9790771,1.8215386,1.7033848,2.356513,2.5238976,2.2613335,1.7591796,1.3259488,1.1946667,0.77456415,0.39056414,0.20348719,0.20020515,0.23302566,0.22646156,0.21661541,0.21661541,0.23630771,0.26256412,0.29538465,0.3249231,0.41682056,0.7253334,1.2570257,1.7099489,1.8445129,1.6213335,1.211077,1.1355898,1.211077,1.3620514,1.5425643,1.7165129,1.463795,1.2931283,1.1257436,0.9321026,0.71548724,0.57764107,0.76800007,1.214359,1.8379488,2.546872,2.9538465,4.3552823,6.2752824,7.975385,8.41518,7.899898,10.292514,13.423591,15.356719,14.362258,12.763899,11.460924,9.324308,7.3025646,8.438154,11.904001,17.237335,23.82113,27.697233,21.546669,15.458463,13.321847,14.306462,16.269129,15.740719,11.10318,7.827693,5.5630774,3.9384618,2.546872,2.0709746,2.0578463,2.1924105,2.3040001,2.359795,2.5435898,2.8980515,3.0129232,2.865231,2.806154,3.620103,4.8082056,5.904411,6.7577443,7.5487185,7.4141545,6.6428723,5.868308,5.802667,7.207385,7.968821,8.01477,7.6012316,7.1909747,7.4896417,7.6931286,7.177847,6.2063594,5.3169236,5.32677,6.124308,5.789539,5.21518,4.8804107,4.844308,4.309334,3.0785644,1.8576412,1.017436,0.5874872,0.65312827,1.1454359,1.3095386,0.97805136,0.5874872,10.056206,8.749949,7.4797955,6.7774363,6.5936418,6.301539,5.654975,5.4843082,5.47118,5.549949,5.904411,6.6002054,7.27959,8.408616,9.40636,8.635077,7.5487185,6.738052,6.3606157,6.49518,7.141744,6.9087186,6.5772314,6.3507695,6.3540516,6.62318,5.7074876,4.8016415,4.201026,4.1550775,4.8377438,5.2512827,4.2207184,2.865231,1.975795,1.9987694,3.4625645,3.501949,3.318154,3.3378465,3.2032824,2.5928206,2.6420515,3.1113849,3.69559,4.013949,4.71959,5.7501545,5.077334,2.92759,1.7558975,1.2307693,0.97805136,0.86974365,0.8730257,1.0666667,0.95835906,0.74830776,0.5284103,0.380718,0.380718,0.32164106,0.2855385,0.32820517,0.47589746,0.7318975,0.7318975,0.7515898,0.7581539,0.72861546,0.65641034,0.42338464,0.27569234,0.17066668,0.0951795,0.04594872,0.032820515,0.03938462,0.052512825,0.06564103,0.09189744,0.09189744,0.055794876,0.02297436,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.0032820515,0.0,0.04266667,0.108307704,0.108307704,0.04594872,0.02297436,0.059076928,0.17394873,0.380718,0.40697438,0.17394873,0.016410258,0.02297436,0.04594872,0.18051283,0.24943592,0.17066668,0.03938462,0.13784617,0.39384618,0.5316923,0.5481026,0.5316923,0.64000005,0.60389745,0.4660513,0.44307697,0.65969235,1.1585642,1.0502565,0.7581539,0.5874872,0.6432821,0.8402052,0.9124103,0.7122052,0.60061544,0.73517954,1.0535386,1.394872,1.5360001,1.1881026,0.51856416,0.15097436,0.06564103,0.108307704,0.24287182,0.39056414,0.4266667,1.4539489,2.0020514,1.3292309,0.029538464,0.029538464,0.06564103,0.07548718,0.04594872,0.0,0.0,0.013128206,0.016410258,0.07548718,0.21661541,0.4135385,0.20348719,0.20676924,0.24943592,0.25271797,0.2297436,0.26584616,0.2100513,0.16738462,0.18051283,0.2297436,0.26584616,0.128,0.029538464,0.029538464,0.029538464,0.029538464,0.029538464,0.036102567,0.055794876,0.09189744,0.15097436,0.17723078,0.16410258,0.12143591,0.06235898,0.098461546,0.39056414,0.8041026,1.1158975,1.0075898,1.2635899,1.2635899,1.2274873,1.2931283,1.5261539,1.3292309,0.86974365,0.5874872,0.65312827,0.94523084,1.2012309,1.339077,1.2964103,1.0601027,0.65641034,0.32820517,0.41025645,0.892718,1.5721027,2.0611284,1.8281027,1.148718,0.5973334,0.42994875,0.56451285,0.4660513,0.40697438,0.3446154,0.31507695,0.4135385,0.7056411,1.2996924,1.9396925,2.3630772,2.28759,2.2383592,1.9068719,1.6705642,1.8149745,2.546872,4.0369234,3.8071797,3.8662567,4.5128207,4.31918,1.1552821,0.4955898,0.6465641,0.8960001,1.4966155,2.1070771,2.103795,1.6311796,1.1323078,1.3259488,2.0709746,3.255795,4.9821544,5.914257,3.2656412,3.1081028,3.945026,4.9296412,5.225026,4.027077,4.2240005,4.57518,4.768821,4.637539,4.1517954,3.4921029,3.5446157,3.8334363,3.8531284,3.0982566,2.7306669,2.5206156,2.2350771,1.8773335,1.6935385,2.1202054,2.612513,3.0523078,3.761231,5.5072823,6.1078978,3.7842054,1.7165129,1.0043077,0.6859488,0.67282057,0.75487185,0.827077,0.81066674,0.64000005,0.51856416,0.37743592,0.23302566,0.101743594,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.009846155,0.016410258,0.02297436,0.04594872,0.04594872,0.01969231,0.0,0.0,0.0,0.013128206,0.016410258,0.009846155,0.0,0.0,0.02297436,0.08533334,0.098461546,0.059076928,0.04594872,0.02297436,0.016410258,0.016410258,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.03938462,0.055794876,0.036102567,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.016410258,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.016410258,0.016410258,0.016410258,0.016410258,0.026256412,0.02297436,0.009846155,0.0032820515,0.016410258,0.016410258,0.032820515,0.068923086,0.108307704,0.108307704,0.0951795,0.08205129,0.0951795,0.16082053,0.32164106,0.28225642,0.33805132,0.3511795,0.26912823,0.12143591,0.049230773,0.07548718,0.15425642,0.22646156,0.21333335,0.1148718,0.08205129,0.06564103,0.04266667,0.029538464,0.006564103,0.0,0.006564103,0.016410258,0.016410258,0.0032820515,0.0,0.01969231,0.04266667,0.029538464,0.01969231,0.006564103,0.006564103,0.026256412,0.07548718,0.026256412,0.07876924,0.17066668,0.24615386,0.25928208,0.11158975,0.13128206,0.16738462,0.15097436,0.09189744,0.128,0.118153855,0.16082053,0.25928208,0.32164106,0.23630771,0.16738462,0.108307704,0.052512825,0.016410258,0.016410258,0.006564103,0.0,0.0,0.0,0.0,0.009846155,0.02297436,0.03938462,0.07548718,0.06564103,0.04266667,0.02297436,0.016410258,0.016410258,0.016410258,0.006564103,0.013128206,0.036102567,0.06235898,0.24287182,0.22646156,0.14112821,0.072205134,0.06235898,0.14769232,0.11158975,0.059076928,0.029538464,0.029538464,0.029538464,0.07548718,0.0951795,0.0951795,0.16738462,0.26584616,0.2986667,0.27569234,0.24943592,0.33476925,0.51856416,0.69251287,0.77128214,0.7089231,0.48902568,0.53825647,0.65969235,0.8533334,1.1552821,1.6311796,1.8773335,2.3302567,2.861949,3.3542566,3.7087183,4.013949,4.31918,4.384821,4.240411,4.164923,4.7261543,4.46359,4.2994876,4.5489235,4.9296412,5.720616,7.706257,8.43159,7.4929237,6.514872,5.100308,3.7743592,3.05559,2.8160002,2.3040001,1.9265642,1.9856411,2.6715899,3.5610259,3.6463592,3.0851285,2.550154,2.2088206,2.1070771,2.166154,1.9593848,1.7624617,1.6147693,1.5425643,1.5425643,1.5425643,1.522872,1.4375386,1.273436,1.0535386,0.73517954,0.7122052,0.6268718,0.40369233,0.24287182,0.4397949,1.1388719,2.2482052,3.2787695,3.3247182,2.7766156,2.3466668,2.2744617,2.6289232,3.31159,4.1550775,4.775385,5.100308,5.156103,5.097026,5.2545643,5.110154,4.673641,4.066462,3.5413337,3.2361028,2.8389745,2.3696413,1.9232821,1.6771283,2.5074873,2.7995899,2.3958976,1.5360001,0.8402052,1.1946667,0.92553854,0.5021539,0.20020515,0.09189744,0.10502565,0.108307704,0.12471796,0.17394873,0.25928208,0.3446154,0.35774362,0.30194873,0.2855385,0.51856416,1.0666667,1.5261539,1.6836925,1.5655385,1.4178462,1.4309745,1.3883078,1.3226668,1.3357949,1.6180514,1.5819489,1.5819489,1.4572309,1.1782565,0.82379496,0.82379496,1.0338463,1.1191796,1.0075898,0.88615394,1.3259488,3.5577438,6.23918,8.303591,8.986258,8.218257,8.2904625,8.94359,9.186462,7.2927184,6.9645133,7.8703594,8.04759,6.961231,5.5072823,10.673231,18.225233,25.225847,29.0199,27.237745,20.62113,15.048206,12.087796,12.688411,17.18154,11.382154,7.506052,5.218462,4.023795,3.2820516,3.3903592,3.9122055,4.069744,3.6168208,2.8225644,2.5304618,2.7142565,2.7798977,2.487795,1.9364104,2.4516926,3.95159,4.7589746,4.827898,5.7665644,6.951385,7.7981544,8.425026,8.976411,9.613129,9.357129,8.329846,6.810257,5.2053337,4.059898,5.756718,7.269744,7.4699492,5.8518977,2.5173335,2.8947694,5.297231,7.6307697,8.615385,7.7981544,5.3202057,3.242667,1.7296412,0.8336411,0.5021539,0.7220513,1.3357949,1.5130258,1.0994873,0.6104616,5.2578464,5.435077,5.681231,6.0980515,6.5969234,6.8988724,6.8988724,7.394462,8.411898,9.337437,8.920616,7.1548724,6.5870776,6.9349747,7.748924,8.41518,8.910769,8.385642,7.578257,6.9809237,6.8496413,5.677949,5.3891287,5.32677,5.175795,4.97559,4.6145644,4.529231,4.6211286,4.9887185,5.937231,7.003898,6.892308,5.8912826,4.4832826,3.318154,3.131077,3.1507695,3.2525132,3.3608208,3.4592824,3.1934361,2.8488207,2.5796926,2.422154,2.3401027,2.6289232,3.0030773,3.170462,2.9472823,2.2547693,1.8379488,1.6377437,1.4539489,1.2438976,1.1158975,0.83035904,0.5973334,0.43323082,0.34133336,0.3314872,0.3117949,0.27241027,0.29210258,0.40369233,0.6104616,0.78769237,0.86317956,0.84348726,0.7417436,0.571077,0.35774362,0.20020515,0.098461546,0.049230773,0.02297436,0.01969231,0.01969231,0.032820515,0.059076928,0.10502565,0.1148718,0.0951795,0.052512825,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.026256412,0.036102567,0.029538464,0.02297436,0.01969231,0.02297436,0.03938462,0.06564103,0.08861539,0.15097436,0.14112821,0.08205129,0.016410258,0.02297436,0.108307704,0.15753847,0.17066668,0.23630771,0.5284103,0.43323082,0.636718,0.9189744,1.0765129,0.9353847,0.48574364,0.48246157,0.56123084,0.574359,0.5874872,0.6826667,0.41682056,0.21333335,0.24943592,0.47261542,0.85005134,1.4834872,1.3850257,0.69251287,0.69907695,1.332513,1.8543591,1.6968206,1.0010257,0.60389745,0.5677949,0.6235898,0.57764107,0.40697438,0.26912823,0.39712822,0.508718,0.44307697,0.26256412,0.26256412,0.41682056,0.45620516,0.44307697,0.45292312,0.5481026,0.32820517,0.256,0.25928208,0.27241027,0.25271797,0.0951795,0.072205134,0.12471796,0.20348719,0.26584616,0.26256412,0.15425642,0.068923086,0.049230773,0.059076928,0.1148718,0.2100513,0.23302566,0.20020515,0.24943592,0.25928208,0.21989745,0.20348719,0.2231795,0.20020515,0.20348719,0.20676924,0.19364104,0.17066668,0.15753847,0.29210258,1.1684103,2.2547693,2.737231,1.4966155,1.5163078,1.6213335,1.8379488,2.103795,2.2580514,0.8730257,0.44964105,0.5415385,0.8205129,1.1060513,1.1946667,1.5556924,1.6278975,1.3850257,1.3161026,1.4736412,1.3062565,1.204513,1.2438976,1.1552821,1.2668719,1.6443079,1.595077,1.2603078,1.6377437,1.785436,1.4703591,1.1684103,0.9321026,0.37415388,0.512,0.8566154,1.3554872,1.9462565,2.556718,3.18359,3.3345644,3.1540515,2.8258464,2.5731285,4.2962055,4.378257,3.8990772,3.3345644,2.5731285,1.4506668,0.9616411,1.1158975,1.7591796,2.5829747,2.802872,1.8740515,1.3161026,1.6508719,2.4024618,3.1376412,3.4527183,3.9351797,4.450462,4.1452312,4.601436,5.2414365,5.2676926,4.4012313,2.8914874,3.0293336,3.3378465,3.3017437,2.9538465,2.8553848,2.481231,2.7667694,3.0752823,2.8127182,1.4506668,2.0118976,2.1924105,2.3171284,2.5665643,2.9997952,3.0654361,2.8882053,2.9669745,3.5052311,4.420923,4.5817437,3.1081028,1.6475899,0.8730257,0.47917953,0.43651286,0.5021539,0.6432821,0.77128214,0.7253334,0.7220513,0.77128214,0.6104616,0.27569234,0.11158975,0.06235898,0.01969231,0.0,0.0,0.0,0.0,0.016410258,0.04266667,0.072205134,0.108307704,0.13456412,0.13784617,0.108307704,0.059076928,0.0,0.0032820515,0.0032820515,0.0032820515,0.0032820515,0.013128206,0.006564103,0.032820515,0.052512825,0.059076928,0.04594872,0.02297436,0.006564103,0.0032820515,0.0032820515,0.0,0.0,0.006564103,0.006564103,0.0,0.0,0.0,0.0,0.0032820515,0.01969231,0.049230773,0.029538464,0.016410258,0.013128206,0.013128206,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.009846155,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.0032820515,0.016410258,0.02297436,0.013128206,0.0032820515,0.006564103,0.0032820515,0.013128206,0.026256412,0.026256412,0.016410258,0.01969231,0.029538464,0.04266667,0.032820515,0.029538464,0.029538464,0.029538464,0.04594872,0.07548718,0.08861539,0.10502565,0.108307704,0.0951795,0.08533334,0.052512825,0.052512825,0.068923086,0.08533334,0.10502565,0.08533334,0.098461546,0.11158975,0.10502565,0.10502565,0.068923086,0.11158975,0.14769232,0.12143591,0.016410258,0.02297436,0.02297436,0.03938462,0.059076928,0.06564103,0.036102567,0.032820515,0.09189744,0.18707694,0.24615386,0.256,0.15425642,0.13456412,0.22646156,0.29538465,0.26584616,0.256,0.21333335,0.14112821,0.07876924,0.1148718,0.19364104,0.32164106,0.42994875,0.39384618,0.27897438,0.19692309,0.15425642,0.13128206,0.07548718,0.055794876,0.036102567,0.013128206,0.0,0.0,0.0,0.0032820515,0.013128206,0.04266667,0.08861539,0.1148718,0.0951795,0.06235898,0.03938462,0.03938462,0.03938462,0.03938462,0.03938462,0.03938462,0.02297436,0.052512825,0.04594872,0.029538464,0.016410258,0.02297436,0.04266667,0.036102567,0.01969231,0.006564103,0.006564103,0.016410258,0.036102567,0.06235898,0.108307704,0.18051283,0.2297436,0.24287182,0.23302566,0.24287182,0.34789747,0.60061544,0.98133343,1.2603078,1.3029745,1.0732309,0.8992821,0.90584624,1.0929232,1.3554872,1.4998976,1.4900514,2.225231,2.793026,2.9833848,3.2689233,3.876103,4.4110775,4.6867695,4.70318,4.630975,4.565334,4.417641,4.125539,4.2436924,5.940513,6.51159,6.957949,6.7872825,6.2851286,6.5280004,5.32677,4.312616,3.6102567,3.2820516,3.318154,2.6453335,2.2022567,1.9528207,1.8149745,1.6443079,1.7755898,1.6640002,1.595077,1.6836925,1.8609232,2.2383592,2.2744617,2.0644104,1.7591796,1.5524104,1.5622566,1.4441026,1.2471796,1.0469744,0.9419488,0.77128214,0.6826667,0.6301539,0.6301539,0.7450257,0.79425645,1.3226668,2.4648206,3.817026,4.460308,3.7349746,2.9538465,2.5304618,2.6945643,3.5052311,4.31918,4.9854364,5.395693,5.5762057,5.671385,5.5663595,5.179077,4.6080003,4.013949,3.626667,3.3969233,3.3345644,3.2754874,3.255795,3.508513,4.2994876,3.7743592,2.5238976,1.2274873,0.6695385,0.72861546,0.51856416,0.25928208,0.07876924,0.01969231,0.029538464,0.03938462,0.04594872,0.055794876,0.11158975,0.24615386,0.3511795,0.380718,0.3708718,0.45620516,1.1355898,1.7690258,2.1234872,2.100513,1.7493335,1.7033848,1.6804104,1.6836925,1.7263591,1.8609232,1.6410258,1.4900514,1.3718976,1.2570257,1.1290257,1.0896411,1.2898463,1.5163078,1.6246156,1.5327181,1.5721027,2.3072822,4.384821,7.1023593,8.402052,7.837539,7.706257,8.411898,8.700719,5.6451287,3.6463592,3.2065644,3.0884104,2.802872,2.5895386,5.4908724,13.269335,23.958977,33.142155,33.939693,26.23672,21.287386,17.795284,14.057027,7.9524107,6.012718,4.457026,3.5774362,3.2820516,3.0851285,3.1277952,3.7710772,4.2371287,4.089436,3.239385,2.281026,2.1431797,2.100513,1.8084104,1.3259488,1.3915899,2.156308,3.0851285,3.948308,4.841026,5.730462,6.619898,7.4896417,8.320001,9.110975,8.835282,7.6012316,5.7107697,3.7973337,2.8258464,3.889231,5.2578464,5.605744,4.857436,4.1911798,5.7107697,6.0324106,5.4153852,4.204308,2.8291285,2.0611284,1.585231,1.2274873,0.90256417,0.61374366,0.84348726,1.4211283,1.6082052,1.2012309,0.53825647,4.673641,4.3651285,4.348718,4.647385,5.106872,5.4186673,5.914257,6.8266673,7.9261546,8.832001,8.996103,7.5552826,7.3091288,7.2664623,7.0925136,7.145026,7.171283,7.056411,6.8365135,6.5378466,6.170257,5.280821,4.972308,5.0149746,5.113436,4.8836927,4.57518,4.4373336,4.263385,4.132103,4.4077954,5.5236926,6.2851286,6.3540516,5.5893335,4.059898,2.8750772,2.3138463,2.15959,2.2613335,2.546872,3.0490258,3.0194874,2.6289232,2.100513,1.719795,2.028308,2.2088206,2.3040001,2.1989746,1.6377437,1.5130258,1.4211283,1.3522053,1.2865642,1.211077,0.9321026,0.58092314,0.33805132,0.24615386,0.2100513,0.18379489,0.18379489,0.2297436,0.33476925,0.50543594,0.6826667,0.77456415,0.77128214,0.67938465,0.512,0.318359,0.16082053,0.068923086,0.032820515,0.016410258,0.006564103,0.006564103,0.013128206,0.03938462,0.08861539,0.1148718,0.10502565,0.06564103,0.01969231,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01969231,0.049230773,0.049230773,0.029538464,0.04594872,0.04266667,0.03938462,0.029538464,0.016410258,0.006564103,0.16738462,0.25271797,0.23630771,0.16082053,0.1148718,0.19692309,0.29210258,0.41682056,0.6170257,0.9747693,0.65969235,0.56123084,0.56451285,0.56123084,0.44964105,0.26584616,0.25271797,0.63343596,1.1881026,1.2373334,0.79097444,0.51856416,0.37415388,0.36430773,0.53825647,0.98133343,1.6607181,1.4572309,0.52512825,0.2986667,0.5677949,0.8172308,0.7811283,0.5513847,0.5874872,0.5874872,0.55794877,0.4660513,0.318359,0.16410258,0.10502565,0.128,0.19692309,0.25928208,0.23958977,0.34133336,0.38728207,0.39384618,0.3708718,0.34789747,0.18379489,0.190359,0.29210258,0.40697438,0.44307697,0.2297436,0.15425642,0.13128206,0.12471796,0.13784617,0.13128206,0.072205134,0.032820515,0.036102567,0.04266667,0.059076928,0.1148718,0.13456412,0.13128206,0.18707694,0.21333335,0.2100513,0.2100513,0.23630771,0.30194873,0.24615386,0.19364104,0.18707694,0.27897438,0.512,0.7384616,1.1913847,1.6836925,1.9035898,1.4145643,1.467077,1.276718,1.1158975,1.1126155,1.270154,0.49230772,0.4135385,0.6432821,0.9616411,1.3095386,1.6640002,1.8346668,1.8838975,1.8740515,1.8642052,1.7493335,1.522872,1.3161026,1.1323078,0.8566154,0.81066674,1.1158975,1.3850257,1.7329233,2.7503593,2.934154,2.6223593,3.0129232,3.4888208,1.6213335,1.014154,1.0436924,1.5392822,2.169436,2.4320002,3.006359,3.2000003,3.131077,2.986667,3.0358977,3.9778464,4.2141542,3.9220517,3.2623591,2.3663592,2.1267693,2.5107694,3.2262566,3.9909747,4.5554876,3.9614363,2.225231,1.2209232,1.4736412,2.166154,2.8324106,3.245949,4.516103,6.439385,7.496206,7.6570263,7.2336416,5.979898,4.2305646,2.8849232,2.7273848,2.678154,2.4648206,2.2711797,2.7602053,2.3335385,2.349949,2.6715899,2.7831798,1.7985642,1.785436,1.9856411,2.356513,2.7076926,2.6847181,3.387077,3.2000003,3.0096412,3.239385,3.876103,3.1934361,2.1333334,1.2406155,0.72861546,0.48246157,0.4266667,0.3708718,0.39712822,0.5481026,0.8205129,1.276718,1.7263591,1.5327181,0.8172308,0.42994875,0.3314872,0.12471796,0.0,0.0,0.0,0.0,0.02297436,0.04266667,0.07548718,0.17723078,0.17066668,0.14112821,0.08861539,0.036102567,0.036102567,0.02297436,0.013128206,0.013128206,0.016410258,0.006564103,0.016410258,0.01969231,0.026256412,0.036102567,0.04594872,0.013128206,0.006564103,0.009846155,0.009846155,0.009846155,0.0032820515,0.0032820515,0.009846155,0.016410258,0.009846155,0.0032820515,0.0,0.006564103,0.02297436,0.052512825,0.072205134,0.07876924,0.055794876,0.02297436,0.016410258,0.016410258,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.0032820515,0.006564103,0.009846155,0.0032820515,0.0,0.0,0.006564103,0.013128206,0.02297436,0.029538464,0.032820515,0.02297436,0.013128206,0.013128206,0.016410258,0.02297436,0.029538464,0.029538464,0.029538464,0.04266667,0.06564103,0.08533334,0.08861539,0.08205129,0.08533334,0.07548718,0.055794876,0.03938462,0.029538464,0.029538464,0.04594872,0.072205134,0.10502565,0.128,0.12143591,0.08533334,0.11158975,0.13456412,0.11158975,0.04266667,0.06235898,0.08205129,0.101743594,0.108307704,0.08533334,0.072205134,0.108307704,0.20676924,0.31507695,0.318359,0.27569234,0.19692309,0.18707694,0.256,0.3052308,0.23302566,0.17394873,0.14769232,0.17066668,0.24943592,0.3249231,0.41025645,0.48246157,0.47589746,0.32164106,0.18379489,0.118153855,0.0951795,0.08861539,0.06564103,0.04594872,0.029538464,0.013128206,0.0032820515,0.009846155,0.009846155,0.0032820515,0.009846155,0.026256412,0.04594872,0.08205129,0.08533334,0.08533334,0.10502565,0.15425642,0.10502565,0.08205129,0.072205134,0.06564103,0.032820515,0.013128206,0.0032820515,0.0,0.0,0.006564103,0.013128206,0.016410258,0.009846155,0.0032820515,0.009846155,0.02297436,0.049230773,0.08205129,0.10502565,0.118153855,0.14112821,0.17394873,0.19692309,0.21661541,0.25928208,0.39712822,0.6498462,0.9485129,1.1946667,1.2471796,1.1979488,1.1749744,1.1848207,1.2800001,1.5458462,1.6344616,2.0676925,2.3827693,2.4549747,2.5271797,2.8750772,3.4625645,4.092718,4.450462,4.1124105,4.854154,5.989744,6.514872,6.3277955,6.2227697,6.3967185,7.1909747,7.7456417,7.79159,7.637334,6.3442054,5.139693,4.1911798,3.5511796,3.1507695,2.3401027,1.6705642,1.2865642,1.2800001,1.6935385,2.7963078,3.4297438,3.5610259,3.383795,3.314872,3.639795,3.5610259,3.1770258,2.6945643,2.4155898,1.9528207,1.3883078,0.97805136,0.8467693,0.97805136,0.8960001,0.69907695,0.5973334,0.69251287,0.97805136,1.1979488,1.9003079,2.9505644,4.0402055,4.71959,4.4045134,3.761231,3.2754874,3.2196925,3.6660516,4.522667,5.366154,5.970052,6.245744,6.235898,5.7403083,5.208616,4.6605134,4.1714873,3.876103,3.9253337,4.2962055,4.7950773,5.3005133,5.7435904,5.7698464,4.571898,2.7241027,1.0043077,0.4135385,0.30851284,0.2100513,0.128,0.06235898,0.0,0.013128206,0.013128206,0.013128206,0.01969231,0.03938462,0.12143591,0.21989745,0.3052308,0.37415388,0.4594872,0.78769237,1.3292309,1.7066668,1.7493335,1.4933335,1.394872,1.4539489,1.5458462,1.6016412,1.6114873,1.4834872,1.463795,1.5261539,1.6147693,1.6443079,1.4703591,1.3587693,1.3095386,1.2931283,1.2438976,1.8051283,3.5807183,5.5236926,7.0104623,7.834257,7.3058467,7.384616,8.411898,9.209436,7.066257,3.4691284,2.2022567,1.9856411,2.0053334,1.9265642,2.7766156,6.6494365,14.742975,25.133951,32.784412,30.920208,26.581335,21.123283,15.274668,9.143796,7.1909747,5.3891287,3.8728209,2.809436,2.4057438,2.605949,3.05559,3.5314875,3.620103,2.7011285,2.1333334,2.2646155,2.422154,2.2153847,1.5327181,1.2406155,1.4605129,2.0545642,2.868513,3.748103,4.857436,6.042257,6.961231,7.4436927,7.4765134,7.0498466,5.973334,4.7622566,3.757949,3.121231,3.4166157,4.6112823,5.5204105,5.805949,5.9536414,6.514872,7.6701546,7.2861543,4.9427695,1.9364104,1.6443079,1.5425643,1.3915899,1.1191796,0.82379496,1.0633847,1.5097437,1.6049232,1.204513,0.58420515,5.868308,5.3005133,4.8705645,5.0149746,5.5138464,5.4941545,5.4186673,5.933949,6.426257,6.7544622,7.2631803,7.1089234,7.53559,7.584821,7.00718,6.2720003,5.7074876,5.543385,5.402257,5.169231,4.9985647,4.8049235,4.670359,4.699898,4.8147697,4.7622566,4.44718,4.2568207,3.9220517,3.383795,2.789744,3.2754874,4.138667,4.9132314,5.182359,4.6145644,3.6693337,2.5600002,1.7985642,1.5786668,1.7887181,2.4943593,2.8389745,2.7536411,2.3302567,1.8379488,1.8281027,1.7755898,1.6180514,1.3489232,1.0272821,1.142154,1.214359,1.2438976,1.2077949,1.0666667,0.81066674,0.4955898,0.26912823,0.17394873,0.14441027,0.12471796,0.15425642,0.21661541,0.31507695,0.45620516,0.5907693,0.65969235,0.6629744,0.60389745,0.49887183,0.30194873,0.14769232,0.052512825,0.016410258,0.009846155,0.0032820515,0.0,0.006564103,0.02297436,0.052512825,0.08205129,0.08533334,0.059076928,0.02297436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.01969231,0.04594872,0.049230773,0.03938462,0.052512825,0.03938462,0.04266667,0.036102567,0.013128206,0.0,0.17723078,0.28882053,0.3249231,0.29210258,0.23302566,0.21989745,0.33476925,0.50543594,0.71548724,1.0043077,0.8730257,0.71548724,0.47917953,0.21661541,0.07548718,0.128,0.08861539,0.5021539,1.1881026,1.2570257,0.67938465,0.51856416,0.5415385,0.6104616,0.69579494,0.9682052,1.3292309,1.1520001,0.53825647,0.3052308,0.21661541,0.14112821,0.08861539,0.1148718,0.3314872,0.3446154,0.28225642,0.22646156,0.2100513,0.21333335,0.12471796,0.1148718,0.15097436,0.19692309,0.21333335,0.3052308,0.30851284,0.26256412,0.20020515,0.128,0.07548718,0.101743594,0.190359,0.30851284,0.39384618,0.26584616,0.21333335,0.16410258,0.11158975,0.11158975,0.14112821,0.08205129,0.052512825,0.07548718,0.10502565,0.0951795,0.055794876,0.03938462,0.06564103,0.12471796,0.15097436,0.17066668,0.16738462,0.17394873,0.26584616,0.27241027,0.28225642,0.34789747,0.5152821,0.8467693,1.6738462,1.9364104,1.7657437,1.4211283,1.3062565,1.2898463,0.8992821,0.5152821,0.38400003,0.60389745,0.36430773,0.4266667,0.5907693,0.764718,0.955077,1.2373334,1.332513,1.4605129,1.6278975,1.6311796,1.3653334,1.2931283,1.2668719,1.2471796,1.2964103,1.5983591,2.172718,2.356513,2.3105643,3.0293336,3.318154,3.4100516,4.1485133,4.781949,2.9571285,2.169436,2.044718,2.412308,2.9078977,2.9505644,3.255795,3.9154875,4.7491283,5.0674877,3.6726158,3.889231,4.161641,4.2371287,4.007385,3.511795,5.146257,5.2742567,4.7950773,4.342154,4.2994876,3.889231,2.789744,2.5074873,3.4166157,4.772103,5.7403083,6.294975,7.174565,8.257642,8.533334,8.198565,7.79159,6.242462,3.9023592,2.5173335,2.2678976,2.2416413,1.9856411,1.6869745,2.156308,2.0545642,2.0775387,2.3335385,2.537026,1.9987694,1.6705642,1.8510771,2.15959,2.3335385,2.2514873,3.0851285,2.8980515,2.487795,2.5009232,3.442872,2.3893335,1.6377437,1.142154,0.80738467,0.512,0.4135385,0.3052308,0.26912823,0.36758977,0.6498462,1.0338463,1.5556924,1.5392822,1.0010257,0.6301539,0.42338464,0.14769232,0.0,0.0,0.0,0.0,0.02297436,0.055794876,0.10502565,0.20676924,0.17066668,0.098461546,0.036102567,0.016410258,0.055794876,0.036102567,0.026256412,0.02297436,0.01969231,0.006564103,0.016410258,0.016410258,0.01969231,0.032820515,0.059076928,0.02297436,0.013128206,0.016410258,0.016410258,0.016410258,0.013128206,0.01969231,0.029538464,0.029538464,0.009846155,0.0032820515,0.0,0.016410258,0.049230773,0.08205129,0.098461546,0.098461546,0.072205134,0.029538464,0.026256412,0.04594872,0.02297436,0.0032820515,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.0032820515,0.006564103,0.013128206,0.009846155,0.0,0.0,0.006564103,0.009846155,0.009846155,0.01969231,0.026256412,0.016410258,0.006564103,0.006564103,0.032820515,0.07548718,0.0951795,0.07548718,0.03938462,0.04266667,0.055794876,0.068923086,0.072205134,0.068923086,0.06235898,0.08205129,0.108307704,0.12143591,0.0951795,0.029538464,0.036102567,0.06235898,0.10502565,0.14441027,0.14112821,0.1148718,0.14441027,0.15097436,0.118153855,0.08533334,0.108307704,0.16082053,0.18707694,0.16082053,0.10502565,0.07548718,0.10502565,0.25271797,0.42338464,0.37743592,0.24287182,0.18707694,0.21333335,0.27241027,0.28225642,0.20676924,0.17066668,0.190359,0.29210258,0.49887183,0.5874872,0.64000005,0.6268718,0.5152821,0.26584616,0.128,0.072205134,0.055794876,0.04594872,0.026256412,0.01969231,0.013128206,0.006564103,0.0032820515,0.009846155,0.009846155,0.036102567,0.06235898,0.06235898,0.032820515,0.055794876,0.06564103,0.08205129,0.1148718,0.18707694,0.15425642,0.118153855,0.101743594,0.108307704,0.0951795,0.08533334,0.055794876,0.026256412,0.009846155,0.006564103,0.009846155,0.013128206,0.016410258,0.01969231,0.02297436,0.029538464,0.0951795,0.16738462,0.19364104,0.13128206,0.17394873,0.21661541,0.22646156,0.20348719,0.20348719,0.25271797,0.37743592,0.5940513,0.8467693,1.0043077,1.1552821,1.276718,1.3029745,1.3128207,1.5097437,1.6705642,1.9035898,2.15959,2.3630772,2.422154,2.4385643,2.868513,3.6069746,4.2240005,3.9844105,4.919795,6.6494365,7.719385,7.5979495,6.675693,6.8496413,8.283898,10.085744,11.057232,9.6754875,8.329846,7.2664623,6.196513,4.9854364,3.636513,2.5435898,1.847795,1.7558975,2.3368206,3.5380516,4.7327185,5.540103,5.720616,5.3431797,4.785231,4.6966157,4.4996924,4.1682053,3.8006158,3.620103,3.1507695,2.2547693,1.5327181,1.2603078,1.3817437,1.4736412,1.1454359,0.8336411,0.74830776,0.86317956,1.2373334,2.0545642,2.9768207,3.8071797,4.4800005,4.57518,4.2338467,3.8367183,3.6562054,3.8859491,4.706462,5.586052,6.2687182,6.5772314,6.422975,5.802667,5.182359,4.604718,4.1156926,3.7710772,4.312616,5.2480006,6.245744,7.0137444,7.2927184,6.363898,4.578462,2.4910772,0.761436,0.17723078,0.068923086,0.049230773,0.052512825,0.04594872,0.006564103,0.009846155,0.0032820515,0.006564103,0.016410258,0.026256412,0.049230773,0.1148718,0.2297436,0.38400003,0.5349744,0.5677949,0.86646163,1.2242053,1.4736412,1.4867693,1.4966155,1.5721027,1.654154,1.6475899,1.4572309,1.3620514,1.3850257,1.4966155,1.719795,2.1464617,2.2121027,1.8773335,1.4605129,1.1815386,1.142154,1.8773335,4.5128207,7.1122055,8.585847,8.700719,7.39118,7.0892315,7.719385,8.39877,7.430565,4.391385,3.2131286,2.6847181,2.2777438,2.1530259,1.9823592,2.7733335,6.9087186,14.8480015,25.114258,29.417028,26.069336,21.458054,17.719797,12.760616,8.306872,5.901129,4.266667,2.9440002,2.294154,2.4155898,2.6486156,2.858667,2.8356924,2.2744617,2.3138463,2.8127182,3.2853336,3.2984617,2.4549747,1.8543591,1.6311796,1.7985642,2.3860514,3.4658465,4.713026,5.986462,6.8266673,6.997334,6.488616,5.504,4.644103,4.1124105,3.8695388,3.6168208,3.7349746,4.5029745,5.297231,5.901129,6.514872,7.4141545,8.342975,8.395488,7.0400004,4.089436,2.8553848,2.4648206,2.1398976,1.5753847,0.9353847,1.2570257,1.7263591,1.9068719,1.591795,0.81394875,6.7840004,6.6560006,6.308103,6.5378466,7.171283,7.0859494,6.2063594,5.986462,5.7403083,5.35959,5.3234878,5.6254363,6.196513,6.665847,6.764308,6.3343596,5.7796926,5.2676926,4.604718,3.9745643,3.9122055,4.07959,4.161641,4.073026,3.9253337,4.020513,3.895795,3.8400004,3.7218463,3.3214362,2.3236926,1.8543591,2.0217438,2.6486156,3.5446157,4.493129,4.713026,3.751385,2.6847181,2.0217438,1.7132308,1.7985642,2.172718,2.487795,2.5107694,2.1333334,1.5819489,1.2242053,0.99774367,0.86646163,0.84348726,1.0502565,1.2471796,1.2800001,1.079795,0.69251287,0.446359,0.30851284,0.21661541,0.15097436,0.15097436,0.17066668,0.21661541,0.27897438,0.35446155,0.446359,0.5415385,0.56451285,0.5481026,0.512,0.47261542,0.26912823,0.13128206,0.04594872,0.0032820515,0.0032820515,0.0,0.0,0.0032820515,0.013128206,0.013128206,0.032820515,0.049230773,0.04266667,0.02297436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.02297436,0.016410258,0.02297436,0.032820515,0.036102567,0.02297436,0.006564103,0.026256412,0.03938462,0.036102567,0.009846155,0.09189744,0.20020515,0.2855385,0.318359,0.29210258,0.17723078,0.32820517,0.49230772,0.58420515,0.7187693,0.955077,0.9485129,0.702359,0.35774362,0.18379489,0.23302566,0.16082053,0.28225642,0.53825647,0.5021539,0.5481026,0.75487185,0.8205129,0.7056411,0.6465641,0.8008206,0.9353847,0.86317956,0.636718,0.5349744,0.4135385,0.2855385,0.17723078,0.098461546,0.06564103,0.08533334,0.07548718,0.08205129,0.14441027,0.2855385,0.15097436,0.10502565,0.12471796,0.18707694,0.26912823,0.36102566,0.28882053,0.2100513,0.20676924,0.26912823,0.23302566,0.16082053,0.0951795,0.06235898,0.08205129,0.128,0.17066668,0.18379489,0.19364104,0.26256412,0.3249231,0.23630771,0.15425642,0.15425642,0.21333335,0.21989745,0.15425642,0.19364104,0.35446155,0.48574364,0.45292312,0.36758977,0.25928208,0.19692309,0.28882053,0.42994875,0.6170257,0.8467693,1.0502565,1.0896411,2.7667694,3.4067695,3.0949745,2.2055387,1.3751796,1.0371283,0.65641034,0.41682056,0.4135385,0.65969235,0.38728207,0.3446154,0.36102566,0.33476925,0.22646156,0.13456412,0.38400003,0.6465641,0.764718,0.761436,0.7220513,0.9517949,1.2077949,1.4736412,1.9790771,2.865231,3.9187696,3.8465643,2.9111798,2.934154,3.4100516,3.7907696,4.2141542,4.417641,3.7349746,3.2886157,3.1442053,3.2886157,3.6824617,4.273231,4.345436,5.169231,6.629744,7.312411,4.4898467,4.516103,4.522667,4.4406157,4.3290257,4.378257,7.4699492,6.5870776,4.4242053,2.7766156,2.553436,3.3805132,4.0434875,5.3366156,7.3616414,9.544206,10.118565,10.33518,9.642668,8.146052,6.6100516,5.920821,6.4656415,5.6451287,3.308308,1.7526156,1.6213335,1.9035898,1.723077,1.1158975,1.0108719,1.4506668,1.7985642,2.0578463,2.103795,1.6705642,1.591795,1.8018463,1.8116925,1.6869745,2.0578463,2.297436,1.9954873,1.5097437,1.4178462,2.5304618,1.8806155,1.5360001,1.2898463,0.97805136,0.4955898,0.33476925,0.256,0.24943592,0.29210258,0.35446155,0.14769232,0.36430773,0.5940513,0.6432821,0.5316923,0.3314872,0.11158975,0.0,0.0,0.0,0.0,0.013128206,0.068923086,0.14769232,0.18379489,0.14441027,0.072205134,0.04266667,0.06235898,0.068923086,0.036102567,0.026256412,0.01969231,0.016410258,0.02297436,0.02297436,0.032820515,0.04266667,0.052512825,0.09189744,0.08205129,0.07548718,0.068923086,0.059076928,0.04266667,0.03938462,0.049230773,0.052512825,0.036102567,0.0032820515,0.0032820515,0.0032820515,0.029538464,0.08861539,0.15097436,0.101743594,0.06564103,0.04266667,0.029538464,0.03938462,0.068923086,0.04266667,0.009846155,0.0,0.0,0.013128206,0.009846155,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016410258,0.029538464,0.026256412,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.049230773,0.118153855,0.14112821,0.101743594,0.032820515,0.013128206,0.013128206,0.006564103,0.006564103,0.013128206,0.013128206,0.052512825,0.14441027,0.20348719,0.18379489,0.06564103,0.052512825,0.08205129,0.12143591,0.14112821,0.14112821,0.128,0.18707694,0.21661541,0.18707694,0.14441027,0.16738462,0.23958977,0.26256412,0.20676924,0.12143591,0.049230773,0.03938462,0.21661541,0.47261542,0.4594872,0.2855385,0.20676924,0.21989745,0.27569234,0.27897438,0.2986667,0.36758977,0.43651286,0.5218462,0.7122052,0.71548724,0.7515898,0.7122052,0.5546667,0.27569234,0.14769232,0.0951795,0.068923086,0.04266667,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.07876924,0.14769232,0.16082053,0.08205129,0.068923086,0.059076928,0.059076928,0.07548718,0.1148718,0.15425642,0.13128206,0.118153855,0.14112821,0.15425642,0.16410258,0.12143591,0.068923086,0.029538464,0.013128206,0.006564103,0.016410258,0.029538464,0.04266667,0.026256412,0.029538464,0.14441027,0.27569234,0.3249231,0.21661541,0.26912823,0.32820517,0.3117949,0.23630771,0.21989745,0.25928208,0.38728207,0.5021539,0.571077,0.6268718,0.92225647,1.2668719,1.4769232,1.4998976,1.4375386,1.5753847,1.8707694,2.284308,2.6847181,2.8553848,2.7503593,2.9243078,3.3608208,3.8564105,4.007385,4.266667,5.408821,6.298257,6.560821,6.5805135,7.387898,9.235693,11.779283,13.157744,9.987283,8.812308,8.349539,7.5946674,6.163693,4.2863593,3.31159,3.0326157,3.4166157,4.3684106,5.737026,6.0980515,6.5247183,6.685539,6.3606157,5.431795,4.8738465,4.6244106,4.4898467,4.394667,4.4012313,4.4045134,3.4789746,2.5140514,1.9889232,1.9692309,2.3433847,2.0742567,1.6869745,1.3587693,0.9288206,1.1388719,1.8116925,2.5993848,3.387077,4.2830772,4.568616,4.4701543,4.197744,4.020513,4.269949,4.97559,5.674667,6.193231,6.4000006,6.1997952,5.7796926,5.169231,4.525949,3.948308,3.4658465,4.650667,6.3179493,7.762052,8.487385,8.192,6.3901544,4.0500517,1.9429746,0.5513847,0.072205134,0.059076928,0.04266667,0.02297436,0.009846155,0.016410258,0.006564103,0.0032820515,0.006564103,0.02297436,0.04594872,0.049230773,0.07876924,0.19692309,0.4135385,0.6826667,0.7187693,0.77456415,1.0994873,1.6180514,1.910154,2.048,1.9954873,1.9003079,1.7624617,1.4572309,1.3653334,1.3456411,1.3686155,1.6180514,2.481231,3.308308,3.2787695,2.8192823,2.2449234,1.7526156,2.0578463,4.092718,7.1154876,9.770667,10.089026,7.50277,6.6461544,6.885744,7.4929237,7.6274877,6.1505647,5.832206,4.886975,3.2032824,2.349949,2.1169233,2.3204105,3.8564105,7.53559,14.089848,20.187899,18.41559,17.253744,17.621334,12.911591,6.997334,4.84759,4.0369234,3.3476925,2.7602053,2.5698464,2.5961027,2.4320002,2.1234872,2.1956925,2.5829747,3.242667,3.945026,4.2338467,3.4330258,2.6486156,2.1398976,2.028308,2.4713848,3.6791797,4.8672824,5.973334,6.669129,6.770872,6.2227697,4.969026,4.2207184,3.754667,3.4658465,3.3608208,3.7842054,4.2830772,4.640821,5.044513,6.088206,8.306872,7.77518,7.532308,7.9294367,6.616616,4.2601027,3.515077,2.986667,2.0808206,0.98461545,1.2832822,1.8576412,2.231795,2.0611284,1.1454359,5.720616,5.464616,5.412103,5.3070774,5.4153852,6.5017443,7.1844106,7.39118,7.128616,6.409847,5.2480006,3.3936412,3.0687182,3.8662567,5.333334,6.957949,6.518154,6.262154,5.8420515,5.1200004,4.1813335,3.6430771,3.4264617,3.255795,3.0785644,3.0687182,3.370667,3.1474874,3.121231,3.2984617,2.9440002,1.9692309,1.3128207,1.0633847,1.3423591,2.3204105,3.4166157,4.0303593,4.092718,3.4822567,2.028308,1.1881026,1.0666667,1.4145643,1.8412309,1.8149745,1.4998976,1.2077949,1.0666667,1.014154,0.79425645,1.0010257,1.1257436,1.083077,0.8402052,0.4135385,0.25271797,0.16738462,0.13784617,0.13784617,0.13784617,0.19692309,0.3052308,0.39712822,0.43323082,0.39712822,0.43323082,0.40697438,0.3708718,0.33805132,0.28882053,0.15425642,0.08533334,0.04266667,0.016410258,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.013128206,0.02297436,0.02297436,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.04594872,0.02297436,0.016410258,0.016410258,0.02297436,0.04594872,0.02297436,0.016410258,0.02297436,0.032820515,0.04594872,0.02297436,0.08861539,0.16738462,0.21989745,0.24287182,0.29210258,0.7089231,0.90256417,0.79097444,0.7778462,0.8402052,0.5349744,0.30851284,0.35446155,0.6104616,0.7089231,0.4955898,0.39056414,0.49230772,0.56451285,1.5163078,2.4516926,1.9692309,0.46276927,0.12143591,0.79425645,1.2537436,1.020718,0.33805132,0.16738462,0.28882053,0.42994875,0.49230772,0.38400003,0.029538464,0.06564103,0.12143591,0.15753847,0.14112821,0.029538464,0.04266667,0.118153855,0.21661541,0.29210258,0.3052308,0.13456412,0.04594872,0.17394873,0.48902568,0.79425645,0.6235898,0.44307697,0.27897438,0.14441027,0.04594872,0.032820515,0.10502565,0.22646156,0.36102566,0.45620516,0.48246157,0.50543594,0.4201026,0.2986667,0.39712822,0.43323082,0.42338464,0.79097444,1.4506668,1.8149745,1.6082052,1.1716924,0.7253334,0.5349744,0.8992821,1.0108719,1.3292309,1.847795,2.1398976,1.3587693,3.1048207,4.125539,4.1878977,3.255795,1.5097437,0.6432821,0.23630771,0.11158975,0.13456412,0.18379489,0.19692309,0.20676924,0.21333335,0.190359,0.09189744,0.16410258,0.4955898,0.6104616,0.41682056,0.19692309,0.39384618,0.955077,1.394872,1.5885129,1.785436,1.9561027,1.9167181,2.1431797,2.8947694,4.2272825,4.7524104,4.1517954,4.2174363,4.8082056,3.8465643,3.0260515,2.7306669,2.865231,3.6627696,5.674667,5.5532312,3.9384618,2.878359,3.4527183,5.7829747,6.0160003,5.0477953,3.436308,2.0118976,1.8773335,1.0732309,0.98133343,1.4867693,2.4943593,3.9220517,5.7042055,7.3025646,8.884514,10.279386,10.985026,7.896616,7.200821,6.931693,6.2063594,5.218462,4.3027697,4.4767184,4.164923,3.0326157,1.9823592,1.7755898,1.7887181,1.6475899,1.2898463,0.9616411,1.1093334,1.4178462,2.1398976,2.793026,2.1825643,1.7920002,1.8937438,1.6935385,1.214359,1.3128207,1.2996924,1.1684103,0.97805136,0.73517954,0.380718,0.6498462,0.8730257,0.90256417,0.7253334,0.45620516,0.2986667,0.17723078,0.14112821,0.23302566,0.48902568,0.098461546,0.04594872,0.0951795,0.1148718,0.09189744,0.45620516,0.21989745,0.0,0.0,0.0,0.0,0.0,0.029538464,0.08533334,0.12143591,0.072205134,0.1148718,0.190359,0.2297436,0.16738462,0.04594872,0.006564103,0.006564103,0.02297436,0.04594872,0.0951795,0.13456412,0.10502565,0.055794876,0.15097436,0.24943592,0.29210258,0.2855385,0.23958977,0.15097436,0.09189744,0.059076928,0.03938462,0.026256412,0.016410258,0.016410258,0.016410258,0.032820515,0.08861539,0.19692309,0.101743594,0.03938462,0.016410258,0.016410258,0.016410258,0.06564103,0.049230773,0.01969231,0.0,0.0,0.013128206,0.02297436,0.02297436,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.02297436,0.026256412,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.016410258,0.009846155,0.0,0.0,0.013128206,0.016410258,0.02297436,0.026256412,0.016410258,0.052512825,0.08861539,0.101743594,0.07876924,0.029538464,0.01969231,0.068923086,0.16738462,0.25271797,0.2297436,0.25271797,0.29538465,0.30851284,0.256,0.12143591,0.049230773,0.07548718,0.18707694,0.3511795,0.5349744,0.48574364,0.41025645,0.35446155,0.3511795,0.4135385,0.508718,0.7187693,0.86974365,0.88287187,0.74830776,0.47917953,0.61374366,0.67282057,0.50543594,0.27569234,0.128,0.09189744,0.06564103,0.02297436,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.026256412,0.06564103,0.17066668,0.26584616,0.16738462,0.0951795,0.059076928,0.059076928,0.07876924,0.09189744,0.09189744,0.101743594,0.118153855,0.13128206,0.108307704,0.108307704,0.098461546,0.072205134,0.036102567,0.0,0.02297436,0.03938462,0.04594872,0.03938462,0.016410258,0.026256412,0.16738462,0.27897438,0.28882053,0.2297436,0.15425642,0.28225642,0.3708718,0.32820517,0.24287182,0.24287182,0.43651286,0.5218462,0.5021539,0.6859488,1.0896411,1.4572309,1.595077,1.5721027,1.6935385,1.9364104,2.2088206,2.5435898,2.806154,2.6847181,2.7470772,2.8356924,2.6289232,2.2613335,2.3335385,2.553436,2.8389745,3.1376412,3.4067695,3.6004105,5.5926156,8.165744,9.997129,9.216001,3.4198978,2.674872,2.7076926,2.9210258,2.868513,2.2580514,3.1967182,4.3585644,5.297231,5.76,5.674667,5.333334,5.7632823,6.0783596,5.8945646,5.3103595,4.565334,4.096,3.8071797,3.6791797,3.754667,3.7776413,3.0227695,2.225231,1.8576412,2.1530259,2.7995899,3.2065644,3.5380516,3.4921029,2.3204105,1.7690258,2.0545642,2.6453335,3.4527183,4.8049235,5.221744,5.2053337,5.0116925,4.854154,4.9296412,5.5762057,6.0028725,6.1078978,5.970052,5.858462,5.7009234,5.3398976,4.841026,4.2830772,3.7842054,5.602462,8.218257,10.292514,10.912822,9.5835905,7.030154,4.1124105,1.8248206,0.5874872,0.24287182,0.21989745,0.15097436,0.08205129,0.03938462,0.016410258,0.016410258,0.016410258,0.016410258,0.02297436,0.04594872,0.059076928,0.06235898,0.14112821,0.39056414,0.9156924,1.1946667,1.1651284,1.3784616,1.8970258,2.28759,2.1530259,1.7558975,1.3161026,1.0404103,1.1126155,1.394872,1.6213335,1.7427694,1.9331284,2.5796926,4.519385,5.802667,6.117744,5.2414365,3.0227695,3.045744,3.170462,4.020513,5.8912826,8.759795,5.6943593,5.927385,8.228104,11.254155,13.548308,10.266257,10.8996935,10.026668,6.2194877,2.044718,1.7624617,2.2613335,3.0293336,3.8367183,4.716308,5.412103,5.8157954,6.0225644,6.038975,5.7829747,5.172513,4.3684106,3.5872824,3.006359,2.7602053,2.481231,2.100513,1.7591796,1.6246156,1.8937438,2.2580514,2.7536411,3.3805132,3.7874875,3.249231,2.5895386,2.15959,2.038154,2.2514873,2.7766156,4.069744,5.110154,5.687795,5.684513,5.0510774,5.464616,4.716308,3.515077,2.409026,1.785436,2.0545642,3.4592824,4.903385,5.868308,6.3934364,6.8955903,7.2927184,7.1122055,6.2884107,5.1889234,4.197744,3.6758976,3.0424619,2.1464617,1.2668719,0.99774367,1.3423591,1.591795,1.5097437,1.3259488,3.511795,4.604718,5.618872,6.442667,7.0892315,7.6964107,7.958975,7.893334,7.6964107,7.3649235,6.7150774,5.648411,5.622154,5.2742567,4.4274874,4.076308,4.076308,4.397949,4.5456414,4.352,3.9975388,3.5577438,3.1770258,2.868513,2.5993848,2.2744617,2.3729234,2.5731285,2.8455386,3.2262566,3.8006158,3.4297438,2.5796926,1.6213335,0.9353847,0.9156924,1.6836925,2.7766156,3.9253337,4.7950773,4.9821544,3.0194874,1.7985642,1.2537436,1.204513,1.3751796,1.4211283,1.6738462,1.9003079,1.9068719,1.5491283,1.1323078,0.8172308,0.64000005,0.60389745,0.6432821,0.6498462,0.50543594,0.32820517,0.20020515,0.16082053,0.25271797,0.30851284,0.32164106,0.29538465,0.24943592,0.256,0.23630771,0.21989745,0.20676924,0.16738462,0.11158975,0.07548718,0.04266667,0.016410258,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.016410258,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.032820515,0.026256412,0.016410258,0.01969231,0.032820515,0.029538464,0.013128206,0.0032820515,0.006564103,0.009846155,0.032820515,0.15753847,0.2986667,0.38728207,0.35446155,0.49230772,1.1257436,1.273436,0.8992821,0.92553854,0.8598975,0.49230772,0.26584616,0.31507695,0.46276927,0.4135385,0.24615386,0.12143591,0.11158975,0.18707694,0.39712822,0.56451285,0.58092314,1.1093334,3.6004105,2.4451284,1.4473847,0.7811283,0.42994875,0.18051283,0.54482055,0.8730257,0.9878975,0.7811283,0.20020515,0.26584616,0.26256412,0.2855385,0.39056414,0.60389745,0.7417436,0.5513847,0.86317956,1.7296412,2.4057438,0.58420515,0.098461546,0.16082053,0.34133336,0.5481026,0.60389745,0.45620516,0.3314872,0.2986667,0.28882053,0.318359,0.4266667,0.4594872,0.4004103,0.36102566,0.33476925,0.33476925,0.24943592,0.12143591,0.14112821,0.2855385,0.44964105,0.58420515,0.67938465,0.7417436,0.65969235,0.5415385,0.45620516,0.5546667,1.0469744,1.0305642,1.083077,1.2996924,1.5983591,1.7362052,2.4484105,2.674872,2.5961027,2.5042052,2.8291285,1.5622566,0.77456415,0.3511795,0.18707694,0.19692309,0.16738462,0.14769232,0.12471796,0.101743594,0.09189744,0.049230773,0.4135385,0.7187693,0.7778462,0.67282057,0.41025645,0.446359,0.60389745,0.8008206,1.0666667,1.5195899,2.4057438,2.5829747,2.4352822,3.8728209,5.277539,4.601436,3.4494362,2.934154,3.698872,3.623385,2.3630772,1.529436,1.529436,1.5622566,1.5885129,1.9364104,3.3444104,5.874872,8.907488,8.192,6.226052,4.013949,2.4681027,2.4024618,2.7667694,3.9647183,5.796103,7.8506675,9.524513,10.016821,10.548513,10.824206,10.505847,9.193027,8.769642,8.838565,8.457847,7.325539,5.7796926,4.640821,3.879385,3.1540515,2.4516926,2.1070771,2.103795,1.4867693,1.0338463,1.0272821,1.2537436,1.4309745,1.4473847,1.4703591,1.5261539,1.5097437,1.657436,1.5130258,1.332513,1.1158975,0.6301539,0.8598975,1.3751796,1.2274873,0.47261542,0.18707694,0.33805132,0.56123084,0.78769237,0.86974365,0.5907693,0.31507695,0.1148718,0.029538464,0.04594872,0.098461546,0.07876924,0.13456412,0.17723078,0.20020515,0.27569234,0.2986667,0.19692309,0.072205134,0.0,0.0,0.0,0.0,0.006564103,0.02297436,0.049230773,0.24287182,0.33476925,0.318359,0.21661541,0.059076928,0.06235898,0.03938462,0.01969231,0.02297436,0.04594872,0.0951795,0.098461546,0.07548718,0.068923086,0.128,0.19692309,0.25271797,0.26584616,0.2297436,0.15097436,0.09189744,0.0951795,0.10502565,0.101743594,0.101743594,0.09189744,0.08861539,0.07876924,0.068923086,0.101743594,0.08205129,0.068923086,0.055794876,0.036102567,0.016410258,0.026256412,0.02297436,0.016410258,0.009846155,0.0,0.013128206,0.009846155,0.0032820515,0.0032820515,0.0,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.006564103,0.0032820515,0.0,0.013128206,0.01969231,0.013128206,0.013128206,0.032820515,0.06564103,0.0951795,0.098461546,0.06235898,0.04266667,0.029538464,0.03938462,0.072205134,0.12143591,0.08533334,0.04594872,0.02297436,0.009846155,0.0,0.0032820515,0.0032820515,0.0032820515,0.006564103,0.0032820515,0.01969231,0.059076928,0.17394873,0.33476925,0.4201026,0.25271797,0.17723078,0.14769232,0.13456412,0.13128206,0.17394873,0.27241027,0.3249231,0.29210258,0.19692309,0.15097436,0.13456412,0.26584616,0.49887183,0.6432821,0.58420515,0.45620516,0.39056414,0.44307697,0.58420515,1.0043077,1.401436,1.3489232,0.9124103,0.6498462,0.508718,0.512,0.43651286,0.256,0.14112821,0.072205134,0.055794876,0.04594872,0.02297436,0.0,0.0,0.0,0.0032820515,0.016410258,0.026256412,0.009846155,0.055794876,0.15097436,0.24287182,0.25271797,0.11158975,0.059076928,0.059076928,0.07876924,0.09189744,0.06235898,0.07876924,0.09189744,0.08861539,0.0951795,0.15425642,0.128,0.08205129,0.052512825,0.072205134,0.128,0.08205129,0.03938462,0.032820515,0.026256412,0.068923086,0.18051283,0.3052308,0.36102566,0.23958977,0.21661541,0.28225642,0.27241027,0.18051283,0.18379489,0.27241027,0.54482055,1.0043077,1.4736412,1.5786668,1.8149745,2.1103592,2.3368206,2.4418464,2.425436,2.4746668,2.5665643,2.681436,2.6157951,1.9790771,1.9200002,2.0020514,2.044718,2.0184617,2.041436,2.9144619,2.989949,2.9505644,3.3575387,4.6276927,7.0859494,8.78277,8.772923,6.875898,3.6758976,3.0949745,2.8192823,2.6715899,2.5961027,2.6486156,3.626667,5.0018463,6.1538467,6.665847,6.3343596,5.865026,6.173539,6.1997952,5.5991797,4.7622566,4.0369234,3.636513,3.131077,2.5042052,2.166154,2.2219489,2.2153847,1.9790771,1.7099489,1.9429746,2.9243078,3.4658465,3.5183592,3.4560003,4.089436,4.388103,4.3651285,4.2929235,4.3618464,4.673641,4.716308,4.594872,4.6145644,5.0149746,5.979898,6.5083084,6.7150774,6.5083084,5.9503593,5.2742567,4.9985647,5.172513,5.5072823,5.914257,6.518154,8.651488,9.957745,10.624001,10.489437,9.081436,5.661539,2.9505644,1.3226668,0.761436,0.8795898,0.69907695,0.47261542,0.26256412,0.11158975,0.026256412,0.026256412,0.01969231,0.016410258,0.01969231,0.032820515,0.04594872,0.04266667,0.072205134,0.18707694,0.4266667,0.69907695,0.9288206,1.3193847,1.8149745,2.1169233,2.3368206,2.1924105,1.8838975,1.6377437,1.7132308,1.9232821,2.0217438,1.8904617,1.6804104,1.8084104,3.564308,4.4767184,4.4832826,3.9023592,3.4494362,3.7349746,3.4133337,3.062154,3.05559,3.570872,2.937436,3.498667,4.532513,6.058667,8.861539,11.047385,9.885539,7.702975,5.6254363,3.5577438,2.9538465,2.5961027,2.8521028,3.570872,4.066462,4.0500517,4.2535386,5.0018463,5.976616,6.196513,5.3924108,4.2469745,3.2623591,2.6978464,2.5895386,2.5435898,2.294154,1.8937438,1.529436,1.5130258,1.7033848,1.9429746,2.3204105,2.6847181,2.6157951,2.103795,1.8116925,1.8313848,2.1300514,2.556718,3.5774362,4.525949,5.139693,5.3792825,5.428513,5.366154,4.923077,4.1452312,3.1409233,2.0775387,2.044718,2.6912823,3.698872,4.841026,5.989744,7.194257,7.506052,6.688821,4.9985647,3.1967182,2.6584618,2.2055387,1.6377437,1.0338463,0.7417436,0.892718,1.591795,2.1300514,2.100513,1.401436,4.086154,4.7950773,5.910975,6.8627696,7.397744,7.5552826,7.5913854,7.5618467,7.529026,7.4075904,6.9809237,6.3901544,6.36718,6.196513,5.5958977,4.70318,4.893539,5.2053337,5.1200004,4.571898,3.9253337,3.2886157,2.9768207,2.861949,2.7208207,2.2219489,1.8379488,1.8281027,2.0184617,2.3696413,2.9702566,3.7251284,3.5971284,2.8717952,1.8510771,0.8566154,0.8598975,1.6344616,2.6518977,3.5807183,4.312616,3.6758976,2.7175386,1.8215386,1.2307693,1.0108719,1.0272821,1.273436,1.6443079,1.9364104,1.8313848,1.3817437,1.0666667,0.86646163,0.79425645,0.90256417,0.88615394,0.6695385,0.44964105,0.34133336,0.38728207,0.43323082,0.40369233,0.3314872,0.24943592,0.17723078,0.14112821,0.118153855,0.108307704,0.10502565,0.08205129,0.068923086,0.052512825,0.032820515,0.016410258,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.013128206,0.016410258,0.016410258,0.013128206,0.009846155,0.009846155,0.0032820515,0.0032820515,0.009846155,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.009846155,0.009846155,0.009846155,0.016410258,0.026256412,0.026256412,0.016410258,0.02297436,0.013128206,0.0032820515,0.0,0.0032820515,0.009846155,0.02297436,0.08861539,0.19692309,0.2986667,0.318359,0.47589746,0.90256417,1.1716924,1.1552821,1.017436,0.7220513,0.36758977,0.23630771,0.34133336,0.41682056,0.3249231,0.20348719,0.10502565,0.055794876,0.06564103,0.38728207,0.48246157,0.47261542,0.7187693,1.8149745,1.5819489,1.3686155,1.2471796,1.1355898,0.82379496,0.571077,0.6235898,0.7220513,0.6859488,0.41682056,0.41025645,0.3446154,0.3249231,0.40369233,0.574359,0.63343596,0.46933338,0.83035904,1.6705642,2.1333334,0.5218462,0.101743594,0.11158975,0.17723078,0.3249231,0.46276927,0.380718,0.318359,0.380718,0.56123084,0.7581539,0.90912825,0.77456415,0.48902568,0.54482055,0.7220513,0.7778462,0.51856416,0.13456412,0.17723078,0.3052308,0.38400003,0.40369233,0.35446155,0.26256412,0.29538465,0.36758977,0.45620516,0.574359,0.79097444,0.7253334,0.98461545,1.5983591,2.3466668,2.7569232,2.100513,1.6640002,1.5622566,1.8740515,2.6289232,2.2416413,1.5458462,0.83035904,0.33476925,0.22646156,0.17394873,0.16410258,0.15753847,0.118153855,0.036102567,0.052512825,0.2231795,0.36758977,0.39712822,0.318359,0.3117949,0.3511795,0.39712822,0.46276927,0.58420515,0.85005134,1.2209232,1.2865642,1.3423591,2.3729234,3.373949,2.5993848,1.7755898,1.7887181,2.6551797,2.8225644,2.0676925,1.8018463,2.0841026,1.6147693,1.7493335,2.7831798,4.4734364,6.170257,6.7971287,5.9536414,4.969026,4.4340515,4.906667,6.9087186,9.061745,11.648001,14.352411,15.937642,14.230975,13.850258,12.950975,11.434668,9.67877,8.4972315,8.28718,8.165744,7.7357955,6.8365135,5.5532312,4.6802053,3.5840003,2.6190772,2.0676925,2.1530259,2.0118976,1.6475899,1.3620514,1.2537436,1.2077949,1.4211283,1.3620514,1.211077,1.1158975,1.204513,1.2438976,1.1290257,1.0732309,1.0371283,0.7318975,0.51856416,0.90584624,0.8763078,0.33476925,0.108307704,0.24615386,0.62030774,0.9485129,1.086359,1.0568206,0.78769237,0.37743592,0.12143591,0.08861539,0.118153855,0.14112821,0.22646156,0.34789747,0.4660513,0.5481026,0.42338464,0.24943592,0.09189744,0.0,0.0,0.0,0.0,0.0,0.006564103,0.029538464,0.24287182,0.33805132,0.3052308,0.17723078,0.03938462,0.16410258,0.24615386,0.25928208,0.20348719,0.08205129,0.190359,0.19364104,0.15097436,0.1148718,0.10502565,0.10502565,0.118153855,0.13128206,0.12471796,0.07876924,0.055794876,0.072205134,0.09189744,0.10502565,0.10502565,0.09189744,0.10502565,0.10502565,0.08861539,0.0951795,0.118153855,0.13456412,0.15425642,0.15753847,0.08861539,0.02297436,0.013128206,0.013128206,0.0032820515,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0032820515,0.006564103,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.0032820515,0.013128206,0.026256412,0.032820515,0.032820515,0.06564103,0.098461546,0.108307704,0.0951795,0.06564103,0.04266667,0.032820515,0.04266667,0.06564103,0.08861539,0.07548718,0.068923086,0.06564103,0.059076928,0.04594872,0.029538464,0.016410258,0.009846155,0.009846155,0.01969231,0.02297436,0.032820515,0.098461546,0.2231795,0.39056414,0.36758977,0.35446155,0.3314872,0.26584616,0.13456412,0.16082053,0.20676924,0.24615386,0.2855385,0.3708718,0.318359,0.23302566,0.26256412,0.42338464,0.58092314,0.45292312,0.43651286,0.43323082,0.43323082,0.48902568,0.7318975,0.93866676,0.8795898,0.6301539,0.571077,0.76800007,0.7450257,0.5481026,0.28225642,0.12471796,0.068923086,0.03938462,0.02297436,0.013128206,0.01969231,0.026256412,0.026256412,0.036102567,0.055794876,0.06564103,0.049230773,0.068923086,0.101743594,0.13128206,0.13784617,0.07548718,0.06564103,0.0951795,0.13456412,0.15425642,0.2297436,0.29210258,0.26256412,0.16082053,0.101743594,0.12143591,0.10502565,0.07876924,0.068923086,0.09189744,0.0951795,0.06564103,0.03938462,0.032820515,0.049230773,0.068923086,0.12471796,0.20348719,0.26584616,0.26256412,0.20676924,0.21333335,0.20348719,0.17066668,0.18707694,0.26584616,0.49887183,0.8336411,1.1355898,1.1782565,1.467077,1.9003079,2.284308,2.5271797,2.6551797,2.6683078,2.7175386,2.6453335,2.3893335,1.9922053,1.9232821,1.9626669,2.0644104,2.2383592,2.537026,3.442872,3.8432825,3.9286156,4.197744,5.4416413,7.2631803,8.195283,7.6274877,5.9536414,4.5522056,4.7491283,5.0116925,4.6145644,3.7874875,3.698872,4.1025643,4.7294364,5.2578464,5.6320004,6.0685134,6.183385,6.301539,5.920821,5.0674877,4.312616,3.9942567,3.8006158,3.4822567,2.9735386,2.4024618,2.4188719,2.1366155,1.6869745,1.5458462,2.5337439,3.945026,4.1156926,3.8629746,3.95159,5.0904617,6.262154,6.560821,6.36718,5.9667697,5.5532312,5.2644105,4.9329233,4.8147697,5.1331286,6.0750775,7.076103,7.39118,7.131898,6.5312824,5.940513,6.0028725,6.7610264,7.6898465,8.536616,9.298052,10.115283,10.049642,9.984001,9.714872,7.939283,4.4701543,2.172718,0.955077,0.574359,0.65312827,0.5152821,0.43323082,0.2855385,0.08861539,0.02297436,0.029538464,0.02297436,0.013128206,0.009846155,0.02297436,0.03938462,0.04266667,0.04594872,0.07876924,0.17723078,0.3708718,0.5677949,0.85005134,1.1979488,1.4802053,1.7493335,1.8018463,1.7558975,1.7362052,1.8904617,2.0841026,2.0644104,1.8084104,1.5425643,1.7263591,3.0490258,3.754667,3.8531284,3.6004105,3.501949,3.5840003,3.5216413,3.3542566,3.0916924,2.7044106,2.422154,2.6354873,2.937436,3.5610259,5.356308,8.402052,8.707283,7.6767187,6.2162056,4.7425647,3.7940516,3.6594875,4.092718,4.768821,5.297231,4.6933336,4.138667,4.1878977,4.7950773,5.3037953,4.7556925,3.9548721,3.2328207,2.7995899,2.7503593,2.8291285,2.809436,2.6912823,2.487795,2.2350771,2.1530259,2.1070771,2.2022567,2.3368206,2.172718,1.6311796,1.4473847,1.591795,1.9790771,2.4484105,3.1376412,4.017231,4.8377438,5.3924108,5.5236926,5.661539,5.618872,5.0543594,3.9876926,2.802872,2.4418464,2.5862565,3.1540515,4.0303593,5.0576415,5.9602056,6.3606157,5.861744,4.4996924,2.7634873,2.03159,1.7427694,1.4441026,1.0305642,0.7384616,0.86317956,1.5360001,2.3991797,2.9407182,2.5009232,6.009436,6.157129,6.4722056,6.5017443,6.2162056,5.986462,6.1341543,6.3474874,6.7249236,7.1647186,7.3747697,6.806975,6.4032826,6.3179493,6.3606157,5.98318,5.730462,6.180103,6.308103,5.7829747,4.97559,4.4406157,3.7382567,3.2131286,2.878359,2.3991797,1.7920002,1.4900514,1.4605129,1.6410258,1.9495386,2.9111798,3.4658465,3.4297438,2.7766156,1.6278975,1.0929232,1.2898463,1.6804104,2.0644104,2.5862565,3.0687182,2.9078977,2.3794873,1.7591796,1.3161026,1.024,0.88287187,0.99774367,1.3128207,1.591795,1.6082052,1.6311796,1.6016412,1.467077,1.1913847,1.0272821,0.82379496,0.636718,0.5152821,0.5218462,0.50543594,0.43323082,0.33476925,0.23630771,0.14112821,0.08861539,0.072205134,0.068923086,0.07548718,0.07548718,0.09189744,0.08533334,0.06564103,0.03938462,0.016410258,0.006564103,0.006564103,0.009846155,0.013128206,0.013128206,0.026256412,0.029538464,0.026256412,0.02297436,0.02297436,0.026256412,0.01969231,0.026256412,0.04594872,0.03938462,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.009846155,0.013128206,0.02297436,0.009846155,0.01969231,0.01969231,0.009846155,0.009846155,0.0032820515,0.0,0.0,0.0032820515,0.016410258,0.009846155,0.026256412,0.08861539,0.18051283,0.24943592,0.43323082,0.67610264,0.9682052,1.1618463,0.9682052,0.60389745,0.3117949,0.21989745,0.29538465,0.36430773,0.34789747,0.29210258,0.2231795,0.15753847,0.13128206,0.47917953,0.54482055,0.43651286,0.26256412,0.13784617,0.702359,1.2077949,1.4769232,1.4276924,1.0568206,0.6268718,0.4660513,0.44964105,0.47261542,0.47261542,0.47589746,0.5481026,0.60389745,0.6104616,0.60389745,0.54482055,0.48246157,0.7056411,1.0962052,1.1388719,0.3117949,0.14441027,0.14441027,0.12471796,0.20020515,0.3446154,0.36430773,0.49887183,0.764718,0.9714873,1.0601027,1.0469744,0.81394875,0.64000005,1.1946667,1.4276924,1.1848207,0.64000005,0.128,0.15753847,0.27569234,0.3249231,0.3052308,0.24615386,0.20020515,0.3314872,0.49887183,0.6498462,0.7187693,0.636718,0.5973334,0.9124103,1.5589745,2.3236926,2.7995899,1.6508719,1.2438976,1.4998976,2.176,2.878359,2.8980515,2.2022567,1.2865642,0.55794877,0.33476925,0.31507695,0.30194873,0.27897438,0.21333335,0.072205134,0.27897438,0.34133336,0.33805132,0.30194873,0.20020515,0.18707694,0.26912823,0.39384618,0.512,0.5874872,0.48246157,0.4135385,0.5021539,0.8008206,1.2832822,1.5655385,0.9682052,0.7220513,1.1158975,1.4834872,1.6180514,1.6705642,2.166154,2.8356924,2.609231,2.665026,3.3312824,4.2141542,4.706462,3.9942567,4.1485133,5.5630774,8.825437,12.987078,15.55036,16.219898,16.836924,18.225233,19.183592,16.505438,15.195899,13.298873,11.1294365,9.373539,9.101129,8.03118,7.276308,6.8266673,6.5050263,5.9569235,5.605744,4.4438977,3.117949,2.162872,1.9823592,1.8609232,1.7788719,1.654154,1.4703591,1.270154,1.657436,1.6738462,1.4572309,1.1749744,0.99774367,0.8598975,0.9321026,1.0043077,0.9485129,0.7089231,0.26256412,0.38400003,0.42994875,0.23630771,0.108307704,0.20676924,0.56123084,0.86646163,1.020718,1.142154,0.9616411,0.5284103,0.21661541,0.13784617,0.13784617,0.1148718,0.2231795,0.3511795,0.5349744,0.9353847,1.0075898,0.6071795,0.19692309,0.0,0.0,0.0,0.0,0.0,0.013128206,0.06235898,0.18707694,0.25928208,0.27241027,0.24287182,0.2100513,0.36430773,0.4955898,0.54482055,0.45292312,0.17394873,0.27569234,0.27569234,0.20348719,0.1148718,0.07876924,0.049230773,0.029538464,0.029538464,0.032820515,0.01969231,0.01969231,0.032820515,0.052512825,0.06564103,0.06564103,0.055794876,0.068923086,0.07876924,0.07548718,0.07548718,0.09189744,0.10502565,0.128,0.14112821,0.08205129,0.016410258,0.006564103,0.006564103,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0,0.006564103,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0032820515,0.009846155,0.016410258,0.026256412,0.04266667,0.055794876,0.052512825,0.06564103,0.07876924,0.07548718,0.055794876,0.04266667,0.029538464,0.02297436,0.029538464,0.032820515,0.026256412,0.03938462,0.055794876,0.06564103,0.06564103,0.052512825,0.04594872,0.04594872,0.049230773,0.06235898,0.07876924,0.068923086,0.03938462,0.029538464,0.08205129,0.23302566,0.3249231,0.37415388,0.38400003,0.3314872,0.19692309,0.20676924,0.2100513,0.21333335,0.23630771,0.30851284,0.26584616,0.20020515,0.19692309,0.26584616,0.36102566,0.28225642,0.35774362,0.4266667,0.4397949,0.45620516,0.5415385,0.5940513,0.60061544,0.574359,0.54482055,0.73517954,0.67610264,0.47589746,0.24287182,0.0951795,0.06235898,0.03938462,0.016410258,0.0032820515,0.02297436,0.036102567,0.03938462,0.04594872,0.059076928,0.06235898,0.06235898,0.098461546,0.12143591,0.1148718,0.08205129,0.072205134,0.13128206,0.21333335,0.28225642,0.30851284,0.39712822,0.41682056,0.35446155,0.23630771,0.15097436,0.108307704,0.09189744,0.09189744,0.0951795,0.09189744,0.055794876,0.052512825,0.055794876,0.052512825,0.06564103,0.06235898,0.06564103,0.08533334,0.118153855,0.17066668,0.128,0.118153855,0.13128206,0.14769232,0.15097436,0.20020515,0.34133336,0.46933338,0.5677949,0.6826667,1.1684103,1.7132308,2.2088206,2.605949,2.9243078,2.8947694,2.9210258,2.8422565,2.6256413,2.3696413,2.3401027,2.359795,2.4713848,2.737231,3.2262566,3.8531284,4.5095387,4.97559,5.353026,6.0750775,6.7249236,6.7610264,6.0619493,5.0477953,4.663795,5.3858466,6.560821,6.7183595,5.8945646,5.6385646,6.373744,6.0160003,5.3924108,4.969026,4.844308,4.9394875,4.9394875,4.634257,4.1517954,3.945026,4.194462,4.210872,4.2469745,4.2469745,3.8465643,3.6660516,3.0129232,2.3958976,2.3204105,3.2820516,4.5554876,4.5489235,4.332308,4.6178465,5.756718,7.069539,7.387898,7.171283,6.8004107,6.5739493,6.3901544,6.038975,5.874872,6.0652313,6.5772314,7.532308,8.201847,8.257642,7.893334,7.8473854,8.054154,8.713847,9.67877,10.65354,11.221334,10.217027,9.416205,9.074872,8.503796,6.0685134,3.186872,1.4703591,0.60389745,0.30851284,0.35446155,0.5481026,0.5481026,0.34133336,0.06564103,0.02297436,0.02297436,0.01969231,0.013128206,0.006564103,0.009846155,0.03938462,0.059076928,0.07548718,0.0951795,0.13456412,0.21661541,0.318359,0.44307697,0.58420515,0.7187693,0.8795898,1.0436924,1.2209232,1.3981539,1.5425643,1.6968206,1.847795,1.847795,1.7952822,2.0086155,3.0654361,4.0467696,4.4110775,4.1189747,3.623385,3.373949,3.515077,3.7152824,3.626667,2.8882053,2.5140514,2.5632823,2.6551797,2.7700515,3.2623591,5.3070774,7.4699492,9.705027,10.679795,7.762052,4.70318,3.8301542,4.2929235,5.3234878,6.2490263,5.366154,4.2962055,3.6758976,3.7087183,4.1682053,3.9089234,3.4724104,3.0326157,2.7241027,2.6289232,2.6584618,2.7076926,2.7437952,2.6880002,2.4057438,2.1103592,1.9593848,1.9298463,1.9068719,1.7033848,1.3161026,1.2504616,1.4408206,1.8281027,2.349949,3.0916924,4.056616,4.969026,5.543385,5.481026,6.088206,6.747898,6.7971287,5.933949,4.197744,2.989949,2.858667,3.2032824,3.6758976,4.1911798,4.522667,4.7458467,4.4701543,3.623385,2.428718,1.8937438,1.8313848,1.7263591,1.4441026,1.2340513,1.1585642,1.4867693,2.3401027,3.2131286,2.9801028,8.280616,8.090257,7.1220517,5.858462,4.7950773,4.450462,4.706462,4.6966157,5.097026,6.0061545,6.951385,6.4623594,5.9634876,5.7731285,5.9634876,6.3442054,5.5236926,6.121026,6.7774363,6.8365135,6.3212314,6.0947695,4.854154,3.6036925,2.802872,2.3630772,1.8773335,1.5195899,1.3522053,1.3587693,1.4342566,1.7329233,2.5140514,3.2098465,3.43959,2.9965131,2.2482052,1.8642052,1.6508719,1.5327181,1.5655385,1.8674873,2.2153847,2.3401027,2.1792822,1.8543591,1.3292309,0.86317956,0.5973334,0.6301539,1.0075898,1.463795,1.7985642,1.9922053,1.913436,1.3128207,1.0962052,0.98133343,0.8566154,0.7122052,0.6301539,0.49230772,0.38728207,0.3117949,0.24615386,0.16738462,0.12471796,0.11158975,0.1148718,0.13128206,0.15425642,0.18379489,0.17723078,0.14441027,0.09189744,0.032820515,0.029538464,0.026256412,0.032820515,0.04594872,0.049230773,0.04266667,0.049230773,0.04594872,0.036102567,0.032820515,0.03938462,0.029538464,0.049230773,0.07876924,0.06564103,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.026256412,0.016410258,0.006564103,0.0,0.0,0.0032820515,0.0032820515,0.0032820515,0.0032820515,0.0032820515,0.013128206,0.0032820515,0.01969231,0.059076928,0.12143591,0.20676924,0.4135385,0.6104616,0.7778462,0.90584624,0.9616411,0.6432821,0.39384618,0.23630771,0.19692309,0.26912823,0.42994875,0.47589746,0.42994875,0.33476925,0.27241027,0.3708718,0.27569234,0.15097436,0.11158975,0.2231795,0.5415385,0.9714873,1.204513,1.1158975,0.7384616,0.636718,0.50543594,0.42338464,0.4266667,0.5284103,0.6498462,0.9124103,1.014154,0.892718,0.7318975,0.6498462,0.6465641,0.65969235,0.6235898,0.45292312,0.20348719,0.19692309,0.20348719,0.16738462,0.17066668,0.28882053,0.44964105,0.86317956,1.3456411,1.3029745,1.0469744,0.81394875,0.6104616,0.7417436,1.7952822,1.8379488,1.1191796,0.40369233,0.06564103,0.08205129,0.2297436,0.34133336,0.318359,0.23630771,0.36758977,0.574359,0.7778462,0.94523084,0.9911796,0.7778462,0.7811283,0.9321026,1.211077,1.5819489,2.0184617,1.2603078,1.4178462,2.28759,3.508513,4.5390773,3.5905645,2.5665643,1.6311796,0.93866676,0.63343596,0.955077,0.9321026,0.7581539,0.5415385,0.32820517,0.62030774,0.65641034,0.60389745,0.54482055,0.45620516,0.20020515,0.2855385,0.56451285,0.8598975,0.95835906,0.47589746,0.44964105,0.62030774,0.8008206,0.8763078,0.77128214,0.6235898,0.6432821,0.7778462,0.71548724,0.7253334,1.270154,2.0873847,2.7963078,2.8750772,2.6322052,2.4418464,2.4582565,2.6551797,2.8356924,4.466872,8.100103,15.195899,22.646156,22.770874,19.495386,16.807386,16.351181,17.404718,16.869745,14.729847,12.393026,10.518975,9.573745,9.83959,8.438154,7.4207187,6.8660517,6.764308,6.994052,6.741334,5.4482055,3.876103,2.5764105,1.8904617,1.8215386,1.8116925,1.8871796,1.9429746,1.7493335,2.1267693,2.1267693,1.8576412,1.529436,1.4408206,1.3226668,1.3423591,1.204513,0.8369231,0.40697438,0.101743594,0.13456412,0.2297436,0.26256412,0.28225642,0.24943592,0.41682056,0.64000005,0.8172308,0.8730257,0.69907695,0.4397949,0.23630771,0.14441027,0.108307704,0.14769232,0.20676924,0.20348719,0.32820517,1.0601027,1.4506668,0.9189744,0.30194873,0.006564103,0.0032820515,0.0,0.0,0.009846155,0.04266667,0.12143591,0.16082053,0.21661541,0.34133336,0.49887183,0.5677949,0.65312827,0.78769237,0.81394875,0.65312827,0.3052308,0.2986667,0.25928208,0.17066668,0.072205134,0.072205134,0.052512825,0.029538464,0.009846155,0.0,0.0,0.0,0.013128206,0.04266667,0.06235898,0.036102567,0.01969231,0.016410258,0.02297436,0.029538464,0.026256412,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.006564103,0.0,0.0,0.029538464,0.04266667,0.052512825,0.059076928,0.049230773,0.029538464,0.026256412,0.029538464,0.026256412,0.016410258,0.013128206,0.013128206,0.013128206,0.009846155,0.0,0.009846155,0.01969231,0.02297436,0.02297436,0.013128206,0.032820515,0.06235898,0.09189744,0.118153855,0.15097436,0.15425642,0.118153855,0.08861539,0.101743594,0.17723078,0.23630771,0.27241027,0.29210258,0.29210258,0.27569234,0.26584616,0.30194873,0.2986667,0.21661541,0.06235898,0.04594872,0.07548718,0.118153855,0.15097436,0.13784617,0.21661541,0.29538465,0.38400003,0.48574364,0.5874872,0.7975385,0.81394875,0.8008206,0.761436,0.5546667,0.43323082,0.30851284,0.18379489,0.08205129,0.026256412,0.036102567,0.03938462,0.02297436,0.0032820515,0.013128206,0.02297436,0.02297436,0.026256412,0.026256412,0.01969231,0.03938462,0.11158975,0.17723078,0.20676924,0.19364104,0.21661541,0.3314872,0.42338464,0.45620516,0.47589746,0.45292312,0.35446155,0.27897438,0.24943592,0.20020515,0.128,0.108307704,0.118153855,0.12471796,0.098461546,0.059076928,0.06235898,0.068923086,0.06564103,0.06564103,0.052512825,0.026256412,0.013128206,0.013128206,0.016410258,0.04266667,0.04594872,0.059076928,0.07876924,0.068923086,0.101743594,0.16082053,0.20348719,0.27569234,0.5152821,1.270154,1.8904617,2.5009232,3.1113849,3.6135387,3.242667,3.2098465,3.2886157,3.242667,2.8422565,2.8389745,2.793026,2.878359,3.1737437,3.6660516,4.0500517,4.8049235,5.671385,6.3376417,6.4623594,5.9470773,5.2480006,4.71959,4.5423594,4.706462,5.2348723,6.426257,7.0465646,6.948103,7.069539,8.792616,7.8539495,6.426257,5.356308,4.1813335,3.892513,3.8400004,3.9844105,4.2535386,4.5489235,5.0182567,5.100308,5.3694363,5.7534366,5.536821,5.0051284,4.33559,4.027077,4.066462,3.945026,4.4734364,4.630975,4.7655387,5.2480006,6.485334,7.3091288,7.1581545,6.669129,6.4754877,7.1909747,7.53559,7.6668725,8.03118,8.63836,9.055181,9.265231,9.882257,10.056206,9.862565,10.305642,10.443488,10.545232,11.0145645,11.657847,11.680821,9.360411,8.441437,7.8834877,6.6461544,3.692308,1.8215386,0.7844103,0.30851284,0.20676924,0.39056414,0.90584624,0.8533334,0.5021539,0.13128206,0.036102567,0.016410258,0.013128206,0.016410258,0.016410258,0.006564103,0.036102567,0.07548718,0.118153855,0.16082053,0.190359,0.18707694,0.23958977,0.27569234,0.26912823,0.24615386,0.3511795,0.57764107,0.8205129,0.97805136,0.9419488,0.9747693,1.3817437,1.8281027,2.2088206,2.6617439,3.892513,5.3037953,5.7009234,4.9132314,3.7973337,3.3050258,3.3509746,3.564308,3.5249233,2.7503593,2.5600002,2.7963078,3.006359,2.9801028,2.7733335,3.5052311,5.8092313,10.282667,13.991385,10.469745,5.4547696,3.1770258,3.0687182,4.2502565,5.5236926,4.919795,4.027077,3.3575387,3.131077,3.2820516,3.114667,2.8291285,2.5731285,2.4057438,2.3204105,2.1924105,2.1169233,2.0644104,1.9889232,1.8379488,1.4802053,1.3751796,1.3423591,1.2996924,1.270154,1.2012309,1.2800001,1.4572309,1.7460514,2.2186668,3.2229745,4.4307694,5.3202057,5.6320004,5.362872,6.2884107,8.349539,9.396514,8.438154,5.6352825,3.3247182,2.9472823,3.259077,3.5872824,3.8465643,3.9909747,3.882667,3.3509746,2.5206156,1.8248206,1.8412309,1.972513,1.9659488,1.8445129,1.9167181,1.7099489,1.657436,2.2186668,3.0194874,2.8389745,10.328616,9.281642,7.315693,5.9963083,5.7665644,5.9503593,5.474462,3.5610259,2.1956925,2.044718,2.4713848,3.3017437,4.397949,5.1364107,5.3792825,5.477744,5.3792825,5.110154,5.156103,5.4416413,5.293949,4.8082056,4.1714873,3.3903592,2.5337439,1.7394873,1.3718976,1.2635899,1.2340513,1.2274873,1.3128207,1.6311796,2.3138463,3.4297438,4.6080003,5.034667,3.9351797,2.930872,2.4155898,2.3466668,2.2121027,1.529436,1.2471796,1.2898463,1.404718,1.1585642,1.0732309,1.0633847,1.024,0.8598975,0.45620516,0.39712822,0.41682056,0.508718,0.6662565,0.88615394,1.079795,1.0010257,0.9156924,0.95835906,1.1290257,0.6892308,0.4135385,0.2986667,0.30194873,0.3511795,0.28882053,0.256,0.24943592,0.26584616,0.28882053,0.28882053,0.25271797,0.20348719,0.15425642,0.108307704,0.08205129,0.06564103,0.07876924,0.108307704,0.12143591,0.098461546,0.08205129,0.068923086,0.059076928,0.04594872,0.02297436,0.006564103,0.01969231,0.04266667,0.029538464,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.016410258,0.006564103,0.0,0.0032820515,0.016410258,0.016410258,0.016410258,0.009846155,0.0,0.0,0.013128206,0.02297436,0.049230773,0.098461546,0.18379489,0.34133336,0.4004103,0.49230772,0.7778462,1.4506668,0.9353847,0.571077,0.3314872,0.20676924,0.18379489,0.5481026,0.7515898,0.7581539,0.5874872,0.32164106,0.47917953,0.35446155,0.16410258,0.03938462,0.016410258,0.052512825,0.48246157,0.82379496,0.8598975,0.64000005,0.17723078,0.16082053,0.40697438,0.761436,1.1126155,1.332513,1.3423591,1.0371283,0.574359,0.36758977,0.48902568,0.45620516,0.4594872,0.52512825,0.48902568,0.32820517,0.1148718,0.06235898,0.14769232,0.12143591,0.21989745,0.574359,1.1355898,1.522872,1.024,0.6695385,0.6432821,0.56451285,0.53825647,1.1585642,0.93866676,0.35446155,0.0,0.059076928,0.28882053,0.43651286,0.49230772,0.41682056,0.34133336,0.5481026,0.8041026,1.0436924,1.2209232,1.2668719,1.083077,1.0469744,1.3226668,1.8051283,2.2613335,2.3335385,1.6738462,2.03159,3.2886157,5.2348723,7.5520005,4.2338467,2.6157951,1.9626669,1.6738462,1.2832822,2.733949,2.7766156,2.166154,1.4408206,0.9156924,0.7581539,0.5349744,0.3249231,0.21333335,0.27569234,0.5907693,0.94523084,1.2504616,1.3850257,1.1913847,0.446359,0.21333335,0.15753847,0.13128206,0.16738462,0.32820517,0.5677949,0.7384616,0.761436,0.64000005,0.60389745,1.2438976,2.0217438,2.484513,2.28759,1.6180514,0.98133343,1.0568206,1.9922053,3.4330258,5.4482055,8.487385,15.425642,22.098053,17.289848,13.124924,13.285745,15.573335,17.821539,17.8839,15.819489,13.033027,10.427077,8.667898,8.178872,8.789334,9.015796,8.057437,6.688821,7.2631803,5.5532312,3.7448208,2.793026,2.7208207,2.6256413,1.8806155,2.097231,2.986667,3.7021542,2.8225644,2.225231,1.7099489,1.5885129,2.1956925,3.9056413,3.9548721,3.006359,1.7165129,0.6859488,0.44307697,0.08861539,0.19364104,0.44307697,0.67282057,0.8533334,0.5973334,0.75487185,0.99774367,1.1158975,1.0075898,0.48246157,0.2855385,0.23302566,0.24287182,0.36758977,0.7089231,0.45620516,0.16082053,0.08205129,0.16738462,0.37415388,0.23630771,0.07548718,0.026256412,0.016410258,0.0032820515,0.0,0.049230773,0.13456412,0.18379489,0.23302566,0.3249231,0.6301539,1.0075898,1.0075898,0.9944616,1.2307693,1.1388719,0.69579494,0.4266667,0.256,0.13128206,0.06564103,0.06235898,0.12143591,0.108307704,0.06235898,0.01969231,0.0,0.0,0.0,0.036102567,0.12143591,0.18379489,0.06235898,0.02297436,0.016410258,0.02297436,0.026256412,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.02297436,0.026256412,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.02297436,0.04266667,0.07548718,0.13784617,0.25928208,0.318359,0.34133336,0.36102566,0.39712822,0.34789747,0.3446154,0.36430773,0.3708718,0.33476925,0.24943592,0.4135385,0.5152821,0.40369233,0.06235898,0.036102567,0.07548718,0.12471796,0.16082053,0.19692309,0.35774362,0.38728207,0.39384618,0.47917953,0.74830776,1.394872,1.2438976,0.90912825,0.67610264,0.51856416,0.446359,0.28225642,0.128,0.03938462,0.016410258,0.016410258,0.006564103,0.0,0.0,0.0,0.0,0.0,0.006564103,0.01969231,0.029538464,0.04266667,0.04594872,0.108307704,0.23958977,0.4135385,0.6301539,0.7975385,0.7187693,0.48902568,0.48902568,0.36758977,0.20676924,0.15097436,0.190359,0.15097436,0.128,0.11158975,0.13128206,0.15753847,0.12143591,0.072205134,0.052512825,0.03938462,0.026256412,0.016410258,0.0032820515,0.0,0.0,0.0032820515,0.016410258,0.052512825,0.052512825,0.03938462,0.032820515,0.04594872,0.059076928,0.08861539,0.13128206,0.19692309,0.32164106,1.3587693,2.231795,3.1573336,4.138667,4.9427695,3.5282054,3.4034874,3.5971284,3.5741541,3.2196925,3.1573336,2.8127182,2.7273848,3.05559,3.5544617,4.1058464,5.2381544,6.2720003,6.744616,6.439385,5.280821,4.8344617,5.395693,6.6100516,7.4765134,7.000616,5.2512827,3.7874875,3.56759,4.95918,6.2884107,5.7534366,5.32677,5.8781543,7.171283,7.9294367,7.7423596,7.8769236,8.346257,7.9195905,7.4797955,7.3419495,7.3682055,7.171283,6.1341543,5.2315903,4.893539,5.3694363,5.8880005,4.6539493,4.457026,4.71959,5.100308,5.8125134,7.643898,8.303591,7.7718983,6.5083084,5.687795,7.200821,8.057437,9.504821,11.500309,13.6697445,15.304206,14.792206,13.718975,12.616206,11.9171295,11.979488,12.42913,12.652308,12.504617,11.815386,10.374565,8.14277,6.951385,5.677949,3.7907696,1.3718976,0.6662565,0.31507695,0.27241027,0.46276927,0.79425645,0.9288206,0.8960001,0.702359,0.39056414,0.06235898,0.013128206,0.009846155,0.02297436,0.029538464,0.029538464,0.029538464,0.03938462,0.06564103,0.10502565,0.15097436,0.190359,0.21661541,0.24615386,0.3314872,0.56451285,0.9419488,1.2570257,1.3292309,1.1257436,0.74830776,0.5152821,0.5874872,1.0305642,2.0644104,4.027077,5.979898,7.0104623,6.629744,5.1265645,3.5413337,2.989949,2.917744,2.9407182,2.8947694,2.8225644,2.8947694,3.1343591,3.446154,3.761231,4.0434875,3.5052311,2.9046156,2.612513,3.3903592,6.3934364,5.1856413,3.4724104,2.1300514,1.7165129,2.4713848,3.0096412,3.1081028,2.937436,2.681436,2.546872,2.2547693,2.100513,2.1300514,2.3302567,2.6256413,2.428718,2.2416413,2.0709746,1.9232821,1.8018463,1.5819489,1.3686155,1.2307693,1.1848207,1.2209232,1.2209232,1.4408206,1.6672822,1.8412309,2.0611284,2.7437952,4.2436924,5.2676926,5.412103,5.142975,5.8256416,10.555078,12.320822,9.4457445,5.5991797,2.9768207,2.0086155,2.2153847,3.1376412,4.332308,5.2611284,5.356308,4.325744,2.6683078,1.6771283,1.4572309,1.6147693,1.8773335,2.0873847,2.1956925,2.1366155,2.156308,2.6289232,3.373949,3.692308,8.109949,7.702975,6.5870776,5.464616,4.955898,5.609026,6.3540516,6.055385,5.1298466,4.007385,3.1540515,3.8400004,4.598154,5.1659493,5.3431797,5.0018463,4.9132314,4.7458467,4.640821,4.667077,4.844308,4.8836927,4.4012313,3.7284105,3.1737437,3.0326157,3.058872,2.3860514,1.5983591,1.1290257,1.2635899,1.8543591,2.0053334,2.1202054,2.4057438,2.861949,3.4527183,3.5347695,3.242667,2.7142565,2.0906668,1.8084104,1.6278975,1.6508719,1.8084104,1.8674873,1.7920002,1.5786668,1.404718,1.3259488,1.2635899,1.2504616,0.86646163,0.5940513,0.60061544,0.761436,0.97805136,1.086359,1.1126155,1.0666667,0.94523084,0.69251287,0.5152821,0.42994875,0.4201026,0.44964105,0.446359,0.44964105,0.45620516,0.46276927,0.44964105,0.4004103,0.32820517,0.256,0.20020515,0.18051283,0.15425642,0.118153855,0.1148718,0.15425642,0.19692309,0.2100513,0.22646156,0.28882053,0.3314872,0.19364104,0.08861539,0.026256412,0.0032820515,0.009846155,0.01969231,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.01969231,0.052512825,0.032820515,0.009846155,0.0,0.006564103,0.026256412,0.016410258,0.016410258,0.013128206,0.009846155,0.0,0.0032820515,0.013128206,0.026256412,0.06235898,0.15753847,0.62030774,0.7384616,0.69907695,0.63343596,0.6301539,0.65641034,0.4594872,0.36102566,0.44964105,0.6104616,0.30194873,0.45292312,0.5513847,0.41682056,0.18707694,0.24615386,0.14769232,0.055794876,0.036102567,0.03938462,0.06564103,0.34133336,0.5415385,0.571077,0.5546667,0.5021539,0.4135385,0.43323082,0.5316923,0.5021539,0.4201026,0.58092314,0.6629744,0.5481026,0.32820517,0.22646156,0.33476925,0.41025645,0.35446155,0.21989745,0.118153855,0.10502565,0.101743594,0.118153855,0.21989745,0.46276927,0.7581539,0.84348726,0.6826667,0.48574364,0.43323082,0.48574364,0.4201026,0.47261542,1.3292309,1.024,0.37743592,0.009846155,0.15097436,0.65641034,0.57764107,0.42338464,0.33476925,0.40369233,0.65969235,0.8960001,1.086359,1.2242053,1.3128207,1.3653334,1.5622566,2.172718,3.18359,4.4996924,5.9602056,4.450462,3.7185643,3.4789746,3.314872,2.6453335,2.412308,2.809436,3.383795,3.764513,3.6857438,4.59159,5.4514875,5.4941545,4.391385,2.2449234,3.1015387,2.4451284,1.7690258,1.7952822,2.4713848,1.9298463,1.4769232,1.1815386,1.020718,0.88615394,0.764718,0.81394875,0.5284103,0.026256412,0.032820515,0.955077,1.3784616,1.5983591,1.6640002,1.3850257,0.7811283,1.2307693,1.6410258,1.5458462,1.1060513,0.5907693,0.37415388,0.7417436,1.7165129,3.0785644,4.821334,6.8463597,9.875693,12.822975,12.809847,12.980514,14.486976,15.530668,15.376411,14.342566,14.135796,14.867694,13.912617,11.1294365,8.874667,7.571693,6.7971287,6.5280004,6.2785645,5.113436,3.748103,2.733949,2.176,2.028308,2.0873847,1.9003079,1.8215386,1.8806155,1.9331284,1.6869745,1.5786668,1.2931283,0.8598975,0.6432821,1.3554872,1.1979488,0.8566154,0.5415385,0.32820517,0.16082053,0.18707694,0.30851284,0.4594872,0.5940513,0.65969235,0.55794877,0.7253334,0.9288206,1.0436924,1.0305642,0.63343596,0.47589746,0.43323082,0.4004103,0.318359,0.318359,0.27897438,0.26912823,0.3249231,0.44964105,1.1060513,0.9747693,0.6071795,0.3117949,0.16082053,0.04266667,0.0032820515,0.009846155,0.029538464,0.049230773,0.059076928,0.07876924,0.13784617,0.21333335,0.21333335,0.2100513,0.25928208,0.23630771,0.13784617,0.08533334,0.06235898,0.029538464,0.013128206,0.013128206,0.02297436,0.02297436,0.013128206,0.0032820515,0.0,0.0,0.0,0.006564103,0.02297436,0.036102567,0.013128206,0.0032820515,0.0032820515,0.0032820515,0.006564103,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.006564103,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.049230773,0.09189744,0.072205134,0.08205129,0.12471796,0.13784617,0.2297436,0.49230772,0.7187693,0.77456415,0.6170257,0.46933338,0.58092314,0.62030774,0.47261542,0.24943592,0.15425642,0.20348719,0.22646156,0.15753847,0.049230773,0.02297436,0.072205134,0.24287182,0.4594872,0.5152821,0.5874872,0.60389745,0.574359,0.56123084,0.6629744,0.9288206,1.0272821,1.0666667,1.0371283,0.8008206,0.67610264,0.49230772,0.23958977,0.006564103,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.009846155,0.01969231,0.026256412,0.02297436,0.006564103,0.009846155,0.02297436,0.055794876,0.101743594,0.15425642,0.2100513,0.28225642,0.30851284,0.29210258,0.28225642,0.24615386,0.190359,0.15097436,0.128,0.09189744,0.06564103,0.052512825,0.04594872,0.04594872,0.049230773,0.07876924,0.068923086,0.06235898,0.06564103,0.06564103,0.013128206,0.006564103,0.02297436,0.036102567,0.03938462,0.026256412,0.04594872,0.07548718,0.108307704,0.118153855,0.08205129,0.101743594,0.20348719,0.40697438,0.73517954,1.3817437,2.1431797,2.9144619,3.4822567,3.515077,2.8127182,2.7700515,3.4002054,4.3027697,4.673641,4.493129,3.8400004,3.4494362,3.498667,3.629949,4.33559,5.3694363,5.398975,4.5029745,4.1682053,4.073026,4.092718,3.7842054,3.436308,4.059898,4.2272825,4.161641,4.6802053,5.658257,6.0324106,6.2490263,6.2687182,6.5280004,7.020308,7.318975,7.4207187,7.3780518,7.509334,8.027898,9.068309,8.257642,7.4469748,6.9152827,6.6625648,6.426257,4.965744,3.826872,3.3411283,3.5380516,4.141949,4.562052,4.854154,5.21518,5.9536414,7.4732313,8.766359,8.592411,7.7456417,7.017026,7.200821,8.008205,9.452309,11.595488,14.296617,17.220924,17.558975,15.504412,13.712411,13.525334,14.992412,14.762668,13.971693,12.652308,10.8767185,8.753231,7.2205133,5.540103,3.7382567,1.9856411,0.60389745,0.3249231,0.19364104,0.19364104,0.29210258,0.4266667,0.318359,0.22646156,0.14769232,0.08205129,0.036102567,0.026256412,0.026256412,0.029538464,0.032820515,0.04266667,0.04266667,0.04594872,0.055794876,0.07548718,0.1148718,0.13456412,0.16410258,0.23302566,0.39384618,0.7220513,1.1027694,1.3128207,1.3587693,1.2406155,0.97805136,1.0010257,1.2832822,1.7526156,2.605949,4.2962055,5.586052,5.832206,5.0051284,3.5905645,2.5993848,2.3827693,2.487795,2.806154,3.1245131,3.1409233,2.9997952,2.92759,2.8914874,2.8258464,2.6289232,2.2580514,1.9528207,1.782154,1.9200002,2.6584618,5.717334,6.3376417,5.2512827,3.7776413,3.8498464,3.2656412,3.0227695,3.0227695,3.0949745,2.9997952,2.5107694,1.9790771,1.5819489,1.4276924,1.5261539,1.6935385,1.8510771,2.0086155,2.166154,2.3368206,2.4681027,2.0906668,1.5786668,1.1848207,1.024,1.2406155,1.6836925,2.0873847,2.409026,2.806154,4.082872,5.0510774,5.412103,5.182359,4.6769233,4.8049235,6.314667,6.6625648,5.280821,3.5741541,2.7667694,2.412308,2.4385643,2.7798977,3.3805132,4.017231,3.9778464,3.308308,2.353231,1.7624617,1.7296412,1.9396925,2.0906668,2.100513,2.1234872,1.9561027,1.6640002,1.8904617,2.5829747,3.0096412,7.141744,7.762052,7.9130263,7.6242056,7.0990777,6.741334,6.554257,6.3277955,5.868308,5.175795,4.4438977,4.562052,5.3431797,5.730462,5.4482055,4.97559,4.969026,4.9493337,5.0116925,5.1659493,5.333334,5.3234878,5.0576415,4.457026,3.69559,3.239385,3.1638978,2.7733335,2.1300514,1.4867693,1.2865642,1.6180514,1.8379488,2.162872,2.5107694,2.5206156,3.1245131,4.2469745,4.57518,3.9056413,3.1770258,2.6945643,2.2646155,1.9331284,1.7165129,1.6246156,1.6246156,1.6902566,1.9429746,2.3433847,2.681436,2.359795,1.7460514,1.339077,1.214359,1.024,0.9944616,1.0896411,1.204513,1.2274873,1.0469744,0.8992821,0.827077,0.7975385,0.7581539,0.6301539,0.56123084,0.508718,0.48246157,0.47261542,0.44307697,0.41682056,0.37415388,0.30851284,0.2297436,0.190359,0.21661541,0.21333335,0.20676924,0.21661541,0.25928208,0.256,0.24287182,0.256,0.25928208,0.14769232,0.07548718,0.032820515,0.01969231,0.01969231,0.02297436,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.032820515,0.02297436,0.013128206,0.009846155,0.009846155,0.013128206,0.02297436,0.02297436,0.01969231,0.013128206,0.0,0.0,0.0032820515,0.016410258,0.055794876,0.16082053,0.53825647,0.6859488,0.65641034,0.5218462,0.3708718,0.47261542,0.35446155,0.39056414,0.63343596,0.827077,0.50543594,0.4266667,0.40697438,0.3511795,0.26256412,0.26256412,0.2231795,0.15753847,0.0951795,0.06564103,0.06564103,0.18707694,0.28225642,0.30851284,0.3249231,0.3511795,0.3314872,0.36758977,0.41682056,0.29538465,0.18051283,0.26584616,0.38728207,0.45292312,0.42994875,0.30194873,0.24943592,0.20676924,0.18051283,0.22646156,0.17723078,0.108307704,0.08533334,0.11158975,0.14441027,0.24943592,0.35774362,0.34133336,0.21989745,0.17723078,0.17066668,0.19692309,0.18379489,0.27897438,0.85005134,0.6695385,0.3052308,0.09189744,0.20348719,0.636718,0.4955898,0.33476925,0.29538465,0.44307697,0.7778462,1.3620514,1.6114873,1.595077,1.6443079,2.3401027,2.5961027,3.242667,4.2502565,5.481026,6.701949,5.989744,5.2315903,4.397949,3.4034874,2.1070771,3.170462,4.535795,5.681231,6.186667,5.733744,6.1374364,6.377026,5.973334,4.7458467,2.8258464,3.3444104,2.7044106,2.172718,2.3729234,3.2787695,3.0490258,2.7175386,2.5107694,2.5304618,2.7306669,2.349949,2.4484105,2.6026669,2.7667694,3.249231,4.1485133,4.5095387,4.562052,4.532513,4.647385,5.293949,4.092718,2.806154,2.1825643,1.9528207,1.8215386,1.6869745,1.8970258,2.5665643,3.5872824,4.965744,6.186667,7.785026,9.941334,12.49477,14.923489,15.520822,15.113848,14.168616,12.780309,12.2617445,12.832822,11.762873,8.950154,6.925129,6.0947695,6.0192823,5.940513,5.3103595,3.8006158,2.809436,2.4713848,2.169436,1.8116925,1.8051283,1.8838975,1.8576412,1.4966155,0.98133343,0.90912825,0.9517949,0.83035904,0.52512825,0.23302566,0.39712822,0.32164106,0.21989745,0.190359,0.24287182,0.29210258,0.42338464,0.508718,0.5415385,0.51856416,0.43651286,0.49230772,0.73517954,1.024,1.1946667,1.0469744,0.7253334,0.57764107,0.5218462,0.4955898,0.46933338,0.34789747,0.38728207,0.45292312,0.47261542,0.446359,0.7089231,0.7187693,0.7089231,0.81066674,1.0666667,0.79097444,0.6892308,0.7318975,0.8369231,0.892718,0.84348726,1.0108719,1.1093334,0.8763078,0.068923086,0.73517954,0.69907695,0.37415388,0.101743594,0.13784617,0.068923086,0.01969231,0.0,0.0032820515,0.01969231,0.16410258,0.13128206,0.049230773,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.009846155,0.01969231,0.029538464,0.036102567,0.036102567,0.013128206,0.013128206,0.013128206,0.016410258,0.04266667,0.068923086,0.06235898,0.07876924,0.13784617,0.21989745,0.23302566,0.42338464,0.62030774,0.69251287,0.54482055,0.50543594,0.5907693,0.58420515,0.43651286,0.24615386,0.26584616,0.29538465,0.28225642,0.21333335,0.128,0.10502565,0.1148718,0.18707694,0.29538465,0.35774362,0.44307697,0.5284103,0.6071795,0.6498462,0.6301539,0.5907693,0.67610264,0.7975385,0.84348726,0.69579494,0.5021539,0.30851284,0.13128206,0.006564103,0.0,0.0,0.006564103,0.009846155,0.009846155,0.01969231,0.029538464,0.052512825,0.06564103,0.06235898,0.04594872,0.059076928,0.07548718,0.098461546,0.11158975,0.101743594,0.10502565,0.13128206,0.16738462,0.19692309,0.19364104,0.17394873,0.15097436,0.128,0.108307704,0.08533334,0.052512825,0.029538464,0.016410258,0.009846155,0.02297436,0.07876924,0.101743594,0.11158975,0.118153855,0.10502565,0.06564103,0.068923086,0.068923086,0.049230773,0.026256412,0.016410258,0.026256412,0.04594872,0.108307704,0.26584616,0.25928208,0.29210258,0.42994875,0.69579494,1.0666667,1.8215386,2.6617439,3.4297438,3.826872,3.3969233,2.9965131,2.9735386,3.3444104,3.9909747,4.650667,4.926359,4.4996924,3.889231,3.4494362,3.3641028,3.8596926,4.4701543,4.516103,3.9745643,3.501949,3.3345644,3.2853336,3.1113849,3.0030773,3.570872,4.2436924,4.588308,5.1856413,5.8945646,5.861744,5.536821,5.586052,5.7534366,5.930667,6.1472826,6.6133337,6.567385,6.75118,7.433847,8.4283085,7.512616,6.810257,6.416411,6.36718,6.6461544,5.4941545,4.637539,4.0402055,3.8990772,4.6539493,6.442667,7.069539,7.128616,7.1089234,7.384616,9.035488,9.7903595,9.29477,8.086975,7.604513,8.612103,9.810052,12.278154,16.098463,20.36513,20.716309,19.236105,17.72636,16.928822,16.544823,15.37313,13.6237955,11.457642,9.045334,6.5903597,5.0576415,3.6726158,2.3368206,1.1716924,0.5021539,0.25928208,0.11158975,0.0951795,0.16082053,0.190359,0.07548718,0.02297436,0.0032820515,0.0032820515,0.02297436,0.036102567,0.055794876,0.07876924,0.0951795,0.09189744,0.068923086,0.049230773,0.036102567,0.04266667,0.07876924,0.1148718,0.16738462,0.21333335,0.28225642,0.4594872,0.7581539,1.0502565,1.3062565,1.4342566,1.276718,1.2800001,1.6705642,2.284308,3.045744,3.95159,4.4438977,4.312616,3.6857438,2.9243078,2.6026669,2.5140514,2.5796926,2.806154,3.131077,3.4297438,3.170462,2.8882053,2.740513,2.6912823,2.5206156,2.1169233,1.7887181,1.5425643,1.4703591,1.7526156,4.194462,6.235898,6.8233852,6.0652313,5.221744,4.0992823,3.2229745,2.8488207,2.8882053,2.9210258,2.6486156,2.1431797,1.6705642,1.394872,1.4145643,1.591795,1.719795,1.8116925,1.9035898,2.0611284,2.294154,2.097231,1.6836925,1.270154,1.0765129,1.3751796,1.9364104,2.553436,3.2032824,4.017231,5.07077,5.5236926,5.4580517,5.0838976,4.7622566,4.8607183,5.2447186,5.1922054,4.46359,3.314872,3.9548721,3.6004105,2.937436,2.5238976,2.7766156,3.2361028,3.1409233,2.6289232,1.9528207,1.463795,1.3522053,1.4178462,1.4736412,1.5163078,1.719795,1.5392822,1.3161026,1.3850257,1.7755898,2.2350771,6.0356927,7.1548724,8.247795,8.953437,9.248821,9.45559,9.025641,7.824411,6.8463597,6.262154,5.425231,4.8607183,5.4153852,6.1046157,6.2818465,5.6320004,5.3858466,5.2414365,5.287385,5.4482055,5.474462,5.4153852,5.4941545,5.2611284,4.630975,3.8859491,3.5840003,3.387077,2.9505644,2.294154,1.8116925,2.0151796,2.3433847,2.6157951,2.7208207,2.612513,2.7798977,3.7710772,4.3290257,4.2174363,4.2141542,3.7448208,3.1803079,2.5764105,2.048,1.7887181,1.6968206,1.7493335,1.972513,2.3958976,3.0687182,3.0391798,2.7864618,2.5993848,2.484513,2.172718,1.4998976,1.2077949,1.1716924,1.2209232,1.1552821,1.0305642,1.014154,1.0305642,0.98461545,0.7581539,0.5513847,0.4266667,0.3708718,0.35446155,0.3314872,0.32820517,0.31507695,0.27897438,0.2297436,0.21333335,0.26912823,0.28882053,0.2855385,0.28225642,0.31507695,0.2986667,0.24287182,0.18051283,0.12471796,0.06564103,0.036102567,0.032820515,0.036102567,0.036102567,0.036102567,0.032820515,0.01969231,0.009846155,0.0032820515,0.0,0.0,0.0,0.0032820515,0.006564103,0.006564103,0.0,0.0,0.0,0.0032820515,0.016410258,0.016410258,0.02297436,0.026256412,0.01969231,0.013128206,0.026256412,0.032820515,0.029538464,0.013128206,0.006564103,0.0,0.0,0.016410258,0.07548718,0.2100513,0.4660513,0.6235898,0.61374366,0.4660513,0.3117949,0.318359,0.29210258,0.36430773,0.54482055,0.7187693,0.6826667,0.6301539,0.51856416,0.38400003,0.33476925,0.31507695,0.29538465,0.26584616,0.21333335,0.13784617,0.13128206,0.18051283,0.21333335,0.21333335,0.24287182,0.27569234,0.29538465,0.3052308,0.3117949,0.3314872,0.40369233,0.508718,0.46933338,0.3314872,0.3708718,0.27897438,0.14112821,0.049230773,0.055794876,0.17723078,0.15753847,0.072205134,0.03938462,0.068923086,0.059076928,0.055794876,0.055794876,0.04266667,0.029538464,0.04266667,0.029538464,0.032820515,0.059076928,0.14112821,0.3314872,0.28225642,0.190359,0.15097436,0.2231795,0.43651286,0.3446154,0.29538465,0.3511795,0.54482055,0.88943595,1.4900514,1.7591796,1.8215386,2.1267693,3.4264617,3.6332312,4.204308,5.0871797,6.124308,7.0367184,6.36718,5.4613338,4.4438977,3.4231799,2.484513,3.8662567,5.280821,6.2687182,6.4590774,5.5696416,5.943795,5.7501545,5.152821,4.3684106,3.6693337,4.1747694,3.9154875,3.5347695,3.4133337,3.6693337,3.4330258,3.249231,3.2984617,3.692308,4.4832826,5.277539,5.4383593,5.280821,5.093744,5.142975,6.5772314,6.3376417,5.7435904,5.5532312,5.9667697,6.685539,5.175795,3.7087183,3.1934361,3.1671798,3.18359,2.9965131,3.1376412,3.761231,4.6605134,5.5696416,6.6822567,8.050873,9.846154,12.373334,14.851283,14.611693,13.436719,12.176412,10.729027,9.757539,9.432616,8.254359,6.298257,5.2512827,5.398975,5.858462,5.5597954,4.3552823,3.0227695,2.3335385,2.353231,2.2711797,1.9068719,1.7263591,1.7296412,1.7296412,1.3161026,0.6662565,0.5316923,0.50543594,0.39712822,0.2855385,0.20676924,0.17066668,0.17394873,0.16738462,0.18051283,0.23630771,0.36102566,0.50543594,0.65312827,0.75487185,0.75487185,0.58420515,0.65969235,0.94523084,1.3193847,1.5097437,1.0962052,0.7844103,0.6859488,0.75487185,0.8467693,0.7253334,0.574359,0.62030774,0.6662565,0.62030774,0.4955898,0.36758977,0.34789747,0.4594872,0.69251287,1.0075898,0.7811283,0.7089231,0.7778462,0.9189744,0.99774367,0.9747693,1.1716924,1.273436,1.024,0.19692309,0.86974365,0.8369231,0.56123084,0.47589746,0.9911796,0.702359,0.47917953,0.318359,0.20020515,0.072205134,0.24943592,0.20348719,0.08533334,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.009846155,0.01969231,0.04266667,0.068923086,0.07876924,0.06235898,0.055794876,0.052512825,0.055794876,0.06564103,0.07548718,0.07876924,0.098461546,0.13456412,0.190359,0.16082053,0.23958977,0.35774362,0.46276927,0.4955898,0.55794877,0.55794877,0.508718,0.4201026,0.31507695,0.37415388,0.42338464,0.36758977,0.23302566,0.14769232,0.13784617,0.14112821,0.16082053,0.20020515,0.27241027,0.39712822,0.5415385,0.7122052,0.8369231,0.74830776,0.6170257,0.6071795,0.60389745,0.54482055,0.39712822,0.24287182,0.1148718,0.036102567,0.006564103,0.0,0.0,0.006564103,0.013128206,0.01969231,0.029538464,0.04266667,0.068923086,0.08861539,0.08861539,0.068923086,0.12471796,0.16082053,0.190359,0.20348719,0.15425642,0.15097436,0.15425642,0.15753847,0.15097436,0.13128206,0.118153855,0.10502565,0.0951795,0.09189744,0.07876924,0.06235898,0.04266667,0.02297436,0.006564103,0.016410258,0.04594872,0.07876924,0.108307704,0.13128206,0.14769232,0.108307704,0.128,0.13128206,0.098461546,0.052512825,0.04266667,0.036102567,0.059076928,0.15425642,0.37415388,0.37415388,0.38400003,0.5218462,0.83035904,1.2438976,2.0841026,2.9669745,3.629949,3.8104618,3.2689233,2.930872,3.0523078,3.2656412,3.5282054,4.1189747,4.97559,5.4843082,5.110154,4.0992823,3.4855387,3.6332312,3.7349746,3.8662567,3.9253337,3.623385,3.2032824,2.9440002,3.0030773,3.5249233,4.644103,6.091488,6.6560006,6.6395903,6.232616,5.533539,4.896821,5.408821,5.76,5.5663595,5.3825645,6.124308,6.163693,6.2687182,6.7774363,7.634052,7.269744,6.626462,6.232616,6.4000006,7.2270775,6.665847,5.684513,4.818052,4.46359,4.886975,7.2237954,8.530052,8.832001,8.562873,8.582564,10.624001,11.680821,11.480617,10.499283,9.961026,10.059488,10.712616,13.157744,17.404718,22.226053,23.138464,22.505028,21.169233,19.475695,17.293129,15.130258,12.547283,9.819899,7.181129,4.8082056,3.3476925,2.3401027,1.5031796,0.8205129,0.5218462,0.2986667,0.128,0.059076928,0.06235898,0.055794876,0.009846155,0.0,0.0032820515,0.009846155,0.026256412,0.052512825,0.08861539,0.128,0.15425642,0.14769232,0.128,0.08205129,0.04266667,0.032820515,0.055794876,0.0951795,0.14769232,0.17066668,0.18051283,0.23958977,0.4135385,0.7089231,1.1027694,1.4539489,1.5261539,1.4473847,1.6246156,2.103795,2.7437952,3.2262566,3.495385,3.4527183,3.4166157,3.6791797,4.4898467,5.139693,4.4898467,3.5347695,3.0194874,3.442872,3.5413337,3.4100516,3.2525132,3.1113849,2.868513,2.9702566,2.5993848,2.0676925,1.6278975,1.4900514,2.484513,4.5423594,5.8223596,5.609026,4.332308,3.3542566,2.612513,2.3204105,2.4484105,2.7142565,2.7437952,2.4943593,2.162872,1.9200002,1.9167181,2.0906668,2.1202054,2.0118976,1.8609232,1.8773335,1.9954873,1.8806155,1.6311796,1.4112822,1.4441026,1.7624617,2.300718,3.0129232,3.895795,4.9920006,5.579488,5.586052,5.2676926,4.84759,4.532513,4.394667,4.322462,4.06318,3.6004105,3.1507695,4.2272825,3.8498464,2.9965131,2.3827693,2.484513,2.6880002,2.5107694,2.0742567,1.5392822,1.1060513,1.0305642,1.014154,0.99774367,1.014154,1.1979488,1.0404103,1.0404103,1.214359,1.5524104,2.0086155,4.7589746,5.5236926,6.741334,8.057437,9.462154,11.300103,11.657847,9.885539,8.362667,7.6603084,6.564103,5.333334,5.211898,6.193231,7.3649235,6.9087186,6.2588725,5.7829747,5.540103,5.431795,5.2053337,5.080616,5.353026,5.5762057,5.4580517,4.8804107,4.4898467,4.1025643,3.636513,3.1573336,2.9013336,3.7776413,3.895795,3.3476925,2.665026,2.8488207,2.6551797,2.6880002,2.9965131,3.5741541,4.348718,4.2994876,3.9384618,3.4330258,2.9505644,2.681436,2.3827693,2.0118976,1.6278975,1.5031796,2.1234872,2.7733335,3.2164104,3.4133337,3.3641028,3.1343591,2.0250258,1.4145643,1.2077949,1.2570257,1.3653334,1.1979488,1.1651284,1.148718,1.0535386,0.7844103,0.44307697,0.27241027,0.21333335,0.20676924,0.2100513,0.19692309,0.19364104,0.19692309,0.21333335,0.256,0.28882053,0.29210258,0.28882053,0.29538465,0.32164106,0.32164106,0.23630771,0.13456412,0.06235898,0.026256412,0.006564103,0.02297436,0.03938462,0.04266667,0.04594872,0.068923086,0.049230773,0.032820515,0.029538464,0.016410258,0.006564103,0.006564103,0.009846155,0.013128206,0.013128206,0.0032820515,0.0,0.0,0.0032820515,0.016410258,0.01969231,0.029538464,0.04266667,0.049230773,0.04266667,0.029538464,0.032820515,0.026256412,0.013128206,0.013128206,0.0032820515,0.0,0.02297436,0.09189744,0.2297436,0.43651286,0.60389745,0.5973334,0.43323082,0.27897438,0.20676924,0.25271797,0.27897438,0.2855385,0.4135385,0.63343596,0.82379496,0.72861546,0.4266667,0.3249231,0.30851284,0.27569234,0.33805132,0.4266667,0.28225642,0.23302566,0.26584616,0.26256412,0.2297436,0.28882053,0.36430773,0.38728207,0.3249231,0.3314872,0.7450257,0.8992821,0.92225647,0.6301539,0.19364104,0.13456412,0.08533334,0.029538464,0.0032820515,0.009846155,0.026256412,0.016410258,0.006564103,0.0032820515,0.006564103,0.02297436,0.032820515,0.036102567,0.02297436,0.0032820515,0.013128206,0.013128206,0.029538464,0.068923086,0.108307704,0.08861539,0.07548718,0.09189744,0.14112821,0.20348719,0.2297436,0.24287182,0.32820517,0.47261542,0.67282057,0.90912825,1.1520001,1.4473847,1.8904617,2.7011285,4.204308,4.4045134,5.0084105,5.917539,6.944821,7.788308,5.933949,4.4045134,3.2689233,2.546872,2.2153847,3.3641028,4.4242053,5.024821,4.8640003,3.7185643,4.2174363,4.2535386,4.1189747,4.1091285,4.5062566,5.464616,5.474462,4.9427695,4.2207184,3.5872824,2.9472823,2.8947694,3.2787695,4.0533338,5.280821,8.024616,8.484103,7.6931286,6.4754877,5.4416413,6.9809237,5.8256416,4.667077,4.6834874,5.540103,5.3005133,4.601436,4.017231,3.7874875,3.7907696,3.7382567,3.4658465,3.7185643,4.637539,5.7632823,6.196513,7.4765134,8.776206,9.80677,10.817642,11.959796,11.943385,11.001437,9.524513,8.0377445,7.138462,6.426257,5.6352825,4.900103,4.7327185,5.3169236,5.4416413,4.772103,3.515077,2.4418464,1.9331284,2.041436,2.1366155,1.9626669,1.6640002,1.4605129,1.2931283,1.0010257,0.6268718,0.41682056,0.24943592,0.08205129,0.072205134,0.17723078,0.15753847,0.14769232,0.16738462,0.17723078,0.17723078,0.20676924,0.36758977,0.63343596,0.9353847,1.1323078,1.0043077,1.0075898,1.2570257,1.5786668,1.6705642,1.1060513,0.8008206,0.7811283,1.0404103,1.2964103,0.99774367,0.88943595,0.9878975,0.9944616,0.8533334,0.7089231,0.49230772,0.27569234,0.13456412,0.07548718,0.07876924,0.07548718,0.098461546,0.13456412,0.17723078,0.22646156,0.2855385,0.3446154,0.37415388,0.36102566,0.3249231,0.34133336,0.36758977,0.4660513,0.83035904,1.7887181,1.3423591,0.9616411,0.67938465,0.44964105,0.14112821,0.18379489,0.15097436,0.07548718,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.032820515,0.07548718,0.10502565,0.118153855,0.11158975,0.108307704,0.118153855,0.13128206,0.15425642,0.15753847,0.14441027,0.118153855,0.059076928,0.049230773,0.068923086,0.14441027,0.2986667,0.5513847,0.7122052,0.6662565,0.5973334,0.56123084,0.49230772,0.42338464,0.44964105,0.39384618,0.26584616,0.27897438,0.22646156,0.23302566,0.28225642,0.35446155,0.4201026,0.5349744,0.7581539,1.0699488,1.339077,1.3062565,1.1158975,0.84348726,0.5677949,0.32164106,0.101743594,0.072205134,0.049230773,0.02297436,0.0,0.0,0.0,0.0,0.006564103,0.01969231,0.029538464,0.03938462,0.059076928,0.07548718,0.08205129,0.068923086,0.15097436,0.2100513,0.24943592,0.26256412,0.21989745,0.2100513,0.20020515,0.17066668,0.118153855,0.072205134,0.072205134,0.06564103,0.068923086,0.07548718,0.068923086,0.08205129,0.07876924,0.052512825,0.016410258,0.013128206,0.0032820515,0.013128206,0.04594872,0.0951795,0.16738462,0.12471796,0.14441027,0.16082053,0.14112821,0.08861539,0.07876924,0.07876924,0.13128206,0.23302566,0.35446155,0.32164106,0.30851284,0.45292312,0.8205129,1.3850257,2.041436,2.681436,3.0326157,3.0030773,2.6880002,2.4385643,2.7667694,3.1442053,3.370667,3.5807183,4.8771286,6.626462,7.0826674,5.973334,4.4996924,4.197744,3.8137438,3.6562054,3.8006158,4.07959,3.639795,3.318154,3.5905645,4.5817437,6.0685134,7.9294367,8.713847,8.372514,7.3025646,6.3310776,5.5729237,6.7577443,7.712821,7.387898,5.8420515,6.170257,6.409847,6.4623594,6.4656415,6.770872,7.4141545,6.8955903,6.409847,6.695385,8.034462,8.057437,6.547693,5.169231,4.7228723,5.152821,6.889026,8.795898,9.869129,10.174359,10.817642,12.983796,14.148924,14.857847,15.126975,14.421334,12.304411,12.09436,14.198155,18.25477,23.168001,24.825438,24.231386,22.33436,19.830154,17.165129,14.464001,11.378873,8.375795,5.7731285,3.7415388,2.612513,1.7690258,1.0994873,0.60389745,0.4004103,0.3052308,0.19364104,0.08533334,0.013128206,0.0032820515,0.0,0.0,0.006564103,0.01969231,0.04266667,0.068923086,0.12143591,0.16410258,0.18379489,0.18707694,0.22646156,0.16082053,0.08861539,0.052512825,0.04594872,0.059076928,0.08861539,0.1148718,0.14112821,0.20348719,0.27569234,0.44307697,0.78769237,1.2504616,1.6475899,1.595077,1.4112822,1.4998976,1.9364104,2.4582565,2.9833848,3.2000003,3.8367183,5.2381544,7.3714876,8.973129,7.6242056,5.211898,3.3509746,3.3969233,4.141949,4.640821,4.7261543,4.352,3.6069746,4.4012313,4.906667,4.3716927,2.9210258,1.5524104,1.6640002,2.5895386,3.1540515,2.8750772,1.9561027,1.5622566,1.5983591,1.8576412,2.228513,2.6912823,2.868513,2.8160002,2.6322052,2.4418464,2.422154,2.6551797,2.681436,2.4582565,2.1267693,2.0118976,1.9922053,1.847795,1.7132308,1.7493335,2.15959,2.556718,3.0162053,3.6627696,4.5489235,5.6385646,5.792821,5.356308,4.775385,4.2601027,3.7710772,3.1540515,2.6223593,2.0939488,1.8215386,2.3893335,3.121231,3.0293336,2.6256413,2.300718,2.3368206,2.2416413,1.9495386,1.5360001,1.1093334,0.827077,0.9321026,0.95835906,0.9124103,0.83035904,0.76800007,0.6465641,0.81394875,1.2176411,1.7099489,2.0545642,4.6244106,4.453744,4.7392826,5.648411,6.7971287,7.24677,7.273026,7.755488,8.602257,9.458873,9.688616,7.785026,6.741334,6.5411286,7.128616,8.421744,7.958975,7.3747697,6.889026,6.439385,5.7074876,4.8771286,4.588308,4.57518,4.6112823,4.5029745,4.3060517,3.698872,3.2098465,3.2820516,4.2568207,7.259898,6.7117953,5.0149746,3.82359,4.0434875,3.370667,3.4592824,3.6430771,3.5544617,3.1277952,3.4691284,3.6463592,3.767795,3.8038976,3.5872824,3.3050258,2.6322052,1.8609232,1.2340513,0.9156924,1.2340513,1.7690258,2.0086155,1.7788719,1.2668719,1.2898463,1.4605129,1.7165129,1.975795,2.1202054,1.8773335,1.7788719,1.585231,1.211077,0.74830776,0.35774362,0.20348719,0.17394873,0.18707694,0.19692309,0.18707694,0.17394873,0.18707694,0.21989745,0.24287182,0.20676924,0.17066668,0.15753847,0.17394873,0.19692309,0.19692309,0.14441027,0.08205129,0.03938462,0.016410258,0.0032820515,0.0,0.013128206,0.032820515,0.04594872,0.059076928,0.052512825,0.068923086,0.101743594,0.07548718,0.03938462,0.029538464,0.01969231,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.03938462,0.01969231,0.055794876,0.128,0.09189744,0.01969231,0.0,0.0,0.0,0.0,0.0,0.0,0.01969231,0.04594872,0.04594872,0.15425642,0.35774362,0.42338464,0.33805132,0.28882053,0.2297436,0.16738462,0.19692309,0.29210258,0.3052308,0.4135385,0.58092314,0.52512825,0.30194873,0.28882053,0.25271797,0.24287182,0.512,0.83035904,0.48902568,0.256,0.16082053,0.118153855,0.0951795,0.108307704,0.23958977,0.39384618,0.49887183,0.8172308,1.9528207,1.4998976,0.62030774,0.06564103,0.0,0.0,0.0,0.0,0.013128206,0.026256412,0.016410258,0.0032820515,0.009846155,0.016410258,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.03938462,0.08861539,0.13784617,0.06564103,0.04594872,0.07548718,0.13128206,0.16738462,0.28882053,0.42994875,0.57764107,0.6892308,0.702359,0.8008206,1.3653334,2.2908719,3.4002054,4.4242053,4.890257,5.901129,7.1089234,8.044309,8.116513,5.333334,3.1638978,1.7558975,1.214359,1.6180514,2.044718,3.2229745,4.2896414,4.4734364,3.0818465,2.802872,3.0523078,3.4855387,3.8104618,3.8006158,4.240411,3.5610259,2.5961027,1.9364104,1.9364104,1.8281027,2.6978464,3.882667,4.9362054,5.6451287,7.463385,8.651488,9.212719,9.114257,8.283898,6.160411,4.532513,4.2830772,5.648411,8.224821,9.284924,7.253334,4.8804107,3.6069746,3.570872,3.754667,3.3411283,3.5249233,4.6276927,6.1046157,6.2752824,6.6822567,7.276308,7.9491286,8.55959,8.756514,9.665642,9.701744,8.490667,6.8660517,5.8912826,4.8114877,4.135385,4.0008206,4.197744,4.4767184,3.82359,3.05559,2.428718,1.6475899,1.2570257,1.4605129,1.585231,1.4309745,1.2964103,1.211077,0.71548724,0.37743592,0.3314872,0.25928208,0.052512825,0.0,0.04266667,0.12143591,0.18379489,0.18379489,0.072205134,0.0,0.0,0.0,0.17066668,0.38728207,0.67610264,0.9682052,1.1126155,1.1749744,1.2996924,1.2996924,1.1290257,0.88615394,0.7253334,0.7220513,0.9189744,1.1815386,1.204513,1.3029745,1.6475899,1.6475899,1.2570257,0.97805136,0.7187693,0.446359,0.190359,0.055794876,0.21333335,0.24943592,0.25928208,0.19364104,0.07876924,0.029538464,0.029538464,0.07548718,0.16738462,0.26256412,0.27569234,0.3117949,0.39384618,0.42338464,0.39712822,0.39712822,0.3117949,0.19692309,0.20348719,0.27569234,0.15097436,0.07876924,0.02297436,0.006564103,0.016410258,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01969231,0.036102567,0.055794876,0.09189744,0.1148718,0.14112821,0.14769232,0.14441027,0.16738462,0.28882053,0.26584616,0.18051283,0.0951795,0.04594872,0.04594872,0.04594872,0.108307704,0.27241027,0.56451285,1.017436,1.0666667,1.017436,0.97805136,0.86974365,0.5284103,0.3708718,0.47261542,0.764718,1.020718,0.71548724,0.6301539,0.61374366,0.5907693,0.58092314,0.5677949,1.0502565,1.8116925,2.540308,2.806154,2.0512822,1.0371283,0.34133336,0.101743594,0.016410258,0.016410258,0.006564103,0.0,0.0,0.0,0.0,0.0,0.006564103,0.01969231,0.029538464,0.029538464,0.03938462,0.052512825,0.068923086,0.108307704,0.118153855,0.13128206,0.13784617,0.14769232,0.18379489,0.18379489,0.14769232,0.1148718,0.098461546,0.06235898,0.049230773,0.06564103,0.07548718,0.08205129,0.108307704,0.118153855,0.12143591,0.08533334,0.02297436,0.0,0.0,0.0,0.006564103,0.032820515,0.108307704,0.14441027,0.1148718,0.06564103,0.026256412,0.016410258,0.06564103,0.13128206,0.19364104,0.20676924,0.12143591,0.108307704,0.21661541,0.45620516,0.92225647,1.8018463,2.0578463,1.8642052,1.7624617,1.9068719,2.0906668,2.297436,2.5862565,3.1081028,3.5314875,3.0654361,4.5817437,6.882462,8.694155,8.933744,6.698667,5.674667,4.821334,4.0336413,3.7152824,4.775385,4.4340515,4.384821,5.5204105,7.1089234,6.7905645,7.059693,7.318975,7.6898465,8.395488,9.750975,9.324308,9.96759,11.211488,11.346052,7.4141545,6.5739493,6.921847,7.4830775,7.0892315,4.378257,5.684513,6.432821,6.688821,6.997334,8.375795,8.976411,8.024616,6.7249236,6.1768208,7.384616,8.3134365,9.816616,11.336206,12.356924,12.406155,13.515489,16.649847,20.233849,22.150566,19.744822,15.058052,13.702565,15.711181,20.41108,26.427078,26.89313,24.644924,21.290668,17.959387,15.333745,13.344822,10.466462,7.4896417,4.9493337,3.1442053,2.1792822,1.4080001,0.81394875,0.4004103,0.16738462,0.18051283,0.14769232,0.10502565,0.06564103,0.016410258,0.0032820515,0.0,0.006564103,0.01969231,0.029538464,0.06564103,0.15097436,0.19364104,0.18707694,0.19692309,0.3446154,0.27241027,0.15425642,0.08205129,0.04594872,0.02297436,0.032820515,0.059076928,0.0951795,0.16738462,0.27897438,0.3249231,0.52512825,0.96492314,1.5885129,1.8182565,1.6738462,1.5786668,1.7263591,2.1070771,2.4713848,2.4549747,3.4855387,5.8223596,8.546462,9.655796,9.511385,7.706257,5.1298466,3.9811285,4.8738465,6.488616,7.496206,7.1844106,5.4613338,5.717334,9.554052,10.299078,6.813539,3.495385,1.9922053,1.6344616,1.6836925,1.7723079,1.9068719,1.9331284,2.1103592,2.412308,2.7634873,3.0818465,3.0818465,2.789744,2.422154,2.1530259,2.1070771,2.2416413,2.3663592,2.3269746,2.1464617,1.9987694,2.1956925,2.3171284,2.3958976,2.5993848,3.2361028,3.9417439,4.457026,4.965744,5.602462,6.4689236,6.2129235,5.159385,3.9942567,3.1737437,2.930872,2.2350771,1.3456411,0.7844103,0.79097444,1.3292309,2.048,2.5862565,2.5665643,2.1530259,2.044718,1.847795,1.4998976,1.0108719,0.58420515,0.5940513,0.67938465,0.7384616,0.7581539,0.7318975,0.67282057,0.5973334,0.6892308,0.94523084,1.211077,1.1749744,9.494975,9.645949,10.003693,9.577026,8.267488,6.882462,6.2818465,6.7544622,8.372514,10.14154,9.980719,7.0826674,6.925129,7.056411,6.764308,7.0925136,7.702975,7.2992826,6.4065647,5.4153852,4.585026,4.2141542,4.46359,4.788513,4.919795,4.8804107,4.5489235,3.817026,3.2820516,3.4166157,4.598154,6.2752824,5.5762057,4.8738465,4.9460516,4.972308,4.378257,3.8400004,3.4100516,2.9833848,2.3236926,2.028308,2.356513,3.0523078,3.9187696,4.781949,4.7360005,3.1442053,2.0118976,1.7788719,1.3554872,1.0371283,0.97805136,1.0010257,0.9747693,0.8041026,0.7384616,0.75487185,0.90912825,1.1651284,1.3883078,1.4867693,1.5688206,1.339077,0.892718,0.7220513,0.6826667,0.6629744,0.56123084,0.39712822,0.32164106,0.25928208,0.22646156,0.21661541,0.2231795,0.256,0.27897438,0.26256412,0.2231795,0.16738462,0.11158975,0.07548718,0.04594872,0.029538464,0.01969231,0.016410258,0.013128206,0.013128206,0.02297436,0.049230773,0.068923086,0.072205134,0.049230773,0.06235898,0.101743594,0.07548718,0.049230773,0.04266667,0.03938462,0.032820515,0.02297436,0.16082053,0.2986667,0.23302566,0.029538464,0.0032820515,0.08533334,0.16082053,0.18707694,0.15097436,0.06564103,0.032820515,0.03938462,0.029538464,0.0,0.0,0.049230773,0.13456412,0.23630771,0.3052308,0.26584616,0.28882053,0.32820517,0.3249231,0.28225642,0.25271797,0.28882053,0.28882053,0.19692309,0.101743594,0.21989745,0.24287182,0.23958977,0.18707694,0.12143591,0.118153855,0.13128206,0.17066668,0.29210258,0.39712822,0.23302566,0.46933338,0.67282057,0.6892308,0.5021539,0.23958977,0.14112821,0.101743594,0.098461546,0.16410258,0.39056414,0.30851284,0.13456412,0.01969231,0.0032820515,0.013128206,0.0032820515,0.006564103,0.01969231,0.026256412,0.0032820515,0.0,0.0032820515,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.016410258,0.026256412,0.02297436,0.029538464,0.04594872,0.07548718,0.13128206,0.23302566,0.44964105,0.6892308,0.80738467,0.60389745,0.56451285,1.1552821,2.0578463,2.858667,3.0326157,3.6036925,4.2207184,4.824616,5.366154,5.8092313,3.5347695,2.048,1.2438976,0.98133343,1.0929232,2.8882053,4.273231,5.0642056,5.074052,4.132103,2.5435898,1.9692309,2.0020514,2.3072822,2.6289232,4.8147697,5.540103,5.1298466,4.2240005,3.8038976,5.9602056,5.7435904,4.6178465,3.7776413,4.1452312,7.5552826,9.028924,9.189744,8.52677,7.394462,6.665847,5.3202057,4.529231,5.037949,7.174565,7.250052,6.8397956,5.930667,4.5489235,2.7634873,2.2547693,2.2121027,2.5009232,2.9965131,3.5774362,4.5095387,5.586052,6.5345645,7.213949,7.6077952,7.6570263,8.772923,9.002667,7.5979495,4.9854364,3.7185643,3.0949745,2.7011285,2.3269746,1.975795,1.9823592,2.8291285,3.1474874,2.4352822,1.0502565,0.84348726,0.6859488,0.52512825,0.36430773,0.25928208,0.48574364,0.3446154,0.18051283,0.12471796,0.101743594,0.01969231,0.0,0.009846155,0.036102567,0.098461546,0.108307704,0.04266667,0.0,0.0,0.0,0.13128206,0.30194873,0.574359,0.90256417,1.1388719,1.083077,1.1848207,1.2964103,1.3357949,1.276718,1.1946667,1.3128207,1.4473847,1.5097437,1.522872,1.6114873,1.7033848,1.6508719,1.4539489,1.2832822,1.1520001,0.86646163,0.58092314,0.3708718,0.23958977,0.108307704,0.14112821,0.15753847,0.10502565,0.055794876,0.07548718,0.14112821,0.25928208,0.380718,0.3708718,0.26256412,0.31507695,0.30194873,0.18051283,0.10502565,0.07548718,0.04594872,0.04594872,0.06564103,0.029538464,0.016410258,0.0032820515,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.013128206,0.006564103,0.0,0.0,0.0,0.0032820515,0.006564103,0.016410258,0.04266667,0.06564103,0.08533334,0.08533334,0.072205134,0.059076928,0.15097436,0.21333335,0.18707694,0.098461546,0.059076928,0.059076928,0.07876924,0.12143591,0.21333335,0.41682056,0.7417436,1.0666667,1.463795,1.7099489,1.2964103,0.8467693,0.63343596,0.7515898,1.0043077,0.88943595,0.67938465,0.60389745,0.6465641,0.71548724,0.65312827,1.0010257,1.5392822,2.0808206,2.3204105,1.8051283,1.1782565,0.6498462,0.3446154,0.21333335,0.03938462,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016410258,0.06564103,0.055794876,0.04266667,0.036102567,0.03938462,0.04594872,0.068923086,0.08205129,0.09189744,0.0951795,0.072205134,0.072205134,0.059076928,0.049230773,0.04266667,0.036102567,0.052512825,0.098461546,0.15425642,0.20020515,0.20348719,0.14769232,0.11158975,0.08533334,0.055794876,0.013128206,0.013128206,0.01969231,0.036102567,0.049230773,0.04594872,0.052512825,0.049230773,0.03938462,0.029538464,0.026256412,0.055794876,0.098461546,0.128,0.13784617,0.12143591,0.108307704,0.19364104,0.43323082,0.88615394,1.6311796,1.9167181,1.6705642,1.3915899,1.4276924,1.9922053,2.162872,2.353231,2.4976413,2.477949,2.1530259,3.5478978,5.034667,6.0783596,6.2752824,5.3694363,4.4701543,4.4274874,4.844308,5.4974365,6.3277955,5.933949,7.0465646,8.704,9.987283,10.013539,9.957745,8.539898,7.171283,6.7249236,7.5520005,8.54318,9.911796,11.477334,12.616206,12.297847,8.769642,7.765334,7.781744,7.8047185,7.322257,7.7981544,8.293744,8.851693,9.511385,10.292514,9.7673855,8.809027,8.237949,8.55959,9.974154,12.015591,11.789129,11.67754,12.570257,13.856822,13.4170265,15.333745,16.928822,16.777847,14.716719,12.724514,13.850258,17.476925,22.472206,27.208208,27.096617,23.168001,19.003078,16.134565,14.076719,11.588924,8.769642,6.193231,4.164923,2.7273848,2.0086155,2.15959,2.0512822,1.4309745,0.92553854,1.3751796,0.8533334,0.28225642,0.052512825,0.0032820515,0.0,0.0,0.006564103,0.01969231,0.04266667,0.068923086,0.11158975,0.12471796,0.108307704,0.101743594,0.16082053,0.12143591,0.06564103,0.029538464,0.02297436,0.016410258,0.026256412,0.049230773,0.07876924,0.0951795,0.108307704,0.16410258,0.33805132,0.6629744,1.148718,1.595077,1.7460514,1.5556924,1.2668719,1.4112822,1.9331284,1.910154,2.0020514,2.5600002,3.6004105,4.585026,5.077334,5.1200004,5.0543594,5.5072823,6.8397956,8.914052,10.010257,9.685334,8.78277,8.845129,10.7848215,11.155693,9.42277,7.9983597,6.7807183,4.824616,3.4330258,3.170462,3.8728209,4.824616,5.149539,4.525949,3.4198978,3.0818465,3.121231,2.9538465,2.5632823,2.1398976,2.0808206,2.1956925,2.2350771,2.1300514,1.975795,2.034872,2.8258464,4.1583595,4.493129,3.8662567,3.892513,4.269949,4.644103,4.893539,5.1331286,5.737026,5.549949,4.535795,3.3411283,2.4516926,2.1956925,1.8543591,1.332513,1.0043077,0.9714873,1.0601027,1.6508719,2.5107694,2.930872,2.7437952,2.300718,2.477949,2.9735386,2.861949,2.048,1.2800001,0.88615394,0.8172308,1.083077,1.3883078,1.1224617,0.9321026,0.9878975,1.204513,1.5327181,1.9561027,9.110975,8.864821,8.795898,8.772923,8.4512825,7.2664623,6.882462,7.4896417,9.088,10.850462,11.145847,8.92718,7.722667,6.8562055,6.2555904,6.4656415,6.4656415,5.8256416,5.0018463,4.457026,4.640821,4.8016415,5.2545643,5.61559,5.477744,4.397949,4.2207184,3.7448208,3.0391798,2.7536411,4.1156926,5.093744,5.0674877,4.9985647,5.1922054,5.3136415,4.6211286,3.8564105,3.255795,2.802872,2.2219489,1.9593848,2.0644104,2.477949,3.242667,4.4964104,5.0215387,4.3684106,3.373949,2.5304618,1.9692309,1.522872,1.1520001,0.86317956,0.65969235,0.5677949,0.5907693,0.6268718,0.6498462,0.6695385,0.702359,0.8336411,0.99774367,1.0305642,0.96492314,1.0272821,0.9517949,0.8402052,0.69579494,0.5546667,0.47917953,0.4135385,0.35774362,0.30851284,0.2986667,0.37743592,0.37743592,0.33805132,0.27569234,0.21333335,0.18379489,0.13456412,0.09189744,0.06235898,0.04594872,0.02297436,0.016410258,0.016410258,0.02297436,0.03938462,0.059076928,0.108307704,0.16738462,0.21989745,0.23302566,0.15097436,0.12471796,0.118153855,0.1148718,0.10502565,0.08533334,0.16082053,0.21989745,0.16410258,0.052512825,0.108307704,0.2231795,0.256,0.20020515,0.0951795,0.04266667,0.026256412,0.029538464,0.01969231,0.0,0.0,0.04594872,0.13456412,0.23302566,0.28882053,0.2100513,0.32820517,0.42338464,0.46933338,0.46933338,0.446359,0.46933338,0.43323082,0.31507695,0.20676924,0.30851284,0.21989745,0.15097436,0.11158975,0.09189744,0.08533334,0.0951795,0.33476925,0.6826667,0.86974365,0.50543594,0.44964105,0.48574364,0.49230772,0.38400003,0.128,0.13784617,0.16738462,0.16738462,0.12471796,0.036102567,0.08533334,0.08533334,0.052512825,0.009846155,0.006564103,0.0,0.0032820515,0.009846155,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.009846155,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.01969231,0.036102567,0.07548718,0.22646156,0.380718,0.51856416,0.5973334,0.5513847,0.98461545,1.591795,2.1530259,2.422154,2.100513,2.3171284,3.0293336,3.876103,4.4865646,4.4734364,2.9997952,1.8642052,1.1881026,1.0732309,1.6016412,2.9407182,4.4045134,5.47118,5.61559,4.3290257,2.7963078,2.3401027,2.4451284,2.678154,2.7011285,3.383795,4.3651285,4.890257,4.6112823,3.6036925,5.175795,4.9920006,4.1682053,3.639795,4.161641,6.514872,6.987488,6.262154,4.9394875,3.5544617,4.07959,3.9942567,3.8498464,4.059898,4.906667,5.9536414,6.5969234,6.688821,6.1768208,5.0904617,3.7776413,3.0752823,2.7142565,2.5238976,2.4320002,3.2623591,4.0303593,4.706462,5.284103,5.786257,5.6385646,6.0652313,6.166975,5.504,4.1058464,3.1638978,2.6289232,2.2547693,1.9396925,1.719795,2.3696413,2.4713848,2.0217438,1.2603078,0.67938465,0.5152821,0.32164106,0.15425642,0.03938462,0.0,0.12143591,0.13456412,0.15425642,0.26584616,0.508718,0.41025645,0.26256412,0.15097436,0.12471796,0.2231795,0.36102566,0.4266667,0.46933338,0.512,0.5415385,0.5513847,0.57764107,0.74830776,1.0699488,1.4276924,1.0929232,0.88287187,0.7778462,0.75487185,0.7778462,0.96492314,1.1060513,1.1552821,1.1388719,1.1454359,1.404718,1.5721027,1.5786668,1.4178462,1.148718,1.0272821,0.7811283,0.5349744,0.34789747,0.20676924,0.13784617,0.118153855,0.09189744,0.052512825,0.032820515,0.04266667,0.108307704,0.21333335,0.3052308,0.31507695,0.16738462,0.17066668,0.18051283,0.16410258,0.16738462,0.13456412,0.072205134,0.02297436,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.016410258,0.009846155,0.0032820515,0.009846155,0.029538464,0.026256412,0.02297436,0.032820515,0.049230773,0.06564103,0.07876924,0.08533334,0.08533334,0.07548718,0.08861539,0.15425642,0.17394873,0.128,0.108307704,0.13456412,0.13784617,0.22646156,0.4201026,0.65641034,0.78769237,0.8566154,0.9714873,1.0666667,0.8992821,0.8402052,0.72861546,0.72861546,0.81066674,0.7253334,0.65969235,0.7811283,1.0765129,1.4244103,1.5786668,1.7690258,1.9528207,1.9528207,1.6410258,0.9353847,0.52512825,0.31507695,0.2297436,0.18707694,0.108307704,0.02297436,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.03938462,0.049230773,0.032820515,0.029538464,0.04266667,0.049230773,0.059076928,0.06564103,0.06235898,0.049230773,0.026256412,0.026256412,0.029538464,0.029538464,0.026256412,0.013128206,0.029538464,0.055794876,0.09189744,0.12143591,0.13784617,0.101743594,0.08533334,0.10502565,0.15425642,0.20676924,0.24287182,0.14769232,0.059076928,0.032820515,0.029538464,0.02297436,0.02297436,0.029538464,0.03938462,0.03938462,0.04266667,0.052512825,0.07548718,0.098461546,0.12143591,0.12471796,0.15097436,0.4135385,0.86974365,1.2471796,1.2274873,1.1651284,1.0502565,1.0404103,1.4736412,1.9561027,2.4352822,2.6190772,2.5271797,2.5009232,3.639795,4.7360005,5.2447186,5.182359,5.1364107,5.3234878,5.756718,6.2030773,6.449231,6.301539,6.0980515,6.8562055,7.4371285,7.4371285,7.174565,6.8496413,6.3540516,5.756718,5.3760004,5.786257,7.056411,8.530052,10.043077,11.414975,12.448821,11.083488,10.131693,9.5606165,9.216001,8.79918,8.67118,8.592411,9.708308,11.684103,12.714667,11.542975,9.537642,8.720411,9.770667,12.048411,14.375385,14.148924,13.052719,12.301129,12.645744,13.092104,15.133539,16.896002,17.237335,15.763694,14.644514,16.728617,21.018257,25.780516,28.566977,26.295797,21.248001,16.672821,13.840411,12.041847,9.970873,7.5487185,5.21518,3.3214362,2.1497438,1.7165129,1.7066668,1.5786668,1.1913847,0.79425645,0.827077,0.45620516,0.13128206,0.01969231,0.0,0.0,0.0,0.0032820515,0.013128206,0.036102567,0.068923086,0.12143591,0.14112821,0.12471796,0.10502565,0.11158975,0.08861539,0.055794876,0.032820515,0.02297436,0.016410258,0.02297436,0.052512825,0.09189744,0.12143591,0.13784617,0.15097436,0.21333335,0.3708718,0.65312827,0.9714873,1.0732309,1.0436924,0.9714873,0.9616411,1.214359,1.4473847,2.044718,2.7864618,2.868513,2.7667694,2.986667,3.5610259,4.6080003,6.3474874,8.316719,9.682052,9.711591,8.513641,7.0400004,7.821129,9.882257,10.154668,8.434873,7.394462,6.189949,3.8104618,2.3105643,2.3269746,3.1113849,4.3027697,5.0642056,5.100308,4.5817437,4.161641,3.7415388,3.239385,2.6880002,2.228513,2.0939488,2.1431797,2.1202054,2.0545642,2.100513,2.546872,3.7743592,5.034667,5.0051284,3.9220517,3.6102567,3.8662567,3.8990772,3.8006158,3.764513,4.089436,4.312616,4.082872,3.2623591,2.172718,1.591795,1.4309745,1.339077,1.273436,1.1815386,0.9747693,1.0502565,1.6246156,2.412308,2.865231,2.162872,1.8904617,2.3958976,2.6157951,2.1989746,1.5130258,1.1552821,0.88943595,1.020718,1.4572309,1.7132308,1.7920002,1.847795,1.8838975,1.972513,2.2514873,6.8529234,6.377026,6.925129,7.834257,8.093539,6.3212314,6.47877,8.195283,10.299078,11.753027,11.651283,10.04636,8.533334,7.3747697,6.803693,7.026872,5.87159,4.9854364,4.240411,3.7907696,4.069744,4.673641,5.910975,6.921847,7.02359,5.7140517,4.59159,3.7448208,2.8947694,2.4615386,3.5478978,4.8082056,4.7983594,4.342154,4.076308,4.4701543,4.516103,4.1583595,3.698872,3.259077,2.7700515,2.5009232,2.3433847,2.3860514,2.6945643,3.3345644,3.7251284,3.7316926,3.1803079,2.3269746,1.8838975,1.7920002,1.4769232,1.0765129,0.72861546,0.5677949,0.58092314,0.5907693,0.54482055,0.4660513,0.43323082,0.5316923,0.6826667,0.86974365,1.0666667,1.2373334,1.1323078,0.93866676,0.7417436,0.5874872,0.49230772,0.44964105,0.380718,0.31507695,0.2986667,0.38400003,0.38400003,0.3708718,0.3446154,0.3249231,0.3249231,0.27569234,0.19692309,0.13128206,0.08533334,0.055794876,0.049230773,0.049230773,0.055794876,0.06564103,0.07548718,0.15097436,0.27241027,0.4201026,0.5513847,0.61374366,0.46276927,0.35446155,0.2855385,0.24943592,0.24287182,0.24287182,0.2231795,0.18379489,0.16410258,0.256,0.38728207,0.36758977,0.24287182,0.098461546,0.049230773,0.04594872,0.059076928,0.06564103,0.052512825,0.01969231,0.055794876,0.10502565,0.16082053,0.190359,0.13128206,0.36102566,0.47261542,0.512,0.52512825,0.5546667,0.63343596,0.5513847,0.4135385,0.32820517,0.4135385,0.26584616,0.17723078,0.12471796,0.098461546,0.08533334,0.072205134,0.41025645,0.85005134,1.0404103,0.5481026,0.3117949,0.22646156,0.22646156,0.21661541,0.06564103,0.13128206,0.17723078,0.17723078,0.13456412,0.06235898,0.09189744,0.08205129,0.049230773,0.006564103,0.0,0.0,0.0,0.0,0.0,0.006564103,0.0,0.0,0.0032820515,0.006564103,0.006564103,0.016410258,0.01969231,0.016410258,0.006564103,0.0,0.0,0.0032820515,0.006564103,0.006564103,0.013128206,0.016410258,0.01969231,0.01969231,0.026256412,0.03938462,0.18707694,0.2986667,0.39384618,0.49887183,0.6432821,0.97805136,1.5392822,2.0939488,2.4188719,2.3072822,2.1136413,2.5698464,3.2787695,3.82359,3.764513,2.8291285,2.0906668,1.6771283,1.7066668,2.3040001,2.737231,3.6857438,4.5423594,4.7294364,3.6824617,2.7011285,2.556718,2.861949,3.0884104,2.5961027,2.3827693,3.4592824,4.4307694,4.6211286,4.056616,4.460308,4.1682053,3.7120004,3.5347695,3.9811285,4.9526157,4.7392826,3.876103,2.868513,2.1891284,2.8914874,3.564308,4.1747694,4.706462,5.146257,6.8299494,7.4043083,7.381334,7.2664623,7.568411,6.1440005,4.568616,3.0654361,1.9167181,1.4867693,1.9167181,2.300718,2.681436,3.0358977,3.2853336,3.1737437,3.2065644,3.249231,3.1770258,2.865231,2.3696413,1.913436,1.5425643,1.3029745,1.2340513,1.9462565,1.6049232,0.9419488,0.43651286,0.32164106,0.28225642,0.21661541,0.14112821,0.072205134,0.04266667,0.055794876,0.1148718,0.16082053,0.3117949,0.8566154,0.47917953,0.26256412,0.16410258,0.16082053,0.25271797,0.33476925,0.4135385,0.62030774,0.955077,1.2800001,1.2209232,1.1093334,1.0929232,1.2471796,1.5425643,1.083077,0.7318975,0.5021539,0.40697438,0.4660513,0.7778462,0.90256417,0.9189744,0.8763078,0.8336411,1.1782565,1.3522053,1.3259488,1.1454359,0.9288206,0.7450257,0.51856416,0.32820517,0.2100513,0.17723078,0.16082053,0.10502565,0.049230773,0.01969231,0.016410258,0.026256412,0.06235898,0.1148718,0.15753847,0.16738462,0.068923086,0.052512825,0.072205134,0.11158975,0.16082053,0.13128206,0.072205134,0.02297436,0.0,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.006564103,0.0,0.0,0.006564103,0.006564103,0.006564103,0.0032820515,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.006564103,0.006564103,0.006564103,0.006564103,0.006564103,0.006564103,0.0032820515,0.0,0.0,0.0,0.006564103,0.009846155,0.006564103,0.0032820515,0.009846155,0.029538464,0.032820515,0.036102567,0.049230773,0.055794876,0.06235898,0.08205129,0.0951795,0.0951795,0.07548718,0.06564103,0.108307704,0.13456412,0.13456412,0.16082053,0.18051283,0.20348719,0.36758977,0.6301539,0.764718,0.7253334,0.6268718,0.53825647,0.512,0.60061544,0.7975385,0.9189744,0.9747693,0.9288206,0.71548724,0.73517954,0.97805136,1.4342566,1.9692309,2.3335385,2.2711797,2.0709746,1.6640002,1.0732309,0.41025645,0.19692309,0.13456412,0.1148718,0.098461546,0.098461546,0.01969231,0.006564103,0.009846155,0.0032820515,0.0,0.0032820515,0.006564103,0.013128206,0.029538464,0.03938462,0.055794876,0.036102567,0.029538464,0.04266667,0.055794876,0.04594872,0.04266667,0.032820515,0.016410258,0.009846155,0.009846155,0.013128206,0.01969231,0.013128206,0.0,0.013128206,0.029538464,0.03938462,0.03938462,0.04594872,0.049230773,0.072205134,0.13456412,0.21661541,0.28225642,0.32164106,0.22646156,0.13784617,0.10502565,0.07876924,0.049230773,0.029538464,0.029538464,0.03938462,0.032820515,0.026256412,0.03938462,0.07876924,0.12471796,0.128,0.13456412,0.15425642,0.35774362,0.6826667,0.827077,0.79425645,0.9288206,1.0436924,1.1848207,1.6443079,1.9790771,2.356513,2.6486156,2.917744,3.4034874,4.338872,4.906667,4.6769233,4.059898,4.3060517,5.2315903,6.1997952,6.8660517,6.7249236,5.1232824,4.6080003,4.8640003,4.9985647,4.7917953,4.709744,4.3290257,4.7425647,5.028103,5.2053337,6.232616,6.7282057,7.1515903,7.837539,8.772923,9.586872,10.246565,10.233437,10.089026,9.852718,9.061745,8.36595,8.169026,9.301334,11.45436,13.184001,12.320822,10.55836,9.705027,10.541949,12.836103,15.471591,16.489027,16.17395,15.025232,13.745232,15.0088215,17.184822,19.423182,20.742565,20.01395,19.86954,22.35077,26.299078,29.824003,30.293335,25.652515,20.263386,15.809642,12.800001,10.594462,9.058462,6.9054365,4.7360005,3.0752823,2.3794873,1.8609232,1.3686155,1.014154,0.76800007,0.46276927,0.18707694,0.04594872,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.009846155,0.029538464,0.06235898,0.1148718,0.14441027,0.14441027,0.14112821,0.118153855,0.0951795,0.068923086,0.049230773,0.029538464,0.02297436,0.026256412,0.052512825,0.09189744,0.12143591,0.16738462,0.190359,0.2231795,0.29210258,0.37743592,0.47261542,0.512,0.6662565,0.8960001,0.955077,0.892718,1.4736412,3.2656412,5.4186673,5.7009234,3.9876926,2.7733335,2.7602053,4.269949,7.250052,10.322052,10.65354,9.403078,7.4371285,5.32677,5.5302567,6.9087186,7.24677,6.2194877,5.3924108,3.761231,1.9232821,1.0108719,1.204513,1.7427694,2.6322052,3.4888208,4.1682053,4.5587697,4.585026,3.9844105,3.2032824,2.5140514,2.0676925,1.8970258,1.8970258,1.8937438,2.0053334,2.3630772,3.121231,4.240411,4.9132314,4.5587697,3.515077,3.0293336,3.249231,3.1277952,2.8160002,2.5435898,2.6322052,3.0982566,3.367385,3.0982566,2.3827693,1.7526156,1.5163078,1.3587693,1.273436,1.211077,1.0699488,1.0404103,1.5163078,2.353231,2.9078977,2.0184617,1.2668719,1.4473847,1.7526156,1.7690258,1.4900514,1.2373334,0.9321026,1.0338463,1.6147693,2.3696413,2.5632823,2.4713848,2.3663592,2.4320002,2.7766156,6.3573337,5.83877,7.197539,8.687591,8.612103,5.333334,4.9460516,7.243488,9.754257,10.998155,10.476309,9.682052,9.38995,9.104411,8.681026,8.320001,6.055385,4.8640003,4.059898,3.3608208,2.8947694,3.7120004,5.9602056,7.9195905,8.664616,8.070564,5.5926156,3.9581542,2.9735386,2.6518977,3.2164104,5.1364107,4.5062566,3.2984617,2.7831798,3.5216413,4.7950773,5.0871797,4.7458467,4.0992823,3.4494362,2.8356924,2.487795,2.3958976,2.3991797,2.169436,1.910154,1.6869745,1.529436,1.4080001,1.2603078,1.522872,1.4244103,1.1684103,0.88943595,0.67282057,0.55794877,0.47589746,0.43651286,0.446359,0.52512825,0.6104616,0.7318975,0.8992821,1.0929232,1.2537436,1.204513,1.0043077,0.7515898,0.52512825,0.38400003,0.36430773,0.29210258,0.23302566,0.2231795,0.26584616,0.30194873,0.36102566,0.4135385,0.4397949,0.446359,0.41025645,0.31507695,0.2100513,0.13456412,0.101743594,0.101743594,0.108307704,0.12471796,0.14769232,0.18051283,0.24615386,0.42338464,0.7515898,1.1782565,1.5524104,1.142154,0.79425645,0.56451285,0.4660513,0.4660513,0.4266667,0.37743592,0.32820517,0.3052308,0.35446155,0.49230772,0.45620516,0.3249231,0.16738462,0.068923086,0.07548718,0.108307704,0.128,0.108307704,0.03938462,0.06564103,0.08533334,0.098461546,0.11158975,0.12471796,0.4266667,0.5349744,0.51856416,0.46276927,0.46276927,0.65969235,0.57764107,0.4266667,0.3511795,0.42994875,0.28225642,0.190359,0.13784617,0.118153855,0.13456412,0.06235898,0.3446154,0.636718,0.67282057,0.26912823,0.20348719,0.17066668,0.16082053,0.15425642,0.098461546,0.07876924,0.04266667,0.01969231,0.01969231,0.052512825,0.029538464,0.02297436,0.01969231,0.013128206,0.0,0.0,0.0,0.0,0.006564103,0.016410258,0.0032820515,0.0,0.006564103,0.016410258,0.016410258,0.036102567,0.036102567,0.02297436,0.006564103,0.0032820515,0.006564103,0.016410258,0.026256412,0.032820515,0.03938462,0.055794876,0.059076928,0.06235898,0.06564103,0.08861539,0.18379489,0.30851284,0.46276927,0.6498462,0.8730257,0.7122052,1.1158975,1.7723079,2.3696413,2.6190772,2.4320002,2.4746668,2.6387694,2.8389745,3.0096412,2.412308,2.3105643,2.5074873,2.8225644,3.0982566,2.7076926,2.5600002,2.5173335,2.4648206,2.3040001,1.8674873,1.9429746,2.409026,2.7963078,2.3072822,2.7700515,4.010667,4.8344617,5.0018463,5.2315903,4.886975,4.1682053,3.4658465,3.006359,2.8521028,3.2656412,3.117949,2.8291285,2.806154,3.43959,3.7021542,4.4438977,5.4514875,6.413129,6.961231,8.218257,8.027898,7.2205133,6.816821,8.01477,7.650462,6.048821,3.82359,1.7296412,0.67282057,0.67282057,0.90912825,1.1979488,1.3292309,1.0896411,1.148718,1.2603078,1.339077,1.3259488,1.1913847,0.9944616,0.7384616,0.47261542,0.27241027,0.23958977,0.318359,0.4135385,0.4660513,0.38728207,0.036102567,0.15097436,0.20348719,0.21661541,0.20348719,0.17723078,0.2231795,0.25928208,0.16410258,0.14769232,0.7450257,0.14769232,0.0,0.036102567,0.101743594,0.13784617,0.04594872,0.04266667,0.380718,1.017436,1.6377437,1.6147693,1.467077,1.3128207,1.2570257,1.3915899,1.0404103,0.82379496,0.69251287,0.6268718,0.6465641,0.80738467,0.88615394,0.9156924,0.92225647,0.9321026,1.1224617,1.0994873,0.9419488,0.7844103,0.8041026,0.5513847,0.30851284,0.15097436,0.10502565,0.15097436,0.118153855,0.07876924,0.04594872,0.029538464,0.01969231,0.03938462,0.032820515,0.029538464,0.036102567,0.026256412,0.006564103,0.0032820515,0.0032820515,0.0032820515,0.013128206,0.013128206,0.0032820515,0.0,0.0032820515,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.009846155,0.013128206,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.016410258,0.0032820515,0.0032820515,0.0,0.006564103,0.013128206,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.013128206,0.016410258,0.01969231,0.01969231,0.026256412,0.01969231,0.013128206,0.006564103,0.0032820515,0.0032820515,0.0032820515,0.006564103,0.016410258,0.01969231,0.01969231,0.026256412,0.036102567,0.04594872,0.049230773,0.052512825,0.08533334,0.1148718,0.118153855,0.08205129,0.08533334,0.09189744,0.10502565,0.13784617,0.2297436,0.2231795,0.30194873,0.48574364,0.65969235,0.5940513,0.48246157,0.46276927,0.4594872,0.48246157,0.6104616,0.7778462,1.1520001,1.3981539,1.3259488,0.8992821,0.98461545,1.1257436,1.4605129,1.9495386,2.3729234,2.228513,1.7887181,1.2668719,0.77128214,0.30851284,0.21333335,0.13128206,0.06235898,0.013128206,0.013128206,0.0032820515,0.013128206,0.02297436,0.016410258,0.016410258,0.04266667,0.049230773,0.055794876,0.068923086,0.07548718,0.07548718,0.049230773,0.029538464,0.029538464,0.03938462,0.016410258,0.013128206,0.006564103,0.0,0.0,0.0032820515,0.0032820515,0.006564103,0.006564103,0.006564103,0.02297436,0.055794876,0.06564103,0.03938462,0.006564103,0.026256412,0.07548718,0.15425642,0.22646156,0.21333335,0.21333335,0.20676924,0.2100513,0.2100513,0.14112821,0.08533334,0.052512825,0.03938462,0.03938462,0.029538464,0.026256412,0.052512825,0.12143591,0.19364104,0.18051283,0.19692309,0.24943592,0.3249231,0.4135385,0.512,0.764718,1.020718,1.273436,1.6311796,2.3138463,2.3040001,2.1858463,2.5632823,3.5610259,4.8114877,5.4514875,5.228308,4.201026,3.0391798,3.0227695,3.8596926,5.152821,6.183385,6.055385,3.6758976,2.737231,2.9604106,3.5741541,4.161641,4.667077,4.7327185,5.35959,5.8125134,6.3343596,8.14277,7.53559,6.6395903,6.442667,6.951385,7.1844106,8.093539,8.759795,9.258667,9.337437,8.41518,7.463385,7.6242056,8.15918,9.084719,11.201642,11.467488,11.369026,11.063796,11.067078,12.232206,14.7790785,17.329231,19.193438,19.64636,17.93641,18.566566,20.115694,22.055386,23.59795,23.699694,25.363695,28.143593,31.031797,32.676105,31.389542,25.5639,20.545643,16.469334,13.184001,10.256411,8.743385,6.564103,4.516103,3.1671798,2.8553848,2.1398976,1.3686155,0.81066674,0.50543594,0.23302566,0.059076928,0.006564103,0.0032820515,0.0,0.0,0.0,0.006564103,0.013128206,0.016410258,0.029538464,0.055794876,0.101743594,0.13784617,0.16082053,0.16082053,0.13784617,0.118153855,0.101743594,0.08533334,0.059076928,0.03938462,0.032820515,0.049230773,0.07548718,0.08533334,0.12143591,0.18379489,0.27897438,0.3708718,0.39712822,0.3511795,0.42994875,0.65969235,0.99774367,1.332513,1.3128207,2.0611284,4.5522056,7.9852314,9.780514,6.928411,3.9548721,2.7831798,4.1156926,7.427283,10.896411,10.541949,8.786052,6.944821,5.208616,4.3060517,4.066462,4.2568207,4.4045134,3.8071797,1.9692309,1.1158975,0.8369231,0.85005134,0.9747693,1.4375386,2.0250258,2.7536411,3.5413337,4.201026,3.82359,3.0227695,2.2613335,1.7723079,1.5753847,1.5589745,1.6344616,1.9462565,2.546872,3.4034874,3.9647183,4.0500517,3.6463592,2.9735386,2.4943593,2.6190772,2.546872,2.225231,1.8346668,1.7690258,2.294154,2.5206156,2.6387694,2.6518977,2.3991797,2.1366155,1.6213335,1.2438976,1.1552821,1.2668719,1.6147693,2.409026,3.1803079,3.3476925,2.2547693,1.2668719,1.0732309,1.1716924,1.270154,1.2865642,1.142154,1.079795,1.3850257,2.0742567,2.8816411,2.8225644,2.5206156,2.481231,2.9571285,3.95159,11.52,10.299078,9.416205,10.55836,12.071385,8.973129,4.637539,3.1442053,3.3772311,4.7261543,7.0957956,9.573745,10.962052,11.608616,11.237744,8.940309,5.681231,3.56759,2.737231,2.8356924,3.006359,3.6660516,5.4875903,7.1548724,7.8506675,7.27959,5.8125134,4.4045134,3.0982566,2.349949,3.0227695,4.4242053,4.0434875,3.69559,4.1682053,5.218462,6.498462,6.6560006,5.8814363,4.5587697,3.2656412,2.1070771,1.4966155,1.4112822,1.7066668,2.1202054,2.1333334,1.6869745,1.4080001,1.4080001,1.2964103,0.9419488,0.7811283,0.71548724,0.67282057,0.6104616,0.47589746,0.40697438,0.4004103,0.4397949,0.48902568,0.52512825,0.7450257,1.0010257,1.204513,1.3259488,1.1815386,0.9353847,0.69579494,0.51856416,0.39712822,0.34789747,0.25271797,0.19692309,0.20348719,0.2297436,0.26584616,0.34789747,0.40369233,0.4201026,0.45620516,0.48246157,0.4135385,0.3117949,0.2100513,0.13784617,0.13784617,0.13784617,0.19364104,0.30194873,0.4135385,0.49887183,0.8467693,1.5195899,2.3236926,2.8225644,2.1398976,1.4375386,0.9485129,0.7220513,0.6268718,0.5152821,0.37743592,0.28225642,0.256,0.3052308,0.40369233,0.41682056,0.33805132,0.19364104,0.04594872,0.02297436,0.02297436,0.02297436,0.016410258,0.016410258,0.0032820515,0.01969231,0.036102567,0.06564103,0.13784617,0.5152821,0.88615394,0.95835906,0.6826667,0.24287182,0.4397949,0.4135385,0.34789747,0.32164106,0.32164106,0.17394873,0.108307704,0.14112821,0.24287182,0.36758977,0.14769232,0.35774362,0.54482055,0.49887183,0.24287182,0.318359,0.23630771,0.118153855,0.036102567,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.052512825,0.08861539,0.0951795,0.06235898,0.0,0.0,0.0,0.006564103,0.016410258,0.016410258,0.0032820515,0.0,0.006564103,0.016410258,0.016410258,0.026256412,0.03938462,0.03938462,0.026256412,0.016410258,0.026256412,0.049230773,0.072205134,0.08861539,0.07548718,0.101743594,0.1148718,0.14769232,0.2100513,0.32164106,0.40697438,0.5284103,0.69251287,0.8960001,1.1290257,1.591795,1.7001027,1.4802053,0.98133343,0.27569234,1.0436924,1.7657437,2.176,2.044718,1.1913847,1.4342566,2.1989746,3.18359,4.086154,4.6244106,3.170462,1.8543591,0.8369231,0.28882053,0.4135385,0.37415388,0.7417436,1.3587693,2.172718,3.2361028,4.027077,4.9854364,5.7140517,5.7435904,4.5456414,3.6069746,3.0687182,2.678154,2.1202054,1.024,1.6213335,1.5786668,1.2537436,1.204513,2.1825643,3.1967182,4.46359,5.6320004,6.045539,4.775385,5.349744,5.1265645,4.4373336,4.023795,5.034667,7.072821,7.584821,6.629744,4.3684106,1.0371283,0.5481026,0.5907693,0.83035904,1.017436,0.9911796,0.8467693,0.7089231,0.5677949,0.4201026,0.27569234,0.22646156,0.19692309,0.108307704,0.07876924,0.39712822,0.41025645,0.4201026,0.446359,0.4135385,0.18379489,0.12143591,0.1148718,0.17723078,0.2986667,0.45620516,0.54482055,0.46276927,0.23958977,0.0,0.0,0.0,0.0,0.036102567,0.08861539,0.07548718,0.101743594,0.21661541,0.4135385,0.636718,0.80738467,0.88287187,0.9189744,0.90584624,0.93866676,1.2209232,1.0732309,0.98133343,1.0075898,1.0502565,0.8533334,0.6826667,0.60389745,0.65312827,0.88287187,1.3587693,1.1520001,0.85005134,0.6498462,0.6301539,0.7778462,0.54482055,0.2855385,0.13456412,0.10502565,0.09189744,0.06564103,0.052512825,0.03938462,0.029538464,0.029538464,0.029538464,0.02297436,0.009846155,0.0032820515,0.016410258,0.016410258,0.02297436,0.01969231,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.016410258,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.016410258,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.02297436,0.029538464,0.029538464,0.06564103,0.07548718,0.059076928,0.026256412,0.016410258,0.016410258,0.016410258,0.03938462,0.07876924,0.09189744,0.09189744,0.055794876,0.036102567,0.049230773,0.06235898,0.072205134,0.13128206,0.20348719,0.26584616,0.28882053,0.20348719,0.14769232,0.15753847,0.23958977,0.3511795,0.4135385,0.508718,0.5218462,0.43651286,0.3511795,0.3249231,0.32164106,0.3314872,0.36758977,0.4266667,0.63343596,1.0633847,1.2635899,1.1946667,1.204513,1.4736412,1.2668719,1.1388719,1.2996924,1.6180514,1.6672822,1.1290257,0.64000005,0.47917953,0.56451285,0.5284103,0.27241027,0.068923086,0.013128206,0.0,0.0,0.0,0.013128206,0.03938462,0.07548718,0.16082053,0.18379489,0.17066668,0.13784617,0.07548718,0.06564103,0.04266667,0.02297436,0.016410258,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.013128206,0.02297436,0.029538464,0.029538464,0.029538464,0.06564103,0.15097436,0.16738462,0.10502565,0.029538464,0.029538464,0.06564103,0.14769232,0.23958977,0.27569234,0.22646156,0.14112821,0.09189744,0.09189744,0.09189744,0.06564103,0.06235898,0.06564103,0.07876924,0.09189744,0.06564103,0.052512825,0.108307704,0.2297436,0.3511795,0.43651286,0.47589746,0.45620516,0.4135385,0.4266667,0.6104616,0.95835906,1.2504616,1.5064616,1.9823592,2.7634873,2.5304618,3.1277952,5.031385,7.3386674,7.1187696,6.1407185,4.9788723,3.9844105,3.2656412,3.5577438,4.023795,4.1058464,3.7218463,3.2951798,3.3444104,3.8498464,4.2601027,4.44718,4.716308,6.117744,7.5421543,8.195283,8.129642,8.241231,7.5552826,7.394462,8.119796,9.45559,10.466462,11.552821,10.86359,9.593436,8.369231,7.2336416,7.0498466,7.325539,7.282872,7.1581545,8.208411,9.6984625,10.630565,11.0145645,10.985026,10.804514,11.195078,14.112822,17.664001,20.502975,21.819078,20.086155,20.056618,20.568617,21.185642,22.186668,26.006977,28.94113,30.660925,31.025232,30.06031,25.678772,21.349745,17.253744,13.61395,10.696206,8.254359,5.8880005,3.895795,2.428718,1.463795,1.404718,0.83035904,0.27569234,0.0,0.0,0.013128206,0.016410258,0.009846155,0.0,0.0,0.0,0.0,0.0,0.006564103,0.029538464,0.06564103,0.15097436,0.21661541,0.2231795,0.13784617,0.16082053,0.17723078,0.19692309,0.20348719,0.16738462,0.068923086,0.04594872,0.052512825,0.072205134,0.12143591,0.06235898,0.055794876,0.13456412,0.3117949,0.58092314,0.60389745,0.7187693,0.86646163,1.1388719,1.785436,2.6157951,2.9604106,4.0402055,6.6428723,11.122872,9.170052,6.055385,4.027077,3.8038976,4.5489235,5.0838976,4.900103,4.460308,4.2436924,4.7458467,5.940513,5.7009234,4.890257,3.882667,2.5632823,2.2088206,1.975795,1.7132308,1.3883078,1.083077,1.6935385,2.2580514,2.8750772,3.6036925,4.4701543,4.1911798,3.4888208,2.6518977,1.9298463,1.5261539,1.5392822,1.6147693,1.8773335,2.3762052,3.0982566,3.2196925,3.0227695,2.6354873,2.2383592,2.028308,1.8838975,1.6804104,1.4736412,1.3062565,1.2209232,2.0873847,2.2678976,2.1398976,2.0578463,2.349949,2.802872,2.6026669,2.0118976,1.4244103,1.3883078,1.9495386,3.190154,4.397949,4.7458467,3.2820516,2.048,1.4933335,1.204513,0.9944616,0.88615394,1.142154,1.6082052,2.1333334,2.5862565,2.868513,2.3302567,2.1136413,2.5009232,3.7087183,5.904411,8.822155,6.705231,6.166975,7.276308,9.26195,10.545232,7.433847,5.4449234,4.965744,5.8092313,7.2303596,10.059488,12.173129,13.078976,12.304411,9.40636,6.633026,4.7458467,3.876103,4.197744,5.910975,5.2414365,4.8344617,5.139693,5.802667,5.677949,5.182359,4.6276927,4.0533338,3.7087183,4.0467696,4.082872,3.820308,3.7907696,4.3749747,5.8157954,6.422975,6.12759,4.857436,3.0982566,1.8609232,1.2209232,0.9714873,1.086359,1.7066668,3.1474874,3.5183592,3.121231,2.3072822,1.4966155,1.1618463,1.014154,0.99774367,1.0633847,1.083077,0.86646163,0.67282057,0.56123084,0.46933338,0.40369233,0.40369233,0.51856416,0.7417436,0.96492314,1.0962052,1.0699488,0.9156924,0.7318975,0.62030774,0.574359,0.48246157,0.36430773,0.21661541,0.18051283,0.26256412,0.3249231,0.40369233,0.508718,0.508718,0.42994875,0.45620516,0.46276927,0.37743592,0.26256412,0.16738462,0.11158975,0.11158975,0.13456412,0.23302566,0.38728207,0.49887183,0.96492314,2.0545642,3.117949,3.6890259,3.5052311,2.609231,1.6902566,1.1290257,0.9682052,0.9321026,0.83035904,0.49887183,0.24943592,0.18707694,0.19692309,0.28225642,0.43651286,0.4135385,0.21989745,0.08205129,0.08861539,0.20020515,0.2100513,0.09189744,0.0032820515,0.0,0.009846155,0.04266667,0.11158975,0.23630771,0.50543594,0.8041026,0.9747693,0.9682052,0.84348726,0.7844103,0.6301539,0.49887183,0.43323082,0.39384618,0.33476925,0.19692309,0.17394873,0.3314872,0.6104616,0.8992821,0.69251287,0.44964105,0.33805132,0.256,0.21333335,0.14441027,0.08861539,0.055794876,0.049230773,0.068923086,0.059076928,0.04266667,0.032820515,0.016410258,0.013128206,0.128,0.19692309,0.16410258,0.072205134,0.032820515,0.016410258,0.009846155,0.006564103,0.016410258,0.0032820515,0.0,0.0,0.0032820515,0.0032820515,0.055794876,0.10502565,0.14112821,0.14441027,0.11158975,0.1148718,0.11158975,0.14112821,0.20676924,0.28225642,0.21989745,0.21989745,0.24615386,0.27241027,0.28225642,0.3117949,0.49887183,0.94523084,1.6869745,2.678154,2.1070771,2.176,2.2153847,1.7460514,0.48246157,0.8402052,1.5721027,2.176,2.2383592,1.4211283,1.1290257,1.782154,2.6518977,3.045744,2.3040001,1.3193847,0.67938465,0.3249231,0.2100513,0.30194873,0.3052308,0.5415385,1.0502565,1.9200002,3.2951798,3.318154,3.1967182,3.0884104,2.7536411,1.5688206,1.204513,1.2438976,1.6311796,2.3171284,3.2820516,3.8006158,3.9154875,3.8137438,3.7940516,4.2338467,4.6211286,4.854154,4.8016415,4.2272825,2.809436,3.8629746,4.630975,4.8147697,4.240411,2.8488207,4.059898,5.2676926,6.045539,5.7042055,3.308308,2.156308,1.972513,2.6912823,3.4002054,2.359795,1.4309745,0.79097444,0.5152821,0.571077,0.82379496,0.7056411,0.60061544,0.6235898,0.764718,0.8960001,0.67610264,0.4397949,0.30194873,0.25271797,0.15753847,0.108307704,0.052512825,0.15753847,0.3314872,0.22646156,0.17394873,0.11158975,0.049230773,0.0,0.0,0.0,0.0,0.006564103,0.03938462,0.12471796,0.29538465,0.5218462,0.6695385,0.67938465,0.57764107,0.571077,0.6695385,0.79425645,0.84348726,0.69579494,0.5284103,0.5218462,0.764718,1.0765129,0.9878975,0.6629744,0.46933338,0.4004103,0.40697438,0.40697438,0.27569234,0.18051283,0.13128206,0.14112821,0.2297436,0.23958977,0.24943592,0.18379489,0.07548718,0.04266667,0.029538464,0.016410258,0.016410258,0.029538464,0.029538464,0.049230773,0.08861539,0.07876924,0.01969231,0.0032820515,0.0032820515,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0032820515,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.009846155,0.01969231,0.036102567,0.055794876,0.06564103,0.06235898,0.03938462,0.049230773,0.036102567,0.04594872,0.0951795,0.16410258,0.14441027,0.12471796,0.101743594,0.08205129,0.08533334,0.21333335,0.27241027,0.26912823,0.20348719,0.08205129,0.06564103,0.068923086,0.098461546,0.15425642,0.21661541,0.28882053,0.42994875,0.5546667,0.60061544,0.5349744,0.49887183,0.46276927,0.4266667,0.4266667,0.53825647,0.55794877,0.7056411,0.8402052,0.90912825,0.9485129,1.8510771,2.0020514,1.7263591,1.4572309,1.7165129,1.7920002,1.3718976,0.74830776,0.22646156,0.13784617,0.12143591,0.06564103,0.02297436,0.0032820515,0.0,0.0,0.0,0.0032820515,0.013128206,0.03938462,0.19364104,0.28225642,0.3052308,0.26912823,0.19692309,0.15753847,0.12143591,0.09189744,0.06564103,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.0032820515,0.01969231,0.055794876,0.09189744,0.09189744,0.08861539,0.11158975,0.13784617,0.15097436,0.128,0.08861539,0.055794876,0.059076928,0.08861539,0.1148718,0.10502565,0.07548718,0.04594872,0.032820515,0.04266667,0.029538464,0.03938462,0.06564103,0.10502565,0.17723078,0.17066668,0.15425642,0.20348719,0.3117949,0.37415388,0.46933338,0.5415385,0.5152821,0.47261542,0.67282057,0.79425645,0.93866676,1.2865642,1.7296412,1.8740515,2.2350771,2.6420515,3.5577438,4.896821,6.0324106,6.340924,6.409847,5.927385,4.8705645,3.498667,3.2623591,4.082872,4.082872,3.121231,2.7700515,2.9571285,3.3805132,3.817026,4.138667,4.2994876,4.824616,5.7501545,7.2861543,8.582564,7.716103,7.5191803,10.673231,13.016617,13.315283,13.275898,12.07795,9.849437,7.4010262,5.290667,3.8038976,3.7284105,3.895795,4.1911798,4.9296412,6.87918,8.89436,8.618668,7.899898,7.7390776,8.28718,9.334154,10.794667,12.806565,15.225437,17.657436,19.098257,19.216412,18.884924,18.835693,19.672617,22.12431,25.3079,28.054977,29.377644,28.471798,24.050873,19.75795,16.022976,12.944411,10.282667,7.643898,4.955898,2.9669745,1.8412309,1.1585642,0.76800007,0.38728207,0.12471796,0.013128206,0.02297436,0.036102567,0.032820515,0.016410258,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.02297436,0.04266667,0.10502565,0.20676924,0.29538465,0.29210258,0.23958977,0.23302566,0.28225642,0.31507695,0.17723078,0.108307704,0.11158975,0.18707694,0.3052308,0.30194873,0.37743592,0.49230772,0.6301539,0.81066674,0.8763078,0.8992821,0.9911796,1.2635899,1.8346668,3.114667,5.277539,6.925129,7.2336416,5.973334,3.8137438,2.477949,1.9396925,2.048,2.5074873,2.986667,3.5183592,4.3585644,5.681231,7.5881033,8.425026,8.832001,8.950154,8.772923,8.178872,8.556309,7.962257,6.8266673,5.792821,5.720616,3.889231,2.9965131,2.7569232,2.8291285,2.7864618,2.7109745,2.6157951,2.425436,2.0906668,1.5983591,1.5425643,1.6311796,1.8445129,2.156308,2.5238976,2.6354873,2.5600002,2.3466668,2.0578463,1.7624617,1.5360001,1.3095386,1.1388719,1.1027694,1.2832822,1.4539489,1.394872,1.3423591,1.5721027,2.412308,2.9604106,2.8455386,2.2514873,1.5688206,1.3751796,1.7132308,3.058872,4.955898,6.114462,4.414359,3.2623591,2.5632823,2.1464617,1.7624617,1.1060513,1.0765129,1.5261539,2.3335385,3.0752823,3.0030773,2.4549747,2.038154,1.9200002,2.428718,4.0500517,5.5663595,4.8344617,4.9132314,5.8125134,7.315693,8.999385,8.631796,8.996103,9.449026,9.655796,9.586872,9.911796,11.378873,12.3306675,11.828514,9.649232,6.5378466,5.093744,5.0871797,6.2490263,8.277334,7.6110773,6.9842057,6.439385,5.805949,4.6933336,4.1813335,3.948308,3.82359,3.7809234,3.9286156,3.5413337,3.3608208,3.511795,4.1222568,5.3169236,5.8814363,5.297231,3.9417439,2.3040001,0.97805136,0.7220513,0.7417436,0.9878975,1.5195899,2.5140514,2.7733335,2.5107694,1.9200002,1.276718,0.94523084,0.9714873,0.99774367,1.0108719,0.9682052,0.79425645,0.6892308,0.6170257,0.54482055,0.46933338,0.43651286,0.446359,0.508718,0.5874872,0.6465641,0.65969235,0.63343596,0.5907693,0.5677949,0.55794877,0.5316923,0.36102566,0.22646156,0.23302566,0.37415388,0.5349744,0.6629744,0.7220513,0.6235898,0.46933338,0.5316923,0.508718,0.41682056,0.2986667,0.20020515,0.18051283,0.25271797,0.34789747,0.48246157,0.761436,1.3686155,2.4516926,3.8629746,5.0477953,5.4482055,4.493129,3.5314875,2.0611284,1.1585642,1.020718,0.9517949,0.7515898,0.40369233,0.16738462,0.10502565,0.11158975,0.21989745,0.38400003,0.3708718,0.18707694,0.072205134,0.055794876,0.11158975,0.13456412,0.09189744,0.026256412,0.026256412,0.068923086,0.2986667,0.6465641,0.8172308,0.8992821,0.96492314,1.0436924,1.1158975,1.1093334,0.9944616,0.827077,0.6892308,0.57764107,0.4135385,0.25928208,0.15097436,0.15425642,0.27569234,0.46933338,0.7515898,0.81394875,0.65641034,0.39712822,0.25928208,0.23630771,0.15425642,0.09189744,0.07876924,0.068923086,0.049230773,0.03938462,0.07876924,0.14441027,0.14441027,0.04266667,0.15425642,0.21989745,0.15425642,0.06564103,0.08205129,0.055794876,0.026256412,0.01969231,0.02297436,0.026256412,0.016410258,0.009846155,0.013128206,0.026256412,0.06564103,0.0951795,0.16082053,0.256,0.32164106,0.21661541,0.20348719,0.23958977,0.29210258,0.3446154,0.29538465,0.26912823,0.26912823,0.28882053,0.32164106,0.35446155,0.4397949,0.7417436,1.3554872,2.297436,2.6978464,2.6584618,2.2744617,1.6147693,0.7187693,0.8205129,1.1552821,1.5622566,1.8806155,1.975795,1.3489232,1.3751796,1.7033848,1.9954873,1.9429746,1.0338463,0.512,0.28225642,0.24615386,0.30194873,0.5481026,0.73517954,0.9419488,1.2832822,1.9003079,1.7887181,1.6278975,1.5589745,1.591795,1.6016412,1.0666667,1.0469744,1.6705642,2.930872,4.6769233,5.3825645,5.5663595,5.3694363,5.034667,4.900103,5.2578464,5.3792825,5.0838976,4.4832826,3.9680004,3.6594875,3.570872,3.8695388,3.9056413,2.1956925,2.6387694,3.4002054,3.9187696,4.059898,4.141949,3.1737437,2.2711797,2.034872,2.300718,2.1333334,1.8806155,1.6246156,1.4080001,1.3915899,1.847795,1.5261539,0.9288206,0.6695385,0.78769237,0.7581539,0.61374366,0.5546667,0.761436,0.99774367,0.5907693,0.29538465,0.25928208,0.38400003,0.4955898,0.3249231,0.3117949,0.47917953,0.51856416,0.36758977,0.21989745,0.101743594,0.029538464,0.0,0.009846155,0.055794876,0.13784617,0.63343596,0.9616411,0.98133343,0.9944616,1.1027694,1.2438976,1.2865642,1.1618463,0.8402052,0.58092314,0.54482055,0.7318975,0.98461545,0.9682052,0.7318975,0.5907693,0.47917953,0.35446155,0.20348719,0.08861539,0.029538464,0.006564103,0.006564103,0.036102567,0.06564103,0.0951795,0.07876924,0.029538464,0.02297436,0.009846155,0.0032820515,0.009846155,0.026256412,0.03938462,0.06564103,0.072205134,0.049230773,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.013128206,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.026256412,0.01969231,0.006564103,0.0032820515,0.009846155,0.016410258,0.013128206,0.026256412,0.036102567,0.049230773,0.08205129,0.07876924,0.049230773,0.052512825,0.0951795,0.13784617,0.11158975,0.09189744,0.108307704,0.14769232,0.15425642,0.20348719,0.19692309,0.15425642,0.0951795,0.03938462,0.055794876,0.055794876,0.07876924,0.15097436,0.27569234,0.37743592,0.39056414,0.44964105,0.571077,0.6629744,0.7515898,0.761436,0.6465641,0.47589746,0.446359,0.45620516,0.57764107,0.6662565,0.75487185,1.020718,2.0250258,2.9505644,3.0260515,2.3630772,1.9790771,1.6968206,1.0666667,0.46933338,0.11158975,0.02297436,0.009846155,0.013128206,0.013128206,0.006564103,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.108307704,0.18051283,0.2100513,0.19692309,0.17394873,0.17723078,0.13784617,0.09189744,0.052512825,0.006564103,0.0,0.0,0.0,0.0,0.0,0.006564103,0.016410258,0.032820515,0.052512825,0.052512825,0.055794876,0.052512825,0.06564103,0.08533334,0.08861539,0.06235898,0.04594872,0.04594872,0.055794876,0.06564103,0.0951795,0.08533334,0.06235898,0.04594872,0.059076928,0.052512825,0.068923086,0.08533334,0.0951795,0.108307704,0.12143591,0.16082053,0.24287182,0.34789747,0.41682056,0.67610264,0.8566154,0.92225647,0.88615394,0.81394875,0.69907695,0.69251287,0.88287187,1.1618463,1.2504616,1.6180514,2.1136413,2.7273848,3.2656412,3.3542566,3.8006158,5.2480006,6.7840004,7.0334363,4.141949,3.767795,4.269949,4.325744,3.629949,2.8947694,3.3214362,3.8465643,4.135385,4.312616,4.97559,5.21518,5.8978467,7.2205133,8.52677,8.326565,8.493949,10.8767185,13.548308,15.199181,15.156514,12.708103,10.128411,8.224821,6.6822567,4.0533338,3.131077,2.9210258,3.6529233,4.827898,5.1987696,5.7009234,5.58277,6.242462,7.702975,8.612103,9.212719,9.90195,11.109744,12.842668,14.667488,16.403694,17.526155,18.75036,20.243694,21.661541,23.341951,25.606565,27.776003,28.918156,27.864618,23.67672,18.70113,14.785643,12.251899,9.895386,7.3091288,4.634257,2.7963078,1.8871796,1.1651284,0.5940513,0.23958977,0.06564103,0.013128206,0.013128206,0.016410258,0.01969231,0.016410258,0.009846155,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.055794876,0.13784617,0.24287182,0.28225642,0.26584616,0.32820517,0.48574364,0.6432821,0.67282057,0.65641034,0.6629744,0.702359,0.7253334,0.636718,0.49230772,0.43323082,0.52512825,0.7515898,0.9714873,1.0568206,1.1355898,1.2964103,1.5885129,2.3072822,3.4067695,4.568616,5.3727183,5.297231,4.8082056,3.3936412,2.1366155,1.6213335,1.9167181,2.5928206,5.0642056,7.6996927,9.478565,9.984001,8.027898,8.635077,9.741129,9.895386,8.274052,7.7718983,6.7905645,5.402257,4.135385,3.9712822,3.249231,2.8980515,2.806154,2.7437952,2.3729234,2.3204105,2.294154,2.1792822,1.913436,1.4900514,1.4539489,1.5491283,1.7263591,1.9429746,2.1431797,2.353231,2.3893335,2.2547693,1.9823592,1.6311796,1.3193847,1.0305642,0.8336411,0.8336411,1.1520001,1.3981539,1.4309745,1.4244103,1.6410258,2.4352822,2.993231,2.9407182,2.3663592,1.6377437,1.3817437,1.657436,2.5042052,3.6693337,4.460308,3.7284105,3.3542566,3.1934361,3.0884104,2.802872,2.0020514,1.6114873,1.6672822,2.2022567,2.989949,3.5478978,3.255795,2.733949,2.2482052,2.1366155,2.8160002,4.890257,5.533539,6.12759,6.7117953,7.64718,9.609847,10.925949,11.759591,11.47077,10.489437,10.328616,10.105436,11.201642,11.969642,11.533129,9.803488,6.885744,5.8814363,6.518154,8.201847,9.997129,9.974154,9.288206,7.8539495,5.8945646,3.9548721,3.1409233,2.861949,2.8389745,2.9078977,2.9997952,2.868513,3.0293336,3.748103,4.818052,5.5663595,5.6943593,4.8049235,3.4002054,1.9167181,0.72861546,0.6301539,0.67282057,0.95835906,1.4441026,1.9298463,2.1300514,1.8182565,1.3981539,1.0732309,0.8467693,0.8960001,0.8992821,0.8533334,0.77456415,0.702359,0.761436,0.7089231,0.63343596,0.571077,0.5284103,0.4397949,0.39712822,0.38400003,0.38728207,0.4135385,0.4266667,0.44964105,0.45292312,0.42994875,0.41025645,0.3314872,0.39056414,0.571077,0.82379496,1.0601027,1.0601027,0.98133343,0.80738467,0.64000005,0.6892308,0.7318975,0.6662565,0.56451285,0.49887183,0.55794877,0.636718,0.79425645,1.079795,1.6607181,2.8422565,4.2436924,5.602462,6.6002054,6.485334,4.0467696,3.242667,2.0086155,1.3193847,1.2537436,0.9944616,0.65641034,0.33476925,0.13784617,0.07876924,0.068923086,0.13784617,0.22646156,0.21661541,0.1148718,0.055794876,0.029538464,0.04594872,0.118153855,0.18707694,0.12471796,0.13128206,0.31507695,0.9517949,1.657436,1.3981539,1.2504616,1.211077,1.1913847,1.1158975,0.9156924,0.83035904,0.83035904,0.7318975,0.5152821,0.32164106,0.16738462,0.118153855,0.14441027,0.2231795,0.32820517,0.46276927,0.6432821,0.6826667,0.5546667,0.4004103,0.3446154,0.256,0.20348719,0.190359,0.15097436,0.09189744,0.07876924,0.13128206,0.21661541,0.27897438,0.2297436,0.28882053,0.26912823,0.15425642,0.06564103,0.101743594,0.072205134,0.04266667,0.03938462,0.04266667,0.049230773,0.036102567,0.026256412,0.026256412,0.04594872,0.07548718,0.08861539,0.14441027,0.24287182,0.33805132,0.26912823,0.30851284,0.37743592,0.42994875,0.4594872,0.4201026,0.3446154,0.3117949,0.35446155,0.44964105,0.512,0.49887183,0.7122052,1.2832822,2.176,2.8455386,2.681436,2.166154,1.6377437,1.2964103,1.142154,1.404718,1.7788719,2.038154,2.034872,1.4900514,1.1913847,1.1323078,1.3062565,1.6935385,1.0469744,0.67282057,0.5546667,0.58420515,0.571077,0.9189744,0.98133343,0.9124103,0.88287187,1.0699488,1.0469744,1.1552821,1.3653334,1.5983591,1.723077,1.394872,1.4900514,2.0611284,2.9735386,3.892513,4.818052,5.2414365,5.142975,4.716308,4.352,4.7458467,5.024821,4.893539,4.535795,4.6080003,3.5347695,2.878359,3.245949,3.820308,2.3827693,2.2186668,2.3991797,2.550154,2.6945643,3.2689233,2.7569232,2.1103592,1.591795,1.4145643,1.7362052,1.8215386,1.6968206,1.4966155,1.4112822,1.7033848,1.5195899,1.1684103,0.8960001,0.75487185,0.5907693,0.53825647,0.58420515,0.9485129,1.3686155,1.086359,0.7778462,0.65312827,0.636718,0.62030774,0.46276927,0.318359,0.574359,0.62030774,0.36758977,0.21989745,0.17723078,0.09189744,0.09189744,0.17723078,0.22646156,0.20020515,0.58420515,0.90584624,1.0404103,1.214359,1.3357949,1.3587693,1.2898463,1.1454359,0.955077,0.7450257,0.65641034,0.65641034,0.6859488,0.6695385,0.6498462,0.5481026,0.40697438,0.26912823,0.19364104,0.24943592,0.18379489,0.0951795,0.03938462,0.029538464,0.016410258,0.009846155,0.009846155,0.016410258,0.032820515,0.006564103,0.0032820515,0.01969231,0.052512825,0.108307704,0.07876924,0.04266667,0.013128206,0.0,0.0,0.0032820515,0.006564103,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.009846155,0.006564103,0.0,0.0,0.0,0.0032820515,0.009846155,0.006564103,0.006564103,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.016410258,0.03938462,0.04266667,0.029538464,0.016410258,0.016410258,0.016410258,0.006564103,0.055794876,0.08205129,0.08205129,0.11158975,0.13456412,0.09189744,0.068923086,0.07876924,0.08205129,0.08861539,0.07548718,0.0951795,0.14112821,0.15097436,0.15425642,0.13128206,0.098461546,0.072205134,0.07548718,0.10502565,0.08861539,0.101743594,0.190359,0.3708718,0.4397949,0.40697438,0.42338464,0.5284103,0.6268718,0.76800007,0.8467693,0.77128214,0.5677949,0.40369233,0.44307697,0.636718,0.80738467,0.92553854,1.1093334,1.5458462,2.3958976,2.6354873,2.1169233,1.5688206,1.211077,0.6695385,0.26912823,0.098461546,0.026256412,0.016410258,0.016410258,0.01969231,0.013128206,0.006564103,0.0,0.0,0.0032820515,0.009846155,0.029538464,0.0951795,0.14769232,0.15425642,0.12471796,0.118153855,0.13128206,0.098461546,0.059076928,0.026256412,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.02297436,0.01969231,0.009846155,0.009846155,0.016410258,0.013128206,0.016410258,0.029538464,0.04594872,0.03938462,0.04594872,0.052512825,0.055794876,0.055794876,0.098461546,0.10502565,0.08861539,0.068923086,0.068923086,0.068923086,0.08861539,0.09189744,0.07548718,0.059076928,0.08861539,0.15425642,0.24287182,0.34789747,0.47261542,0.88943595,1.3095386,1.4572309,1.273436,0.8992821,0.5973334,0.5021539,0.571077,0.77128214,1.086359,1.595077,1.8116925,1.9331284,1.9626669,1.7165129,2.356513,3.9712822,5.9569235,6.9021544,4.598154,4.1485133,4.568616,5.074052,5.0871797,4.2338467,4.315898,4.3684106,4.263385,4.2174363,4.7983594,5.208616,6.0652313,7.2336416,8.356103,8.881231,8.539898,9.07159,10.587898,12.314258,12.563693,10.699488,9.094564,8.3134365,7.683283,5.3037953,4.2601027,4.135385,4.713026,5.3169236,4.8082056,3.8662567,3.6824617,4.969026,7.259898,8.897642,8.982975,9.409642,10.279386,11.244308,11.500309,12.1698475,13.879796,16.873028,20.378258,22.59036,25.294771,27.549541,29.108515,29.410463,27.56595,22.898874,17.483488,13.453129,11.162257,9.199591,6.9021544,4.516103,2.8521028,1.9889232,1.2406155,0.6301539,0.22646156,0.04594872,0.029538464,0.036102567,0.04594872,0.04594872,0.036102567,0.01969231,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.006564103,0.029538464,0.07548718,0.14112821,0.2297436,0.29538465,0.41025645,0.5907693,0.7778462,0.86646163,0.8795898,0.8763078,0.86646163,0.8008206,0.636718,0.39712822,0.25271797,0.27569234,0.43323082,0.64000005,0.73517954,0.8008206,0.892718,1.0535386,1.3161026,1.4178462,2.0939488,3.5314875,5.35959,6.6428723,5.3037953,4.2896414,4.5062566,4.7917953,4.2502565,6.1407185,8.129642,8.864821,7.965539,5.9963083,6.665847,7.79159,7.90318,6.242462,6.2720003,6.51159,5.907693,4.578462,3.7874875,3.2951798,2.9833848,2.8816411,2.8389745,2.5337439,2.284308,2.1333334,1.9790771,1.7788719,1.5130258,1.4867693,1.5589745,1.6738462,1.7755898,1.8182565,2.0217438,2.103795,2.03159,1.8182565,1.5392822,1.276718,0.9878975,0.7450257,0.65969235,0.86317956,1.2012309,1.3981539,1.5130258,1.719795,2.28759,2.8192823,2.789744,2.3171284,1.7066668,1.4441026,1.6082052,1.972513,2.3926156,2.7733335,3.045744,3.5216413,3.8662567,3.9811285,3.8038976,3.3247182,2.733949,2.3466668,2.5107694,3.2098465,4.056616,3.9253337,3.3509746,2.7536411,2.4418464,2.6223593,6.8496413,7.499488,8.457847,9.229129,10.240001,12.849232,13.915898,12.941129,10.568206,8.362667,8.789334,10.105436,11.260718,11.661129,11.017847,9.373539,7.643898,6.931693,7.2992826,8.408616,9.524513,9.921641,9.035488,7.351795,5.402257,3.751385,2.6847181,2.1464617,1.9364104,1.9364104,2.0808206,2.422154,3.0720003,4.466872,6.091488,6.4656415,5.924103,4.824616,3.2853336,1.7362052,0.90912825,0.8205129,0.75487185,1.0765129,1.7132308,2.1792822,2.4024618,1.8970258,1.3554872,1.0633847,0.9124103,0.86974365,0.88943595,1.0502565,1.3193847,1.5458462,1.6410258,1.1323078,0.7220513,0.6268718,0.5874872,0.49230772,0.4660513,0.446359,0.41682056,0.38728207,0.32820517,0.318359,0.3052308,0.27241027,0.24287182,0.380718,0.7220513,1.1388719,1.5064616,1.7165129,1.467077,1.2373334,1.0568206,0.9616411,0.9911796,1.1552821,1.1520001,1.1191796,1.1585642,1.332513,1.3883078,1.5786668,2.0611284,2.9735386,4.4340515,5.802667,6.672411,7.00718,6.058667,2.3794873,1.8543591,1.5655385,1.5425643,1.5491283,1.083077,0.6432821,0.34133336,0.17066668,0.101743594,0.06564103,0.07548718,0.072205134,0.06564103,0.055794876,0.06564103,0.13456412,0.21661541,0.33805132,0.44307697,0.39384618,0.36430773,0.636718,1.4769232,2.2777438,1.5524104,1.3029745,1.3357949,1.3193847,1.0765129,0.6170257,0.5316923,0.6695385,0.60389745,0.318359,0.21661541,0.17066668,0.14769232,0.16410258,0.21989745,0.3117949,0.32820517,0.32820517,0.49887183,0.7581539,0.7778462,0.64000005,0.512,0.44307697,0.4004103,0.27897438,0.20348719,0.21333335,0.23958977,0.26912823,0.34789747,0.41025645,0.38728207,0.28882053,0.16082053,0.07876924,0.07548718,0.055794876,0.04266667,0.049230773,0.06564103,0.072205134,0.068923086,0.06235898,0.055794876,0.072205134,0.118153855,0.12471796,0.13456412,0.16082053,0.20020515,0.27241027,0.37415388,0.47589746,0.5513847,0.5874872,0.5349744,0.446359,0.43323082,0.5284103,0.69579494,0.8041026,0.761436,0.9714873,1.5753847,2.4615386,2.5304618,2.422154,2.284308,2.2153847,2.2547693,2.0644104,2.5337439,2.8980515,2.6157951,1.3915899,1.214359,1.0765129,0.9944616,0.97805136,1.017436,0.90584624,0.8336411,0.8533334,0.90584624,0.81066674,1.020718,0.95835906,0.8369231,0.8467693,1.1618463,1.1749744,1.3653334,1.6114873,1.6443079,1.0469744,1.2996924,1.6836925,2.048,2.1464617,1.6443079,2.4385643,3.0194874,3.2000003,3.0326157,2.8127182,3.1081028,3.4330258,3.4756925,3.2820516,3.242667,2.6256413,2.3269746,2.8553848,3.5478978,2.5435898,2.0742567,1.9790771,2.3040001,2.5632823,1.7394873,1.5360001,1.8806155,1.9626669,1.6705642,1.591795,1.3817437,1.0371283,0.81066674,0.7450257,0.6662565,0.8205129,1.2471796,1.2438976,0.82379496,0.7056411,0.7844103,0.702359,0.79097444,1.0601027,1.2012309,1.0699488,0.8598975,0.7515898,0.75487185,0.7187693,0.32820517,0.3446154,0.24943592,0.0,0.0,0.18379489,0.15425642,0.20020515,0.36758977,0.47261542,0.4594872,0.446359,0.5481026,0.7581539,0.96492314,0.97805136,0.85005134,0.761436,0.76800007,0.80738467,0.77456415,0.6629744,0.49887183,0.34789747,0.30194873,0.44307697,0.34133336,0.18379489,0.09189744,0.12143591,0.37743592,0.3249231,0.18707694,0.09189744,0.07876924,0.03938462,0.01969231,0.016410258,0.029538464,0.049230773,0.013128206,0.013128206,0.04594872,0.098461546,0.16738462,0.072205134,0.026256412,0.006564103,0.0,0.0,0.009846155,0.013128206,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01969231,0.08205129,0.18051283,0.10502565,0.02297436,0.0,0.0,0.0,0.0,0.009846155,0.02297436,0.013128206,0.016410258,0.009846155,0.006564103,0.006564103,0.0032820515,0.0032820515,0.0032820515,0.0032820515,0.0,0.0,0.0,0.006564103,0.016410258,0.026256412,0.029538464,0.06564103,0.07548718,0.068923086,0.055794876,0.032820515,0.032820515,0.14112821,0.20348719,0.18051283,0.12143591,0.190359,0.15425642,0.108307704,0.08533334,0.06564103,0.098461546,0.0951795,0.08205129,0.07876924,0.08205129,0.12143591,0.13784617,0.13456412,0.12471796,0.118153855,0.15097436,0.13128206,0.14112821,0.2297436,0.42338464,0.42994875,0.4660513,0.5349744,0.5874872,0.52512825,0.58092314,0.67610264,0.7253334,0.6892308,0.55794877,0.58420515,0.7581539,1.0010257,1.1618463,1.0272821,0.73517954,0.77128214,0.8533334,0.83035904,0.67610264,0.5481026,0.38728207,0.23630771,0.118153855,0.055794876,0.04594872,0.036102567,0.029538464,0.01969231,0.016410258,0.0032820515,0.0032820515,0.009846155,0.026256412,0.072205134,0.15425642,0.21333335,0.21333335,0.16410258,0.14441027,0.12143591,0.07548718,0.032820515,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.026256412,0.03938462,0.026256412,0.0,0.0,0.0,0.0,0.006564103,0.01969231,0.03938462,0.04594872,0.055794876,0.059076928,0.049230773,0.04266667,0.072205134,0.0951795,0.0951795,0.07548718,0.068923086,0.07548718,0.08205129,0.07548718,0.068923086,0.09189744,0.14441027,0.20348719,0.26584616,0.35774362,0.5152821,0.9878975,1.6278975,1.8445129,1.5163078,0.99774367,0.64000005,0.49887183,0.571077,0.8566154,1.3817437,1.972513,1.9232821,1.7033848,1.595077,1.6968206,2.5993848,3.3575387,4.069744,4.604718,4.585026,4.325744,5.208616,6.2720003,6.698667,5.8223596,4.97559,4.1550775,3.6594875,3.5347695,3.5774362,4.309334,5.6451287,7.0465646,8.1066675,8.553026,7.131898,6.426257,6.2162056,6.3868723,6.8988724,6.6625648,6.413129,6.5280004,6.701949,5.9503593,5.4974365,5.5893335,5.481026,5.146257,5.284103,4.1156926,3.3345644,3.8596926,5.7501545,8.198565,8.349539,8.789334,9.458873,9.757539,8.562873,7.955693,9.396514,13.272616,18.33354,21.697643,25.45231,28.425848,30.080002,29.833849,27.076925,21.625437,16.416822,12.507898,10.095591,8.500513,6.5312824,4.450462,2.8324106,1.8313848,1.1782565,0.63343596,0.21661541,0.036102567,0.055794876,0.098461546,0.13128206,0.12471796,0.08861539,0.03938462,0.02297436,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.032820515,0.06564103,0.15425642,0.28225642,0.40697438,0.508718,0.5973334,0.6104616,0.6268718,0.65641034,0.65641034,0.5513847,0.36102566,0.20348719,0.11158975,0.07548718,0.06564103,0.0951795,0.118153855,0.15425642,0.23958977,0.42338464,0.64000005,0.761436,1.2373334,2.3072822,3.9811285,5.7764106,5.3858466,6.009436,7.9819493,8.789334,6.994052,6.229334,5.395693,4.194462,3.131077,4.204308,5.35959,6.0783596,6.0783596,5.3234878,6.7282057,8.556309,8.87795,7.6077952,6.488616,4.7950773,3.4166157,2.7634873,2.7142565,2.612513,2.1497438,1.913436,1.8313848,1.8182565,1.7985642,1.7690258,1.7788719,1.7526156,1.6607181,1.5097437,1.5721027,1.6443079,1.6344616,1.529436,1.4145643,1.3423591,1.1224617,0.8402052,0.61374366,0.574359,0.764718,1.0732309,1.3915899,1.7099489,2.1136413,2.5829747,2.5337439,2.1858463,1.7624617,1.4933335,1.522872,1.7394873,2.044718,2.4746668,3.1934361,3.9975388,4.4012313,4.4373336,4.2929235,4.325744,3.8564105,3.3345644,3.308308,3.7940516,4.2830772,4.2207184,3.7251284,3.2295387,3.0194874,3.2361028,8.421744,7.2861543,8.743385,11.32636,13.640206,14.372104,14.106257,12.977232,11.204924,9.193027,7.506052,7.88677,8.162462,8.12636,7.765334,7.2631803,7.250052,6.6625648,5.5696416,4.384821,3.8596926,3.4592824,3.43959,4.056616,4.923077,5.0215387,3.751385,2.865231,2.359795,2.228513,2.4713848,2.861949,3.6102567,4.7261543,5.796103,5.9667697,5.8453336,5.0543594,3.442872,1.6311796,1.0075898,1.0436924,1.1093334,1.6311796,2.5206156,3.1442053,2.9965131,2.4943593,1.8510771,1.2898463,1.020718,0.99774367,1.2209232,2.228513,3.7940516,4.9296412,4.57518,2.3335385,0.764718,0.5481026,0.48902568,0.46276927,0.47589746,0.45620516,0.4004103,0.3511795,0.30194873,0.28225642,0.26256412,0.28225642,0.4266667,0.7187693,1.1585642,1.5983591,1.8970258,1.9232821,1.6049232,1.3883078,1.3161026,1.3817437,1.5425643,1.723077,1.8051283,1.9331284,2.162872,2.4549747,2.674872,2.8882053,3.373949,4.240411,5.3858466,6.7544622,6.554257,5.4383593,3.7710772,1.6475899,1.2570257,1.332513,1.4178462,1.2898463,0.9616411,0.5218462,0.28225642,0.16738462,0.11158975,0.07548718,0.17394873,0.18051283,0.13784617,0.10502565,0.15097436,0.5316923,0.77128214,0.8467693,0.8467693,0.9911796,0.7975385,0.67282057,0.67938465,0.7975385,0.9321026,0.9911796,1.0896411,1.1946667,1.2274873,1.0666667,0.8369231,0.5940513,0.42994875,0.36430773,0.3511795,0.26584616,0.190359,0.17066668,0.21333335,0.27569234,0.21333335,0.21661541,0.5218462,1.0601027,1.4506668,1.3883078,1.0633847,0.78769237,0.62030774,0.3511795,0.26584616,0.35446155,0.46276927,0.48246157,0.33476925,0.16410258,0.07548718,0.04594872,0.04266667,0.029538464,0.01969231,0.02297436,0.036102567,0.052512825,0.07548718,0.11158975,0.14112821,0.14769232,0.14769232,0.18379489,0.256,0.18379489,0.15097436,0.21333335,0.27569234,0.2855385,0.30851284,0.3511795,0.40697438,0.44307697,0.41682056,0.47589746,0.6235898,0.84348726,1.0994873,1.2931283,1.2242053,1.0962052,1.0699488,1.2668719,2.2416413,2.6978464,2.917744,3.0982566,3.3411283,3.95159,4.096,3.5872824,2.356513,0.4266667,0.46276927,0.51856416,0.58092314,0.636718,0.6859488,0.9682052,0.9911796,0.74830776,0.39712822,0.27569234,0.24943592,0.36430773,0.57764107,0.7975385,0.86974365,0.73517954,0.53825647,0.256,0.14441027,0.7187693,0.8041026,0.82379496,0.8369231,0.827077,0.7187693,0.48574364,0.36430773,0.43651286,0.60389745,0.58092314,0.7384616,0.88943595,0.9124103,0.7778462,0.5349744,0.42338464,0.50543594,0.892718,1.4080001,1.6016412,1.3718976,1.1552821,1.6082052,2.3368206,1.9232821,1.6311796,1.7493335,1.6278975,1.2274873,1.1290257,1.1913847,1.214359,1.1848207,1.0929232,0.94523084,0.8369231,1.0272821,0.9485129,0.7056411,1.083077,1.7296412,1.4539489,1.014154,0.7253334,0.45620516,0.09189744,0.2100513,0.636718,1.1585642,1.5261539,1.2340513,0.69251287,0.2297436,0.0,0.0,0.18379489,0.14769232,0.07876924,0.068923086,0.108307704,0.27897438,0.34789747,0.39056414,0.45292312,0.5481026,0.574359,0.65312827,0.71548724,0.7122052,0.6268718,0.6498462,0.53825647,0.43323082,0.4004103,0.4135385,0.43651286,0.37743592,0.26912823,0.14769232,0.06235898,0.02297436,0.016410258,0.026256412,0.055794876,0.09189744,0.029538464,0.006564103,0.0,0.0,0.0,0.013128206,0.032820515,0.068923086,0.0951795,0.04594872,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.02297436,0.01969231,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.0951795,0.4135385,0.8992821,0.5284103,0.118153855,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02297436,0.029538464,0.029538464,0.026256412,0.016410258,0.016410258,0.016410258,0.009846155,0.0,0.0,0.0,0.0,0.0,0.006564103,0.029538464,0.1148718,0.17394873,0.21661541,0.21661541,0.108307704,0.108307704,0.19692309,0.27897438,0.26912823,0.12143591,0.17066668,0.17394873,0.18707694,0.19692309,0.13784617,0.11158975,0.08861539,0.07548718,0.08205129,0.108307704,0.108307704,0.108307704,0.0951795,0.08205129,0.108307704,0.118153855,0.13128206,0.15097436,0.21661541,0.4135385,0.49887183,0.53825647,0.65969235,0.79425645,0.67282057,0.56123084,0.5349744,0.62030774,0.79097444,0.9616411,0.88943595,0.7220513,0.6695385,0.73517954,0.74830776,0.69907695,0.67610264,0.67610264,0.65312827,0.51856416,0.3117949,0.16738462,0.08861539,0.06564103,0.09189744,0.09189744,0.06564103,0.04594872,0.03938462,0.016410258,0.0032820515,0.01969231,0.02297436,0.02297436,0.06235898,0.12143591,0.19364104,0.25928208,0.31507695,0.3511795,0.33805132,0.19692309,0.068923086,0.013128206,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.07548718,0.06564103,0.026256412,0.0,0.0,0.0,0.0,0.006564103,0.016410258,0.016410258,0.03938462,0.06564103,0.07548718,0.06564103,0.029538464,0.029538464,0.03938462,0.059076928,0.08205129,0.108307704,0.13128206,0.09189744,0.06564103,0.09189744,0.15097436,0.27569234,0.37743592,0.4266667,0.44307697,0.5021539,0.9189744,1.3883078,1.7362052,1.7558975,1.204513,0.827077,0.6695385,0.7778462,1.0404103,1.1749744,1.6738462,1.9561027,1.8084104,1.5491283,2.0151796,2.868513,3.6496413,3.9975388,3.9844105,4.1189747,5.07077,6.6822567,7.5552826,7.030154,5.1889234,3.4921029,2.5074873,2.1792822,2.3696413,2.868513,3.6004105,5.3398976,6.87918,7.4797955,6.882462,5.149539,4.2305646,3.7284105,3.6791797,4.532513,4.568616,4.027077,4.352,5.402257,5.4613338,4.6080003,3.6332312,3.1409233,3.3542566,4.135385,4.1583595,3.2229745,3.5511796,5.4908724,7.4929237,8.579283,9.005949,9.242257,9.160206,8.024616,6.695385,7.4436927,11.270565,17.352207,23.04,23.102362,25.094566,27.431387,28.383183,26.0759,21.316925,16.794258,13.010053,10.282667,8.743385,6.764308,4.5489235,2.6322052,1.3489232,0.82379496,0.39712822,0.12471796,0.026256412,0.06235898,0.12143591,0.19692309,0.21333335,0.17066668,0.0951795,0.04594872,0.02297436,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.026256412,0.12143591,0.23302566,0.29210258,0.24287182,0.3052308,0.42994875,0.62030774,0.761436,0.6268718,0.3446154,0.14769232,0.04266667,0.01969231,0.029538464,0.029538464,0.029538464,0.04266667,0.068923086,0.108307704,0.16738462,0.24615386,0.33805132,0.44307697,0.56451285,0.6498462,1.4966155,2.8192823,4.6276927,7.200821,8.533334,7.683283,5.346462,2.9472823,2.6551797,5.1331286,8.041026,10.043077,10.328616,8.621949,8.060719,7.7259493,6.9087186,6.048821,6.744616,5.7435904,3.5052311,2.1530259,2.0873847,2.0151796,1.7591796,1.6016412,1.6705642,1.9429746,2.2744617,2.3236926,2.2350771,1.9593848,1.5721027,1.2668719,1.2307693,1.2931283,1.3128207,1.2570257,1.2209232,1.3423591,1.1618463,0.8566154,0.5973334,0.5481026,0.6235898,0.99774367,1.4933335,1.9692309,2.3335385,2.674872,2.5435898,2.1464617,1.6869745,1.3587693,1.4572309,1.910154,2.6354873,3.436308,3.9975388,4.069744,3.9351797,3.7382567,3.629949,3.7382567,3.7874875,3.8728209,3.9351797,4.0008206,4.197744,4.4767184,4.33559,3.9581542,3.636513,3.7842054,5.664821,6.3343596,6.8004107,8.536616,11.260718,12.921437,12.914873,11.588924,9.7214365,7.8834877,6.432821,5.835488,4.8640003,4.3749747,4.4964104,4.637539,4.266667,3.3805132,2.5042052,1.9593848,1.8838975,1.8904617,3.0424619,4.7917953,6.5411286,7.643898,8.172308,6.806975,5.405539,4.844308,5.0116925,4.2994876,3.9056413,4.4406157,6.2490263,9.409642,10.262975,8.421744,5.3103595,2.4024618,1.214359,1.7493335,2.7208207,3.948308,5.152821,5.9503593,4.585026,3.4100516,2.537026,2.0841026,2.156308,2.1924105,3.3312824,5.7107697,8.03118,7.565129,4.827898,2.1169233,0.65969235,0.512,0.5481026,0.50543594,0.49887183,0.58092314,0.6662565,0.508718,0.4135385,0.3708718,0.380718,0.4955898,0.8172308,1.3062565,1.8838975,2.2744617,2.353231,2.1431797,1.8642052,1.7165129,1.6869745,1.7493335,1.8576412,2.100513,2.4451284,2.7306669,2.8882053,2.9571285,3.0194874,3.3444104,3.8695388,4.594872,5.605744,6.5936418,5.5072823,4.0533338,2.9078977,1.719795,1.4080001,1.4309745,1.3357949,0.9878975,0.571077,0.30851284,0.26584616,0.25928208,0.190359,0.07548718,0.055794876,0.13456412,0.2100513,0.27569234,0.43323082,1.4867693,1.3456411,0.77456415,0.3249231,0.3446154,0.5316923,0.6071795,0.7056411,0.90912825,1.2471796,1.3489232,1.3620514,1.2800001,1.0765129,0.71548724,0.6104616,0.508718,0.42338464,0.33805132,0.2297436,0.28882053,0.31507695,0.27241027,0.21333335,0.27569234,0.3314872,0.37743592,0.46276927,0.7220513,1.3751796,1.6475899,1.6836925,1.5819489,1.3850257,1.0469744,0.98133343,1.0371283,0.9878975,0.7450257,0.38400003,0.15425642,0.08861539,0.07876924,0.06564103,0.055794876,0.052512825,0.052512825,0.052512825,0.052512825,0.07548718,0.09189744,0.1148718,0.16738462,0.2231795,0.21989745,0.14769232,0.118153855,0.12143591,0.14441027,0.17723078,0.21989745,0.28225642,0.34133336,0.37415388,0.380718,0.33805132,0.4201026,0.60389745,0.86974365,1.1848207,1.4375386,2.0644104,2.2613335,1.8379488,1.1946667,1.7493335,1.8642052,1.9823592,2.3072822,2.806154,2.6912823,2.6978464,2.4418464,1.7132308,0.48902568,1.0896411,1.1257436,0.9485129,0.8533334,1.0765129,0.9682052,1.0043077,0.97805136,0.8008206,0.48246157,0.5940513,0.6695385,0.65641034,0.512,0.17394873,0.30194873,0.4266667,0.5677949,0.67938465,0.65641034,0.4594872,0.29210258,0.19692309,0.16410258,0.14441027,0.098461546,0.072205134,0.08861539,0.12143591,0.1148718,0.14769232,0.39712822,0.69579494,0.9189744,0.99774367,0.8008206,0.54482055,0.7187693,1.1520001,1.0043077,0.9878975,1.3751796,1.7887181,1.9954873,1.9232821,1.7066668,1.4736412,1.4834872,1.6278975,1.4211283,1.1126155,1.0962052,1.1388719,1.1093334,0.98133343,0.88287187,1.1585642,1.4342566,1.5425643,1.5097437,1.2209232,0.9124103,0.51856416,0.14441027,0.09189744,0.19364104,0.34133336,0.49230772,0.5349744,0.3052308,0.65641034,0.512,0.28882053,0.20348719,0.28225642,0.56123084,0.512,0.36102566,0.26584616,0.30194873,0.7844103,0.90584624,0.83035904,0.7089231,0.65969235,0.7417436,0.8205129,0.8336411,0.71548724,0.40697438,0.42994875,0.4135385,0.39056414,0.40697438,0.49887183,0.5415385,0.4594872,0.2986667,0.14769232,0.108307704,0.101743594,0.07876924,0.04266667,0.013128206,0.029538464,0.01969231,0.006564103,0.0,0.013128206,0.06235898,0.072205134,0.06564103,0.049230773,0.029538464,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02297436,0.0951795,0.19364104,0.12471796,0.04266667,0.013128206,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.016410258,0.029538464,0.026256412,0.016410258,0.016410258,0.009846155,0.0,0.0,0.0,0.0,0.0,0.009846155,0.04266667,0.098461546,0.12143591,0.14769232,0.17723078,0.15425642,0.118153855,0.08205129,0.068923086,0.072205134,0.072205134,0.13128206,0.20348719,0.26584616,0.27569234,0.18707694,0.12143591,0.14112821,0.190359,0.23958977,0.25271797,0.21333335,0.14441027,0.108307704,0.118153855,0.14441027,0.14441027,0.14112821,0.2855385,0.574359,0.8402052,0.88615394,0.7975385,0.76800007,0.84348726,0.9288206,1.0633847,1.0075898,0.88943595,0.77456415,0.67938465,0.5973334,0.6498462,0.83035904,1.0633847,1.211077,0.85005134,0.62030774,0.50543594,0.47917953,0.48246157,0.3249231,0.20020515,0.12471796,0.09189744,0.06564103,0.055794876,0.049230773,0.03938462,0.032820515,0.026256412,0.026256412,0.01969231,0.02297436,0.036102567,0.072205134,0.10502565,0.118153855,0.11158975,0.098461546,0.108307704,0.2231795,0.24615386,0.16410258,0.04594872,0.02297436,0.013128206,0.0032820515,0.0,0.0032820515,0.016410258,0.016410258,0.013128206,0.006564103,0.0,0.0,0.0,0.0,0.009846155,0.026256412,0.026256412,0.04266667,0.08533334,0.12143591,0.12143591,0.055794876,0.026256412,0.026256412,0.03938462,0.08205129,0.20348719,0.28882053,0.18051283,0.10502565,0.13784617,0.23958977,0.3708718,0.50543594,0.6071795,0.67282057,0.7220513,0.86646163,1.1126155,1.270154,1.2307693,0.9747693,0.5349744,0.38400003,0.43651286,0.6432821,0.9911796,2.0184617,2.169436,1.910154,1.6508719,1.7329233,2.3433847,2.6617439,2.9078977,3.308308,4.096,5.586052,6.048821,5.7698464,4.893539,3.442872,2.7798977,2.6289232,2.7766156,2.9669745,2.8816411,2.9702566,3.5216413,4.1846156,4.6080003,4.4406157,3.8596926,3.6890259,3.8038976,3.9909747,3.9581542,3.4855387,3.1343591,3.2098465,3.7743592,4.6572313,4.6244106,4.197744,3.6496413,3.3378465,3.7185643,4.056616,4.2896414,4.6080003,5.0838976,5.661539,6.678975,8.165744,9.340718,9.508103,8.050873,7.6176414,8.743385,11.296822,15.14995,20.184616,24.97313,29.200413,31.93436,32.141132,28.70154,23.05313,18.372925,14.749539,11.98277,9.586872,6.925129,4.4734364,2.550154,1.276718,0.5546667,0.3511795,0.21661541,0.12143591,0.06235898,0.08533334,0.13784617,0.23958977,0.25271797,0.15425642,0.04594872,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.03938462,0.08205129,0.11158975,0.12143591,0.12471796,0.13128206,0.15097436,0.16082053,0.12471796,0.07876924,0.04266667,0.01969231,0.016410258,0.01969231,0.029538464,0.03938462,0.049230773,0.06235898,0.068923086,0.08205129,0.10502565,0.15425642,0.24287182,0.39384618,0.6268718,1.5819489,3.4034874,5.83877,8.228104,8.746667,8.04759,6.49518,4.4865646,2.4352822,2.1103592,2.428718,2.7798977,2.7766156,2.2482052,2.1464617,2.3040001,2.6518977,2.9965131,3.0096412,2.3991797,1.6672822,1.3423591,1.4736412,1.6344616,1.8379488,2.0676925,2.4188719,2.793026,2.9078977,2.7241027,2.487795,2.162872,1.7755898,1.401436,1.1782565,1.1158975,1.0502565,0.9419488,0.86646163,0.9288206,0.90256417,0.827077,0.7515898,0.7318975,0.8533334,1.404718,2.044718,2.5829747,2.9702566,3.0391798,2.8947694,2.6420515,2.349949,2.028308,1.7952822,2.0939488,2.6847181,3.3411283,3.8629746,4.201026,4.1583595,3.9712822,3.8334363,3.8859491,4.1091285,4.0336413,3.7973337,3.5971284,3.69559,4.1911798,4.4406157,4.2535386,3.5872824,2.550154,7.463385,8.3823595,8.546462,8.753231,9.019077,8.612103,8.89436,8.411898,7.0859494,5.546667,5.1298466,4.3684106,3.4297438,3.1376412,3.4002054,3.2131286,3.0293336,3.18359,4.516103,6.157129,5.5269747,4.785231,5.1364107,6.2720003,7.4075904,7.2861543,6.665847,5.3169236,4.460308,4.2371287,3.7218463,2.4943593,2.28759,4.164923,7.5487185,10.223591,11.657847,9.819899,6.76759,4.0500517,2.6683078,3.2164104,4.338872,5.156103,5.3136415,4.9788723,3.7448208,3.511795,3.318154,2.8160002,2.2580514,2.4385643,5.037949,7.9491286,9.366975,7.77518,5.146257,2.665026,1.0043077,0.36758977,0.46276927,0.42338464,0.50543594,0.6826667,0.827077,0.7220513,0.77456415,0.7844103,0.81066674,0.99774367,1.585231,2.041436,2.3663592,2.4484105,2.28759,2.0053334,1.8084104,1.7362052,1.782154,1.9364104,2.166154,2.5271797,2.8980515,3.0851285,3.0884104,3.1015387,3.3214362,3.7874875,4.266667,4.6933336,5.149539,5.2414365,4.1813335,3.2295387,2.7175386,2.0512822,1.6180514,1.404718,1.1224617,0.7187693,0.39056414,0.2231795,0.18379489,0.25928208,0.35446155,0.2855385,0.12143591,0.3708718,0.6695385,0.8533334,0.9714873,1.3489232,1.3095386,1.0962052,0.90256417,0.86974365,0.86646163,0.8533334,0.88943595,1.0272821,1.2996924,1.6377437,1.3554872,0.98133343,0.80738467,0.88287187,0.9485129,0.74830776,0.5021539,0.37415388,0.48246157,0.380718,0.39056414,0.41682056,0.42338464,0.40369233,0.4135385,0.41682056,0.40369233,0.45292312,0.7253334,1.1618463,1.467077,1.6049232,1.5458462,1.2570257,1.2242053,1.3357949,1.4867693,1.3817437,0.54482055,0.190359,0.101743594,0.10502565,0.10502565,0.07876924,0.06564103,0.055794876,0.052512825,0.059076928,0.07548718,0.11158975,0.16082053,0.19364104,0.20348719,0.19364104,0.14769232,0.15097436,0.14112821,0.1148718,0.12471796,0.17394873,0.26256412,0.30851284,0.30194873,0.30194873,0.318359,0.380718,0.5021539,0.6662565,0.8205129,0.8763078,1.3161026,1.6311796,1.6410258,1.4966155,1.7788719,1.7952822,1.782154,1.847795,1.9561027,1.5819489,1.4211283,1.339077,1.2668719,1.1979488,1.9889232,2.0939488,1.7920002,1.2931283,0.761436,0.761436,0.86317956,0.94523084,0.892718,0.5973334,0.8533334,0.8795898,0.76800007,0.7417436,1.1454359,1.2373334,1.1257436,0.8795898,0.6071795,0.4660513,0.37415388,0.27569234,0.13456412,0.0,0.0,0.0,0.059076928,0.14441027,0.16738462,0.0,0.0,0.15425642,0.32820517,0.46276927,0.5546667,0.60061544,0.67938465,0.6170257,0.43323082,0.34133336,0.35774362,0.9288206,1.3587693,1.3817437,1.1913847,0.77456415,0.88615394,1.1191796,1.1913847,0.9353847,0.50543594,0.7778462,1.1716924,1.4309745,1.6311796,1.8510771,1.7788719,1.595077,1.3620514,1.024,0.58420515,0.34789747,0.15753847,0.0,0.0,0.08861539,0.15097436,0.18051283,0.28225642,0.6498462,0.48902568,0.6301539,0.892718,1.0371283,0.79097444,0.69251287,0.5021539,0.33476925,0.28225642,0.4135385,0.8369231,0.93866676,0.8730257,0.83035904,1.0436924,1.0666667,1.0075898,0.8795898,0.7220513,0.5973334,0.61374366,0.67282057,0.827077,1.0043077,1.014154,0.7778462,0.42338464,0.17394873,0.098461546,0.13128206,0.14441027,0.098461546,0.055794876,0.04266667,0.068923086,0.06235898,0.036102567,0.009846155,0.006564103,0.03938462,0.04594872,0.032820515,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.006564103,0.016410258,0.02297436,0.02297436,0.016410258,0.009846155,0.0032820515,0.0032820515,0.009846155,0.009846155,0.009846155,0.009846155,0.016410258,0.032820515,0.03938462,0.04266667,0.026256412,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.01969231,0.03938462,0.049230773,0.06235898,0.13456412,0.36102566,1.2635899,1.5425643,1.5064616,1.3292309,1.0502565,0.69907695,0.47261542,0.3511795,0.32164106,0.36430773,0.44307697,0.43323082,0.3708718,0.30194873,0.26256412,0.27897438,0.23302566,0.17394873,0.15753847,0.22646156,0.23302566,0.22646156,0.3052308,0.49887183,0.77128214,0.8172308,0.7318975,0.6071795,0.51856416,0.5349744,0.6695385,0.6892308,0.58092314,0.41682056,0.35446155,0.4660513,0.7056411,0.9124103,1.0043077,0.9616411,0.6465641,0.41025645,0.30194873,0.30851284,0.35446155,0.28882053,0.17394873,0.118153855,0.12471796,0.08861539,0.04594872,0.036102567,0.03938462,0.04266667,0.049230773,0.06235898,0.059076928,0.055794876,0.06235898,0.08533334,0.108307704,0.101743594,0.072205134,0.04266667,0.026256412,0.08533334,0.118153855,0.101743594,0.06564103,0.08533334,0.04266667,0.02297436,0.029538464,0.049230773,0.068923086,0.036102567,0.016410258,0.006564103,0.0032820515,0.009846155,0.009846155,0.013128206,0.02297436,0.026256412,0.013128206,0.032820515,0.06564103,0.0951795,0.098461546,0.068923086,0.049230773,0.06235898,0.11158975,0.23302566,0.5021539,0.446359,0.27569234,0.16738462,0.190359,0.31507695,0.47917953,0.6235898,0.6892308,0.6662565,0.61374366,0.636718,0.761436,0.92553854,0.9944616,0.761436,0.41025645,0.27569234,0.49230772,0.90256417,1.0666667,1.6968206,2.356513,2.3302567,1.8904617,2.294154,3.0424619,2.484513,2.2547693,2.9571285,4.1714873,5.7009234,5.8092313,4.9952826,3.7185643,2.3926156,2.0053334,2.2547693,2.5600002,2.6354873,2.4910772,2.6584618,2.7602053,3.0358977,3.4822567,3.8662567,3.9089234,3.9975388,4.1878977,4.4045134,4.4274874,3.6693337,3.2361028,3.0358977,3.045744,3.3214362,3.7251284,4.1124105,4.3716927,4.4406157,4.3027697,4.886975,5.2053337,5.1364107,4.772103,4.4438977,4.630975,5.658257,7.026872,7.899898,7.0859494,6.987488,7.686565,9.091283,11.933539,17.785437,25.11754,31.422361,34.92103,34.648617,30.457438,24.746668,19.666052,16.25272,13.99795,10.857026,7.565129,4.7228723,2.6617439,1.4966155,1.1388719,1.0568206,0.5218462,0.14112821,0.07876924,0.07548718,0.0951795,0.15097436,0.14769232,0.08205129,0.01969231,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.009846155,0.0032820515,0.006564103,0.016410258,0.026256412,0.036102567,0.03938462,0.03938462,0.032820515,0.02297436,0.009846155,0.013128206,0.016410258,0.01969231,0.029538464,0.04266667,0.03938462,0.04266667,0.052512825,0.06235898,0.06235898,0.052512825,0.06235898,0.07876924,0.118153855,0.19692309,0.34789747,0.9485129,2.1169233,3.5905645,4.7491283,5.467898,5.914257,6.1078978,5.6418467,3.6791797,2.1497438,1.0502565,0.5546667,0.512,0.46276927,0.51856416,0.6892308,1.020718,1.3522053,1.2865642,1.1257436,1.1158975,1.2603078,1.5163078,1.7788719,2.0611284,2.3105643,2.5928206,2.8389745,2.8553848,2.6912823,2.612513,2.3893335,1.9954873,1.5885129,1.2832822,1.1651284,1.083077,0.98461545,0.90584624,0.88943595,1.0010257,1.1323078,1.2373334,1.3259488,1.4408206,1.9593848,2.4943593,2.8225644,2.8980515,2.5764105,2.537026,2.5862565,2.5928206,2.4713848,2.0676925,1.9626669,2.1234872,2.5173335,3.1343591,3.4789746,3.5840003,3.6004105,3.6758976,3.9318976,4.20759,4.092718,3.7087183,3.2984617,3.239385,3.6791797,4.0500517,4.1485133,3.6824617,2.2711797,8.021334,8.493949,8.625232,8.4053335,7.7981544,6.7249236,6.2884107,6.7085133,6.452513,5.35959,4.630975,3.3312824,2.6847181,2.9505644,3.8859491,4.7392826,5.677949,6.9809237,9.271795,11.411694,10.518975,8.228104,6.8266673,6.363898,6.3212314,5.6352825,4.7622566,3.9876926,3.6463592,3.508513,2.789744,1.5983591,1.5688206,3.5413337,6.4722056,7.433847,8.713847,8.310155,6.4557953,4.2994876,3.9122055,4.578462,5.47118,5.930667,5.6352825,4.588308,3.7382567,3.8695388,4.023795,3.9778464,4.2601027,5.5302567,8.310155,9.813334,9.012513,6.6527185,4.6539493,2.5632823,1.014154,0.3249231,0.48246157,0.6104616,0.6104616,0.65641034,0.764718,0.79097444,0.9156924,0.98461545,1.1355898,1.5130258,2.2547693,2.487795,2.4976413,2.3236926,2.044718,1.7920002,1.7329233,1.7657437,1.8970258,2.1070771,2.356513,2.7306669,3.0720003,3.255795,3.2984617,3.370667,3.6693337,4.07959,4.4045134,4.466872,4.1156926,3.6824617,3.0523078,2.6617439,2.484513,2.0644104,1.6213335,1.2898463,0.9288206,0.56123084,0.3708718,0.24287182,0.17394873,0.34133336,0.5907693,0.446359,0.4004103,1.0305642,1.3751796,1.273436,1.3292309,1.2438976,1.0896411,1.1257436,1.3653334,1.5721027,1.5655385,1.2242053,1.024,1.1060513,1.2865642,1.6311796,1.4178462,1.0896411,0.92553854,1.0404103,0.98461545,0.74830776,0.49887183,0.39056414,0.5316923,0.37743592,0.36430773,0.42994875,0.508718,0.512,0.4955898,0.40369233,0.29538465,0.21989745,0.21989745,0.6498462,1.0371283,1.2996924,1.3423591,1.0732309,1.0075898,1.086359,1.2865642,1.2964103,0.49887183,0.18707694,0.08861539,0.08205129,0.08205129,0.06235898,0.052512825,0.049230773,0.059076928,0.07876924,0.101743594,0.12471796,0.15097436,0.15753847,0.15097436,0.15097436,0.16410258,0.20348719,0.18051283,0.101743594,0.08861539,0.11158975,0.17723078,0.2231795,0.24615386,0.29538465,0.36102566,0.36430773,0.4201026,0.5349744,0.6301539,0.63343596,0.76800007,0.9419488,1.1323078,1.3784616,1.7493335,2.1530259,2.481231,2.6223593,2.481231,1.4342566,0.9124103,0.7581539,0.8795898,1.2537436,1.9659488,2.1267693,1.8937438,1.3883078,0.702359,0.69907695,0.8041026,0.9517949,1.014154,0.82379496,0.9156924,0.8008206,0.60389745,0.5907693,1.1454359,1.1585642,0.96492314,0.62030774,0.28225642,0.2100513,0.22646156,0.21333335,0.12143591,0.055794876,0.27569234,0.33476925,0.35446155,0.36102566,0.31507695,0.10502565,0.068923086,0.068923086,0.14769232,0.26256412,0.256,0.27241027,0.5513847,0.48902568,0.1148718,0.09189744,0.10502565,0.571077,0.90912825,0.8992821,0.65312827,0.2297436,0.57764107,0.9124103,0.9288206,0.827077,0.67938465,1.0404103,1.4342566,1.6672822,1.8346668,1.9495386,1.6443079,1.2307693,0.8566154,0.5284103,0.21661541,0.055794876,0.0,0.009846155,0.04266667,0.08205129,0.07548718,0.03938462,0.17394873,0.8763078,0.4266667,0.53825647,0.85005134,1.0272821,0.7417436,0.51856416,0.3314872,0.2231795,0.29538465,0.702359,0.9878975,1.0371283,0.92225647,0.8402052,1.0929232,1.0502565,0.90584624,0.7384616,0.6432821,0.7318975,0.81394875,0.88943595,1.0896411,1.3226668,1.276718,0.9156924,0.42338464,0.14769232,0.14112821,0.15425642,0.12471796,0.072205134,0.04266667,0.052512825,0.08861539,0.0951795,0.06564103,0.029538464,0.013128206,0.009846155,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.009846155,0.013128206,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.026256412,0.04594872,0.059076928,0.04266667,0.02297436,0.016410258,0.026256412,0.03938462,0.072205134,0.068923086,0.055794876,0.049230773,0.04594872,0.059076928,0.03938462,0.026256412,0.01969231,0.006564103,0.006564103,0.006564103,0.0032820515,0.0,0.0,0.0,0.006564103,0.009846155,0.06564103,0.29210258,1.2176411,1.5589745,1.5983591,1.522872,1.4342566,1.0765129,0.69907695,0.46933338,0.45620516,0.61374366,0.76800007,0.7220513,0.5284103,0.2986667,0.21989745,0.2855385,0.318359,0.29538465,0.26912823,0.34133336,0.39712822,0.40369233,0.4201026,0.48574364,0.61374366,0.56451285,0.49230772,0.37415388,0.23302566,0.16738462,0.22646156,0.28225642,0.24943592,0.16410258,0.18379489,0.37743592,0.62030774,0.761436,0.7417436,0.5940513,0.4266667,0.36758977,0.39056414,0.43323082,0.38400003,0.26584616,0.13456412,0.08205129,0.098461546,0.07548718,0.059076928,0.06235898,0.07876924,0.10502565,0.15097436,0.13784617,0.101743594,0.072205134,0.06564103,0.09189744,0.1148718,0.1148718,0.10502565,0.09189744,0.07548718,0.07548718,0.07876924,0.07876924,0.08533334,0.108307704,0.059076928,0.03938462,0.049230773,0.07548718,0.0951795,0.055794876,0.02297436,0.006564103,0.009846155,0.026256412,0.04594872,0.06235898,0.055794876,0.036102567,0.013128206,0.026256412,0.059076928,0.08205129,0.07876924,0.068923086,0.06235898,0.08861539,0.16410258,0.3117949,0.56451285,0.43651286,0.29538465,0.318359,0.5677949,1.0043077,1.0075898,0.9517949,0.81394875,0.6268718,0.4660513,0.49887183,0.571077,0.7056411,0.83035904,0.77128214,0.46276927,0.31507695,0.52512825,0.94523084,1.1093334,1.3095386,2.0020514,2.2646155,2.0808206,2.349949,2.9735386,2.556718,2.4057438,3.0293336,4.128821,5.106872,5.0510774,4.141949,2.8291285,1.8313848,1.7263591,2.1792822,2.5961027,2.7306669,2.6847181,2.7109745,2.537026,2.740513,3.4067695,4.1222568,4.388103,4.4406157,4.4274874,4.4340515,4.4767184,3.9614363,3.6660516,3.4100516,3.1540515,3.0030773,3.7251284,4.71959,5.546667,5.904411,5.61559,6.242462,6.3967185,5.979898,5.0609236,3.876103,3.31159,3.5872824,4.601436,5.87159,6.5444107,6.770872,6.928411,7.6307697,10.075898,16.022976,24.77949,31.442053,34.85539,34.773335,31.88513,26.948925,22.022566,18.484514,15.9573345,12.281437,8.402052,5.1265645,2.8717952,1.6902566,1.2800001,1.1848207,0.5874872,0.15097436,0.072205134,0.068923086,0.07548718,0.08205129,0.06564103,0.032820515,0.013128206,0.006564103,0.0032820515,0.0,0.0,0.006564103,0.0,0.0,0.0032820515,0.009846155,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.006564103,0.02297436,0.029538464,0.026256412,0.016410258,0.016410258,0.016410258,0.02297436,0.04266667,0.06564103,0.06564103,0.068923086,0.07548718,0.08533334,0.08533334,0.08205129,0.098461546,0.1148718,0.12471796,0.14112821,0.18051283,0.380718,0.764718,1.2242053,1.5064616,2.5173335,3.892513,5.4449234,6.4689236,5.76,3.5314875,1.5097437,0.446359,0.35774362,0.4955898,0.571077,0.571077,0.5874872,0.636718,0.67282057,0.81394875,1.1355898,1.5195899,1.975795,2.6387694,3.1442053,3.242667,3.2196925,3.1803079,3.0687182,2.793026,2.6486156,2.412308,2.0512822,1.7066668,1.4145643,1.2373334,1.1388719,1.0896411,1.0699488,1.079795,1.2931283,1.6114873,1.9561027,2.284308,2.412308,2.6256413,2.8127182,2.8914874,2.8324106,2.2416413,2.0775387,2.1202054,2.1924105,2.1924105,1.8970258,1.6869745,1.6771283,1.9462565,2.546872,2.789744,3.0851285,3.3805132,3.6036925,3.6758976,3.751385,3.6594875,3.3247182,2.8389745,2.4713848,2.6026669,2.8356924,3.1474874,3.2065644,2.3630772,5.8978467,5.924103,5.9930263,6.442667,7.062975,7.0892315,5.8945646,6.951385,7.755488,7.072821,4.962462,2.868513,2.4385643,3.515077,5.7829747,8.753231,10.952206,12.356924,13.269335,13.548308,12.612924,9.078155,6.3442054,4.565334,3.767795,3.8301542,4.201026,4.3060517,4.1222568,3.7448208,3.3772311,2.5107694,2.353231,2.8980515,3.5380516,3.0818465,3.8301542,5.179077,4.827898,3.4691284,4.8049235,5.5630774,6.0225644,6.3376417,6.2851286,5.2709746,4.7392826,4.604718,4.9296412,5.9569235,8.090257,10.108719,11.221334,10.28595,7.6603084,5.228308,3.6693337,2.041436,0.90256417,0.48574364,0.7187693,1.0666667,0.79097444,0.53825647,0.56451285,0.7318975,0.8369231,0.92553854,1.2307693,1.8018463,2.481231,2.4910772,2.294154,2.03159,1.7985642,1.6311796,1.6902566,1.8740515,2.097231,2.294154,2.425436,2.6715899,3.0391798,3.4100516,3.7021542,3.892513,3.9975388,4.082872,4.1025643,3.8400004,2.9210258,2.5698464,2.356513,2.1989746,2.0118976,1.7033848,1.4605129,1.2373334,0.9714873,0.702359,0.5874872,0.4201026,0.2986667,0.446359,0.7187693,0.6071795,0.8467693,1.6869745,1.8445129,1.3259488,1.4375386,1.4998976,1.0633847,0.98133343,1.3981539,1.7624617,1.8970258,1.2635899,0.9156924,1.1158975,1.3128207,1.4244103,1.529436,1.463795,1.211077,0.92225647,0.6268718,0.5218462,0.48246157,0.4397949,0.38728207,0.32820517,0.32820517,0.37415388,0.45292312,0.5415385,0.512,0.3446154,0.16082053,0.055794876,0.09189744,0.35446155,0.65312827,0.90584624,1.0010257,0.8008206,0.6301539,0.56451285,0.571077,0.5415385,0.28882053,0.17394873,0.108307704,0.068923086,0.049230773,0.04594872,0.049230773,0.06564103,0.08533334,0.108307704,0.13128206,0.118153855,0.08205129,0.072205134,0.0951795,0.108307704,0.15097436,0.2231795,0.20348719,0.10502565,0.07548718,0.08205129,0.1148718,0.17394873,0.25271797,0.36430773,0.4594872,0.46933338,0.512,0.6170257,0.73517954,0.82379496,0.90912825,0.9189744,0.9124103,1.0962052,1.8051283,2.7667694,3.5347695,3.8301542,3.5446157,1.9068719,1.1224617,0.77128214,0.61374366,0.5973334,1.0896411,1.3128207,1.3653334,1.3357949,1.3161026,0.9156924,0.86974365,1.0272821,1.1749744,1.0338463,0.761436,0.48902568,0.23630771,0.049230773,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.108307704,0.5481026,0.69251287,0.63343596,0.48574364,0.33805132,0.24943592,0.17723078,0.06235898,0.15753847,0.380718,0.31507695,0.08205129,0.21989745,0.3446154,0.32820517,0.31507695,0.37415388,0.57764107,0.7417436,0.81066674,0.84348726,0.8467693,0.9189744,1.0108719,1.1257436,1.3226668,1.5097437,1.6771283,1.719795,1.585231,1.2898463,1.0699488,0.827077,0.61374366,0.4397949,0.31507695,0.18379489,0.09189744,0.029538464,0.02297436,0.12143591,0.2100513,0.20676924,0.12471796,0.12143591,0.49887183,0.33476925,0.21989745,0.18379489,0.20348719,0.2100513,0.2100513,0.20020515,0.22646156,0.42338464,1.0108719,1.1946667,1.214359,1.020718,0.75487185,0.75487185,0.69907695,0.5973334,0.5349744,0.56451285,0.7253334,0.88615394,0.90584624,0.9878975,1.1257436,1.1060513,0.8763078,0.4594872,0.22646156,0.21661541,0.15425642,0.06235898,0.02297436,0.013128206,0.02297436,0.052512825,0.07876924,0.06235898,0.03938462,0.01969231,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.026256412,0.03938462,0.036102567,0.026256412,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.026256412,0.059076928,0.098461546,0.08205129,0.055794876,0.03938462,0.03938462,0.06564103,0.15097436,0.14441027,0.11158975,0.07876924,0.055794876,0.055794876,0.049230773,0.049230773,0.04594872,0.016410258,0.013128206,0.013128206,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.01969231,0.1148718,0.256,0.47917953,0.892718,0.9189744,0.764718,0.65641034,0.702359,0.8730257,1.0469744,1.020718,0.7581539,0.37415388,0.16410258,0.21989745,0.34789747,0.42994875,0.45292312,0.47917953,0.5481026,0.5349744,0.5316923,0.5415385,0.4660513,0.30194873,0.23302566,0.19364104,0.14441027,0.07548718,0.07876924,0.11158975,0.128,0.13128206,0.16410258,0.27241027,0.3708718,0.4266667,0.4266667,0.36758977,0.30851284,0.4397949,0.6071795,0.6662565,0.49887183,0.26256412,0.13456412,0.072205134,0.049230773,0.03938462,0.07548718,0.0951795,0.12471796,0.17394873,0.26584616,0.2100513,0.13784617,0.07548718,0.049230773,0.07876924,0.101743594,0.12471796,0.14441027,0.15753847,0.15425642,0.16082053,0.17066668,0.16082053,0.12471796,0.08205129,0.049230773,0.049230773,0.06564103,0.07876924,0.07548718,0.055794876,0.02297436,0.009846155,0.02297436,0.04594872,0.08861539,0.108307704,0.09189744,0.059076928,0.04594872,0.04266667,0.07876924,0.09189744,0.072205134,0.049230773,0.052512825,0.08861539,0.19692309,0.3511795,0.45292312,0.35774362,0.3314872,0.571077,1.1093334,1.8281027,1.5589745,1.2077949,0.86317956,0.57764107,0.37743592,0.46276927,0.5513847,0.58420515,0.6170257,0.8369231,0.62030774,0.47589746,0.48246157,0.65969235,0.97805136,1.0535386,1.3784616,1.847795,2.1497438,1.7624617,2.169436,2.740513,3.1573336,3.4855387,4.164923,4.453744,4.1156926,3.2164104,2.1825643,1.8018463,2.2121027,2.7437952,3.2032824,3.4921029,3.6332312,3.2623591,2.8717952,3.0687182,3.8629746,4.647385,4.962462,4.9362054,4.6802053,4.3290257,4.059898,4.010667,3.9909747,3.879385,3.754667,3.9056413,4.9427695,6.163693,7.000616,7.256616,7.128616,7.5454364,7.3682055,6.5969234,5.3037953,3.626667,2.8947694,2.865231,3.4691284,4.70318,6.636308,7.2927184,7.27959,8.024616,10.555078,15.507693,24.214975,29.518772,31.88185,32.17067,31.648823,28.419285,24.65149,21.106873,17.723078,13.610668,9.143796,5.4908724,3.0293336,1.6640002,0.83035904,0.69579494,0.4201026,0.17066668,0.04594872,0.06564103,0.07876924,0.07876924,0.06564103,0.04266667,0.026256412,0.016410258,0.006564103,0.0032820515,0.0032820515,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.006564103,0.006564103,0.0032820515,0.006564103,0.036102567,0.059076928,0.06235898,0.029538464,0.01969231,0.013128206,0.02297436,0.049230773,0.06564103,0.07876924,0.0951795,0.11158975,0.12471796,0.13128206,0.15097436,0.190359,0.23302566,0.25928208,0.26256412,0.24615386,0.2231795,0.20676924,0.23302566,0.35774362,1.2274873,2.6683078,4.4110775,5.9667697,6.619898,4.6966157,2.3236926,0.86974365,0.7450257,1.4342566,1.4539489,1.0305642,0.69907695,0.62030774,0.5907693,0.77128214,1.2307693,1.785436,2.4746668,3.5544617,4.2601027,4.2207184,3.9154875,3.620103,3.4002054,2.9440002,2.5600002,2.2383592,1.9692309,1.7493335,1.4998976,1.2471796,1.0994873,1.079795,1.1257436,1.2274873,1.4867693,1.9200002,2.481231,3.0654361,3.2065644,3.0162053,2.8521028,2.8717952,3.0490258,2.4451284,1.910154,1.6311796,1.5885129,1.5425643,1.4900514,1.4703591,1.5688206,1.8281027,2.2383592,2.4385643,2.92759,3.4724104,3.764513,3.4231799,3.0490258,2.8882053,2.665026,2.228513,1.5458462,1.3456411,1.3718976,1.7427694,2.2908719,2.5665643,4.0434875,4.1156926,3.9351797,4.3060517,4.8672824,4.073026,5.024821,6.820103,7.706257,7.0137444,5.156103,3.436308,3.498667,5.717334,9.350565,12.57354,14.194873,13.568001,11.851488,9.7673855,7.584821,4.9952826,3.0391798,2.0151796,1.913436,2.425436,2.9144619,3.639795,4.066462,4.013949,3.6463592,2.865231,3.045744,3.2525132,2.9965131,2.228513,3.131077,3.9351797,4.1780515,4.4734364,6.5017443,6.488616,6.2916927,5.8157954,4.965744,3.6463592,3.817026,4.8771286,6.7807183,9.028924,10.666668,9.67877,7.9294367,6.4623594,5.5072823,4.4701543,3.7152824,2.9768207,1.8576412,0.81394875,1.1454359,1.3751796,0.90256417,0.4955898,0.48902568,0.79425645,1.024,1.0568206,1.2504616,1.6640002,2.028308,2.176,1.910154,1.654154,1.5589745,1.5097437,1.4998976,1.8707694,2.231795,2.412308,2.487795,2.546872,3.0293336,3.629949,4.138667,4.457026,4.089436,3.639795,3.170462,2.7142565,2.2744617,2.2383592,2.0709746,1.8412309,1.6049232,1.4342566,1.4966155,1.5392822,1.5425643,1.463795,1.2209232,0.8795898,0.53825647,0.2986667,0.38728207,1.1454359,1.3161026,1.3489232,1.2274873,1.1552821,1.5721027,1.6311796,1.5556924,1.5819489,1.5819489,1.0666667,0.60389745,0.23302566,0.41025645,1.020718,1.3718976,1.4473847,1.2996924,1.014154,0.702359,0.51856416,0.5546667,0.6662565,0.7384616,0.72861546,0.65641034,0.508718,0.49887183,0.53825647,0.5513847,0.5021539,0.30851284,0.15753847,0.07876924,0.06564103,0.09189744,0.04266667,0.19692309,0.45620516,0.7384616,0.94523084,0.6892308,0.49887183,0.380718,0.3249231,0.28882053,0.28882053,0.28882053,0.25271797,0.19364104,0.16738462,0.14441027,0.128,0.128,0.13128206,0.108307704,0.0951795,0.072205134,0.049230773,0.036102567,0.06235898,0.12143591,0.19364104,0.19364104,0.13784617,0.13784617,0.2100513,0.32164106,0.36430773,0.3511795,0.4135385,0.5940513,0.86974365,0.98461545,0.892718,0.74830776,0.6498462,0.94523084,1.2570257,1.5097437,1.9364104,2.802872,3.6069746,3.7054362,2.9735386,1.8018463,1.5064616,1.2865642,1.0436924,0.7450257,0.4266667,0.6826667,1.142154,1.6475899,2.1070771,2.487795,1.3161026,0.892718,0.92553854,1.0338463,0.7778462,0.48574364,0.26584616,0.101743594,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.12143591,0.23630771,0.25928208,0.21333335,0.21333335,0.190359,0.072205134,0.036102567,0.0951795,0.108307704,0.118153855,0.15097436,0.27897438,0.48574364,0.65641034,0.81394875,0.761436,0.8533334,1.2438976,1.8904617,2.7963078,2.0611284,1.3456411,1.332513,1.723077,1.4441026,1.4998976,1.463795,1.1191796,0.47261542,0.7778462,0.73517954,0.508718,0.23958977,0.04594872,0.2297436,0.256,0.14769232,0.036102567,0.18379489,0.23302566,0.26256412,0.21989745,0.15425642,0.2297436,0.25271797,0.17723078,0.108307704,0.101743594,0.13784617,0.18707694,0.28882053,0.49887183,0.72861546,0.7778462,0.81394875,0.9156924,0.82379496,0.58420515,0.5349744,0.54482055,0.55794877,0.6301539,0.761436,0.88615394,0.94523084,0.86974365,0.8205129,0.8369231,0.82379496,0.702359,0.38728207,0.14441027,0.059076928,0.04594872,0.02297436,0.006564103,0.006564103,0.016410258,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.03938462,0.07548718,0.08861539,0.06564103,0.026256412,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06235898,0.08533334,0.072205134,0.03938462,0.016410258,0.101743594,0.14112821,0.14112821,0.1148718,0.09189744,0.055794876,0.036102567,0.029538464,0.026256412,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.029538464,0.10502565,0.20348719,0.29538465,0.35774362,0.380718,0.35774362,0.7187693,0.9682052,0.9944616,1.0666667,1.4966155,1.591795,1.3423591,0.8008206,0.09189744,0.07876924,0.26912823,0.4955898,0.636718,0.6268718,0.47917953,0.3314872,0.2231795,0.16082053,0.13784617,0.08861539,0.08533334,0.108307704,0.12471796,0.07548718,0.08861539,0.101743594,0.11158975,0.1148718,0.09189744,0.14112821,0.18051283,0.19692309,0.19692309,0.18379489,0.18379489,0.2297436,0.30194873,0.3511795,0.28882053,0.23958977,0.2100513,0.17394873,0.12471796,0.07548718,0.052512825,0.036102567,0.055794876,0.108307704,0.16738462,0.18051283,0.14769232,0.10502565,0.06564103,0.029538464,0.04266667,0.09189744,0.12143591,0.118153855,0.108307704,0.13128206,0.21989745,0.26256412,0.20348719,0.04594872,0.02297436,0.06235898,0.1148718,0.13784617,0.07548718,0.06564103,0.04266667,0.02297436,0.02297436,0.04594872,0.068923086,0.07548718,0.07548718,0.08205129,0.108307704,0.0951795,0.08205129,0.052512825,0.013128206,0.0,0.02297436,0.08533334,0.3117949,0.6235898,0.7318975,0.5973334,0.636718,0.88287187,1.1815386,1.204513,0.9353847,0.6235898,0.43323082,0.36758977,0.24287182,0.26912823,0.47589746,0.48902568,0.3249231,0.39712822,0.7384616,0.7318975,0.6826667,0.69907695,0.6859488,0.7122052,1.5589745,2.176,2.1267693,1.6016412,2.665026,3.3312824,3.7415388,4.141949,4.896821,5.362872,4.598154,3.3247182,2.349949,2.5928206,3.4231799,3.8498464,3.9417439,4.023795,4.6834874,4.5390773,4.31918,4.2338467,4.4996924,5.356308,5.904411,6.0324106,5.6976414,5.07077,4.5456414,4.2535386,4.007385,3.9581542,4.2240005,4.8836927,6.2129235,7.397744,8.129642,8.3134365,8.057437,8.03118,6.698667,5.044513,3.7120004,2.989949,2.8553848,3.2164104,4.1550775,5.4153852,6.3934364,7.2369237,7.7292314,9.494975,12.944411,17.302977,22.698668,26.466463,27.831797,27.280413,26.535387,26.10872,24.638361,22.46236,19.383797,14.647796,9.508103,5.605744,2.9144619,1.3554872,0.79425645,0.8533334,0.5021539,0.16082053,0.029538464,0.09189744,0.10502565,0.08861539,0.06564103,0.03938462,0.016410258,0.016410258,0.016410258,0.016410258,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.02297436,0.029538464,0.026256412,0.016410258,0.03938462,0.101743594,0.17394873,0.20020515,0.09189744,0.029538464,0.006564103,0.013128206,0.029538464,0.029538464,0.04266667,0.072205134,0.10502565,0.13128206,0.16738462,0.21661541,0.29210258,0.37743592,0.446359,0.45620516,0.43323082,0.4004103,0.33805132,0.27241027,0.25928208,0.45620516,0.98133343,1.5458462,2.0906668,2.7634873,4.2272825,2.9440002,1.5458462,1.7263591,4.240411,4.096,2.546872,1.4933335,1.2996924,0.82379496,0.7515898,1.1454359,1.7920002,2.481231,3.006359,3.006359,3.0326157,2.9046156,2.6683078,2.5928206,2.412308,2.2383592,2.0906668,1.9692309,1.847795,1.529436,1.2406155,1.014154,0.88287187,0.86974365,0.9419488,1.1355898,1.5130258,2.0512822,2.6256413,2.6617439,2.412308,2.3663592,2.7175386,3.4034874,3.0720003,2.2022567,1.7624617,1.8576412,1.723077,1.6147693,1.5491283,1.5327181,1.5786668,1.723077,2.1530259,2.7634873,3.4527183,3.9844105,3.9975388,3.058872,2.484513,2.1234872,1.7657437,1.1454359,1.0108719,1.1520001,1.4178462,1.9068719,2.9440002,5.7403083,5.648411,5.664821,5.914257,6.3967185,6.99077,7.650462,8.3823595,8.667898,7.8670774,5.2315903,3.5478978,3.0358977,3.69559,5.2578464,7.200821,7.643898,7.584821,8.306872,9.31118,8.316719,6.626462,4.673641,3.8104618,4.1682053,4.673641,5.277539,5.6451287,5.031385,3.9286156,4.0500517,5.034667,5.832206,6.7840004,7.433847,6.5378466,4.6867695,4.125539,4.525949,5.5269747,6.744616,6.3310776,6.1538467,5.8781543,5.3924108,4.8049235,4.5390773,5.3169236,6.3442054,6.931693,6.5280004,5.5991797,4.9854364,4.6244106,4.3060517,3.6758976,3.3312824,3.7284105,4.525949,4.7589746,2.8422565,2.097231,1.4539489,0.8566154,0.5284103,0.9517949,0.9878975,0.8533334,0.90256417,1.1782565,1.4178462,1.5261539,1.522872,1.5524104,1.6705642,1.8281027,1.9232821,1.9626669,2.0939488,2.3401027,2.609231,2.9636924,3.43959,3.7973337,3.9056413,3.7349746,3.2032824,2.7142565,2.3466668,2.1103592,1.9429746,1.8084104,1.6869745,1.5195899,1.332513,1.2406155,1.6114873,1.8740515,1.9856411,1.8773335,1.4276924,0.8041026,0.6235898,0.74830776,1.0305642,1.3259488,1.3423591,1.211077,1.0699488,1.1355898,1.7066668,1.7755898,1.5622566,1.3784616,1.3193847,1.276718,1.270154,1.3423591,1.4309745,1.394872,1.0075898,0.9714873,1.2406155,1.3587693,1.1815386,0.8598975,0.702359,0.83035904,0.8960001,0.8205129,0.764718,0.6695385,0.4955898,0.4004103,0.40369233,0.39384618,0.29538465,0.2231795,0.17066668,0.14112821,0.1148718,0.049230773,0.16738462,0.3446154,0.50543594,0.60389745,0.47589746,0.38728207,0.3117949,0.21661541,0.08205129,0.21989745,0.26912823,0.24615386,0.18379489,0.13128206,0.118153855,0.10502565,0.07876924,0.049230773,0.04594872,0.06235898,0.072205134,0.072205134,0.06564103,0.06235898,0.072205134,0.0951795,0.108307704,0.21333335,0.61374366,0.75487185,0.6104616,0.44307697,0.36430773,0.33805132,0.38400003,0.4660513,0.6629744,0.88287187,0.8336411,0.6465641,0.9353847,1.276718,1.5097437,1.7296412,2.0217438,2.2482052,2.3072822,2.166154,1.8740515,1.5031796,1.4473847,1.401436,1.2242053,0.9288206,0.9485129,1.4966155,1.9954873,2.028308,1.3029745,1.0994873,0.8533334,0.6301539,0.52512825,0.67938465,0.38728207,0.14441027,0.01969231,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06235898,0.0951795,0.08205129,0.04266667,0.04266667,0.07548718,0.08533334,0.059076928,0.01969231,0.02297436,0.02297436,0.13128206,0.24943592,0.36430773,0.5349744,0.83035904,0.7089231,0.7187693,1.0043077,1.3292309,0.74830776,0.574359,0.5973334,0.7384616,1.0404103,1.1224617,1.0929232,0.9353847,0.6432821,0.23958977,0.18379489,0.14769232,0.101743594,0.049230773,0.009846155,0.13456412,0.16082053,0.0951795,0.006564103,0.036102567,0.20348719,0.31507695,0.35774362,0.36430773,0.38728207,0.4201026,0.44964105,0.5284103,0.62030774,0.5874872,0.5316923,0.62030774,0.81066674,0.9353847,0.7417436,0.61374366,0.71548724,0.81394875,0.78769237,0.6301539,0.3708718,0.26912823,0.2855385,0.37415388,0.50543594,0.65641034,0.69579494,0.6432821,0.5218462,0.3708718,0.36758977,0.23630771,0.1148718,0.059076928,0.059076928,0.032820515,0.01969231,0.013128206,0.013128206,0.0032820515,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.01969231,0.026256412,0.016410258,0.026256412,0.026256412,0.02297436,0.01969231,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.013128206,0.0032820515,0.0,0.0,0.0,0.013128206,0.02297436,0.032820515,0.029538464,0.016410258,0.04266667,0.10502565,0.190359,0.26256412,0.23958977,0.1148718,0.06564103,0.04594872,0.026256412,0.016410258,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.013128206,0.07548718,0.22646156,0.16082053,0.08861539,0.059076928,0.07548718,0.08861539,0.12143591,0.36430773,0.6498462,0.8205129,0.7253334,1.1355898,1.5261539,1.6968206,1.4112822,0.41025645,0.12471796,0.10502565,0.2100513,0.32820517,0.39384618,0.43323082,0.43651286,0.36102566,0.24287182,0.19692309,0.19692309,0.25928208,0.2986667,0.28882053,0.25928208,0.28225642,0.34133336,0.34789747,0.28882053,0.22646156,0.18707694,0.20348719,0.22646156,0.23958977,0.256,0.18707694,0.14441027,0.118153855,0.108307704,0.0951795,0.0951795,0.12143591,0.13128206,0.11158975,0.052512825,0.036102567,0.02297436,0.01969231,0.02297436,0.04594872,0.08861539,0.098461546,0.098461546,0.0951795,0.06564103,0.07876924,0.12143591,0.12143591,0.07876924,0.059076928,0.101743594,0.15097436,0.16410258,0.128,0.059076928,0.04266667,0.07876924,0.20676924,0.34133336,0.27241027,0.13128206,0.0951795,0.07548718,0.059076928,0.08205129,0.108307704,0.098461546,0.098461546,0.1148718,0.118153855,0.108307704,0.0951795,0.08205129,0.072205134,0.049230773,0.032820515,0.098461546,0.31507695,0.6662565,1.0502565,1.0929232,1.0502565,1.0469744,1.079795,1.0469744,0.67938465,0.47261542,0.39712822,0.36430773,0.23302566,0.45292312,0.5021539,0.45620516,0.45620516,0.71548724,0.8205129,0.7778462,0.6170257,0.4594872,0.5152821,0.571077,0.9189744,1.6869745,2.4582565,2.2744617,2.281026,2.612513,3.6857438,5.21518,6.2162056,6.183385,4.8705645,3.7940516,3.6168208,4.1452312,4.535795,4.516103,4.4406157,4.5587697,5.0018463,5.4908724,5.428513,5.2348723,5.277539,5.868308,6.6428723,6.242462,5.349744,4.5095387,4.132103,4.3651285,4.3684106,4.3060517,4.46359,5.2480006,7.076103,8.474257,9.353847,9.908514,10.607591,8.864821,6.633026,4.8771286,4.092718,4.309334,4.2830772,4.0303593,3.889231,4.4307694,6.491898,8.231385,9.728001,11.963078,15.793232,21.930668,25.488413,26.436926,25.760822,24.658052,24.556309,24.6679,24.083694,22.416412,19.373951,14.795488,9.819899,5.651693,2.8225644,1.3423591,0.6826667,0.44307697,0.24287182,0.11158975,0.06564103,0.1148718,0.15753847,0.15753847,0.14769232,0.14769232,0.16082053,0.17066668,0.16082053,0.12471796,0.07876924,0.036102567,0.016410258,0.013128206,0.02297436,0.032820515,0.02297436,0.026256412,0.036102567,0.04266667,0.04266667,0.03938462,0.101743594,0.14441027,0.15425642,0.13456412,0.10502565,0.08205129,0.04594872,0.026256412,0.036102567,0.055794876,0.10502565,0.15425642,0.20020515,0.24615386,0.30194873,0.3511795,0.38400003,0.41025645,0.42994875,0.4201026,0.40697438,0.39056414,0.35774362,0.3117949,0.27241027,0.26256412,0.37743592,0.50543594,0.60389745,0.69907695,0.9419488,0.7417436,1.0765129,2.4188719,4.71959,3.7021542,2.2744617,1.2832822,0.9288206,0.77456415,0.761436,0.9124103,1.2274873,1.6278975,1.9692309,1.9396925,1.7985642,1.5524104,1.2964103,1.214359,1.3456411,1.4309745,1.5688206,1.7329233,1.7985642,1.6640002,1.5031796,1.2340513,0.9156924,0.74830776,0.85005134,1.079795,1.5261539,2.1398976,2.733949,2.556718,2.2547693,2.1924105,2.4615386,2.8914874,3.0194874,2.7700515,2.3204105,1.8838975,1.7132308,1.5524104,1.4998976,1.5786668,1.7263591,1.785436,1.910154,2.166154,2.5862565,3.0851285,3.4494362,3.1540515,2.4681027,1.8609232,1.4933335,1.2406155,0.9911796,0.9124103,0.97805136,1.1881026,1.5524104,5.605744,5.221744,5.024821,5.0510774,5.35959,6.0258465,6.738052,8.280616,9.468719,9.5835905,8.362667,7.4371285,6.76759,6.5345645,6.7905645,7.4699492,8.218257,8.736821,9.353847,9.622975,8.333129,6.1440005,4.8147697,4.8082056,6.0028725,7.6964107,8.65477,8.011488,5.622154,3.1376412,4.0041027,5.1167183,6.1768208,7.7948723,9.304616,8.749949,6.7314878,5.333334,5.612308,6.9349747,6.997334,6.088206,5.3431797,4.893539,4.785231,4.969026,5.1232824,5.179077,5.3169236,5.4186673,5.0543594,4.525949,4.0402055,3.7021542,3.5741541,3.6726158,4.8640003,5.156103,5.293949,5.179077,3.8498464,2.4024618,1.5622566,1.017436,0.7318975,0.9189744,1.0469744,0.9747693,0.9288206,1.024,1.276718,1.3653334,1.4473847,1.5556924,1.6672822,1.7066668,1.7329233,1.7690258,1.9987694,2.3630772,2.5862565,2.8947694,3.2065644,3.31159,3.1638978,2.878359,2.4057438,1.9265642,1.6278975,1.5392822,1.5130258,1.4572309,1.3193847,1.1520001,1.0929232,1.3653334,2.166154,2.356513,2.284308,2.0841026,1.6640002,0.892718,1.0469744,1.3357949,1.332513,0.9419488,0.7220513,0.955077,1.3226668,1.6213335,1.7755898,1.6508719,1.7165129,1.9167181,1.9856411,1.463795,1.3554872,1.5163078,1.8215386,1.9265642,1.2635899,1.1946667,1.3817437,1.467077,1.2964103,0.9288206,0.72861546,0.7187693,0.69251287,0.60389745,0.5546667,0.5218462,0.47917953,0.43651286,0.39056414,0.34789747,0.27569234,0.2297436,0.23958977,0.26912823,0.23958977,0.12471796,0.26256412,0.39384618,0.4135385,0.36430773,0.23630771,0.190359,0.17066668,0.14441027,0.0951795,0.19364104,0.23958977,0.23630771,0.18379489,0.0951795,0.10502565,0.118153855,0.13456412,0.15425642,0.20348719,0.13456412,0.07548718,0.049230773,0.052512825,0.068923086,0.068923086,0.07548718,0.0951795,0.17066668,0.35774362,0.47917953,0.47261542,0.39056414,0.29538465,0.23958977,0.3446154,0.60389745,0.82379496,0.8960001,0.79097444,0.65641034,0.9714873,1.3423591,1.6443079,2.0250258,2.5600002,2.7667694,2.8192823,2.7766156,2.5796926,1.9626669,1.9265642,1.9528207,1.7657437,1.3554872,0.8992821,1.0994873,1.5064616,1.7887181,1.7493335,1.1618463,0.761436,0.5218462,0.43323082,0.49230772,0.190359,0.04594872,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01969231,0.052512825,0.04266667,0.0,0.0,0.01969231,0.036102567,0.026256412,0.0,0.0,0.02297436,0.06235898,0.098461546,0.14112821,0.23958977,0.34133336,0.5415385,0.702359,0.7089231,0.47589746,0.16738462,0.26584616,0.446359,0.56451285,0.6301539,0.58420515,0.47917953,0.34789747,0.2100513,0.072205134,0.013128206,0.0,0.108307704,0.24615386,0.128,0.17066668,0.20020515,0.14112821,0.04266667,0.072205134,0.3117949,0.5907693,0.7515898,0.7253334,0.5546667,0.41682056,0.38400003,0.5874872,0.90584624,0.95835906,0.9616411,1.401436,1.5064616,1.1191796,0.6859488,0.60389745,0.72861546,0.7778462,0.636718,0.380718,0.19692309,0.101743594,0.07876924,0.11158975,0.16410258,0.2855385,0.2855385,0.23958977,0.17723078,0.11158975,0.13128206,0.098461546,0.055794876,0.032820515,0.032820515,0.016410258,0.009846155,0.006564103,0.0032820515,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.009846155,0.0,0.013128206,0.01969231,0.02297436,0.016410258,0.0,0.006564103,0.009846155,0.009846155,0.013128206,0.02297436,0.016410258,0.013128206,0.009846155,0.009846155,0.009846155,0.009846155,0.006564103,0.013128206,0.029538464,0.068923086,0.04594872,0.049230773,0.08533334,0.13128206,0.13784617,0.07876924,0.06235898,0.059076928,0.052512825,0.032820515,0.01969231,0.006564103,0.0,0.0032820515,0.009846155,0.009846155,0.0032820515,0.006564103,0.40697438,1.9593848,1.8838975,0.7844103,0.04266667,0.009846155,0.006564103,0.026256412,0.12143591,0.29210258,0.48574364,0.6235898,1.0994873,1.6180514,1.7329233,1.3128207,0.52512825,0.18707694,0.12471796,0.15097436,0.17394873,0.20676924,0.40369233,0.4594872,0.40697438,0.2986667,0.20348719,0.19364104,0.23958977,0.28225642,0.2986667,0.3052308,0.3446154,0.35774362,0.318359,0.24615386,0.18707694,0.17723078,0.20676924,0.24615386,0.27241027,0.28225642,0.21333335,0.15097436,0.1148718,0.101743594,0.06564103,0.055794876,0.06564103,0.072205134,0.06235898,0.036102567,0.032820515,0.026256412,0.02297436,0.01969231,0.02297436,0.04266667,0.052512825,0.06564103,0.08205129,0.0951795,0.13456412,0.27241027,0.3117949,0.21333335,0.06564103,0.08205129,0.14441027,0.16738462,0.128,0.04266667,0.029538464,0.07548718,0.27897438,0.67282057,1.1979488,0.77128214,0.512,0.36430773,0.29210258,0.26584616,0.20348719,0.16738462,0.17394873,0.19692309,0.15753847,0.108307704,0.08861539,0.14769232,0.22646156,0.14441027,0.10502565,0.16738462,0.33476925,0.5940513,0.9353847,1.0601027,1.0469744,0.9485129,0.8960001,1.079795,1.1158975,0.6662565,0.33476925,0.28882053,0.26584616,0.37415388,0.36758977,0.3511795,0.40369233,0.5907693,0.6629744,0.60389745,0.4660513,0.3511795,0.41025645,0.65969235,0.8336411,1.2012309,1.6968206,1.9298463,2.2055387,2.9078977,4.076308,5.395693,6.180103,5.5236926,4.5587697,4.1780515,4.4964104,4.8607183,4.827898,4.5062566,4.082872,3.889231,4.4045134,4.9985647,5.284103,5.3727183,5.467898,5.858462,6.2129235,5.730462,4.972308,4.3716927,4.210872,4.571898,4.7917953,4.84759,5.0182567,5.87159,7.9195905,9.278359,10.361437,11.349334,12.179693,10.666668,8.254359,6.1308722,4.9788723,4.969026,5.1232824,4.457026,3.876103,4.266667,6.488616,8.323282,9.068309,9.885539,12.465232,19.02277,22.511591,23.555285,22.944822,21.979898,22.478771,22.820105,22.646156,21.477745,18.884924,14.519796,9.90195,5.8453336,2.934154,1.3095386,0.65641034,0.43323082,0.30194873,0.20020515,0.12143591,0.11158975,0.14769232,0.16738462,0.20348719,0.26256412,0.35446155,0.47589746,0.52512825,0.5218462,0.47261542,0.40369233,0.27569234,0.16082053,0.08533334,0.052512825,0.049230773,0.026256412,0.026256412,0.02297436,0.01969231,0.01969231,0.055794876,0.072205134,0.07548718,0.08861539,0.14441027,0.108307704,0.06564103,0.036102567,0.03938462,0.068923086,0.13128206,0.19364104,0.26256412,0.32820517,0.39056414,0.43323082,0.45620516,0.47917953,0.49230772,0.4660513,0.41682056,0.380718,0.35446155,0.33805132,0.3117949,0.27897438,0.26584616,0.25271797,0.2231795,0.18379489,0.13784617,0.14769232,0.4594872,1.1782565,2.2744617,2.3138463,3.170462,3.7120004,3.3312824,1.9265642,1.0994873,0.81394875,0.88287187,1.1520001,1.4802053,1.3259488,1.1749744,1.0436924,0.94523084,0.88943595,0.9124103,0.9485129,1.0666667,1.3817437,2.03159,2.0118976,1.847795,1.7427694,1.6049232,1.0469744,0.8795898,1.0075898,1.394872,1.8773335,2.166154,2.097231,2.0841026,2.3794873,2.8750772,3.1081028,3.0916924,2.7766156,2.3827693,2.0742567,1.9659488,1.8248206,1.6147693,1.5458462,1.657436,1.8084104,1.9167181,2.0709746,2.28759,2.5337439,2.7437952,2.609231,2.100513,1.5721027,1.1979488,0.96492314,0.80738467,0.7318975,0.74830776,0.8336411,0.9485129,5.2414365,4.972308,4.7655387,4.647385,4.5029745,4.0434875,4.5095387,6.1374364,7.8014364,9.321027,11.474052,11.979488,11.07036,9.734565,8.625232,8.073847,8.300308,8.241231,7.9261546,7.3353853,6.419693,5.0543594,4.240411,4.535795,5.901129,7.709539,8.251078,6.9382567,4.332308,2.0841026,2.930872,4.6834874,5.8190775,7.0990777,8.2904625,8.169026,8.080411,7.2992826,7.259898,7.762052,6.997334,6.012718,5.152821,4.6572313,4.585026,4.8147697,5.1659493,4.9362054,4.6572313,4.535795,4.450462,4.132103,3.620103,3.4100516,3.6069746,3.9089234,5.540103,6.5805135,6.87918,6.3967185,5.2053337,2.737231,1.5261539,1.0732309,0.9944616,1.0469744,1.1158975,1.1126155,1.1060513,1.1815386,1.4473847,1.5064616,1.5130258,1.5097437,1.5031796,1.4441026,1.5491283,1.6836925,1.9331284,2.231795,2.3663592,2.9078977,3.239385,3.2000003,2.8389745,2.4024618,1.9561027,1.4834872,1.148718,1.024,1.1158975,1.1716924,1.1716924,1.3850257,1.8281027,2.231795,2.8488207,2.868513,2.5731285,2.172718,1.8149745,1.2307693,1.204513,1.401436,1.5031796,1.1881026,0.80738467,1.0502565,1.4933335,1.8313848,1.847795,1.8970258,2.228513,2.5074873,2.3696413,1.4342566,1.6869745,1.7624617,1.8313848,1.8018463,1.3292309,1.2242053,1.214359,1.1848207,1.0929232,0.9517949,0.7515898,0.6104616,0.508718,0.4397949,0.38400003,0.3708718,0.40369233,0.4266667,0.40369233,0.318359,0.23302566,0.19692309,0.27897438,0.41682056,0.380718,0.2297436,0.30851284,0.38400003,0.35774362,0.25271797,0.118153855,0.07548718,0.09189744,0.13456412,0.16738462,0.14769232,0.17723078,0.19364104,0.16082053,0.07548718,0.0951795,0.15097436,0.20676924,0.24943592,0.26584616,0.16410258,0.0951795,0.07876924,0.11158975,0.17394873,0.16410258,0.14441027,0.12471796,0.1148718,0.0951795,0.20348719,0.3249231,0.33476925,0.24287182,0.21989745,0.34789747,0.6170257,0.77456415,0.7811283,0.80738467,0.9321026,1.3259488,2.0250258,2.8849232,3.5774362,3.9647183,3.8400004,3.6627696,3.5938463,3.495385,3.1015387,3.0949745,3.0358977,2.7109745,2.1300514,1.3915899,1.1355898,1.2504616,1.6738462,2.3827693,1.3915899,0.8205129,0.55794877,0.46276927,0.3708718,0.07548718,0.0,0.06235898,0.128,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.026256412,0.026256412,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02297436,0.009846155,0.0,0.006564103,0.036102567,0.1148718,0.380718,0.51856416,0.39384618,0.055794876,0.13784617,0.28882053,0.42994875,0.49230772,0.41682056,0.31507695,0.24943592,0.2231795,0.26256412,0.41025645,0.47261542,0.44307697,0.41682056,0.43323082,0.48902568,0.55794877,0.5415385,0.43651286,0.3117949,0.3117949,0.4397949,0.60061544,0.702359,0.67282057,0.48902568,0.3052308,0.36102566,0.6465641,1.0436924,1.3193847,1.6771283,2.0086155,1.8379488,1.2176411,0.73517954,0.702359,0.764718,0.7187693,0.508718,0.23958977,0.15097436,0.07548718,0.026256412,0.0,0.0,0.052512825,0.026256412,0.0,0.0032820515,0.016410258,0.02297436,0.02297436,0.01969231,0.013128206,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.01969231,0.026256412,0.02297436,0.006564103,0.0,0.006564103,0.01969231,0.055794876,0.128,0.23302566,0.11158975,0.04266667,0.01969231,0.029538464,0.03938462,0.07876924,0.07876924,0.055794876,0.16738462,0.72861546,0.83035904,0.7417436,0.446359,0.118153855,0.118153855,0.14441027,0.08205129,0.049230773,0.059076928,0.04594872,0.02297436,0.006564103,0.0,0.0032820515,0.016410258,0.016410258,0.009846155,0.0032820515,0.40697438,2.038154,2.294154,1.0994873,0.17723078,0.049230773,0.029538464,0.009846155,0.032820515,0.12143591,0.3117949,0.6301539,1.2274873,1.7755898,1.9232821,1.591795,0.9714873,0.48902568,0.26256412,0.16738462,0.128,0.098461546,0.27241027,0.3314872,0.31507695,0.24615386,0.15097436,0.14441027,0.17723078,0.21661541,0.23958977,0.24943592,0.27569234,0.23958977,0.18707694,0.13456412,0.101743594,0.12143591,0.15097436,0.190359,0.2231795,0.2231795,0.15753847,0.12471796,0.118153855,0.12143591,0.08861539,0.06564103,0.055794876,0.049230773,0.04266667,0.04266667,0.032820515,0.032820515,0.03938462,0.04266667,0.049230773,0.03938462,0.032820515,0.036102567,0.049230773,0.068923086,0.14441027,0.33476925,0.47589746,0.446359,0.16082053,0.11158975,0.18379489,0.25271797,0.23958977,0.10502565,0.03938462,0.06564103,0.27241027,0.702359,1.3522053,1.0502565,0.88615394,0.7056411,0.49230772,0.33805132,0.3249231,0.37743592,0.4201026,0.39384618,0.28225642,0.17723078,0.16082053,0.24287182,0.3314872,0.2231795,0.23302566,0.38400003,0.64000005,0.96492314,1.3456411,1.2668719,1.079795,0.8402052,0.7450257,1.1290257,1.2504616,0.7844103,0.4660513,0.4594872,0.3511795,0.318359,0.3511795,0.43651286,0.51856416,0.52512825,0.49230772,0.39056414,0.28882053,0.26584616,0.43323082,0.8369231,0.86646163,0.90912825,1.148718,1.5556924,2.0020514,2.806154,3.9122055,5.106872,6.052103,5.1856413,4.394667,4.059898,4.1124105,4.0500517,4.1222568,3.882667,3.4494362,3.170462,3.6168208,4.8705645,5.6287184,5.7698464,5.5663595,5.674667,5.7731285,5.5236926,5.106872,4.7360005,4.670359,4.8705645,5.044513,5.146257,5.3431797,5.9930263,7.719385,9.173334,11.145847,13.354668,14.444309,13.302155,10.387693,7.6077952,5.940513,5.431795,5.4482055,4.886975,4.391385,4.5587697,5.943795,7.574975,7.8112826,7.936001,9.6525135,15.090873,21.333336,23.64718,23.2599,21.746874,21.051079,20.614565,20.450462,19.98113,18.310566,14.208001,9.977437,6.232616,3.3444104,1.522872,0.81394875,0.5677949,0.4266667,0.30851284,0.2100513,0.18051283,0.18051283,0.17394873,0.2100513,0.29538465,0.4201026,0.636718,0.82379496,0.9288206,0.9353847,0.8533334,0.65969235,0.48246157,0.3511795,0.26256412,0.19692309,0.07548718,0.026256412,0.013128206,0.006564103,0.013128206,0.029538464,0.036102567,0.04594872,0.072205134,0.12471796,0.101743594,0.07548718,0.068923086,0.08861539,0.14441027,0.2297436,0.32820517,0.42994875,0.508718,0.49887183,0.47261542,0.446359,0.43651286,0.4397949,0.4135385,0.34789747,0.2986667,0.27569234,0.26912823,0.256,0.24943592,0.24287182,0.22646156,0.20676924,0.190359,0.190359,0.26256412,0.3249231,0.4004103,0.58420515,1.1323078,2.6223593,3.6496413,3.4592824,1.9495386,0.96492314,0.61374366,0.6301539,0.8336411,1.1191796,0.94523084,0.8402052,0.8172308,0.8598975,0.9353847,0.85005134,0.76800007,0.7581539,0.9878975,1.7263591,1.9068719,1.8937438,1.8740515,1.7591796,1.1815386,0.9156924,1.0436924,1.3292309,1.595077,1.7099489,1.7263591,1.8281027,2.2186668,2.7536411,2.9440002,2.861949,2.3958976,2.0611284,2.0250258,2.1070771,2.0709746,1.785436,1.5819489,1.595077,1.7788719,1.9265642,2.156308,2.349949,2.4615386,2.5304618,2.1530259,1.7263591,1.3423591,1.0601027,0.892718,0.84348726,0.8008206,0.77456415,0.761436,0.761436,5.113436,5.3037953,5.5532312,5.605744,5.074052,3.43959,3.4756925,4.2994876,5.5007186,7.50277,11.546257,12.826258,11.772718,9.856001,8.060719,6.872616,5.723898,4.417641,3.4592824,3.121231,3.4297438,4.279795,4.132103,4.1878977,4.7327185,5.149539,4.7983594,3.757949,2.7864618,2.4024618,2.8717952,5.8486156,7.2631803,7.427283,6.9349747,6.675693,8.51036,8.89436,8.444718,7.6143594,6.7150774,6.114462,5.8256416,5.658257,5.4908724,5.280821,5.4153852,5.3792825,5.0543594,4.5062566,4.007385,3.5249233,3.131077,3.3214362,3.882667,3.892513,5.0116925,7.4108725,9.002667,8.694155,6.4032826,3.062154,1.4834872,1.0666667,1.204513,1.276718,1.1257436,1.1126155,1.2077949,1.3718976,1.5688206,1.585231,1.4736412,1.3653334,1.3226668,1.3226668,1.522872,1.6869745,1.8412309,2.0217438,2.2514873,3.2853336,4.092718,4.384821,4.1091285,3.4756925,2.6978464,2.034872,1.4703591,1.1716924,1.5097437,1.5556924,1.654154,2.2088206,3.0391798,3.383795,3.4330258,3.3247182,2.8488207,2.2088206,2.0184617,1.8904617,1.3817437,1.2865642,1.6640002,1.847795,1.4933335,1.4966155,1.6147693,1.7427694,1.910154,2.2646155,2.553436,2.5206156,2.103795,1.4178462,2.2482052,2.1956925,1.7329233,1.2603078,1.1191796,0.8795898,0.7253334,0.65641034,0.69907695,0.88943595,0.7089231,0.5415385,0.446359,0.41025645,0.36758977,0.3314872,0.31507695,0.36102566,0.41682056,0.30851284,0.20676924,0.14441027,0.256,0.44964105,0.4135385,0.27897438,0.23958977,0.24615386,0.256,0.20676924,0.118153855,0.07548718,0.09189744,0.14441027,0.18707694,0.0951795,0.108307704,0.13128206,0.12471796,0.08861539,0.101743594,0.17723078,0.24615386,0.26256412,0.19692309,0.16410258,0.15425642,0.17723078,0.2297436,0.3117949,0.28225642,0.23302566,0.16738462,0.098461546,0.07548718,0.19364104,0.34133336,0.4201026,0.45292312,0.56123084,0.5940513,0.56451285,0.5316923,0.6071795,0.9419488,1.4834872,2.103795,3.5905645,5.546667,6.36718,5.6976414,4.9427695,4.345436,4.007385,3.892513,4.056616,4.073026,3.8728209,3.43959,2.8127182,2.0808206,1.529436,1.3095386,1.5589745,2.3991797,1.6049232,1.0601027,0.7187693,0.5152821,0.3708718,0.15425642,0.098461546,0.20020515,0.28882053,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.02297436,0.23302566,0.26912823,0.23630771,0.190359,0.13128206,0.20020515,0.31507695,0.4201026,0.46276927,0.39712822,0.42994875,0.4955898,0.61374366,0.7975385,1.0305642,1.1388719,1.083077,0.7778462,0.49887183,0.88615394,1.0272821,0.88287187,0.6892308,0.571077,0.5415385,0.50543594,0.39384618,0.31507695,0.28882053,0.25271797,0.2100513,0.4955898,0.82379496,1.1290257,1.5753847,2.2482052,2.0250258,1.5130258,1.0502565,0.7187693,0.6892308,0.65641034,0.5907693,0.48902568,0.35446155,0.18707694,0.108307704,0.052512825,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.013128206,0.013128206,0.013128206,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0,0.0,0.0032820515,0.013128206,0.02297436,0.02297436,0.013128206,0.0,0.0,0.0032820515,0.02297436,0.0951795,0.24615386,0.48902568,0.27897438,0.13128206,0.06235898,0.06235898,0.10502565,0.21661541,0.22646156,0.17723078,0.38400003,1.4572309,1.7624617,1.6443079,1.1585642,0.65312827,0.764718,0.46933338,0.17066668,0.032820515,0.059076928,0.06564103,0.032820515,0.013128206,0.0032820515,0.006564103,0.01969231,0.01969231,0.016410258,0.009846155,0.07548718,0.37743592,1.0535386,0.8205129,0.4266667,0.21333335,0.13128206,0.101743594,0.118153855,0.17066668,0.30194873,0.5907693,1.1848207,1.6246156,1.9429746,2.0578463,1.7591796,1.3489232,0.7778462,0.38400003,0.23302566,0.1148718,0.15097436,0.190359,0.19364104,0.15753847,0.09189744,0.098461546,0.14769232,0.17723078,0.17394873,0.15097436,0.14112821,0.098461546,0.06564103,0.055794876,0.04266667,0.055794876,0.06235898,0.08205129,0.101743594,0.101743594,0.03938462,0.049230773,0.068923086,0.07876924,0.08861539,0.06564103,0.052512825,0.052512825,0.059076928,0.06235898,0.03938462,0.036102567,0.04266667,0.052512825,0.06564103,0.04594872,0.032820515,0.026256412,0.01969231,0.02297436,0.098461546,0.24287182,0.45292312,0.5677949,0.28225642,0.16738462,0.23630771,0.35446155,0.40369233,0.26912823,0.12471796,0.108307704,0.23302566,0.45292312,0.65969235,0.78769237,0.9616411,0.90256417,0.60061544,0.3117949,0.4135385,0.60061544,0.7089231,0.67610264,0.52512825,0.4004103,0.39056414,0.38728207,0.33805132,0.23958977,0.3249231,0.6235898,1.0502565,1.5524104,2.0939488,1.8018463,1.3817437,0.98133343,0.78769237,1.0338463,0.8533334,0.69907695,0.7187693,0.764718,0.4135385,0.3249231,0.4266667,0.5940513,0.6826667,0.54482055,0.35446155,0.21989745,0.14112821,0.2100513,0.5940513,1.014154,0.8960001,0.8566154,1.1027694,1.4441026,1.719795,2.2908719,3.1770258,4.2962055,5.4843082,4.9362054,4.0008206,3.1770258,2.6453335,2.284308,2.8192823,3.3312824,3.5905645,3.748103,4.3290257,6.370462,7.2369237,6.9120007,5.937231,5.4153852,5.730462,5.9536414,5.910975,5.6352825,5.3694363,5.290667,5.2315903,5.293949,5.4875903,5.737026,6.633026,7.9786673,10.581334,13.83713,15.721026,14.667488,11.503591,8.54318,6.7840004,5.8847184,5.408821,5.152821,4.8836927,4.716308,5.110154,6.675693,7.4732313,8.4283085,10.489437,14.608412,23.512617,26.574772,26.052925,23.69313,20.719591,18.481232,18.080822,18.28431,17.51631,13.856822,10.092308,6.701949,3.876103,1.8838975,1.0568206,0.7056411,0.5349744,0.4135385,0.32164106,0.36102566,0.34789747,0.2986667,0.26912823,0.28882053,0.3511795,0.55794877,0.8402052,1.0568206,1.1388719,1.1027694,0.94523084,0.7975385,0.65312827,0.5021539,0.33476925,0.13128206,0.04266667,0.01969231,0.029538464,0.04266667,0.068923086,0.09189744,0.101743594,0.0951795,0.07548718,0.08533334,0.098461546,0.12471796,0.17066668,0.256,0.37743592,0.5021539,0.62030774,0.67282057,0.574359,0.45292312,0.3511795,0.28882053,0.26256412,0.24615386,0.20348719,0.17066668,0.15097436,0.13784617,0.12143591,0.12143591,0.14441027,0.15753847,0.16082053,0.17394873,0.22646156,0.40369233,0.5284103,0.5481026,0.51856416,0.5513847,0.702359,0.8795898,0.9353847,0.6662565,0.3511795,0.28882053,0.380718,0.5513847,0.7581539,0.67282057,0.61374366,0.62030774,0.7220513,0.94523084,0.90584624,0.78769237,0.67282057,0.6859488,0.97805136,1.3357949,1.529436,1.4736412,1.2635899,1.1749744,1.1027694,1.2176411,1.3259488,1.394872,1.5458462,1.5753847,1.6049232,1.7887181,2.1169233,2.3860514,2.4484105,1.9922053,1.6607181,1.7099489,1.9790771,2.0939488,1.9068719,1.7001027,1.6344616,1.7558975,1.8707694,2.1924105,2.5074873,2.7011285,2.740513,2.03159,1.5655385,1.3062565,1.1979488,1.1651284,1.1716924,1.1158975,1.024,0.90256417,0.74830776,4.578462,4.8836927,5.976616,6.7807183,6.806975,6.1505647,6.4295387,7.817847,8.562873,7.8080006,5.5991797,4.391385,4.1813335,4.5587697,5.0051284,4.8836927,3.7842054,2.6847181,1.9035898,1.7099489,2.3204105,4.1747694,6.0652313,6.6100516,5.733744,4.6834874,4.5489235,4.9460516,5.76,6.9349747,8.4972315,11.270565,13.784616,13.453129,10.65354,8.713847,8.763078,8.113232,7.2960005,6.6527185,6.3474874,6.189949,6.5805135,7.1056414,7.4797955,7.5520005,7.7718983,7.5979495,6.921847,5.72718,4.1058464,3.249231,2.8816411,2.8882053,3.0720003,3.1573336,5.3431797,7.1548724,8.41518,8.320001,5.402257,2.861949,1.404718,1.0075898,1.214359,1.1290257,1.0075898,0.9682052,1.0043077,1.0666667,1.0666667,1.0568206,1.017436,1.1618463,1.4572309,1.6016412,1.3456411,1.3653334,1.6311796,2.1431797,2.8980515,4.010667,5.979898,7.6734366,8.395488,7.9195905,6.0750775,4.673641,3.5971284,3.1573336,4.073026,3.817026,3.4133337,2.9571285,2.7864618,3.495385,3.7874875,3.6594875,2.9702566,2.2383592,2.6387694,2.934154,2.7503593,2.3401027,1.847795,1.2964103,1.1881026,1.847795,2.2416413,2.0939488,1.8609232,1.6311796,1.3981539,1.3915899,1.6640002,2.0906668,2.1891284,2.048,1.8215386,1.5721027,1.2668719,0.7056411,0.41025645,0.3117949,0.33805132,0.4135385,0.3511795,0.30851284,0.30851284,0.34133336,0.36758977,0.34133336,0.36430773,0.42994875,0.47917953,0.380718,0.25928208,0.128,0.10502565,0.16738462,0.16738462,0.14441027,0.09189744,0.06235898,0.06235898,0.06235898,0.098461546,0.07876924,0.06235898,0.06564103,0.07548718,0.11158975,0.11158975,0.11158975,0.12471796,0.13784617,0.15097436,0.190359,0.21989745,0.23302566,0.24287182,0.28225642,0.28882053,0.27897438,0.26256412,0.27569234,0.22646156,0.19692309,0.17066668,0.13784617,0.07548718,0.17394873,0.41682056,0.827077,1.3193847,1.7099489,1.6344616,1.2340513,0.8008206,0.6498462,1.1126155,2.0545642,3.249231,6.009436,9.271795,9.613129,7.1483083,6.38359,5.4941545,3.9909747,2.7470772,2.8816411,2.7503593,2.546872,2.349949,2.1070771,1.4211283,0.93866676,0.7450257,0.9353847,1.6180514,1.5556924,1.3489232,1.0305642,0.6892308,0.45620516,0.4955898,0.48574364,0.3708718,0.17066668,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02297436,0.108307704,0.0951795,0.19364104,0.29538465,0.30194873,0.108307704,0.3511795,0.5415385,0.6498462,0.67610264,0.64000005,0.6662565,0.8008206,1.1060513,1.3620514,1.0666667,0.9714873,0.9747693,0.81394875,0.60389745,0.82379496,0.8467693,0.43323082,0.15425642,0.18707694,0.32164106,0.49230772,0.56123084,0.48246157,0.31507695,0.2297436,0.30194873,0.64000005,0.98133343,1.2340513,1.463795,1.6114873,1.2274873,0.71548724,0.32820517,0.16738462,0.2297436,0.25271797,0.29538465,0.39056414,0.5481026,0.108307704,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.016410258,0.016410258,0.009846155,0.0,0.0,0.0,0.0,0.006564103,0.016410258,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.013128206,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.006564103,0.006564103,0.072205134,0.3052308,0.37743592,0.3249231,0.19692309,0.10502565,0.21333335,0.38400003,0.380718,0.3708718,0.446359,0.64000005,0.85005134,0.90912825,1.3620514,2.2055387,2.9144619,1.1946667,0.36102566,0.098461546,0.11158975,0.13784617,0.07548718,0.04266667,0.02297436,0.01969231,0.029538464,0.029538464,0.02297436,0.009846155,0.0,0.0,0.4397949,0.71548724,0.78769237,0.65641034,0.3511795,0.4004103,0.38400003,0.26256412,0.15097436,0.33476925,0.46933338,0.48574364,0.6695385,1.2438976,2.3794873,3.1737437,2.2646155,1.1946667,0.6301539,0.33476925,0.3708718,0.3708718,0.3249231,0.23958977,0.15097436,0.09189744,0.12143591,0.15753847,0.15097436,0.09189744,0.07876924,0.06564103,0.055794876,0.04266667,0.029538464,0.04266667,0.036102567,0.02297436,0.016410258,0.016410258,0.0032820515,0.009846155,0.016410258,0.016410258,0.016410258,0.0032820515,0.0,0.01969231,0.049230773,0.06235898,0.049230773,0.01969231,0.0,0.0032820515,0.016410258,0.016410258,0.02297436,0.029538464,0.032820515,0.04594872,0.032820515,0.08533334,0.15097436,0.2100513,0.25928208,0.16082053,0.2297436,0.36430773,0.47589746,0.48902568,0.35446155,0.3117949,0.3249231,0.37743592,0.48902568,0.5481026,0.6465641,0.7384616,0.7253334,0.45620516,0.38400003,0.47589746,0.6826667,0.892718,0.9156924,0.8795898,0.8336411,0.6268718,0.31507695,0.16738462,0.20348719,0.52512825,0.9353847,1.3620514,1.8609232,2.0578463,1.9495386,1.657436,1.2307693,0.65641034,0.43651286,0.574359,0.7384616,0.69251287,0.28882053,0.19364104,0.23958977,0.31507695,0.3249231,0.2297436,0.108307704,0.07548718,0.101743594,0.27897438,0.8402052,1.1684103,1.142154,0.94523084,0.8467693,1.1749744,1.9200002,2.7175386,2.8488207,2.4451284,2.5173335,2.5173335,1.8937438,1.4244103,1.3587693,1.4178462,1.8838975,4.1878977,6.055385,7.174565,9.199591,10.226872,9.915077,8.631796,6.803693,4.9132314,5.7665644,6.669129,7.1876926,7.0531287,6.1505647,5.85518,5.8092313,5.927385,6.0783596,6.1046157,5.9930263,5.9667697,6.436103,7.906462,10.971898,10.689642,9.69518,8.602257,7.5552826,6.226052,5.211898,4.5029745,3.9876926,3.9286156,4.9296412,6.941539,9.028924,11.32636,14.546052,20.004105,24.582565,26.2039,26.134975,24.769644,21.622156,17.227488,16.587488,16.745028,15.835898,13.075693,10.121847,6.9776416,4.082872,1.9364104,1.0666667,0.82379496,0.7187693,0.571077,0.446359,0.64000005,0.7253334,0.7384616,0.6170257,0.4135385,0.28882053,0.3511795,0.45620516,0.58092314,0.69907695,0.80738467,0.80738467,0.7089231,0.4955898,0.23958977,0.09189744,0.04266667,0.029538464,0.04266667,0.06564103,0.09189744,0.128,0.17394873,0.19692309,0.18707694,0.13784617,0.13784617,0.15425642,0.18051283,0.21989745,0.3052308,0.4135385,0.48902568,0.512,0.48902568,0.4266667,0.318359,0.25271797,0.20348719,0.16082053,0.13784617,0.11158975,0.108307704,0.101743594,0.08533334,0.06235898,0.06235898,0.06235898,0.06235898,0.06564103,0.07548718,0.101743594,0.108307704,0.12471796,0.15425642,0.15425642,0.16410258,0.15097436,0.11158975,0.06564103,0.029538464,0.029538464,0.029538464,0.09189744,0.256,0.5481026,0.47589746,0.44964105,0.49887183,0.6170257,0.761436,0.8467693,0.8041026,0.7089231,0.6629744,0.80738467,0.9321026,0.9353847,0.92225647,1.0765129,1.6640002,1.8346668,1.4834872,1.1782565,1.142154,1.2504616,1.4572309,1.719795,1.9659488,2.2022567,2.5337439,2.5074873,2.1070771,1.6804104,1.4769232,1.6475899,1.8445129,1.8740515,1.7887181,1.7165129,1.8773335,1.8773335,2.0512822,2.4352822,2.789744,2.5928206,2.03159,1.7263591,1.6475899,1.654154,1.4966155,1.5688206,1.4966155,1.3718976,1.1881026,0.80738467,5.687795,6.560821,6.872616,7.062975,7.515898,8.5661545,9.304616,10.532104,10.617436,9.547488,8.920616,6.8430777,6.698667,7.752206,9.045334,9.409642,8.077128,7.0826674,6.482052,6.488616,7.4699492,8.018052,7.4207187,6.235898,5.0674877,4.57518,6.7840004,8.937026,10.390975,10.509129,8.681026,9.577026,10.84718,11.369026,11.109744,11.142565,11.113027,10.791386,9.777231,8.572719,8.582564,8.950154,9.133949,8.776206,7.9819493,7.3321033,6.567385,6.11118,5.408821,4.381539,3.4330258,3.9844105,4.1780515,4.269949,4.31918,4.2207184,6.1013336,6.875898,6.9776416,6.5411286,5.402257,3.5446157,2.2580514,1.5721027,1.3193847,1.1158975,0.955077,0.8467693,0.7975385,0.9419488,1.5556924,1.6902566,1.6508719,1.9035898,2.3893335,2.5042052,2.3171284,2.6518977,3.623385,5.037949,6.3901544,7.578257,7.6734366,6.810257,5.2578464,3.4166157,2.4516926,1.9987694,2.225231,3.2131286,4.9788723,6.0685134,6.11118,5.5762057,4.9132314,4.5554876,3.8432825,3.5741541,3.3903592,3.1770258,3.0424619,3.1803079,3.1245131,2.6880002,2.1858463,2.4549747,2.3762052,2.1333334,1.975795,1.9889232,2.1169233,2.0118976,1.4769232,1.214359,1.3423591,1.3718976,1.2438976,1.3259488,1.3883078,1.3489232,1.2800001,1.1651284,0.9321026,0.71548724,0.5907693,0.54482055,0.40697438,0.27897438,0.22646156,0.28882053,0.48902568,0.45292312,0.4135385,0.37743592,0.34789747,0.30851284,0.24615386,0.18707694,0.15753847,0.15097436,0.13128206,0.12471796,0.12471796,0.108307704,0.08205129,0.072205134,0.08205129,0.15097436,0.15097436,0.08533334,0.08861539,0.10502565,0.108307704,0.12143591,0.15097436,0.17394873,0.20676924,0.2297436,0.26256412,0.318359,0.37743592,0.33805132,0.3052308,0.28882053,0.28225642,0.27569234,0.24615386,0.2986667,0.41682056,0.5677949,0.7220513,1.2012309,1.723077,2.2613335,2.4320002,1.5130258,1.1093334,1.0043077,1.1651284,1.6377437,2.5435898,3.3444104,3.8465643,4.4832826,4.9854364,4.4012313,3.1376412,3.3050258,3.8367183,4.263385,4.6867695,5.35959,4.0008206,2.802872,2.6322052,3.0326157,1.8904617,1.2438976,1.1257436,1.585231,2.678154,1.9528207,1.4572309,1.1191796,0.8566154,0.5546667,0.5349744,0.62030774,0.7581539,0.69907695,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.036102567,0.1148718,0.256,0.49887183,0.5546667,0.5218462,0.4201026,0.28882053,0.18051283,0.101743594,0.108307704,0.36102566,0.6465641,0.39712822,0.380718,0.50543594,0.7450257,0.93866676,0.81066674,0.65641034,0.5415385,0.76800007,1.1716924,1.1158975,0.7220513,0.508718,0.46276927,0.5513847,0.73517954,0.92553854,0.7515898,0.56451285,0.48902568,0.42338464,0.4201026,0.512,0.58092314,0.57764107,0.52512825,0.4660513,0.36758977,0.26912823,0.17394873,0.032820515,0.04594872,0.049230773,0.17066668,0.30194873,0.108307704,0.02297436,0.029538464,0.029538464,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.016410258,0.016410258,0.006564103,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.006564103,0.006564103,0.0032820515,0.013128206,0.04266667,0.029538464,0.013128206,0.032820515,0.108307704,0.15425642,0.25271797,0.54482055,0.94523084,1.1520001,1.2077949,1.1684103,1.0929232,1.0962052,1.3620514,2.1267693,2.0184617,1.6672822,1.9954873,4.194462,2.2613335,0.77128214,0.10502565,0.108307704,0.11158975,0.08205129,0.055794876,0.036102567,0.029538464,0.04266667,0.04266667,0.03938462,0.029538464,0.009846155,0.0,0.128,0.2855385,0.45620516,0.56123084,0.4594872,0.2855385,0.16082053,0.0951795,0.0951795,0.190359,0.3511795,0.45620516,0.5546667,0.7450257,1.148718,1.8051283,1.8346668,1.6016412,1.2570257,0.7384616,0.6662565,0.52512825,0.3446154,0.18051283,0.10502565,0.101743594,0.13128206,0.15425642,0.14441027,0.10502565,0.08205129,0.06564103,0.049230773,0.032820515,0.029538464,0.032820515,0.02297436,0.026256412,0.03938462,0.03938462,0.016410258,0.013128206,0.016410258,0.016410258,0.016410258,0.0032820515,0.0,0.013128206,0.04266667,0.072205134,0.072205134,0.055794876,0.029538464,0.0,0.0032820515,0.0032820515,0.013128206,0.01969231,0.026256412,0.059076928,0.055794876,0.059076928,0.06235898,0.07548718,0.12471796,0.17394873,0.23302566,0.31507695,0.4004103,0.45292312,0.5316923,0.65312827,0.7778462,0.8402052,0.7450257,0.56123084,0.52512825,0.5907693,0.7056411,0.78769237,0.8992821,0.6859488,0.5316923,0.60389745,0.84348726,0.7187693,0.76800007,0.9156924,1.0929232,1.2307693,0.9944616,1.017436,1.1913847,1.394872,1.4966155,1.5064616,1.3522053,1.1454359,0.90256417,0.5349744,0.3446154,0.29210258,0.30851284,0.31507695,0.20348719,0.20348719,0.24943592,0.33476925,0.38400003,0.2297436,0.098461546,0.072205134,0.16082053,0.36102566,0.6695385,0.8795898,0.9124103,1.1224617,1.6180514,2.2613335,2.156308,2.0545642,2.2514873,2.9210258,4.1156926,3.5314875,2.8488207,2.1300514,1.5031796,1.1749744,1.2865642,2.1924105,3.3280003,4.4767184,5.7698464,7.4797955,8.717129,7.752206,5.225026,4.132103,4.128821,4.6605134,5.5302567,6.4065647,6.8332314,7.4469748,7.210667,6.8430777,6.626462,6.3967185,6.091488,5.540103,5.32677,5.861744,7.381334,8.635077,8.805744,8.914052,9.245539,9.350565,7.1154876,5.5138464,5.0149746,5.1626673,4.562052,5.8256416,8.815591,12.563693,16.498873,20.43077,24.549746,27.542976,28.504618,26.985027,22.977642,18.474669,16.656412,16.817232,17.414566,16.091898,11.907283,7.9130263,5.832206,5.428513,4.4734364,1.9626669,0.84348726,0.56451285,0.75487185,1.214359,1.2603078,1.0075898,0.65641034,0.36102566,0.2297436,0.20348719,0.26584616,0.34789747,0.39712822,0.3708718,0.32164106,0.24287182,0.14441027,0.049230773,0.01969231,0.009846155,0.013128206,0.026256412,0.04594872,0.07876924,0.10502565,0.128,0.13784617,0.13456412,0.12471796,0.14441027,0.15425642,0.15753847,0.16738462,0.18379489,0.21333335,0.23302566,0.23302566,0.21661541,0.19692309,0.16410258,0.14769232,0.12471796,0.09189744,0.07548718,0.06235898,0.049230773,0.04594872,0.04266667,0.036102567,0.04594872,0.055794876,0.06564103,0.08205129,0.12471796,0.17723078,0.2231795,0.23958977,0.2297436,0.190359,0.16082053,0.12143591,0.08205129,0.049230773,0.04266667,0.11158975,0.2100513,0.256,0.24287182,0.23302566,0.21661541,0.2855385,0.4266667,0.6104616,0.77456415,0.81066674,0.78769237,0.702359,0.6104616,0.60061544,0.67610264,0.7253334,0.81066674,1.0075898,1.4178462,2.0578463,2.2121027,1.6869745,0.892718,0.8369231,0.92553854,1.1881026,1.6377437,2.1366155,2.3860514,2.2547693,1.9462565,1.6508719,1.5064616,1.5983591,1.7263591,1.7460514,1.6902566,1.6246156,1.657436,1.7755898,2.0512822,2.2055387,2.1267693,1.8740515,1.595077,1.4572309,1.401436,1.3587693,1.2406155,1.0765129,0.9747693,0.90256417,0.83035904,0.73517954,8.054154,8.136206,8.339693,8.602257,8.523488,7.3485136,9.537642,11.405129,11.923694,11.0145645,9.567181,8.457847,8.933744,10.31877,11.631591,11.579078,11.175385,11.703795,11.395283,10.20718,9.829744,9.829744,8.743385,7.351795,6.3934364,6.550975,9.032206,10.834052,11.401847,10.469745,8.067283,8.87795,10.676514,12.386462,13.210258,12.629334,12.681848,12.714667,12.458668,11.808822,10.824206,10.066052,9.235693,8.192,7.0137444,6.0160003,5.149539,4.6080003,4.2830772,4.056616,3.7874875,4.066462,3.9581542,3.9876926,4.332308,4.8147697,6.160411,5.9569235,5.4613338,5.1331286,4.650667,2.674872,1.9922053,1.7394873,1.4506668,1.0601027,1.4802053,1.7558975,1.8904617,1.9593848,2.1267693,2.1300514,2.1136413,2.3335385,2.986667,4.2338467,3.9220517,3.43959,3.3312824,4.023795,5.8256416,6.564103,5.7534366,4.345436,2.9604106,1.9035898,1.8248206,2.3729234,3.2984617,4.5554876,6.2916927,8.283898,8.615385,7.9130263,6.7085133,5.425231,4.893539,4.466872,4.2174363,4.2305646,4.6080003,4.2141542,4.1813335,4.1452312,3.8104618,2.937436,2.609231,2.3630772,2.3696413,2.5206156,2.4484105,2.2219489,1.7887181,1.529436,1.4867693,1.3554872,1.1716924,1.1454359,1.1126155,1.0305642,0.9517949,0.892718,0.71548724,0.5218462,0.37415388,0.2855385,0.25928208,0.20348719,0.17723078,0.21661541,0.3446154,0.49887183,0.446359,0.32820517,0.26256412,0.35446155,0.26912823,0.24287182,0.25271797,0.25928208,0.21333335,0.20676924,0.20348719,0.18379489,0.15753847,0.15753847,0.15753847,0.18379489,0.16738462,0.118153855,0.118153855,0.13784617,0.18051283,0.20676924,0.20676924,0.2100513,0.21661541,0.21661541,0.23630771,0.27569234,0.32164106,0.27569234,0.26256412,0.30851284,0.4266667,0.60389745,0.8205129,1.1520001,1.5524104,1.9954873,2.4582565,2.28759,2.0709746,1.8707694,1.5753847,0.92553854,0.9124103,1.1552821,1.4211283,1.7985642,2.6880002,3.7284105,4.71959,4.9985647,4.6605134,4.5522056,4.263385,3.2328207,2.550154,2.605949,3.1048207,4.1058464,3.4034874,2.540308,2.1989746,2.166154,1.5261539,1.083077,1.0436924,1.5261539,2.5698464,1.5983591,1.0469744,0.79425645,0.67282057,0.45292312,0.26256412,0.26256412,0.44964105,0.571077,0.13784617,0.09189744,0.07548718,0.072205134,0.059076928,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0951795,0.18707694,0.27569234,0.47589746,0.31507695,0.24287182,0.29210258,0.42338464,0.5284103,0.40697438,0.30851284,0.41025645,0.65312827,0.7581539,0.8730257,0.9353847,1.0568206,1.2471796,1.4244103,1.4441026,1.1191796,1.0962052,1.3784616,1.3095386,0.9189744,0.6629744,0.56451285,0.60061544,0.702359,0.64000005,0.46276927,0.35774362,0.39056414,0.49230772,0.446359,0.4201026,0.39384618,0.36102566,0.3249231,0.24615386,0.19364104,0.13784617,0.07876924,0.04594872,0.009846155,0.0,0.055794876,0.11158975,0.0,0.0,0.013128206,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.006564103,0.006564103,0.0032820515,0.0,0.0,0.0,0.0,0.006564103,0.009846155,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.029538464,0.04594872,0.04594872,0.016410258,0.029538464,0.04266667,0.04594872,0.052512825,0.08861539,0.06564103,0.03938462,0.03938462,0.068923086,0.13456412,0.24943592,0.44307697,0.67610264,0.81066674,0.98133343,1.1355898,1.2964103,1.4834872,1.7066668,2.2580514,2.4155898,2.3302567,2.5271797,3.9023592,2.8816411,1.5031796,0.88287187,0.9189744,0.3249231,0.13456412,0.07876924,0.06235898,0.049230773,0.04594872,0.04594872,0.055794876,0.052512825,0.029538464,0.009846155,0.02297436,0.13128206,0.3511795,0.6268718,0.86317956,0.49887183,0.23630771,0.08861539,0.049230773,0.07876924,0.21333335,0.4004103,0.7318975,1.1027694,1.204513,1.3653334,1.4441026,1.4933335,1.4408206,1.0962052,0.84348726,0.54482055,0.28882053,0.13128206,0.072205134,0.108307704,0.17723078,0.20348719,0.16082053,0.08861539,0.08533334,0.072205134,0.055794876,0.04594872,0.03938462,0.026256412,0.016410258,0.02297436,0.036102567,0.026256412,0.009846155,0.013128206,0.016410258,0.013128206,0.006564103,0.0,0.0,0.0032820515,0.02297436,0.059076928,0.072205134,0.072205134,0.049230773,0.016410258,0.009846155,0.009846155,0.006564103,0.006564103,0.013128206,0.032820515,0.055794876,0.14112821,0.20020515,0.20676924,0.18379489,0.2100513,0.28225642,0.3446154,0.3708718,0.36102566,0.37743592,0.4660513,0.5874872,0.67938465,0.6432821,0.5907693,0.58420515,0.5973334,0.63343596,0.7220513,0.86646163,0.79425645,0.57764107,0.41025645,0.5874872,0.6071795,0.6235898,0.65969235,0.7811283,1.083077,1.3128207,1.6738462,2.041436,2.2646155,2.162872,1.8116925,1.3259488,0.90256417,0.6235898,0.47589746,0.30851284,0.20348719,0.16410258,0.18379489,0.256,0.54482055,0.65312827,0.5874872,0.4135385,0.256,0.15097436,0.11158975,0.16082053,0.27569234,0.38728207,0.5940513,0.82379496,1.0765129,1.3850257,1.8182565,1.9265642,1.8313848,2.15959,2.9144619,3.4822567,2.7864618,2.0841026,1.5195899,1.1716924,1.0666667,1.3128207,1.8084104,2.3762052,2.9013336,3.3378465,4.069744,5.4974365,6.226052,5.83877,4.9362054,4.2896414,3.9909747,4.273231,5.179077,6.564103,7.8834877,8.333129,9.130668,9.947898,8.923898,7.381334,5.8190775,5.0904617,5.398975,6.2916927,7.4732313,7.768616,8.096821,8.5891285,8.585847,7.4371285,6.7085133,6.3179493,5.930667,4.9296412,5.979898,9.429334,13.466257,17.24718,20.896822,25.911797,29.272617,29.705849,26.985027,21.943796,18.871796,17.178257,16.820515,16.810667,15.225437,11.529847,7.817847,5.428513,4.378257,3.367385,1.6443079,0.6826667,0.36758977,0.5415385,0.9911796,1.1454359,0.8008206,0.42338464,0.22646156,0.15753847,0.13128206,0.128,0.13456412,0.13456412,0.10502565,0.07876924,0.052512825,0.02297436,0.0,0.0,0.006564103,0.013128206,0.016410258,0.026256412,0.03938462,0.055794876,0.068923086,0.07876924,0.08861539,0.0951795,0.11158975,0.1148718,0.12471796,0.13128206,0.1148718,0.1148718,0.11158975,0.11158975,0.10502565,0.101743594,0.11158975,0.118153855,0.11158975,0.08861539,0.068923086,0.049230773,0.036102567,0.02297436,0.013128206,0.02297436,0.026256412,0.036102567,0.049230773,0.06564103,0.101743594,0.15425642,0.20020515,0.21661541,0.20676924,0.18051283,0.15097436,0.118153855,0.08861539,0.068923086,0.055794876,0.0951795,0.15753847,0.20020515,0.2100513,0.19692309,0.22646156,0.3249231,0.4660513,0.6104616,0.7220513,0.75487185,0.69251287,0.5874872,0.48574364,0.42994875,0.49887183,0.6104616,0.7122052,0.79425645,0.88287187,1.1716924,1.3161026,1.211077,0.9321026,0.76800007,0.88287187,1.1224617,1.522872,1.9232821,1.9922053,1.847795,1.6147693,1.4244103,1.3554872,1.4145643,1.4933335,1.5163078,1.4572309,1.3522053,1.3095386,1.3686155,1.522872,1.5786668,1.4966155,1.3718976,1.2964103,1.270154,1.2931283,1.339077,1.3686155,1.1618463,0.9517949,0.7844103,0.6826667,0.6432821,8.388924,8.12636,8.487385,8.536616,7.781744,6.183385,9.780514,11.52,11.995898,11.539693,10.213744,9.83959,10.043077,10.689642,11.369026,11.437949,10.59118,10.729027,10.118565,8.674462,7.9261546,7.8834877,7.3780518,6.7971287,6.698667,7.8047185,10.052924,11.661129,12.058257,11.418258,10.673231,11.72677,12.681848,13.312001,13.384206,12.645744,13.8075905,13.942155,13.610668,12.790154,10.873437,8.6580515,7.0137444,5.799385,4.9460516,4.4406157,3.7973337,3.4067695,3.3936412,3.6332312,3.7251284,3.6693337,3.5380516,3.7776413,4.309334,4.5029745,4.772103,4.06318,3.5282054,3.442872,3.1934361,1.8937438,1.8510771,2.1792822,2.3204105,2.028308,2.2088206,2.6387694,2.9604106,3.0293336,2.9210258,2.9702566,3.318154,3.8104618,4.5554876,5.924103,5.3398976,4.1911798,3.1113849,2.8488207,4.269949,4.46359,3.6069746,2.4681027,1.6771283,1.7099489,2.284308,3.308308,4.325744,5.2676926,6.4590774,8.1755905,8.792616,8.375795,7.2303596,5.8945646,5.4514875,5.031385,4.969026,5.405539,6.2752824,5.8453336,5.5236926,5.280821,4.8049235,3.4756925,3.0785644,2.8553848,2.809436,2.8291285,2.6912823,2.6026669,2.428718,2.2121027,2.0118976,1.9298463,1.7066668,1.4342566,1.1027694,0.78769237,0.67282057,0.58420515,0.4201026,0.27897438,0.20020515,0.14769232,0.18707694,0.20020515,0.190359,0.17394873,0.18051283,0.35774362,0.33805132,0.25928208,0.2297436,0.34789747,0.26256412,0.24615386,0.27241027,0.29210258,0.256,0.25271797,0.23958977,0.21333335,0.190359,0.20020515,0.21661541,0.21661541,0.19692309,0.17394873,0.18051283,0.21989745,0.3052308,0.32164106,0.26912823,0.24615386,0.256,0.26584616,0.28225642,0.30194873,0.30194873,0.24615386,0.28225642,0.45620516,0.7811283,1.2340513,1.7001027,2.1497438,2.5764105,2.9833848,3.373949,3.0982566,2.5140514,1.7296412,0.9616411,0.5415385,0.7515898,1.1651284,1.5622566,1.8740515,2.162872,3.5216413,5.477744,5.792821,4.706462,4.9329233,5.2381544,3.6463592,2.2547693,1.8970258,2.1202054,2.9571285,3.045744,2.6683078,2.044718,1.3554872,1.1388719,0.9682052,1.0404103,1.4539489,2.228513,1.2373334,0.6892308,0.47261542,0.4004103,0.23958977,0.049230773,0.0,0.13456412,0.2986667,0.13784617,0.09189744,0.07548718,0.072205134,0.059076928,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.032820515,0.036102567,0.006564103,0.0,0.0,0.03938462,0.190359,0.49230772,0.56451285,0.446359,0.33805132,0.5907693,0.48574364,0.40369233,0.32820517,0.40697438,0.9321026,1.2373334,1.4473847,1.4802053,1.4572309,1.7099489,1.8248206,1.723077,1.8248206,2.1202054,2.1530259,1.7165129,1.2471796,1.083077,1.2077949,1.2537436,1.014154,0.5973334,0.3511795,0.35446155,0.4135385,0.31507695,0.23302566,0.20348719,0.256,0.42338464,0.34789747,0.28882053,0.26256412,0.28882053,0.380718,0.3249231,0.2231795,0.10502565,0.02297436,0.04594872,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.006564103,0.016410258,0.01969231,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.01969231,0.009846155,0.0,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.009846155,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.036102567,0.068923086,0.08861539,0.068923086,0.07548718,0.08533334,0.08205129,0.08861539,0.14112821,0.13128206,0.09189744,0.07548718,0.17394873,0.2100513,0.2100513,0.2297436,0.318359,0.4955898,0.8402052,1.2537436,1.6377437,1.9429746,2.176,2.487795,2.6551797,2.8225644,3.0916924,3.5249233,2.8816411,3.3050258,3.8301542,3.3575387,0.6301539,0.21333335,0.118153855,0.128,0.12143591,0.068923086,0.055794876,0.055794876,0.049230773,0.032820515,0.009846155,0.0032820515,0.108307704,0.44964105,0.9353847,1.2537436,0.8992821,0.5284103,0.24615386,0.098461546,0.049230773,0.12471796,0.28225642,0.64000005,1.2438976,2.0545642,4.1714873,3.5478978,2.425436,1.8937438,1.8707694,1.1585642,0.6268718,0.29210258,0.13784617,0.108307704,0.2231795,0.31507695,0.32164106,0.23302566,0.108307704,0.08533334,0.068923086,0.059076928,0.052512825,0.04594872,0.029538464,0.01969231,0.01969231,0.02297436,0.016410258,0.0032820515,0.009846155,0.013128206,0.006564103,0.0,0.0,0.0032820515,0.006564103,0.013128206,0.032820515,0.04266667,0.04594872,0.036102567,0.016410258,0.009846155,0.029538464,0.032820515,0.026256412,0.01969231,0.02297436,0.049230773,0.14769232,0.2297436,0.25271797,0.20676924,0.2100513,0.27897438,0.31507695,0.29538465,0.26912823,0.25271797,0.29538465,0.37743592,0.4660513,0.49230772,0.50543594,0.5349744,0.5284103,0.49230772,0.49230772,0.5677949,0.60061544,0.48246157,0.3052308,0.38400003,0.5152821,0.57764107,0.6170257,0.7056411,0.9485129,1.6475899,2.3302567,2.7700515,2.8455386,2.5173335,1.9561027,1.3292309,0.9189744,0.761436,0.64000005,0.41025645,0.2855385,0.24287182,0.2986667,0.53825647,1.0699488,1.0601027,0.76800007,0.43323082,0.26912823,0.21333335,0.18707694,0.21333335,0.29210258,0.36758977,0.5513847,1.0010257,1.4375386,1.6672822,1.5819489,2.2744617,2.740513,3.2164104,3.5544617,3.2262566,2.409026,1.6147693,1.404718,1.654154,1.5688206,1.6082052,1.910154,2.0611284,1.9954873,1.9790771,2.1103592,3.0227695,4.266667,5.1659493,4.8016415,4.325744,3.7776413,3.6430771,4.240411,5.717334,8.231385,9.058462,9.577026,9.9282055,8.986258,7.210667,5.6320004,4.926359,5.3070774,6.5378466,7.1680007,7.0957956,7.1581545,7.4075904,7.1187696,7.177847,7.7325134,8.027898,7.860513,7.5585647,8.493949,10.889847,13.761642,16.918976,20.955898,27.825233,31.593027,31.757132,28.612925,23.273027,21.943796,20.676924,19.48554,17.91672,15.041642,11.221334,7.716103,5.093744,3.4166157,2.2416413,1.4211283,0.7844103,0.446359,0.45620516,0.81394875,0.94523084,0.54482055,0.2100513,0.13456412,0.1148718,0.1148718,0.072205134,0.032820515,0.013128206,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0,0.013128206,0.016410258,0.016410258,0.013128206,0.009846155,0.016410258,0.02297436,0.029538464,0.04266667,0.06564103,0.08205129,0.08861539,0.08861539,0.08205129,0.072205134,0.06564103,0.06564103,0.06564103,0.06564103,0.07548718,0.10502565,0.11158975,0.10502565,0.098461546,0.08205129,0.06235898,0.04594872,0.026256412,0.013128206,0.016410258,0.009846155,0.013128206,0.02297436,0.032820515,0.059076928,0.09189744,0.12471796,0.15097436,0.17066668,0.18707694,0.190359,0.19364104,0.20020515,0.2231795,0.256,0.32164106,0.39384618,0.47917953,0.571077,0.636718,0.6826667,0.7220513,0.7450257,0.7515898,0.761436,0.78769237,0.7089231,0.58092314,0.44964105,0.3446154,0.38400003,0.47589746,0.5349744,0.5284103,0.45620516,0.4594872,0.5152821,0.6892308,0.8763078,0.77456415,0.96492314,1.2340513,1.5819489,1.8576412,1.7657437,1.5983591,1.3915899,1.2438976,1.1848207,1.1815386,1.2077949,1.2471796,1.2209232,1.142154,1.0765129,1.0535386,1.0896411,1.1257436,1.1355898,1.142154,1.1520001,1.1881026,1.2307693,1.2603078,1.2504616,1.1158975,0.9419488,0.79425645,0.6859488,0.6071795,7.269744,7.834257,8.684308,8.533334,7.532308,7.269744,10.312206,10.627283,10.187488,9.977437,9.987283,9.586872,8.917334,8.470975,8.556309,9.301334,7.177847,5.481026,4.348718,3.8367183,3.9286156,4.2371287,4.5817437,5.0018463,5.7665644,7.384616,9.747693,12.081232,13.610668,14.401642,15.37313,15.91795,14.70359,12.832822,11.385437,11.418258,13.528616,13.46954,12.2847185,10.594462,8.595693,5.868308,4.138667,3.2361028,3.0326157,3.4297438,3.121231,2.8389745,2.7503593,2.868513,3.0358977,3.2000003,3.4231799,3.8728209,4.1583595,3.308308,2.7076926,2.172718,1.9429746,1.9593848,1.8543591,1.8445129,2.0841026,2.5895386,3.1376412,3.255795,2.8160002,3.2787695,3.882667,4.1846156,4.0467696,3.9548721,4.5456414,5.2644105,5.792821,6.048821,5.362872,4.420923,3.3641028,2.6026669,2.7995899,2.7733335,2.4352822,1.8149745,1.3718976,1.9790771,3.0851285,4.2240005,5.113436,5.609026,5.7074876,6.091488,6.803693,7.2894363,7.2205133,6.521436,5.8814363,5.7140517,5.910975,6.377026,7.0498466,7.072821,6.4623594,5.58277,4.706462,4.0041027,3.7874875,3.43959,3.0851285,2.865231,2.930872,3.1409233,3.1770258,2.9669745,2.6256413,2.4451284,2.1792822,1.8018463,1.3456411,0.92553854,0.75487185,0.60389745,0.37743592,0.24615386,0.24287182,0.28225642,0.2986667,0.2855385,0.24943592,0.19364104,0.13128206,0.13784617,0.17394873,0.21989745,0.256,0.28225642,0.26256412,0.24615386,0.24615386,0.25271797,0.26256412,0.28225642,0.26912823,0.23630771,0.20348719,0.19692309,0.21333335,0.24287182,0.27241027,0.28882053,0.2855385,0.3249231,0.39712822,0.39384618,0.32164106,0.30194873,0.34133336,0.38728207,0.43323082,0.4660513,0.4660513,0.43651286,0.5874872,0.92225647,1.4211283,2.0578463,2.7208207,2.9965131,3.0490258,2.989949,2.8750772,3.249231,2.9702566,2.1530259,1.1323078,0.47917953,0.5316923,0.955077,1.7033848,2.2777438,1.7033848,2.92759,5.2315903,5.6385646,4.2535386,4.276513,4.5456414,3.5216413,2.6518977,2.4615386,2.553436,2.8849232,3.1573336,2.937436,2.1792822,1.214359,1.0305642,1.0108719,1.1388719,1.401436,1.7887181,0.94523084,0.47589746,0.26584616,0.18051283,0.06564103,0.013128206,0.0,0.068923086,0.15097436,0.059076928,0.049230773,0.01969231,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.01969231,0.04266667,0.072205134,0.072205134,0.052512825,0.04266667,0.036102567,0.098461546,0.37743592,1.1290257,1.2471796,1.0075898,0.7778462,1.017436,1.1618463,1.1290257,0.8566154,0.69579494,1.394872,2.0939488,2.7109745,2.9046156,2.7437952,2.6912823,2.487795,2.2088206,2.3105643,2.5764105,2.1464617,1.083077,0.6859488,0.65312827,0.76800007,0.8795898,0.8041026,0.33805132,0.036102567,0.04594872,0.13456412,0.2100513,0.2100513,0.17394873,0.16410258,0.28225642,0.20020515,0.14112821,0.12471796,0.190359,0.3708718,0.32820517,0.19364104,0.06564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.013128206,0.032820515,0.036102567,0.02297436,0.0,0.0,0.0,0.006564103,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.029538464,0.036102567,0.02297436,0.0032820515,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.032820515,0.072205134,0.098461546,0.108307704,0.10502565,0.09189744,0.07876924,0.09189744,0.15097436,0.16410258,0.17394873,0.23630771,0.4397949,0.35446155,0.21661541,0.20348719,0.380718,0.7056411,1.0666667,1.5589745,2.0053334,2.3991797,2.9046156,3.1967182,3.1507695,3.2525132,3.5052311,3.4100516,2.425436,4.640821,6.373744,5.4416413,1.1520001,0.47917953,0.22646156,0.190359,0.20020515,0.108307704,0.068923086,0.03938462,0.026256412,0.02297436,0.0,0.0,0.0951795,0.5677949,1.2504616,1.5195899,1.1913847,0.8402052,0.5546667,0.34789747,0.17723078,0.15097436,0.16738462,0.28225642,0.84348726,2.4976413,6.9382567,5.7435904,3.3772311,2.1858463,2.4024618,1.3686155,0.69579494,0.32164106,0.17066668,0.17723078,0.36758977,0.48246157,0.46276927,0.3249231,0.15097436,0.08861539,0.068923086,0.059076928,0.049230773,0.04594872,0.049230773,0.032820515,0.02297436,0.01969231,0.01969231,0.006564103,0.009846155,0.006564103,0.0,0.0,0.0032820515,0.016410258,0.029538464,0.036102567,0.02297436,0.0032820515,0.0032820515,0.0032820515,0.0,0.0,0.03938462,0.059076928,0.055794876,0.04594872,0.04266667,0.06235898,0.08861539,0.118153855,0.14769232,0.15097436,0.17394873,0.2100513,0.2100513,0.18707694,0.24287182,0.30194873,0.34789747,0.37743592,0.4004103,0.4397949,0.38728207,0.40697438,0.41682056,0.38728207,0.3249231,0.3117949,0.27569234,0.25928208,0.28225642,0.35446155,0.508718,0.75487185,0.97805136,1.1224617,1.1618463,2.028308,2.7109745,2.9505644,2.6945643,2.1103592,1.5556924,1.1585642,1.1191796,1.2603078,1.0436924,0.65312827,0.44964105,0.38400003,0.49887183,0.92225647,1.5688206,1.4441026,1.017436,0.6071795,0.40369233,0.40369233,0.45292312,0.512,0.5874872,0.71548724,0.85005134,1.339077,2.038154,2.5796926,2.3663592,3.7120004,4.824616,5.366154,5.172513,4.263385,3.1048207,2.15959,2.1070771,2.5993848,2.2646155,1.9626669,2.1169233,2.1497438,1.972513,1.9790771,2.2383592,2.409026,2.7700515,3.2656412,3.4921029,3.511795,3.4494362,3.6627696,4.273231,5.156103,8.503796,8.937026,7.8736415,6.665847,6.6100516,5.8945646,5.3136415,5.0215387,5.353026,6.8365135,7.131898,6.813539,6.616616,6.701949,6.6461544,7.243488,8.553026,9.498257,9.882257,10.381129,11.142565,11.818667,13.078976,15.619284,20.161642,28.425848,33.29313,34.425438,32.15754,27.477335,26.177643,24.74995,22.741335,19.820309,15.78995,11.444513,8.011488,5.5630774,3.8629746,2.3696413,1.6771283,1.214359,0.90912825,0.78769237,0.93866676,0.83035904,0.39384618,0.12143591,0.118153855,0.108307704,0.1148718,0.07548718,0.036102567,0.013128206,0.0,0.0,0.006564103,0.006564103,0.0,0.0,0.009846155,0.013128206,0.013128206,0.009846155,0.0,0.0,0.0,0.0,0.009846155,0.03938462,0.06235898,0.07548718,0.06235898,0.036102567,0.04266667,0.049230773,0.052512825,0.052512825,0.052512825,0.072205134,0.101743594,0.09189744,0.07876924,0.07876924,0.07548718,0.068923086,0.055794876,0.03938462,0.029538464,0.01969231,0.009846155,0.006564103,0.006564103,0.009846155,0.029538464,0.04266667,0.068923086,0.1148718,0.17723078,0.25928208,0.32164106,0.3708718,0.42338464,0.5021539,0.6301539,0.77128214,0.9156924,1.0568206,1.1913847,1.2865642,1.3161026,1.2603078,1.1355898,0.98461545,0.88943595,0.8795898,0.81066674,0.6662565,0.47917953,0.318359,0.3052308,0.3117949,0.32164106,0.32164106,0.2986667,0.35774362,0.4135385,0.53825647,0.7056411,0.77128214,1.020718,1.3357949,1.6640002,1.8576412,1.6705642,1.467077,1.2996924,1.2012309,1.1454359,1.0601027,1.0108719,1.0305642,1.0469744,1.0305642,0.98461545,0.93866676,0.96492314,1.0338463,1.1191796,1.1848207,1.1881026,1.1979488,1.1585642,1.0371283,0.8402052,0.79425645,0.7844103,0.7778462,0.7384616,0.64000005,9.124104,11.369026,13.571283,14.815181,14.299898,11.323078,9.015796,7.1581545,5.691077,4.713026,4.457026,4.309334,4.1452312,4.457026,5.1889234,5.737026,5.1265645,4.453744,3.9876926,3.7809234,3.6463592,4.7589746,5.5302567,5.986462,6.189949,6.226052,9.143796,12.373334,15.300924,16.938667,15.898257,14.470565,13.033027,11.539693,10.282667,9.90195,9.573745,9.225847,8.303591,6.9382567,5.937231,4.8377438,3.8301542,3.3280003,3.4067695,3.7842054,4.0533338,3.2689233,2.537026,2.3762052,2.7306669,3.3050258,3.2918978,2.986667,2.4910772,1.7099489,2.2711797,2.5764105,2.550154,2.3302567,2.2580514,2.15959,1.9429746,1.6935385,1.6311796,2.1202054,3.0490258,4.3060517,5.717334,6.560821,5.586052,3.9614363,3.4264617,3.1573336,2.789744,2.412308,2.3991797,2.678154,2.5337439,1.723077,0.5021539,1.017436,1.273436,1.4506668,1.8051283,2.6847181,4.663795,6.419693,7.762052,8.024616,6.0717955,5.0116925,5.093744,6.875898,9.084719,8.621949,8.402052,8.713847,8.027898,6.51159,6.012718,6.0717955,6.0160003,5.4580517,4.493129,3.6627696,3.564308,3.4592824,3.3903592,3.3936412,3.4789746,3.4658465,3.4822567,3.3345644,2.8225644,1.723077,1.5163078,1.529436,1.7296412,1.8642052,1.4506668,0.98461545,0.5940513,0.3708718,0.3446154,0.5021539,0.5284103,0.37743592,0.2855385,0.28882053,0.2297436,0.16738462,0.25271797,0.3249231,0.3314872,0.32164106,0.40697438,0.380718,0.3446154,0.34789747,0.39712822,0.446359,0.4397949,0.39712822,0.32820517,0.24287182,0.19692309,0.2297436,0.3708718,0.51856416,0.45620516,0.39712822,0.33476925,0.3249231,0.36430773,0.4135385,0.4594872,0.49887183,0.5874872,0.7220513,0.86974365,1.0535386,1.4998976,1.972513,2.3991797,2.8980515,3.826872,3.692308,3.0752823,2.349949,1.6771283,2.2777438,2.2153847,1.6902566,0.9682052,0.380718,0.35774362,0.892718,2.0742567,3.0818465,2.166154,2.03159,2.5862565,3.8367183,5.142975,5.2020516,4.457026,3.3575387,2.4976413,2.0775387,1.9068719,1.9922053,2.0873847,1.972513,1.6049232,1.1290257,0.98133343,0.90912825,0.84348726,0.7384616,0.58092314,0.1148718,0.0,0.0,0.029538464,0.15097436,0.029538464,0.0,0.055794876,0.16738462,0.28882053,0.23958977,0.09189744,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.072205134,0.101743594,0.08861539,0.049230773,0.0,0.18379489,0.2100513,0.17394873,0.108307704,0.0,0.7318975,1.3653334,1.847795,2.0053334,1.5425643,1.4441026,1.6114873,2.0873847,2.5173335,2.1530259,1.9922053,2.172718,2.6847181,3.1081028,2.5928206,1.6672822,1.4441026,1.2373334,0.827077,0.47261542,0.38728207,0.40369233,0.39056414,0.3052308,0.18379489,0.29210258,0.256,0.17723078,0.13456412,0.18379489,0.17066668,0.15097436,0.08205129,0.03938462,0.19692309,0.17394873,0.11158975,0.04594872,0.026256412,0.13784617,0.12471796,0.049230773,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.036102567,0.036102567,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02297436,0.049230773,0.098461546,0.13456412,0.06235898,0.013128206,0.01969231,0.02297436,0.01969231,0.029538464,0.029538464,0.029538464,0.29210258,0.7318975,0.9156924,0.63343596,0.5284103,0.6071795,0.8402052,1.1454359,1.0962052,1.1552821,1.5360001,2.356513,3.6627696,3.892513,4.161641,4.3651285,4.1156926,2.7634873,1.9922053,1.6902566,1.9396925,2.3958976,2.2744617,1.2603078,0.5021539,0.15425642,0.13128206,0.108307704,0.059076928,0.026256412,0.016410258,0.013128206,0.0,0.0,0.0,0.34133336,1.0305642,1.7394873,0.9353847,0.85005134,0.9747693,0.94523084,0.58092314,0.34789747,0.22646156,0.21333335,0.33476925,0.64000005,0.77456415,0.79097444,0.74830776,0.7417436,0.8992821,0.7187693,0.39712822,0.17723078,0.128,0.15097436,0.27569234,0.49887183,0.5218462,0.3249231,0.15097436,0.128,0.0951795,0.068923086,0.059076928,0.04594872,0.059076928,0.06235898,0.055794876,0.04266667,0.029538464,0.01969231,0.006564103,0.0,0.0,0.0,0.013128206,0.04266667,0.09189744,0.12143591,0.06235898,0.013128206,0.009846155,0.009846155,0.0,0.0,0.0,0.009846155,0.026256412,0.055794876,0.09189744,0.14112821,0.14441027,0.13128206,0.128,0.15097436,0.16410258,0.14112821,0.128,0.18379489,0.36758977,0.46276927,0.48902568,0.4135385,0.34133336,0.48902568,0.52512825,0.54482055,0.5481026,0.5349744,0.47261542,0.44964105,0.36102566,0.29210258,0.318359,0.48902568,0.7811283,1.2209232,1.3686155,1.211077,1.1749744,2.041436,2.422154,2.4155898,2.0709746,1.3883078,0.86317956,0.9517949,1.3357949,1.6672822,1.5556924,0.9714873,0.5481026,0.34789747,0.46933338,1.0666667,1.7624617,2.156308,1.8937438,1.2209232,0.97805136,1.0371283,1.2438976,1.3259488,1.2504616,1.2504616,1.4473847,1.5327181,1.9298463,2.806154,4.073026,6.2227697,7.4929237,7.8506675,7.2894363,5.8125134,4.1780515,3.117949,2.4352822,2.0217438,1.8609232,2.3138463,2.793026,3.2984617,3.7251284,3.8596926,3.5905645,3.1409233,3.31159,3.7710772,3.0523078,2.3302567,2.7569232,4.141949,5.7435904,6.2555904,7.6603084,7.197539,6.5870776,6.5017443,6.560821,6.744616,6.7249236,6.5739493,6.2851286,5.799385,6.2490263,6.4557953,6.5017443,6.6592827,7.3550773,8.441437,9.45559,9.29477,8.198565,7.722667,8.4053335,9.426052,10.916103,13.446565,18.034874,24.786053,31.727592,35.232822,34.349953,30.821747,24.999386,22.06195,19.705437,16.804104,13.397334,10.906258,8.516924,6.088206,3.7251284,1.785436,1.6377437,1.5392822,1.5130258,1.4408206,1.0371283,0.5874872,0.21661541,0.07548718,0.118153855,0.108307704,0.0951795,0.072205134,0.04266667,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.016410258,0.016410258,0.026256412,0.03938462,0.04594872,0.04266667,0.029538464,0.055794876,0.07876924,0.07876924,0.06235898,0.06235898,0.06235898,0.04266667,0.029538464,0.026256412,0.016410258,0.026256412,0.03938462,0.04594872,0.04266667,0.029538464,0.029538464,0.03938462,0.03938462,0.029538464,0.029538464,0.04266667,0.09189744,0.17066668,0.28225642,0.44307697,0.5513847,0.6432821,0.7187693,0.8008206,0.94523084,1.079795,1.204513,1.3095386,1.3850257,1.4342566,1.4211283,1.3718976,1.2635899,1.1093334,0.9616411,0.8763078,0.77128214,0.5874872,0.36758977,0.24287182,0.23302566,0.24615386,0.27241027,0.2986667,0.33476925,0.43323082,0.512,0.63343596,0.7844103,0.86974365,1.0896411,1.3357949,1.4900514,1.4605129,1.204513,1.0699488,1.1191796,1.2537436,1.3522053,1.2668719,1.1191796,0.98133343,0.8960001,0.86317956,0.8402052,0.85005134,0.9288206,1.1060513,1.3292309,1.463795,1.4408206,1.2603078,1.0272821,0.81394875,0.65641034,0.62030774,0.6301539,0.6662565,0.702359,0.702359,7.90318,8.910769,10.610872,11.9860525,12.2847185,11.004719,9.780514,8.822155,7.4075904,5.799385,5.2611284,5.3103595,4.6802053,3.876103,3.4822567,4.1878977,4.466872,4.269949,3.9909747,3.8400004,3.8432825,4.1222568,4.460308,4.6539493,4.890257,5.737026,8.254359,10.095591,11.027693,10.981745,10.052924,10.325335,9.750975,9.074872,8.710565,8.743385,8.054154,7.2927184,6.38359,5.5958977,5.533539,5.536821,5.3858466,5.172513,5.0576415,5.2480006,4.7950773,3.9548721,3.692308,4.1189747,4.4996924,4.5489235,4.309334,3.636513,2.6617439,1.782154,2.1398976,2.3105643,2.297436,2.1497438,1.9790771,1.7723079,1.5425643,1.3850257,1.404718,1.719795,2.2547693,2.8816411,3.4494362,3.6857438,3.1671798,2.8127182,2.7076926,2.5173335,2.166154,1.8379488,1.6311796,1.6640002,1.5524104,1.1881026,0.74830776,0.8205129,0.8566154,0.96492314,1.2635899,1.8806155,3.446154,4.6867695,5.533539,5.7403083,4.850872,4.785231,4.9493337,5.540103,6.117744,5.5926156,5.7829747,6.2785645,6.698667,6.7774363,6.36718,5.8518977,5.333334,5.179077,5.0182567,3.761231,2.5206156,2.5961027,2.9243078,3.1015387,3.3936412,3.6660516,3.1803079,2.4582565,1.7920002,1.2603078,1.5524104,1.5327181,1.3686155,1.1552821,0.92553854,0.764718,0.54482055,0.2986667,0.1148718,0.13784617,0.16082053,0.16738462,0.23630771,0.38400003,0.54482055,0.60389745,0.51856416,0.4594872,0.46276927,0.42994875,0.34133336,0.36758977,0.36430773,0.28882053,0.20020515,0.21989745,0.43323082,0.64000005,0.67938465,0.4266667,0.29210258,0.26584616,0.3314872,0.42994875,0.446359,0.45292312,0.52512825,0.72861546,1.014154,1.2176411,1.3751796,1.4769232,1.5721027,1.7099489,1.9429746,2.2449234,2.5698464,2.9210258,3.242667,3.4133337,3.3247182,2.9571285,2.6157951,2.4484105,2.4713848,3.0884104,3.1573336,2.9243078,2.6322052,2.5042052,2.3040001,2.3105643,2.5698464,2.9210258,3.0227695,2.9078977,2.9669745,3.698872,4.598154,4.141949,3.4166157,3.0293336,2.8980515,2.802872,2.409026,1.6836925,1.6705642,1.5622566,1.1060513,0.5907693,0.7187693,0.7581539,0.7056411,0.5513847,0.27569234,0.26912823,0.2231795,0.20020515,0.22646156,0.2986667,0.23630771,0.17723078,0.098461546,0.07876924,0.27897438,0.3249231,0.25271797,0.118153855,0.0,0.0,0.128,0.14441027,0.108307704,0.059076928,0.0,0.013128206,0.101743594,0.17723078,0.2100513,0.21989745,0.2855385,0.34133336,0.41682056,0.5481026,0.76800007,1.5885129,2.0217438,2.0086155,1.657436,1.273436,1.2537436,1.3751796,1.5327181,1.6344616,1.5885129,1.5589745,1.5655385,1.6475899,1.7066668,1.4966155,1.1158975,1.014154,0.99774367,0.94523084,0.827077,0.47917953,0.20676924,0.07876924,0.06235898,0.036102567,0.28225642,0.318359,0.2231795,0.118153855,0.15753847,0.059076928,0.029538464,0.016410258,0.006564103,0.03938462,0.036102567,0.02297436,0.009846155,0.006564103,0.026256412,0.026256412,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.0032820515,0.0,0.0,0.02297436,0.049230773,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.016410258,0.029538464,0.08205129,0.15097436,0.14769232,0.118153855,0.068923086,0.052512825,0.0951795,0.22646156,0.4004103,0.39384618,0.45620516,0.67610264,0.97805136,0.93866676,0.84348726,0.8730257,1.2307693,2.1333334,1.7526156,1.4900514,1.6607181,2.1267693,2.2711797,2.4648206,2.6420515,2.9636924,3.2951798,3.190154,3.0162053,2.4746668,2.0512822,1.9232821,1.9692309,2.1366155,1.1027694,0.30194873,0.15097436,0.059076928,0.049230773,0.036102567,0.026256412,0.02297436,0.013128206,0.0032820515,0.052512825,0.2855385,0.7253334,1.2865642,1.1355898,1.3062565,1.5458462,1.5360001,0.88615394,0.47589746,0.47261542,0.44964105,0.31507695,0.2855385,0.380718,0.5349744,0.6235898,0.63343596,0.65641034,0.5218462,0.33805132,0.22646156,0.25271797,0.43323082,0.380718,0.3314872,0.26912823,0.20348719,0.190359,0.20348719,0.20348719,0.16738462,0.12143591,0.118153855,0.24943592,0.43323082,0.4004103,0.16082053,0.04266667,0.029538464,0.009846155,0.0032820515,0.009846155,0.0,0.0032820515,0.009846155,0.01969231,0.02297436,0.013128206,0.0032820515,0.0032820515,0.006564103,0.013128206,0.013128206,0.0032820515,0.009846155,0.026256412,0.06564103,0.14112821,0.2100513,0.2231795,0.21661541,0.21333335,0.23958977,0.2100513,0.14112821,0.098461546,0.11158975,0.15753847,0.22646156,0.21333335,0.190359,0.20348719,0.29210258,0.38728207,0.3708718,0.32164106,0.30194873,0.33805132,0.42338464,0.4266667,0.38400003,0.4201026,0.7581539,1.273436,1.9593848,2.8882053,3.5807183,3.006359,2.3105643,1.9922053,1.7329233,1.4441026,1.2800001,1.5163078,1.9692309,2.2088206,2.03159,1.4834872,0.9353847,0.5481026,0.39056414,0.54482055,1.0929232,1.8281027,1.9593848,1.6935385,1.2537436,0.90256417,1.1290257,1.4441026,1.591795,1.5819489,1.6902566,2.169436,3.249231,4.273231,5.044513,5.796103,7.00718,7.4043083,6.7840004,5.467898,4.325744,4.240411,3.6890259,3.3411283,3.4198978,3.692308,3.4034874,3.0358977,2.8980515,3.0687182,3.4100516,2.858667,2.422154,2.2744617,2.3302567,2.2350771,2.169436,3.1015387,5.179077,7.2237954,6.7183595,6.3376417,5.8223596,5.874872,6.2851286,5.927385,5.5729237,5.98318,6.5050263,6.813539,6.921847,7.24677,7.381334,7.712821,8.169026,8.2215395,8.116513,8.218257,8.1755905,8.064001,8.379078,8.274052,8.109949,8.602257,10.410667,14.129231,19.951591,25.790361,31.215591,35.14749,35.876106,31.996721,26.840618,21.546669,16.981335,13.751796,11.349334,8.418462,5.7107697,3.6594875,2.3827693,1.847795,1.4572309,1.0666667,0.67282057,0.4135385,0.23630771,0.098461546,0.04594872,0.06235898,0.068923086,0.068923086,0.06235898,0.055794876,0.04594872,0.02297436,0.02297436,0.016410258,0.013128206,0.009846155,0.0,0.0,0.006564103,0.013128206,0.009846155,0.0,0.0,0.006564103,0.029538464,0.072205134,0.16082053,0.28225642,0.32820517,0.3249231,0.27569234,0.17723078,0.17066668,0.1148718,0.08205129,0.08205129,0.072205134,0.052512825,0.03938462,0.026256412,0.01969231,0.026256412,0.03938462,0.13128206,0.17723078,0.13456412,0.055794876,0.06564103,0.09189744,0.1148718,0.128,0.128,0.15097436,0.2231795,0.3511795,0.51856416,0.6859488,0.7581539,0.7450257,0.72861546,0.7811283,0.95835906,1.142154,1.3226668,1.4703591,1.5819489,1.6902566,1.7362052,1.7460514,1.6968206,1.595077,1.4998976,1.4900514,1.2537436,0.98133343,0.7318975,0.4135385,0.42338464,0.48574364,0.574359,0.65312827,0.6892308,0.7089231,0.7253334,0.7844103,0.8763078,0.9419488,1.142154,1.3718976,1.4736412,1.3850257,1.1191796,1.0633847,1.4178462,1.9561027,2.300718,1.913436,1.3751796,1.1618463,1.0568206,0.9747693,0.9485129,1.020718,0.90584624,0.79097444,0.7581539,0.8041026,0.9485129,1.0371283,0.9714873,0.76800007,0.571077,0.52512825,0.56123084,0.6301539,0.7056411,0.761436,8.257642,8.910769,10.538668,12.219078,13.223386,13.02318,12.839386,14.221129,14.631386,13.397334,11.733335,9.882257,8.89436,7.958975,6.76759,5.4843082,4.460308,4.0303593,4.0041027,4.132103,4.1025643,3.817026,3.82359,4.135385,4.7261543,5.543385,6.810257,8.04759,8.920616,9.176616,8.644924,8.710565,8.684308,8.54318,8.4053335,8.553026,7.972103,7.2894363,6.892308,6.892308,7.0990777,6.764308,6.770872,6.7938466,6.5247183,5.651693,5.113436,4.9854364,5.3891287,5.7698464,4.906667,4.338872,3.9056413,3.0654361,2.0118976,1.6738462,2.0217438,2.1497438,2.1924105,2.1792822,2.034872,1.6705642,1.3686155,1.1585642,1.0896411,1.2340513,1.8182565,2.156308,2.3368206,2.422154,2.4451284,2.225231,1.9429746,1.5425643,1.1257436,0.9616411,0.82379496,0.79097444,0.8533334,0.93866676,0.9288206,0.9124103,0.8336411,0.82379496,0.99774367,1.467077,2.4418464,2.917744,3.3312824,3.7842054,4.0336413,4.2994876,4.450462,4.522667,4.4406157,4.0500517,4.562052,4.8344617,4.916513,5.080616,5.805949,6.2720003,6.6034875,6.7774363,6.816821,6.7971287,6.193231,5.6385646,4.8607183,4.007385,3.6463592,3.8498464,3.2656412,2.6420515,2.294154,2.0873847,1.8871796,1.9659488,1.9659488,1.7493335,1.3981539,0.90912825,0.62030774,0.44307697,0.3117949,0.17394873,0.24287182,0.318359,0.34133336,0.380718,0.6432821,0.9189744,1.1782565,1.1552821,0.8598975,0.5677949,0.380718,0.5415385,0.60389745,0.47917953,0.4004103,0.5513847,0.77128214,0.9353847,0.93866676,0.7187693,0.48246157,0.4004103,0.41025645,0.4594872,0.49887183,0.65969235,0.8467693,1.0962052,1.4834872,2.1234872,2.4910772,2.6486156,2.5698464,2.4057438,2.487795,2.809436,3.259077,3.876103,4.394667,4.2535386,3.0916924,2.5993848,2.4976413,2.6322052,2.9801028,3.7349746,4.0336413,4.161641,4.332308,4.6933336,4.069744,3.5183592,3.1507695,3.318154,4.6080003,4.5489235,4.2174363,4.4242053,4.965744,4.644103,4.2535386,4.2174363,4.394667,4.391385,3.5577438,1.9200002,1.4112822,1.142154,0.7581539,0.42994875,0.67610264,0.6629744,0.5481026,0.40697438,0.22646156,0.15097436,0.11158975,0.101743594,0.108307704,0.13456412,0.1148718,0.08861539,0.04266667,0.02297436,0.108307704,0.13784617,0.35774362,0.2986667,0.0,0.0,0.13784617,0.108307704,0.055794876,0.029538464,0.0,0.0,0.12143591,0.2855385,0.45292312,0.6301539,0.49887183,0.56123084,0.71548724,0.8533334,0.84348726,1.0404103,1.0994873,0.99774367,0.8041026,0.65641034,0.72861546,0.8730257,0.99774367,1.0732309,1.1388719,1.1454359,1.0436924,0.955077,0.8960001,0.8008206,0.6301539,0.5316923,0.48574364,0.44964105,0.36758977,0.20020515,0.06235898,0.0,0.0,0.0,0.18707694,0.2297436,0.15425642,0.04594872,0.06235898,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0,0.013128206,0.02297436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.009846155,0.013128206,0.013128206,0.006564103,0.0,0.0,0.006564103,0.009846155,0.009846155,0.016410258,0.02297436,0.049230773,0.0951795,0.14441027,0.18707694,0.27241027,0.24943592,0.23302566,0.3117949,0.55794877,0.6892308,0.6662565,0.5973334,0.7122052,1.3489232,1.467077,1.1191796,0.8566154,0.98133343,1.5195899,1.6213335,2.0873847,2.3466668,2.2777438,2.1956925,2.8356924,2.6978464,2.7831798,3.3608208,3.9548721,3.3969233,2.5829747,1.8018463,1.3226668,1.4145643,2.9407182,3.0720003,1.9889232,0.5349744,0.21989745,0.18379489,0.2100513,0.18379489,0.101743594,0.06235898,0.026256412,0.08205129,0.7122052,1.6344616,1.8149745,1.1388719,1.2865642,1.6804104,1.8937438,1.657436,1.014154,0.827077,0.65969235,0.3708718,0.1148718,0.12143591,0.20348719,0.28225642,0.32820517,0.36758977,0.36758977,0.3314872,0.24615386,0.20020515,0.38400003,0.36758977,0.28882053,0.2297436,0.2231795,0.26256412,0.26584616,0.23302566,0.17723078,0.12471796,0.118153855,0.20348719,0.30851284,0.28225642,0.13784617,0.036102567,0.03938462,0.02297436,0.013128206,0.013128206,0.0,0.006564103,0.01969231,0.029538464,0.029538464,0.009846155,0.0032820515,0.0,0.0032820515,0.006564103,0.006564103,0.009846155,0.03938462,0.08861539,0.14441027,0.21661541,0.27569234,0.23630771,0.18707694,0.18051283,0.20348719,0.22646156,0.17394873,0.13456412,0.13456412,0.15097436,0.18379489,0.13784617,0.09189744,0.08533334,0.14441027,0.19364104,0.20348719,0.21333335,0.2855385,0.46933338,0.5513847,0.4594872,0.38728207,0.50543594,0.9714873,1.7624617,2.9078977,3.9187696,4.201026,3.0227695,1.9167181,2.0775387,2.428718,2.353231,1.7001027,2.1924105,2.4648206,2.2678976,1.6935385,1.1815386,0.8402052,0.61374366,0.5349744,0.73517954,1.4572309,2.0545642,2.2482052,2.2383592,2.1234872,1.9298463,1.6246156,1.9528207,2.2088206,2.156308,2.0118976,2.5895386,3.2065644,3.7448208,4.2174363,4.7524104,5.0838976,4.9394875,4.4734364,4.0467696,4.197744,5.293949,5.5762057,5.605744,5.85518,6.685539,6.416411,5.98318,5.3792825,4.7261543,4.276513,3.5872824,2.9604106,2.4648206,2.1431797,1.9922053,2.353231,2.9571285,4.3651285,6.380308,8.064001,7.7981544,7.0400004,6.5312824,6.5280004,6.810257,6.449231,6.436103,6.6100516,6.961231,7.640616,8.644924,9.176616,9.639385,9.984001,9.7214365,10.358154,10.71918,10.256411,9.091283,8.01477,7.4896417,7.5552826,8.507077,10.571488,13.922462,19.02277,24.280617,29.718977,34.71426,38.009438,34.73395,29.88308,24.146053,18.54031,14.424617,11.670976,8.769642,6.2818465,4.5489235,3.69559,2.7076926,1.6016412,0.81394875,0.44307697,0.23302566,0.12143591,0.055794876,0.029538464,0.032820515,0.052512825,0.059076928,0.06235898,0.072205134,0.098461546,0.14112821,0.0951795,0.059076928,0.036102567,0.01969231,0.0,0.006564103,0.013128206,0.01969231,0.02297436,0.01969231,0.026256412,0.052512825,0.13456412,0.28225642,0.46276927,0.64000005,0.7122052,0.7450257,0.72861546,0.5973334,0.32820517,0.20020515,0.118153855,0.049230773,0.029538464,0.01969231,0.01969231,0.026256412,0.04266667,0.08533334,0.2297436,0.28225642,0.2297436,0.15097436,0.20676924,0.23302566,0.256,0.29538465,0.33476925,0.33476925,0.33805132,0.40697438,0.56451285,0.7811283,0.95835906,1.0272821,0.955077,0.86646163,0.8467693,0.9353847,1.086359,1.2373334,1.3718976,1.5031796,1.6640002,1.8412309,1.9561027,1.9561027,1.8313848,1.6147693,1.4736412,1.2570257,1.0404103,0.8402052,0.61374366,0.5973334,0.6432821,0.7253334,0.81394875,0.8795898,0.92225647,0.9714873,1.020718,1.0699488,1.1093334,1.2012309,1.657436,2.0841026,2.162872,1.6311796,1.6311796,1.7493335,1.9232821,2.1792822,2.6617439,1.8510771,1.3554872,1.1749744,1.1946667,1.1782565,1.1618463,1.0568206,0.92225647,0.8336411,0.88943595,1.014154,1.083077,1.020718,0.8763078,0.81394875,0.88943595,0.8763078,0.81394875,0.76800007,0.84348726,8.2445135,8.635077,9.888822,11.424822,12.616206,12.809847,12.924719,14.834873,16.65313,17.112617,15.553642,13.492514,12.796719,12.304411,11.047385,8.234667,5.0838976,4.2436924,4.4012313,4.6769233,4.630975,3.8990772,3.82359,4.3716927,5.356308,6.439385,6.0258465,6.186667,6.636308,7.00718,6.8397956,7.197539,7.9097443,8.260923,8.234667,8.480822,8.093539,7.3616414,7.2960005,7.9425645,8.372514,8.185436,8.342975,8.411898,7.958975,6.5312824,5.579488,5.5171285,5.8486156,5.858462,4.601436,3.5610259,2.9407182,2.284308,1.6935385,1.8445129,2.1333334,2.1825643,2.0841026,1.9987694,2.1530259,1.9331284,1.5360001,1.2077949,1.0732309,1.1290257,1.6180514,1.7526156,1.7493335,1.7723079,1.9265642,1.6705642,1.5163078,1.3423591,1.1618463,1.1257436,0.9911796,0.77456415,0.6301539,0.6235898,0.7515898,0.9911796,1.2406155,1.522872,1.8018463,1.9922053,2.425436,2.6026669,2.7864618,3.1376412,3.7218463,4.1025643,4.378257,4.4340515,4.2994876,4.1485133,4.9526157,4.9788723,4.8804107,5.4416413,7.574975,7.529026,7.7292314,7.893334,8.277334,9.665642,9.472001,8.5661545,7.453539,6.3868723,5.356308,4.8114877,3.8596926,3.3805132,3.4560003,3.373949,2.8127182,2.7273848,2.6190772,2.294154,1.8543591,1.5491283,1.1323078,0.7778462,0.5415385,0.35774362,0.4201026,0.44307697,0.35774362,0.2986667,0.5940513,0.9353847,1.3226668,1.3850257,1.1257436,0.90912825,0.72861546,0.7187693,0.827077,0.9682052,1.0469744,1.1585642,1.2012309,1.273436,1.3620514,1.3357949,0.9321026,0.636718,0.45292312,0.38400003,0.42338464,0.7384616,1.1257436,1.6114873,2.3335385,3.570872,4.2240005,4.352,3.7316926,2.7700515,2.5173335,2.6978464,3.1277952,3.8465643,4.568616,4.6769233,3.8104618,3.3641028,3.1770258,3.1376412,3.190154,3.308308,3.69559,4.2962055,5.100308,6.1407185,5.0510774,4.1058464,3.4133337,3.3805132,4.7360005,4.8049235,4.4964104,4.3552823,4.562052,4.9362054,4.8836927,4.44718,4.6178465,5.1922054,4.778667,3.314872,2.1431797,1.4309745,1.1651284,1.1323078,1.1848207,1.0338463,0.83035904,0.6432821,0.46276927,0.58092314,0.5677949,0.40369233,0.16738462,0.0,0.0,0.032820515,0.068923086,0.101743594,0.14769232,0.15097436,0.35446155,0.34789747,0.128,0.098461546,0.09189744,0.036102567,0.0,0.006564103,0.036102567,0.04266667,0.15425642,0.30194873,0.44964105,0.5874872,0.6071795,0.7450257,0.892718,0.9189744,0.6465641,0.42994875,0.28882053,0.22646156,0.23630771,0.31507695,0.42338464,0.49230772,0.5415385,0.58420515,0.6268718,0.636718,0.56123084,0.50543594,0.5021539,0.48246157,0.3314872,0.23958977,0.17394873,0.101743594,0.0,0.0,0.0,0.0,0.0,0.0,0.072205134,0.098461546,0.059076928,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.009846155,0.013128206,0.013128206,0.006564103,0.0,0.013128206,0.049230773,0.072205134,0.06564103,0.016410258,0.072205134,0.15097436,0.23958977,0.3314872,0.44307697,0.43651286,0.32820517,0.29210258,0.42338464,0.7220513,0.8172308,0.74830776,0.75487185,1.1093334,2.1103592,2.674872,1.913436,1.2406155,1.2077949,1.4769232,1.6738462,2.0742567,2.2121027,2.2022567,2.7536411,3.370667,3.1606157,3.0424619,3.3050258,3.6069746,3.0129232,2.353231,1.5097437,0.8205129,1.079795,2.6256413,3.245949,2.5961027,1.2077949,0.48246157,0.27897438,0.25928208,0.23302566,0.15425642,0.12143591,0.07876924,0.101743594,0.77128214,1.8871796,2.4943593,1.4408206,1.3161026,1.585231,1.8576412,1.8642052,1.4506668,1.2931283,0.9944616,0.53825647,0.256,0.19364104,0.098461546,0.068923086,0.118153855,0.18379489,0.25271797,0.27897438,0.21333335,0.12471796,0.20020515,0.23958977,0.23958977,0.23630771,0.24287182,0.24287182,0.22646156,0.18707694,0.14112821,0.10502565,0.08205129,0.098461546,0.108307704,0.10502565,0.08205129,0.036102567,0.032820515,0.02297436,0.013128206,0.006564103,0.0,0.006564103,0.02297436,0.036102567,0.036102567,0.016410258,0.006564103,0.006564103,0.006564103,0.006564103,0.013128206,0.02297436,0.068923086,0.128,0.19364104,0.25928208,0.27569234,0.20348719,0.15097436,0.15425642,0.19364104,0.2231795,0.17723078,0.19364104,0.27569234,0.2986667,0.2297436,0.13456412,0.055794876,0.02297436,0.059076928,0.068923086,0.1148718,0.19692309,0.3314872,0.5546667,0.5677949,0.46933338,0.4594872,0.71548724,1.3981539,2.1825643,3.1376412,3.7874875,3.7185643,2.5961027,1.8215386,2.284308,2.7963078,2.793026,2.3466668,2.9965131,3.045744,2.4943593,1.6410258,1.083077,1.2964103,1.3292309,1.273436,1.2668719,1.4998976,1.9396925,2.477949,3.0982566,3.501949,3.0884104,2.868513,3.3641028,3.7087183,3.4658465,2.6322052,2.7044106,2.9472823,3.0523078,3.0523078,3.3280003,3.446154,3.4822567,3.370667,3.2623591,3.5282054,4.886975,5.5105643,5.87159,6.498462,7.962257,8.395488,7.9950776,6.774154,5.2742567,4.562052,4.2929235,3.8498464,3.1081028,2.294154,2.0053334,2.428718,2.8127182,3.7251284,5.622154,8.854975,10.256411,9.235693,7.7981544,7.000616,6.944821,6.363898,6.1046157,6.1997952,6.803693,8.172308,10.230155,11.021129,10.962052,10.496001,10.092308,11.30995,12.25518,11.88759,10.171078,8.073847,7.125334,7.056411,8.2445135,10.722463,14.185027,19.203283,24.982977,30.480413,35.088413,38.63959,36.562054,32.643284,27.24431,21.083899,15.225437,11.969642,9.120821,6.8529234,5.3103595,4.588308,3.3411283,1.9265642,1.0699488,0.79425645,0.4201026,0.17066668,0.06235898,0.032820515,0.059076928,0.15425642,0.26584616,0.23302566,0.17066668,0.13784617,0.14769232,0.098461546,0.07876924,0.068923086,0.052512825,0.02297436,0.032820515,0.029538464,0.032820515,0.04266667,0.049230773,0.08205129,0.128,0.2231795,0.37415388,0.5907693,0.9189744,1.273436,1.3292309,1.0994873,0.9156924,0.5874872,0.43323082,0.28882053,0.12471796,0.036102567,0.032820515,0.04266667,0.06564103,0.0951795,0.14112821,0.3052308,0.33476925,0.29210258,0.26912823,0.41025645,0.4397949,0.446359,0.46276927,0.48902568,0.48902568,0.4955898,0.5546667,0.6826667,0.85005134,0.9878975,1.0568206,0.9944616,0.8992821,0.84348726,0.8467693,0.9124103,0.9878975,1.086359,1.2340513,1.4572309,1.7952822,2.0118976,2.0545642,1.8970258,1.522872,1.2504616,1.0502565,0.8992821,0.7778462,0.6859488,0.6662565,0.69251287,0.7581539,0.8402052,0.9156924,0.97805136,1.0469744,1.1290257,1.2274873,1.332513,1.4178462,1.6968206,1.9167181,1.8674873,1.404718,1.5195899,1.6311796,1.7394873,1.9954873,2.6912823,2.0020514,1.463795,1.2603078,1.3292309,1.3554872,1.332513,1.3029745,1.2373334,1.1782565,1.2406155,1.332513,1.2537436,1.1454359,1.1093334,1.204513,1.4178462,1.4244103,1.2964103,1.1257436,1.020718,7.9786673,8.04759,8.162462,8.832001,9.83959,10.259693,10.157949,10.650257,12.406155,14.477129,14.309745,14.083283,13.804309,13.338258,12.3766165,10.423796,6.6100516,5.536821,5.398975,5.293949,5.2348723,4.44718,4.5489235,5.1626673,6.1538467,7.6176414,6.3343596,5.3070774,4.706462,4.5587697,4.7327185,6.564103,7.6996927,8.03118,7.9327188,8.274052,7.8802056,6.9842057,6.9054365,7.8080006,8.697436,9.321027,9.632821,9.40636,8.602257,7.3616414,5.858462,5.228308,4.8607183,4.457026,4.023795,3.2656412,2.609231,2.281026,2.3335385,2.6683078,2.9243078,2.917744,2.5928206,2.2547693,2.553436,2.5796926,2.1464617,1.7723079,1.6410258,1.585231,1.7362052,1.7329233,1.6311796,1.5130258,1.4769232,1.4276924,1.6804104,1.972513,2.1234872,2.0545642,1.723077,1.2471796,0.69907695,0.3117949,0.44307697,1.2996924,2.1333334,2.8422565,3.2196925,2.937436,2.8882053,3.1606157,3.4067695,3.5380516,3.7185643,4.197744,4.7458467,5.093744,5.2512827,5.536821,6.5706673,6.5411286,6.6822567,7.7948723,10.256411,8.720411,7.8834877,7.8834877,8.910769,11.221334,11.0375395,10.374565,9.872411,9.55077,8.822155,7.4469748,5.930667,5.2348723,5.287385,5.0018463,4.322462,3.6004105,2.9013336,2.300718,1.8904617,2.162872,1.8215386,1.2668719,0.78769237,0.5513847,0.508718,0.4266667,0.2986667,0.23302566,0.43323082,0.64000005,0.827077,0.9616411,1.0633847,1.204513,1.1323078,0.8566154,0.9747693,1.4703591,1.7132308,1.6836925,1.591795,1.6705642,1.9298463,2.1464617,1.7657437,1.2406155,0.77456415,0.49887183,0.44964105,0.77456415,1.4211283,2.3302567,3.5282054,5.1167183,6.0324106,6.1374364,5.037949,3.3805132,2.8356924,2.6945643,2.7536411,3.131077,3.8006158,4.6145644,5.221744,5.031385,4.4406157,3.7120004,2.9440002,2.0676925,2.5665643,3.7185643,5.100308,6.6034875,4.97559,3.9647183,3.4330258,3.2918978,3.5249233,3.5544617,3.5183592,3.4231799,3.5577438,4.519385,4.6178465,3.629949,3.5183592,4.4832826,4.9821544,4.7622566,3.508513,2.487795,2.1333334,2.0512822,1.6836925,1.7001027,1.8707694,2.044718,2.15959,2.0020514,1.6016412,1.0272821,0.44964105,0.13128206,0.08861539,0.098461546,0.16410258,0.26584616,0.34789747,0.34789747,0.25928208,0.24615386,0.3052308,0.24943592,0.08533334,0.01969231,0.0,0.013128206,0.072205134,0.14441027,0.24615386,0.3117949,0.29210258,0.17066668,0.5218462,0.72861546,0.79097444,0.69579494,0.4135385,0.25271797,0.15753847,0.1148718,0.14112821,0.30851284,0.38400003,0.32164106,0.23958977,0.18707694,0.15753847,0.14769232,0.16082053,0.21333335,0.29210258,0.34133336,0.18707694,0.13784617,0.12471796,0.08861539,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.0032820515,0.0032820515,0.0,0.0032820515,0.049230773,0.1148718,0.14441027,0.12471796,0.08533334,0.2231795,0.37415388,0.6170257,0.90912825,1.079795,0.80738467,0.49230772,0.35446155,0.4594872,0.7122052,0.9321026,0.81394875,0.9485129,1.595077,2.6912823,3.570872,2.681436,1.9232821,1.9987694,2.428718,2.0939488,1.5721027,1.4834872,2.1070771,3.3969233,3.5282054,3.4560003,3.170462,2.7503593,2.349949,2.4713848,2.6420515,2.038154,0.98461545,0.9353847,1.4900514,1.8281027,2.1333334,2.0906668,0.8730257,0.36102566,0.20348719,0.18707694,0.19692309,0.2231795,0.190359,0.14441027,0.36758977,1.1126155,2.609231,1.9856411,1.5786668,1.4572309,1.5064616,1.4342566,1.654154,1.6475899,1.2340513,0.6432821,0.512,0.5940513,0.35774362,0.14441027,0.08861539,0.128,0.17394873,0.17723078,0.14112821,0.0951795,0.08533334,0.13784617,0.21989745,0.25928208,0.23958977,0.18051283,0.16410258,0.14112821,0.118153855,0.09189744,0.049230773,0.03938462,0.036102567,0.03938462,0.04594872,0.04594872,0.02297436,0.016410258,0.013128206,0.009846155,0.02297436,0.029538464,0.032820515,0.029538464,0.016410258,0.016410258,0.013128206,0.013128206,0.016410258,0.02297436,0.036102567,0.04594872,0.072205134,0.108307704,0.15425642,0.21661541,0.19364104,0.15097436,0.13128206,0.14441027,0.190359,0.18051283,0.14112821,0.23630771,0.4397949,0.50543594,0.34133336,0.19692309,0.09189744,0.032820515,0.03938462,0.055794876,0.1148718,0.20676924,0.3249231,0.4594872,0.4266667,0.45620516,0.60389745,1.0010257,1.8445129,2.353231,2.5271797,2.6289232,2.6289232,2.1989746,2.0709746,2.3893335,2.5731285,2.5961027,2.9833848,3.7284105,3.7809234,3.114667,2.0644104,1.3095386,1.9167181,2.1202054,2.0939488,1.913436,1.5425643,2.1136413,3.249231,4.571898,5.3169236,4.312616,4.2535386,4.8607183,5.3398976,5.10359,3.761231,2.865231,2.9407182,2.9046156,2.550154,2.550154,2.930872,3.4560003,3.4592824,2.8553848,2.1530259,2.9669745,3.4888208,4.1485133,5.2611284,7.0400004,8.329846,7.8145647,6.1505647,4.450462,4.2863593,4.6802053,4.5522056,3.6168208,2.3663592,2.0644104,2.5435898,3.2229745,4.20759,5.8157954,8.549745,11.323078,10.371283,8.631796,7.3583593,6.11118,5.179077,5.149539,5.609026,6.51159,8.1755905,10.568206,11.254155,10.656821,9.636104,9.4916935,11.0145645,12.484924,12.694975,11.378873,9.216001,7.7357955,6.8430777,7.4863596,9.905231,13.61395,19.042463,25.974155,32.518566,37.3399,39.66031,38.262157,33.96595,28.409437,22.340925,15.638975,12.281437,9.40636,7.138462,5.5663595,4.7491283,3.5052311,2.3236926,1.6377437,1.3357949,0.761436,0.31507695,0.101743594,0.04266667,0.10502565,0.28882053,0.51856416,0.48246157,0.33805132,0.18379489,0.06564103,0.04594872,0.07548718,0.108307704,0.1148718,0.08533334,0.072205134,0.055794876,0.052512825,0.06564103,0.07548718,0.16082053,0.24943592,0.3249231,0.47589746,0.88615394,1.3883078,1.9593848,1.9265642,1.4244103,1.3686155,1.332513,1.0502565,0.67938465,0.33805132,0.10502565,0.09189744,0.1148718,0.14769232,0.17723078,0.20348719,0.26256412,0.318359,0.38728207,0.4660513,0.5546667,0.56451285,0.54482055,0.5152821,0.4955898,0.4955898,0.52512825,0.571077,0.6268718,0.6892308,0.7581539,0.81394875,0.79425645,0.75487185,0.7253334,0.71548724,0.69579494,0.69251287,0.7450257,0.892718,1.1618463,1.6246156,1.9035898,1.9692309,1.7952822,1.3653334,1.0732309,0.8566154,0.7187693,0.6432821,0.6071795,0.60061544,0.6235898,0.6859488,0.77456415,0.8467693,0.90256417,0.9517949,1.0666667,1.2603078,1.4867693,1.6607181,1.4703591,1.0732309,0.6892308,0.5973334,0.85005134,1.2438976,1.7165129,2.100513,2.1333334,1.8346668,1.5130258,1.3193847,1.2931283,1.3686155,1.467077,1.529436,1.5425643,1.522872,1.5425643,1.5753847,1.3718976,1.2340513,1.276718,1.4178462,1.6869745,1.8084104,1.7952822,1.6640002,1.404718,9.6295395,9.810052,7.834257,7.003898,8.172308,9.734565,10.052924,10.167795,10.450052,10.965334,11.490462,12.064821,10.725744,8.326565,6.8496413,9.399796,9.6065645,8.67118,7.076103,5.5991797,5.293949,5.5630774,5.986462,6.1768208,6.2129235,6.6527185,7.3714876,7.059693,6.5444107,6.491898,7.3682055,10.811078,10.564924,9.117539,8.103385,8.283898,7.4929237,6.9645133,6.892308,7.4896417,9.002667,9.540924,9.353847,8.316719,6.774154,5.5532312,4.6867695,4.332308,3.7907696,3.1671798,3.387077,4.6802053,4.4274874,4.0008206,4.0336413,4.4242053,5.0838976,5.293949,5.1364107,4.6769233,3.9811285,3.5807183,3.2853336,3.1277952,2.9636924,2.487795,2.4746668,2.6190772,2.5009232,2.2088206,2.3204105,2.5632823,2.5600002,2.425436,2.1989746,1.847795,1.1749744,0.7515898,0.512,0.47917953,0.74830776,2.6387694,3.570872,3.826872,3.5446157,2.7175386,2.044718,1.9396925,2.5829747,3.4888208,3.5249233,4.0008206,4.8147697,5.5171285,6.170257,7.3550773,8.4283085,8.579283,8.326565,8.011488,7.765334,7.8506675,7.506052,7.7948723,9.330873,12.2847185,13.371078,13.082257,12.196103,11.848206,13.53518,12.754052,11.283693,9.849437,8.687591,7.5520005,6.11118,4.269949,2.865231,2.1333334,1.6935385,1.595077,1.8642052,1.8576412,1.394872,0.74830776,0.47917953,0.4201026,0.4266667,0.3708718,0.15097436,0.21333335,0.34789747,0.5316923,0.7056411,0.7778462,0.8992821,1.0305642,1.1848207,1.3456411,1.4802053,1.6738462,1.9265642,2.156308,2.3762052,2.6715899,3.0720003,2.733949,2.166154,1.6443079,1.204513,1.2176411,1.9987694,3.18359,4.4340515,5.4482055,6.413129,6.7544622,6.3212314,5.4580517,5.0215387,4.4110775,3.754667,3.314872,3.4658465,4.699898,6.12759,6.413129,5.421949,3.6036925,1.9692309,1.4309745,2.6617439,4.315898,5.6287184,6.409847,3.882667,3.2787695,3.7842054,4.2929235,3.4034874,2.7208207,2.556718,3.117949,3.9942567,4.164923,4.164923,4.056616,3.367385,2.4648206,2.5632823,3.4297438,3.9844105,3.7120004,2.6486156,1.404718,0.7318975,1.9298463,3.8498464,5.8223596,7.6274877,4.493129,2.3433847,1.086359,0.58420515,0.65641034,0.44964105,0.15753847,0.12143591,0.2986667,0.27569234,0.22646156,0.16738462,0.18051283,0.24943592,0.27569234,0.23958977,0.09189744,0.0,0.0,0.0,0.3052308,0.508718,0.5874872,0.49887183,0.18379489,0.28225642,0.31507695,0.25928208,0.16738462,0.16738462,0.15425642,0.13456412,0.10502565,0.08861539,0.13784617,0.17394873,0.18379489,0.17723078,0.15753847,0.12143591,0.02297436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.026256412,0.02297436,0.009846155,0.0032820515,0.016410258,0.101743594,0.14112821,0.09189744,0.072205134,0.36758977,0.574359,0.761436,1.3193847,2.044718,2.166154,1.8248206,1.3456411,0.9321026,0.7220513,0.80738467,1.4178462,1.3062565,1.1716924,1.3620514,1.8609232,1.7165129,1.7788719,2.0118976,2.4155898,3.0523078,2.2580514,1.7033848,2.0086155,3.006359,3.7382567,3.8596926,3.5807183,2.793026,1.9462565,2.044718,3.0949745,4.821334,4.785231,2.7076926,0.47261542,1.1946667,2.3991797,3.245949,3.1081028,1.5556924,0.65312827,0.36430773,0.3314872,0.3708718,0.44307697,0.42994875,0.27241027,0.16082053,0.43651286,1.5721027,2.156308,1.9364104,1.4802053,1.1782565,1.2504616,1.8609232,1.4473847,0.77456415,0.34133336,0.36758977,1.1093334,0.9682052,0.48574364,0.09189744,0.09189744,0.128,0.128,0.098461546,0.098461546,0.24287182,0.36758977,0.43323082,0.39056414,0.28882053,0.28882053,0.31507695,0.256,0.18379489,0.12143591,0.06235898,0.06235898,0.052512825,0.04594872,0.04594872,0.04594872,0.02297436,0.016410258,0.02297436,0.049230773,0.12143591,0.14769232,0.13456412,0.07876924,0.016410258,0.016410258,0.0032820515,0.0,0.01969231,0.049230773,0.06235898,0.06235898,0.032820515,0.016410258,0.02297436,0.04594872,0.068923086,0.08533334,0.07876924,0.055794876,0.029538464,0.04266667,0.101743594,0.21661541,0.39712822,0.64000005,0.5907693,0.44307697,0.24615386,0.08861539,0.07548718,0.11158975,0.14112821,0.15753847,0.18051283,0.2297436,0.30194873,0.42994875,0.6859488,1.0994873,1.6475899,2.0020514,1.7427694,1.394872,1.2603078,1.4178462,1.7985642,2.3236926,2.92759,3.4133337,3.4494362,3.8990772,4.1780515,3.5872824,2.359795,1.6640002,1.332513,1.2406155,1.4572309,2.0053334,2.8849232,4.33559,6.3212314,7.6635904,7.7292314,6.422975,4.2272825,4.1911798,5.0510774,5.7403083,5.3858466,3.7743592,2.5764105,2.0020514,1.9659488,2.0742567,2.2088206,2.3171284,2.281026,2.0578463,1.6771283,1.8871796,2.7995899,3.817026,4.7589746,5.8453336,7.1614366,6.557539,5.612308,5.179077,5.3858466,5.6418467,4.8640003,3.6069746,2.4681027,2.0906668,3.4592824,4.7983594,5.674667,6.2916927,7.4765134,8.001641,8.004924,7.712821,7.1483083,6.1341543,5.6320004,5.8912826,6.193231,6.3573337,6.7610264,7.003898,7.384616,7.9885135,8.854975,9.980719,13.397334,15.458463,15.606155,13.952001,11.290257,9.363693,8.093539,7.972103,9.426052,12.832822,18.435284,25.632822,34.1399,41.57703,43.457645,38.02585,30.083284,23.023592,18.179283,14.8480015,12.599796,9.961026,7.506052,5.664821,4.699898,3.6135387,2.609231,1.8149745,1.2635899,0.88615394,0.50543594,0.19364104,0.04594872,0.068923086,0.16738462,0.28882053,0.4397949,0.446359,0.2986667,0.15097436,0.09189744,0.11158975,0.15425642,0.18379489,0.18379489,0.108307704,0.06564103,0.059076928,0.07548718,0.07548718,0.25928208,0.4594872,0.6432821,1.079795,2.349949,2.7634873,2.6026669,2.2055387,2.0644104,2.8225644,3.2754874,2.425436,1.3522053,0.5907693,0.15097436,0.14112821,0.19364104,0.25928208,0.31507695,0.3511795,0.4004103,0.4397949,0.47589746,0.50543594,0.51856416,0.46933338,0.4201026,0.3708718,0.33476925,0.33476925,0.33476925,0.3446154,0.380718,0.4397949,0.48902568,0.52512825,0.5152821,0.5152821,0.54482055,0.58092314,0.5907693,0.55794877,0.55794877,0.6498462,0.86974365,1.3226668,1.5885129,1.6278975,1.4605129,1.204513,1.020718,0.8402052,0.67938465,0.55794877,0.47261542,0.43651286,0.446359,0.51856416,0.636718,0.74830776,0.8336411,0.892718,0.98133343,1.1323078,1.3259488,1.522872,1.4244103,1.1684103,0.9156924,0.8533334,1.086359,1.4473847,1.8806155,2.1956925,2.0611284,1.8904617,1.6344616,1.3489232,1.1388719,1.1749744,1.3587693,1.5688206,1.7033848,1.7132308,1.6016412,1.3817437,1.2176411,1.0962052,1.017436,0.9911796,1.1618463,1.3981539,1.6607181,1.9167181,2.1366155,14.132514,13.5548725,12.317539,11.201642,10.742155,11.1983595,11.447796,11.503591,11.569232,11.871181,12.649027,13.466257,12.517745,10.440206,8.192,7.030154,6.4295387,6.308103,6.3540516,6.5312824,7.076103,7.384616,7.387898,6.8955903,6.370462,6.9087186,7.5913854,7.9261546,7.2303596,6.11118,6.442667,7.6964107,8.054154,7.77518,7.276308,7.125334,7.076103,7.003898,6.994052,7.128616,7.4896417,7.8703594,7.394462,6.2227697,4.972308,4.7360005,5.579488,6.311385,6.547693,6.2129235,5.536821,5.031385,4.273231,3.95159,4.2962055,5.0477953,5.366154,4.634257,3.882667,3.5938463,3.6890259,4.896821,4.164923,3.2000003,3.062154,4.1583595,3.9220517,4.0303593,4.263385,4.493129,4.699898,4.71959,4.601436,4.414359,4.2207184,4.092718,4.279795,5.3005133,5.5072823,4.9329233,5.287385,7.2205133,6.183385,4.768821,4.2207184,4.4373336,3.131077,2.7602053,3.2525132,4.2830772,5.2578464,5.3136415,5.504,5.7764106,5.9963083,5.9503593,5.805949,5.618872,6.183385,7.3649235,8.096821,8.756514,9.478565,9.708308,9.42277,9.133949,10.397539,11.191795,10.692924,8.881231,6.554257,7.8506675,9.291488,10.952206,12.455385,12.960821,11.510155,9.219283,6.491898,3.9680004,2.5238976,2.0644104,2.2219489,2.484513,2.5140514,2.1398976,1.3226668,1.0108719,1.0338463,1.2373334,1.4966155,1.214359,1.1618463,1.2077949,1.2307693,1.1191796,1.2406155,1.3653334,1.4736412,1.529436,1.467077,1.4276924,1.4375386,1.6114873,1.9265642,2.231795,2.4582565,2.3827693,2.176,1.9528207,1.7657437,1.8379488,2.2744617,2.8914874,3.56759,4.240411,4.7458467,4.781949,4.420923,4.1058464,4.640821,4.9985647,5.1265645,4.7983594,4.1813335,3.8334363,3.495385,2.8291285,2.2711797,2.103795,2.4681027,3.7185643,4.6834874,5.333334,5.6418467,5.602462,4.571898,3.6496413,2.865231,2.1956925,1.6082052,1.6968206,2.0775387,2.7241027,3.3050258,3.2131286,3.18359,3.3247182,4.141949,5.0018463,4.1124105,2.605949,3.0162053,4.1222568,5.221744,6.114462,6.340924,6.9710774,7.3747697,7.1548724,6.1407185,3.9318976,2.225231,1.014154,0.35774362,0.4135385,0.54482055,0.5973334,0.39056414,0.08533334,0.17723078,0.256,0.318359,0.38728207,0.446359,0.4201026,0.26584616,0.20020515,0.15425642,0.08861539,0.0,0.06235898,0.101743594,0.118153855,0.128,0.17066668,0.17066668,0.15097436,0.0951795,0.032820515,0.032820515,0.029538464,0.026256412,0.01969231,0.016410258,0.026256412,0.036102567,0.036102567,0.036102567,0.032820515,0.02297436,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.02297436,0.055794876,0.13128206,0.25928208,0.26584616,0.16082053,0.059076928,0.052512825,0.20676924,0.40369233,0.4660513,0.72861546,1.2373334,1.7394873,2.2186668,2.048,1.6508719,1.3423591,1.3095386,1.332513,1.5655385,2.0742567,2.6157951,2.6190772,2.8914874,3.0391798,2.6847181,2.034872,1.8806155,1.8970258,2.356513,2.6518977,2.5961027,2.4188719,2.6486156,2.7995899,2.5829747,2.0873847,1.7755898,3.255795,3.82359,3.318154,2.028308,0.69251287,1.6672822,2.8553848,3.511795,3.387077,2.7175386,2.1169233,0.9944616,0.37743592,0.41682056,0.39384618,0.256,0.5021539,0.6432821,0.6629744,1.0469744,2.540308,2.8324106,2.477949,1.8149745,0.9714873,0.86646163,0.6498462,0.4660513,0.5152821,1.0371283,1.1881026,0.7975385,0.3446154,0.08861539,0.07876924,0.12471796,0.21661541,0.23302566,0.17723078,0.14769232,0.2100513,0.20348719,0.18051283,0.17394873,0.19364104,0.19692309,0.17066668,0.13128206,0.08861539,0.036102567,0.04594872,0.06235898,0.068923086,0.068923086,0.068923086,0.06564103,0.049230773,0.036102567,0.036102567,0.06235898,0.10502565,0.11158975,0.13128206,0.17066668,0.2100513,0.09189744,0.04594872,0.04594872,0.059076928,0.06235898,0.06235898,0.03938462,0.016410258,0.009846155,0.032820515,0.059076928,0.08205129,0.08533334,0.07548718,0.09189744,0.08533334,0.101743594,0.16738462,0.26584616,0.3249231,0.19692309,0.17394873,0.15425642,0.108307704,0.07548718,0.07548718,0.07548718,0.0951795,0.13784617,0.21661541,0.27897438,0.5021539,1.0305642,1.654154,1.782154,1.7263591,1.5556924,1.5130258,1.7001027,2.0545642,2.3729234,2.605949,2.6715899,2.5731285,2.3860514,3.0227695,2.7634873,2.15959,1.7526156,2.041436,2.0742567,1.9692309,1.8379488,1.8084104,2.0545642,2.8717952,3.882667,4.70318,4.8311796,3.639795,3.2984617,4.348718,5.477744,5.8420515,5.0576415,3.515077,3.1081028,3.0424619,3.006359,3.1737437,2.986667,2.7634873,2.3696413,1.847795,1.4211283,1.5425643,2.0512822,2.8750772,3.82359,4.598154,5.0084105,4.630975,4.3290257,4.46359,4.886975,4.713026,4.3027697,4.1583595,4.70318,6.2785645,8.044309,8.664616,8.267488,7.0498466,5.2545643,4.6080003,4.663795,5.3169236,6.2752824,7.0498466,6.5870776,5.927385,5.5532312,5.8945646,7.322257,9.058462,9.301334,9.856001,11.044104,11.687386,12.95754,14.257232,15.058052,14.92677,13.525334,12.133744,11.753027,12.2157955,13.525334,15.849027,20.240412,26.453335,34.116924,41.41949,45.105236,39.11549,29.814156,22.498463,18.635489,15.858873,12.773745,9.8592825,7.6931286,6.3934364,5.61559,4.381539,3.0720003,1.9003079,1.0535386,0.6662565,0.36430773,0.20348719,0.20676924,0.30851284,0.33805132,0.26584616,0.21989745,0.21661541,0.23630771,0.22646156,0.23302566,0.24287182,0.27569234,0.32820517,0.37743592,0.38400003,0.32820517,0.25271797,0.19692309,0.18707694,0.36102566,0.86646163,1.585231,2.228513,2.3368206,3.4756925,4.161641,4.1583595,3.8301542,4.1156926,4.1583595,4.0434875,3.69559,2.8225644,0.90912825,0.26256412,0.12471796,0.16410258,0.20348719,0.2297436,0.24943592,0.27241027,0.30194873,0.3249231,0.34789747,0.37743592,0.40697438,0.43651286,0.446359,0.41025645,0.380718,0.3511795,0.36102566,0.39384618,0.40369233,0.39056414,0.3708718,0.35446155,0.36102566,0.39712822,0.44964105,0.46933338,0.4594872,0.4594872,0.5513847,0.77128214,0.9419488,0.99774367,0.90912825,0.69251287,0.636718,0.56451285,0.51856416,0.4955898,0.44964105,0.42994875,0.446359,0.508718,0.6268718,0.7844103,0.97805136,1.1946667,1.3915899,1.5261539,1.5360001,1.4867693,1.3128207,1.1290257,1.0436924,1.148718,1.3489232,1.657436,1.9561027,2.0939488,1.9003079,1.7887181,1.595077,1.3522053,1.1257436,1.017436,1.2077949,1.5031796,1.7624617,1.913436,1.9200002,1.8740515,1.7690258,1.6278975,1.5097437,1.5031796,1.7723079,2.1070771,2.4549747,2.7011285,2.6354873,15.340309,15.832617,15.330462,14.099693,12.714667,12.068104,12.156719,12.235488,12.35036,12.681848,13.561437,14.119386,13.328411,11.851488,10.144821,8.480822,7.066257,6.442667,6.518154,6.997334,7.3682055,6.7610264,6.5969234,6.298257,5.805949,5.5893335,5.543385,5.5926156,5.221744,4.7228723,5.2020516,5.691077,5.8945646,5.901129,5.733744,5.3727183,5.4974365,5.72718,6.1078978,6.5870776,6.9809237,7.6110773,8.848411,8.914052,7.765334,7.0957956,7.6996927,8.064001,8.149334,7.899898,7.253334,5.832206,4.821334,4.6244106,5.110154,5.6254363,6.186667,6.294975,6.3376417,6.2851286,5.684513,5.3037953,5.1232824,4.844308,4.6802053,5.356308,5.4941545,5.467898,5.6320004,6.012718,6.301539,6.2720003,6.308103,6.2720003,6.38359,7.2270775,6.875898,6.449231,6.242462,6.445949,7.1483083,7.9228725,6.678975,5.3037953,4.604718,4.31918,3.0818465,2.9013336,3.5446157,4.821334,6.5706673,7.781744,7.8539495,7.1581545,6.166975,5.4547696,4.84759,4.7392826,5.668103,7.3025646,8.41518,9.485129,10.788103,11.030975,10.112,9.124104,9.465437,10.049642,9.435898,7.240206,4.128821,4.2929235,6.2752824,9.137232,11.9171295,13.643488,12.301129,10.187488,7.899898,6.186667,5.9634876,5.412103,4.6900516,3.892513,3.2229745,2.989949,2.6617439,2.0611284,1.5753847,1.3883078,1.5097437,1.8412309,1.9790771,1.9331284,1.7132308,1.332513,1.2373334,1.214359,1.276718,1.3357949,1.2176411,1.0404103,0.9517949,1.1355898,1.5721027,2.038154,2.3466668,2.3466668,2.2055387,2.041436,1.9364104,1.9987694,2.0578463,2.2219489,2.540308,3.0030773,3.3345644,3.56759,3.6463592,3.5840003,3.4494362,3.879385,4.2568207,4.2272825,3.8432825,3.5872824,3.0424619,2.1398976,1.7427694,2.1366155,3.0227695,4.450462,5.1626673,5.431795,5.3924108,5.044513,4.0500517,3.05559,2.156308,1.4998976,1.2865642,1.5261539,1.8773335,2.2580514,2.4746668,2.2350771,2.550154,3.1245131,3.5216413,3.5774362,3.3936412,3.2131286,3.7842054,4.420923,4.923077,5.58277,6.774154,6.232616,5.333334,4.8771286,5.0904617,4.007385,2.868513,1.7460514,0.92553854,0.8992821,0.79097444,0.6268718,0.32164106,0.013128206,0.06235898,0.10502565,0.14112821,0.19692309,0.256,0.256,0.16738462,0.1148718,0.07548718,0.04266667,0.0,0.0,0.0,0.0,0.01969231,0.10502565,0.0951795,0.059076928,0.02297436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01969231,0.03938462,0.01969231,0.016410258,0.02297436,0.07876924,0.16410258,0.2297436,0.15753847,0.09189744,0.055794876,0.07876924,0.18707694,0.446359,0.54482055,0.7187693,1.1716924,2.0545642,2.6584618,2.6945643,2.3433847,1.8576412,1.5885129,1.8838975,2.7175386,3.0949745,2.8488207,2.6518977,3.0818465,3.6791797,3.620103,2.878359,2.2449234,2.8455386,3.0194874,2.793026,2.3236926,1.8970258,2.1169233,2.3105643,2.3236926,2.169436,2.0118976,3.1803079,3.698872,3.2164104,2.1530259,1.7099489,2.4155898,3.1770258,3.9614363,4.5062566,4.325744,2.4451284,1.0568206,0.43651286,0.4135385,0.36430773,0.23630771,0.40697438,0.9321026,1.591795,1.8674873,2.4549747,2.481231,2.169436,1.6147693,0.79097444,0.4135385,0.318359,0.47589746,0.8467693,1.3620514,1.3161026,0.82379496,0.36430773,0.14769232,0.12143591,0.19364104,0.33476925,0.5218462,0.65641034,0.5513847,0.43323082,0.3052308,0.18707694,0.11158975,0.12143591,0.14441027,0.15753847,0.13456412,0.07876924,0.02297436,0.01969231,0.036102567,0.049230773,0.049230773,0.049230773,0.049230773,0.04594872,0.04266667,0.049230773,0.08205129,0.14441027,0.18379489,0.21661541,0.24287182,0.23302566,0.128,0.07876924,0.068923086,0.0951795,0.16082053,0.18379489,0.18051283,0.13128206,0.06564103,0.06564103,0.1148718,0.098461546,0.072205134,0.059076928,0.068923086,0.06564103,0.08533334,0.12471796,0.16410258,0.16082053,0.08861539,0.11158975,0.12143591,0.08205129,0.03938462,0.036102567,0.04594872,0.098461546,0.19692309,0.29538465,0.37743592,0.52512825,0.97805136,1.6246156,1.972513,1.5261539,1.2307693,1.2438976,1.5983591,2.1858463,2.2416413,2.1792822,1.972513,1.6672822,1.3718976,1.9593848,2.1300514,2.0118976,1.9922053,2.7503593,3.6102567,3.387077,2.6551797,1.9331284,1.6804104,1.8346668,2.3630772,3.062154,3.498667,2.989949,3.4724104,4.7458467,5.868308,6.009436,4.4438977,3.3936412,3.4855387,3.5905645,3.3969233,3.4133337,3.2820516,3.006359,2.5238976,2.0151796,1.8970258,1.9167181,2.2383592,2.8225644,3.5347695,4.1517954,4.3552823,3.9318976,3.4067695,3.117949,3.2131286,3.1245131,3.2000003,3.8137438,5.4186673,8.549745,11.237744,11.730052,10.085744,7.138462,4.4898467,3.8038976,4.1124105,5.3202057,7.0531287,8.67118,7.6176414,6.196513,5.3398976,5.4153852,6.242462,7.273026,7.686565,8.205129,8.92718,9.350565,10.134975,11.283693,12.432411,13.321847,13.781334,14.194873,14.838155,16.000002,17.611488,19.22954,22.081642,26.978464,33.631184,40.697437,45.810875,39.51262,30.503387,23.112207,18.825848,16.269129,13.37436,10.732308,8.388924,6.5280004,5.4974365,4.4012313,3.2131286,2.1202054,1.3062565,0.9321026,0.57764107,0.33476925,0.29210258,0.40697438,0.49887183,0.42338464,0.32820517,0.29210258,0.33476925,0.41682056,0.44307697,0.44964105,0.44307697,0.46933338,0.6104616,0.72861546,0.65312827,0.47261542,0.3446154,0.46933338,1.0371283,2.103795,3.4560003,4.5423594,4.466872,3.882667,4.391385,5.044513,5.228308,4.650667,3.7316926,2.986667,2.409026,1.7526156,0.5415385,0.15097436,0.06235898,0.08533334,0.118153855,0.14441027,0.16410258,0.18707694,0.20020515,0.2100513,0.23958977,0.27569234,0.31507695,0.3511795,0.37415388,0.36430773,0.33476925,0.31507695,0.3249231,0.35446155,0.36430773,0.3249231,0.29210258,0.26256412,0.24943592,0.27897438,0.318359,0.3511795,0.36102566,0.36102566,0.41025645,0.5021539,0.5907693,0.61374366,0.5513847,0.41682056,0.3708718,0.3446154,0.3446154,0.37415388,0.42338464,0.46276927,0.512,0.5677949,0.63343596,0.7384616,0.9156924,1.1323078,1.3522053,1.5163078,1.5589745,1.4998976,1.3489232,1.214359,1.1684103,1.2471796,1.4145643,1.591795,1.7132308,1.7296412,1.6311796,1.7920002,1.7755898,1.5130258,1.1388719,0.97805136,1.1290257,1.3718976,1.6869745,1.9954873,2.162872,2.2514873,2.2153847,2.1530259,2.1366155,2.2186668,2.5042052,2.7766156,2.9472823,2.9604106,2.7995899,15.579899,16.475899,16.502155,15.589745,14.145642,13.046155,12.970668,13.6467705,14.14236,14.093129,13.702565,12.980514,12.475078,12.173129,11.802258,10.824206,9.314463,8.434873,8.664616,9.524513,9.5835905,8.753231,8.454565,8.306872,8.004924,7.3058467,6.442667,5.861744,5.4449234,5.3037953,5.7403083,5.7074876,5.464616,5.3103595,5.2742567,5.1200004,5.2480006,5.4875903,5.9503593,6.744616,7.958975,8.644924,9.777231,9.872411,8.815591,7.890052,7.9491286,8.224821,8.300308,8.077128,7.748924,7.6209235,7.181129,6.9021544,6.820103,6.557539,7.0957956,7.430565,7.2861543,6.7577443,6.301539,5.3103595,5.293949,5.152821,4.7983594,5.1659493,5.8781543,5.7042055,5.717334,6.3573337,7.4240007,8.986258,9.511385,9.334154,8.871386,8.635077,7.2992826,5.901129,5.5565133,6.3343596,7.269744,7.177847,6.2916927,5.4547696,5.041231,4.9460516,4.70318,4.8344617,5.58277,6.961231,8.736821,10.348309,9.508103,7.6701546,6.0192823,5.47118,4.3585644,4.414359,5.6320004,7.463385,8.845129,9.747693,10.857026,10.880001,9.833026,9.058462,8.87795,9.26195,8.592411,6.564103,4.164923,3.3575387,3.9154875,5.4153852,7.325539,9.032206,8.704,7.9425645,7.2927184,7.3682055,8.845129,9.53436,9.173334,7.453539,5.172513,4.2305646,3.7842054,2.9440002,2.15959,1.7165129,1.7362052,2.5238976,2.8291285,2.7076926,2.2613335,1.6311796,1.3751796,1.4211283,1.6475899,1.8281027,1.6508719,1.5655385,1.5097437,1.5360001,1.8051283,2.5993848,3.2196925,3.4789746,3.3444104,2.9702566,2.6912823,2.5304618,2.169436,1.8674873,1.782154,1.9462565,2.5271797,3.0293336,3.3411283,3.259077,2.484513,2.7864618,3.1967182,3.4625645,3.498667,3.3805132,2.9801028,2.3171284,2.3368206,3.1507695,4.020513,4.896821,5.159385,4.9985647,4.5587697,3.9154875,2.8455386,2.0151796,1.4441026,1.1913847,1.3489232,1.4145643,1.5983591,1.8346668,1.9495386,1.6475899,1.9035898,2.3991797,2.4976413,2.5764105,4.0041027,5.654975,5.8781543,5.182359,4.273231,4.0500517,5.9602056,5.031385,3.6463592,3.1803079,3.9811285,3.9253337,3.2787695,2.225231,1.2176411,0.9747693,0.69907695,0.446359,0.21661541,0.059076928,0.072205134,0.072205134,0.029538464,0.032820515,0.0951795,0.14112821,0.18051283,0.16410258,0.15425642,0.17066668,0.190359,0.03938462,0.0,0.0,0.006564103,0.036102567,0.036102567,0.013128206,0.013128206,0.02297436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.052512825,0.08205129,0.06235898,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.029538464,0.118153855,0.15425642,0.1148718,0.049230773,0.06564103,0.13128206,0.2297436,0.3117949,0.28225642,0.23630771,0.256,0.30194873,0.36102566,0.44307697,0.7417436,0.9747693,1.2471796,1.7657437,2.8160002,3.249231,3.0523078,2.5304618,2.0086155,1.8149745,2.7470772,4.020513,4.1813335,3.1671798,2.3269746,3.2328207,4.397949,4.9296412,4.5062566,3.4067695,3.6660516,3.3805132,2.9669745,2.5731285,2.0939488,1.9232821,1.8182565,2.0217438,2.428718,2.5895386,2.930872,3.242667,2.9472823,2.2678976,2.2350771,2.5862565,3.2295387,4.1485133,4.8640003,4.4045134,2.4648206,1.0929232,0.48246157,0.4397949,0.4004103,0.30194873,0.27897438,1.1027694,2.3335385,2.3138463,1.9823592,1.8149745,1.5885129,1.1913847,0.6432821,0.26256412,0.21333335,0.42994875,0.7811283,1.079795,1.0994873,0.77456415,0.43323082,0.26584616,0.3249231,0.36102566,0.4201026,0.6170257,0.8467693,0.77128214,0.5940513,0.48902568,0.40697438,0.35774362,0.39056414,0.42338464,0.36758977,0.24615386,0.118153855,0.04594872,0.029538464,0.032820515,0.036102567,0.032820515,0.02297436,0.02297436,0.026256412,0.032820515,0.052512825,0.108307704,0.190359,0.23958977,0.24615386,0.2100513,0.15097436,0.0951795,0.108307704,0.13784617,0.16082053,0.17394873,0.190359,0.20020515,0.16082053,0.101743594,0.108307704,0.15097436,0.12471796,0.08533334,0.06564103,0.06564103,0.055794876,0.06564103,0.08533334,0.10502565,0.11158975,0.16082053,0.23302566,0.24287182,0.17066668,0.06564103,0.055794876,0.06564103,0.1148718,0.18707694,0.24615386,0.3052308,0.4397949,0.88287187,1.4834872,1.6968206,1.1651284,0.79097444,0.86646163,1.3883078,2.0250258,1.9954873,1.7952822,1.5031796,1.204513,1.020718,1.332513,1.9987694,2.4910772,2.6683078,2.7864618,3.7448208,3.6332312,2.937436,2.1464617,1.7723079,1.463795,1.522872,1.9987694,2.6256413,2.8192823,3.495385,4.716308,5.5597954,5.3070774,3.4560003,2.7798977,3.190154,3.6069746,3.5741541,3.2656412,2.930872,2.477949,2.038154,1.9429746,2.7273848,3.0490258,3.255795,3.5249233,3.826872,3.948308,3.7284105,2.993231,2.2744617,1.8937438,1.9790771,2.3827693,2.9538465,3.9975388,5.937231,9.3078985,11.493745,11.608616,9.915077,7.2927184,5.2447186,4.9854364,5.622154,6.954667,8.628513,10.154668,9.124104,7.138462,5.789539,5.586052,5.9503593,6.6822567,6.885744,6.918565,7.0400004,7.4207187,8.572719,10.177642,11.940104,13.51877,14.513232,15.2155905,15.927796,17.240616,19.137642,20.982155,23.785027,28.2519,34.254772,40.592415,44.996925,38.944824,30.447592,23.017027,18.189129,15.537232,13.298873,11.1294365,8.822155,6.6002054,5.1167183,3.9811285,2.9735386,2.2088206,1.6935385,1.3259488,0.8467693,0.42994875,0.27897438,0.39384618,0.58092314,0.61374366,0.5907693,0.5546667,0.5415385,0.571077,0.67938465,0.7122052,0.6859488,0.6629744,0.7581539,0.9156924,0.8763078,0.71548724,0.57764107,0.69579494,1.5195899,3.062154,4.824616,6.12759,6.11118,4.57518,4.6080003,5.2742567,5.691077,5.0116925,3.7743592,2.3893335,1.2832822,0.5973334,0.2100513,0.12143591,0.101743594,0.12143591,0.15425642,0.18051283,0.16410258,0.15097436,0.13784617,0.13456412,0.15425642,0.17066668,0.190359,0.21333335,0.23958977,0.27241027,0.27241027,0.27897438,0.28882053,0.29210258,0.27241027,0.23630771,0.2100513,0.18707694,0.18707694,0.24615386,0.30194873,0.3511795,0.37415388,0.3708718,0.37743592,0.39384618,0.39384618,0.3708718,0.32820517,0.27241027,0.22646156,0.21661541,0.23302566,0.27897438,0.3708718,0.49230772,0.5907693,0.6629744,0.7089231,0.7450257,0.86317956,1.0535386,1.2931283,1.5195899,1.6508719,1.6508719,1.5524104,1.4309745,1.332513,1.2964103,1.3620514,1.3883078,1.3784616,1.3456411,1.3226668,1.4933335,1.5327181,1.3554872,1.0633847,0.94523084,1.0666667,1.2668719,1.5622566,1.9068719,2.1891284,2.3893335,2.5304618,2.6322052,2.7142565,2.806154,3.0030773,3.1803079,3.2262566,3.1409233,3.0293336,14.808617,14.759386,14.87754,14.592001,13.827283,13.016617,12.685129,13.74195,14.575591,14.263796,12.557129,10.840616,10.939077,11.874462,12.698257,12.4685135,11.664412,10.932513,11.336206,12.521027,12.708103,12.911591,12.816411,12.711386,12.511181,11.766154,10.322052,9.088,8.155898,7.683283,7.893334,7.634052,7.322257,7.02359,6.8529234,6.9743595,7.1154876,6.941539,6.961231,7.7423596,9.924924,10.066052,9.170052,8.027898,7.1548724,6.7905645,6.7872825,7.506052,8.119796,8.306872,8.231385,9.911796,10.226872,9.613129,8.536616,7.4863596,7.77518,7.532308,6.4557953,5.2644105,5.681231,5.5630774,5.2020516,4.663795,4.325744,4.890257,5.691077,5.366154,5.3169236,6.173539,7.7981544,10.843898,11.769437,11.542975,10.555078,8.605539,7.0465646,5.986462,5.674667,6.058667,6.764308,6.550975,6.2129235,6.1538467,6.5247183,7.2369237,8.116513,8.480822,9.15036,10.223591,11.093334,11.513436,9.147078,6.5411286,5.100308,5.097026,3.9253337,4.132103,5.346462,6.99077,8.283898,8.769642,9.340718,9.209436,8.4512825,8.008205,8.021334,8.454565,7.955693,6.370462,4.7655387,4.0041027,2.989949,2.4155898,2.5238976,3.1277952,3.515077,4.325744,5.287385,6.4754877,8.320001,10.354873,11.224616,9.731283,6.7150774,5.0543594,4.017231,3.1540515,2.4451284,2.0020514,2.0676925,2.7470772,3.0916924,2.9801028,2.4582565,1.7526156,1.467077,1.8084104,2.349949,2.7011285,2.5173335,2.9144619,3.0982566,2.9440002,2.7831798,3.4198978,4.31918,5.0871797,5.211898,4.7261543,4.2305646,3.7316926,3.0523078,2.3794873,1.8707694,1.6443079,2.4418464,2.993231,3.2262566,3.05559,2.3762052,2.4516926,2.6683078,2.9669745,3.1376412,2.8356924,2.6289232,2.553436,3.2032824,4.384821,5.1167183,5.353026,4.9920006,4.204308,3.1934361,2.2121027,1.522872,1.1651284,0.98133343,0.98461545,1.3522053,1.083077,1.211077,1.6771283,2.0742567,1.654154,1.4375386,1.401436,1.7001027,2.793026,5.4514875,7.8014364,7.4863596,5.756718,3.8334363,2.9046156,4.8672824,4.5029745,3.5774362,3.0227695,2.9440002,3.2656412,2.8389745,1.9167181,0.97805136,0.73517954,0.508718,0.318359,0.23958977,0.25271797,0.24287182,0.18707694,0.10502565,0.08205129,0.128,0.18379489,0.3052308,0.36102566,0.38728207,0.41025645,0.42994875,0.11158975,0.03938462,0.055794876,0.055794876,0.0,0.0,0.0,0.029538464,0.059076928,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.101743594,0.17066668,0.13784617,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.059076928,0.318359,0.42338464,0.2855385,0.06564103,0.15097436,0.32164106,0.4955898,0.5874872,0.48246157,0.5284103,0.62030774,0.71548724,0.8041026,0.9124103,1.2176411,1.5688206,2.0118976,2.6223593,3.501949,3.636513,3.0654361,2.412308,2.048,2.1103592,3.5872824,4.844308,4.919795,3.7809234,2.3269746,4.210872,6.1440005,6.7872825,5.8781543,4.240411,3.626667,3.4067695,3.4691284,3.511795,3.0358977,1.9561027,1.401436,1.719795,2.5829747,3.0096412,2.8225644,2.6223593,2.3269746,2.041436,2.0676925,2.3236926,3.2032824,4.1846156,4.5456414,3.3805132,2.477949,1.204513,0.571077,0.6695385,0.6629744,0.5481026,0.3446154,1.0404103,2.15959,1.7493335,1.4998976,1.4933335,1.2996924,0.86317956,0.48902568,0.3117949,0.40697438,0.72861546,1.0436924,0.9288206,0.7581539,0.6662565,0.5316923,0.41025645,0.5218462,0.46933338,0.4594872,0.5677949,0.7056411,0.64000005,0.52512825,0.5284103,0.58420515,0.6826667,0.86974365,0.90256417,0.7220513,0.51856416,0.36430773,0.2297436,0.128,0.09189744,0.08205129,0.068923086,0.04266667,0.03938462,0.02297436,0.01969231,0.04266667,0.09189744,0.18051283,0.21989745,0.19364104,0.12143591,0.06564103,0.03938462,0.13456412,0.25928208,0.3052308,0.16738462,0.108307704,0.09189744,0.11158975,0.15753847,0.22646156,0.25928208,0.2231795,0.16738462,0.128,0.13784617,0.10502565,0.08205129,0.072205134,0.07876924,0.10502565,0.28225642,0.44964105,0.5021539,0.41025645,0.2231795,0.17394873,0.16410258,0.15753847,0.14112821,0.118153855,0.0951795,0.26912823,0.72861546,1.1782565,0.9353847,0.63343596,0.4004103,0.6235898,1.2274873,1.6607181,1.7132308,1.5589745,1.3357949,1.1979488,1.3226668,1.4834872,2.4451284,3.2295387,3.2229745,2.166154,2.540308,2.7044106,2.5731285,2.2219489,1.910154,1.4703591,1.1093334,1.1782565,1.6804104,2.2547693,2.8225644,3.8400004,4.266667,3.7251284,2.4910772,2.1136413,2.6912823,3.5183592,3.9811285,3.5511796,2.7208207,1.8215386,1.3029745,1.6377437,3.31159,3.9056413,4.013949,4.07959,4.0369234,3.308308,2.4943593,1.5819489,1.0896411,1.1749744,1.6344616,2.5895386,3.639795,4.886975,6.49518,8.700719,9.091283,8.956718,8.641642,8.237949,7.5881033,7.893334,8.717129,9.724719,10.745437,11.798975,11.188514,8.825437,6.8660517,6.193231,6.426257,7.4863596,7.2631803,6.961231,7.171283,7.8736415,9.31118,11.221334,13.436719,15.409232,16.210052,15.724309,15.776822,16.705643,18.58954,21.215181,25.416206,30.624823,36.867287,42.578056,44.596516,39.171284,30.516516,22.852924,17.88718,14.811898,12.78359,10.939077,9.028924,7.0400004,5.1954875,3.7349746,2.7766156,2.3236926,2.1366155,1.723077,1.0896411,0.49887183,0.26256412,0.39056414,0.61374366,0.7450257,0.79425645,0.761436,0.67938465,0.5874872,0.79097444,0.88287187,0.9124103,0.92225647,0.9485129,1.0502565,1.1224617,1.1454359,1.1093334,0.99774367,1.7296412,3.2984617,4.97559,6.189949,6.5050263,5.9963083,5.8978467,5.868308,5.681231,5.2348723,4.2863593,2.8324106,1.463795,0.571077,0.3446154,0.27897438,0.25928208,0.26256412,0.27897438,0.2986667,0.21989745,0.13128206,0.08205129,0.07876924,0.08205129,0.08533334,0.09189744,0.11158975,0.14769232,0.20348719,0.23630771,0.256,0.24943592,0.2100513,0.14112821,0.128,0.118153855,0.12143591,0.15753847,0.26584616,0.36102566,0.43323082,0.446359,0.40369233,0.36758977,0.32820517,0.25928208,0.2100513,0.190359,0.18379489,0.16738462,0.16738462,0.18707694,0.2297436,0.29210258,0.49887183,0.6465641,0.74830776,0.79425645,0.7581539,0.83035904,1.024,1.3161026,1.6246156,1.8051283,1.8510771,1.8346668,1.7329233,1.5753847,1.4309745,1.3456411,1.2570257,1.1848207,1.1388719,1.0994873,1.014154,0.9616411,0.9353847,0.92553854,0.8960001,1.0010257,1.1881026,1.4408206,1.7427694,2.0578463,2.3368206,2.674872,2.934154,3.0720003,3.1343591,3.2229745,3.3312824,3.4067695,3.4560003,3.5544617,10.620719,9.399796,8.910769,9.015796,9.291488,9.048616,8.083693,7.2303596,7.5421543,8.822155,9.6295395,10.325335,11.369026,12.245335,12.786873,13.154463,13.3251295,11.884309,10.535385,10.253129,11.290257,13.282462,14.565744,15.140103,14.930053,13.794462,12.035283,10.197334,8.907488,8.549745,9.245539,10.345026,11.21477,11.264001,10.597744,10.023385,10.20718,9.055181,8.310155,8.996103,11.414975,10.167795,8.933744,7.785026,7.1680007,7.890052,8.218257,8.704,10.125129,11.867898,11.9171295,11.185231,10.59118,9.53436,8.146052,7.27959,8.04759,8.4512825,8.54318,8.329846,7.781744,6.8430777,6.744616,7.3485136,8.100103,8.024616,7.4896417,6.9349747,6.9087186,7.1515903,6.5772314,6.038975,6.3540516,7.4469748,8.973129,10.315488,10.778257,9.649232,8.2215395,7.240206,6.8955903,6.764308,7.6176414,9.222565,10.676514,10.420513,10.725744,11.234463,11.690667,11.762873,11.030975,9.324308,6.5050263,4.2371287,3.1540515,2.8980515,3.9253337,4.381539,4.522667,4.5095387,4.4242053,5.3037953,6.117744,6.8266673,7.2992826,7.325539,7.3353853,7.2664623,6.9382567,6.0619493,4.240411,2.861949,3.3969233,4.397949,4.923077,4.532513,2.1267693,2.2678976,2.8947694,2.8521028,1.8609232,1.8379488,2.0611284,2.481231,2.8947694,2.930872,2.7208207,2.3302567,1.6475899,0.92225647,0.761436,1.020718,1.4966155,1.6410258,1.3489232,0.94523084,0.65312827,1.1749744,1.847795,2.284308,2.3958976,3.8367183,4.634257,4.8114877,4.312616,3.006359,3.639795,4.9427695,5.9503593,6.242462,5.9503593,5.366154,4.788513,4.1583595,3.5249233,3.0358977,2.9636924,3.1737437,3.3936412,3.4625645,3.3411283,2.5961027,2.0808206,1.782154,1.6869745,1.785436,2.409026,3.259077,4.1452312,4.8738465,5.2644105,5.1167183,4.240411,2.9801028,1.7001027,0.74830776,0.67610264,1.2242053,1.4802053,1.339077,1.5097437,0.75487185,1.0305642,2.1103592,3.058872,2.228513,1.8740515,1.6935385,1.3751796,1.4211283,3.1442053,4.9854364,5.402257,4.2469745,2.1858463,0.67282057,1.4900514,1.6016412,1.7132308,2.1267693,2.7634873,1.9692309,1.2931283,0.8041026,0.74830776,1.5425643,1.1881026,0.5415385,0.39384618,0.6826667,0.48902568,0.20676924,0.23958977,0.2855385,0.256,0.24287182,0.318359,0.380718,0.4004103,0.35774362,0.25928208,0.18707694,0.20348719,0.27897438,0.28225642,0.0,0.0,0.0,0.02297436,0.049230773,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02297436,0.049230773,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.4135385,0.74830776,0.67610264,0.029538464,0.21333335,0.44307697,0.6859488,0.81066674,0.58092314,0.6170257,0.761436,0.8960001,1.0338463,1.3259488,1.6804104,1.972513,2.428718,3.0030773,3.3575387,3.0030773,2.8947694,2.8422565,2.733949,2.5632823,4.076308,4.6834874,4.525949,3.9745643,3.629949,6.806975,10.115283,9.419488,5.3398976,3.2656412,2.7273848,3.318154,4.342154,5.100308,4.8672824,2.3401027,1.5064616,1.4998976,1.8379488,2.412308,3.4231799,3.4034874,2.5304618,1.6180514,2.1070771,2.789744,3.6463592,4.716308,5.3234878,4.089436,2.2580514,1.0305642,0.8467693,1.3587693,1.4178462,1.2373334,0.7515898,0.45292312,0.47917953,0.6268718,1.6738462,1.8838975,1.4080001,0.65969235,0.3052308,0.5973334,1.2931283,2.5862565,3.6496413,2.6256413,1.148718,0.81394875,0.72861546,0.508718,0.28882053,0.16738462,0.4955898,0.8041026,0.8369231,0.51856416,0.33476925,0.22646156,0.20676924,0.39384618,0.9911796,1.0535386,0.93866676,0.9878975,1.1093334,0.7778462,0.37415388,0.256,0.22646156,0.190359,0.15097436,0.128,0.08533334,0.049230773,0.029538464,0.029538464,0.09189744,0.1148718,0.10502565,0.07548718,0.07548718,0.101743594,0.18051283,0.4004103,0.62030774,0.47261542,0.21661541,0.12471796,0.19692309,0.38400003,0.58092314,0.702359,0.5481026,0.36102566,0.27241027,0.32164106,0.25928208,0.19692309,0.12471796,0.055794876,0.029538464,0.2855385,0.5973334,0.761436,0.7220513,0.56451285,0.41682056,0.35446155,0.3249231,0.28882053,0.2297436,0.108307704,0.0951795,0.12471796,0.15425642,0.15425642,0.16410258,0.36102566,0.702359,1.024,1.0371283,0.96492314,0.90912825,0.93866676,1.1388719,1.6016412,2.4681027,3.9122055,4.125539,2.9604106,1.9232821,2.3269746,2.4549747,2.3269746,1.9364104,1.2504616,1.0568206,0.85005134,0.6859488,0.7187693,1.204513,1.595077,1.9331284,2.097231,2.172718,2.4418464,2.9046156,3.4527183,4.2436924,5.0904617,5.431795,4.4077954,2.878359,1.7985642,1.723077,2.8225644,2.3827693,2.428718,2.8258464,2.8947694,1.404718,0.84348726,0.6826667,0.7384616,0.96492314,1.463795,2.428718,4.017231,5.4153852,6.2588725,6.636308,6.1505647,7.463385,9.235693,10.676514,11.58236,12.6063595,13.174155,13.3940525,13.7386675,15.044924,13.5548725,10.95877,8.237949,6.1472826,5.218462,5.0477953,5.1987696,6.373744,8.39877,10.194052,10.791386,11.332924,12.425847,14.418053,17.394873,17.112617,17.319386,18.021746,19.46913,22.15713,27.283695,33.765747,41.64267,48.416824,49.027287,43.982773,34.162876,25.770668,20.78195,16.938667,13.433437,11.395283,9.826463,8.185436,6.377026,4.6080003,3.5347695,3.0523078,2.809436,2.2121027,1.4309745,0.7318975,0.46933338,0.61374366,0.74830776,0.77128214,0.6695385,0.5415385,0.45292312,0.4266667,0.52512825,0.67610264,0.8960001,1.1946667,1.5721027,1.595077,1.7952822,2.1070771,2.281026,1.8773335,2.2678976,3.0227695,3.895795,4.9920006,6.774154,8.421744,9.137232,8.470975,6.698667,4.8049235,3.4888208,2.3433847,1.4572309,0.88287187,0.6268718,0.5415385,0.46276927,0.39056414,0.33476925,0.33476925,0.22646156,0.07876924,0.006564103,0.02297436,0.04594872,0.059076928,0.098461546,0.14769232,0.19364104,0.2297436,0.23958977,0.22646156,0.19692309,0.15097436,0.09189744,0.07876924,0.08533334,0.098461546,0.13128206,0.2297436,0.31507695,0.36430773,0.3511795,0.29210258,0.24287182,0.20676924,0.15097436,0.1148718,0.108307704,0.12143591,0.13456412,0.128,0.13456412,0.17066668,0.24287182,0.49887183,0.67282057,0.761436,0.7318975,0.5481026,0.6235898,0.81394875,1.1815386,1.595077,1.7558975,1.8412309,1.9790771,2.0184617,1.9200002,1.785436,1.6016412,1.4736412,1.3653334,1.2570257,1.1585642,0.9878975,0.892718,0.8598975,0.8730257,0.88615394,0.92225647,1.0305642,1.3259488,1.7394873,2.044718,2.3138463,2.5895386,2.8488207,3.0720003,3.2820516,3.4264617,3.4921029,3.626667,3.9220517,4.4110775,13.804309,12.527591,11.0145645,9.544206,8.326565,7.4863596,7.1187696,7.3419495,8.155898,9.386667,10.689642,11.474052,11.930258,11.897437,12.018872,13.764924,14.647796,14.168616,12.36677,10.089026,8.996103,9.337437,10.66995,11.956513,12.688411,12.891898,12.852514,13.594257,14.815181,16.039387,16.607182,15.2155905,14.326155,14.319591,15.100719,16.128002,17.142155,17.792002,17.204514,15.724309,14.930053,13.712411,12.763899,11.575796,10.049642,8.474257,9.028924,9.403078,9.780514,9.974154,9.426052,8.910769,8.523488,8.090257,7.5421543,6.8988724,6.5280004,6.196513,6.235898,6.554257,6.6592827,6.304821,6.426257,6.944821,7.6242056,8.086975,7.8145647,7.6964107,7.77518,7.860513,7.5421543,8.379078,9.29477,9.058462,7.88677,7.433847,7.194257,6.416411,5.6254363,5.044513,4.6145644,4.276513,4.2502565,4.9526157,6.4623594,8.530052,9.186462,9.898667,10.7158985,11.890873,13.863386,13.453129,11.480617,8.933744,6.7216415,5.6943593,5.5762057,5.7042055,5.927385,6.160411,6.377026,6.7282057,6.518154,6.3474874,6.5870776,7.3714876,6.1440005,5.8518977,6.5444107,7.1483083,5.474462,3.764513,2.5140514,2.3433847,2.878359,2.7503593,2.0250258,3.0752823,4.1714873,4.453744,3.9253337,2.806154,2.2711797,2.228513,2.5928206,3.2820516,2.7142565,2.1825643,1.7099489,1.332513,1.1060513,0.84348726,0.5677949,0.4955898,0.6071795,0.65312827,0.69251287,1.3029745,1.7690258,1.847795,1.7723079,3.3214362,4.089436,4.309334,4.128821,3.6036925,4.522667,5.8880005,7.394462,8.4283085,8.086975,7.24677,6.232616,4.97559,3.7120004,2.9997952,3.0424619,3.114667,3.242667,3.4231799,3.623385,3.3575387,2.930872,2.5435898,2.3729234,2.5796926,3.1507695,3.7054362,3.9417439,3.9056413,3.9942567,4.082872,4.066462,3.4100516,2.2186668,1.2373334,0.79097444,0.6170257,0.51856416,0.4594872,0.58420515,0.49887183,0.85005134,1.4736412,1.8838975,1.2865642,1.5688206,1.8773335,1.2996924,0.41682056,1.2865642,2.0578463,2.481231,2.1989746,1.4539489,1.1224617,2.0086155,1.9692309,1.6114873,1.2537436,0.9321026,1.017436,0.9124103,0.64000005,0.38728207,0.5284103,0.58420515,0.60389745,0.6268718,0.60061544,0.36758977,0.16410258,0.190359,0.2297436,0.20348719,0.17066668,0.16738462,0.21661541,0.2855385,0.33805132,0.35774362,0.30194873,0.24615386,0.19364104,0.13784617,0.06235898,0.06235898,0.07548718,0.055794876,0.009846155,0.0,0.0,0.029538464,0.029538464,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.0032820515,0.006564103,0.006564103,0.0,0.0,0.0,0.0,0.0,0.013128206,0.06235898,0.08205129,0.32164106,0.67610264,0.86974365,0.45620516,0.54482055,0.80738467,1.0010257,1.020718,0.88615394,0.8533334,0.99774367,1.0535386,0.99774367,1.0469744,1.585231,2.162872,2.6518977,2.9669745,3.0752823,2.9571285,3.0096412,3.2295387,3.511795,3.6726158,3.7907696,3.501949,2.8521028,2.28759,2.6190772,4.1124105,5.1889234,4.8049235,3.3280003,2.5206156,2.8127182,2.9965131,2.986667,2.7864618,2.487795,1.8149745,1.6147693,1.719795,2.048,2.5829747,3.058872,3.0490258,2.6289232,2.1267693,2.1169233,2.3138463,3.0194874,3.6824617,3.895795,3.4067695,1.8182565,0.8730257,0.5284103,0.6662565,1.0896411,0.96492314,0.71548724,0.44964105,0.34133336,0.61374366,1.1848207,1.6738462,1.5360001,0.955077,0.8533334,1.6049232,1.4802053,1.5983591,2.2022567,2.6617439,2.0906668,1.8313848,1.522872,1.1290257,0.9485129,0.9156924,1.014154,1.0075898,0.81066674,0.4955898,0.28225642,0.20020515,0.22646156,0.34789747,0.56451285,0.6268718,0.5940513,0.53825647,0.47261542,0.33805132,0.69907695,1.0633847,1.4080001,1.5360001,1.079795,0.69579494,0.38728207,0.23302566,0.2231795,0.26256412,0.3052308,0.27897438,0.2100513,0.12471796,0.07548718,0.09189744,0.16082053,0.3117949,0.49887183,0.5940513,0.56451285,0.571077,0.5874872,0.57764107,0.51856416,0.4266667,0.36758977,0.3446154,0.34133336,0.3314872,0.3511795,0.45620516,0.44964105,0.2986667,0.128,0.14112821,0.17723078,0.24943592,0.37743592,0.60061544,0.8369231,0.88943595,0.7417436,0.48246157,0.31507695,0.19364104,0.15097436,0.15097436,0.16082053,0.14112821,0.17066668,0.29210258,0.4135385,0.48902568,0.5021539,0.6629744,0.6071795,0.5677949,0.76800007,1.4080001,2.3138463,2.9243078,2.5665643,1.6869745,1.8609232,2.176,1.8346668,1.585231,1.6016412,1.4966155,1.3981539,1.2176411,1.1060513,1.1158975,1.1946667,1.6607181,1.7624617,1.6771283,1.6705642,2.0742567,2.2547693,2.4976413,2.7831798,2.9801028,2.8324106,2.3138463,1.8412309,1.8576412,2.3696413,2.9801028,2.7076926,2.172718,1.7493335,1.4736412,1.0502565,0.81066674,0.74830776,0.9156924,1.6049232,3.3444104,4.788513,5.6943593,5.6320004,4.9526157,4.7950773,5.1659493,6.806975,9.248821,11.562668,12.337232,11.001437,10.551796,10.9686165,12.028719,13.334975,12.911591,11.336206,8.470975,5.1954875,3.387077,4.0467696,5.4449234,7.2369237,9.416205,12.304411,14.083283,12.704822,11.605334,12.422565,14.989129,18.927591,20.086155,20.43077,21.523693,24.51036,28.944412,33.920002,39.233643,43.85149,45.925747,41.196312,33.352207,25.93149,20.476719,16.534975,13.636924,12.035283,10.564924,8.694155,6.5247183,4.6178465,3.6562054,3.3312824,3.3247182,3.31159,2.7733335,2.3926156,2.172718,1.9790771,1.529436,1.1913847,1.014154,0.9288206,0.8730257,0.76800007,0.7384616,0.8960001,1.6443079,3.0096412,4.647385,5.07077,4.785231,4.31918,3.9286156,3.5872824,2.8816411,2.6190772,3.121231,4.84759,8.39877,11.385437,12.074668,9.527796,5.0576415,2.2186668,2.041436,1.6607181,1.1913847,0.7811283,0.61374366,0.48902568,0.50543594,0.5677949,0.5546667,0.3117949,0.2100513,0.15425642,0.13456412,0.12471796,0.068923086,0.032820515,0.04594872,0.09189744,0.14769232,0.20348719,0.21661541,0.18707694,0.14112821,0.10502565,0.09189744,0.07876924,0.09189744,0.118153855,0.15425642,0.19364104,0.21989745,0.2231795,0.20676924,0.17723078,0.15753847,0.13128206,0.0951795,0.07548718,0.08861539,0.108307704,0.16082053,0.2231795,0.28225642,0.33805132,0.39056414,0.44307697,0.49230772,0.5021539,0.47261542,0.4135385,0.46933338,0.61374366,0.93866676,1.3193847,1.401436,1.3784616,1.5425643,1.7690258,2.034872,2.409026,2.92759,2.9833848,2.7109745,2.169436,1.3292309,1.1191796,0.99774367,0.8992821,0.82379496,0.8369231,0.90256417,1.0338463,1.3357949,1.7985642,2.28759,2.6453335,2.9669745,3.1934361,3.318154,3.3772311,3.515077,3.751385,4.056616,4.384821,4.6769233,13.824001,13.190565,12.09436,10.663385,9.245539,8.43159,7.8769236,7.9294367,8.674462,9.90195,11.113027,11.30995,11.296822,10.889847,10.410667,10.70277,11.0605135,10.840616,9.826463,8.487385,7.9458466,7.8506675,8.280616,9.110975,10.029949,10.532104,10.9226675,11.723488,12.852514,14.027489,14.775796,13.965129,13.495796,13.574565,14.263796,15.504412,16.239592,16.708925,16.177233,14.890668,14.096412,13.334975,12.373334,11.158976,9.83959,8.766359,9.032206,9.209436,9.258667,9.104411,8.612103,7.972103,7.2237954,6.51159,5.9470773,5.6254363,5.674667,5.786257,6.11118,6.6002054,7.000616,7.1876926,7.3714876,7.6701546,8.080411,8.457847,8.39877,8.021334,7.860513,8.001641,8.109949,8.854975,9.353847,8.933744,7.6110773,6.1013336,5.284103,4.5423594,3.7973337,3.170462,2.989949,3.515077,4.8311796,6.4065647,8.067283,9.961026,10.604308,11.460924,12.314258,13.144616,14.122667,13.548308,12.202667,10.345026,8.664616,8.280616,8.293744,8.454565,8.234667,7.899898,8.523488,9.452309,7.709539,5.917539,5.284103,5.5729237,4.394667,4.1124105,4.598154,5.139693,4.46359,3.6660516,2.9144619,2.7470772,2.9965131,2.7798977,2.8849232,4.1124105,5.356308,6.0160003,5.9963083,5.031385,4.027077,3.2032824,2.6420515,2.3105643,1.847795,1.4408206,1.083077,0.7975385,0.64000005,0.5218462,0.39384618,0.40369233,0.5415385,0.63343596,0.72861546,1.0535386,1.273436,1.3489232,1.5261539,2.7634873,3.6660516,4.2272825,4.4406157,4.3027697,5.028103,5.976616,7.1187696,8.329846,9.38995,8.802463,7.269744,5.3005133,3.5610259,2.8816411,3.1442053,3.3345644,3.9056413,4.857436,5.717334,4.8672824,4.706462,5.2545643,6.6560006,9.16677,9.964309,9.429334,7.194257,4.384821,3.6135387,3.2164104,2.865231,2.3368206,1.6344616,0.98133343,0.51856416,0.40369233,0.4135385,0.45292312,0.52512825,0.79425645,1.0666667,1.2832822,1.3981539,1.3718976,1.2406155,0.99774367,0.512,0.06564103,0.32820517,0.5284103,0.9714873,1.1881026,1.1224617,1.1093334,1.1552821,1.3095386,1.3784616,1.2570257,0.9321026,0.90584624,0.764718,0.512,0.29210258,0.38400003,0.5284103,0.64000005,0.5973334,0.4201026,0.26256412,0.20348719,0.3052308,0.38728207,0.380718,0.33476925,0.318359,0.29210258,0.28225642,0.31507695,0.4004103,0.35774362,0.28882053,0.2100513,0.14769232,0.13128206,0.15425642,0.2100513,0.20020515,0.13128206,0.108307704,0.08861539,0.049230773,0.013128206,0.0,0.0,0.0,0.0,0.009846155,0.02297436,0.0,0.04266667,0.06564103,0.04266667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.0,0.009846155,0.009846155,0.0032820515,0.009846155,0.0032820515,0.026256412,0.026256412,0.029538464,0.15097436,0.21661541,0.3708718,0.702359,1.024,0.86646163,0.58420515,0.6662565,0.9911796,1.2931283,1.1618463,0.94523084,1.0699488,1.2307693,1.2668719,1.1520001,1.4211283,2.0545642,2.868513,3.4822567,3.2820516,2.92759,2.4976413,2.3171284,2.422154,2.5796926,2.5895386,2.1924105,1.8937438,1.9626669,2.4582565,3.05559,2.930872,2.2055387,1.3357949,1.079795,1.3751796,1.5622566,1.6246156,1.5819489,1.5064616,1.5064616,1.6016412,1.8773335,2.3368206,2.8980515,3.3575387,3.3050258,2.92759,2.4155898,1.975795,1.9232821,2.3072822,2.7733335,2.9472823,2.428718,1.5786668,1.2373334,1.1716924,1.3193847,1.7952822,1.7296412,1.1355898,0.5415385,0.256,0.3708718,0.574359,1.0075898,1.3193847,1.5753847,2.2547693,2.3105643,2.169436,2.6289232,3.626667,4.2436924,3.7874875,2.917744,1.9593848,1.2242053,0.9944616,1.0633847,0.97805136,0.892718,0.8566154,0.80738467,0.508718,0.45292312,0.5513847,0.6662565,0.61374366,0.55794877,0.4660513,0.36430773,0.31507695,0.4135385,0.8008206,1.0568206,1.5163078,2.0841026,2.2449234,1.9298463,1.4900514,1.2373334,1.2340513,1.2898463,1.2898463,1.1027694,0.72861546,0.32820517,0.23302566,0.26584616,0.3511795,0.41025645,0.446359,0.5152821,0.58420515,0.6662565,0.7122052,0.69251287,0.6235898,0.41025645,0.3117949,0.28225642,0.28225642,0.27241027,0.36758977,0.5218462,0.61374366,0.63343596,0.67282057,0.6104616,0.36102566,0.18379489,0.20020515,0.41025645,0.67938465,0.7515898,0.69579494,0.5907693,0.5284103,0.38400003,0.29538465,0.2231795,0.190359,0.27569234,0.43651286,0.5513847,0.56123084,0.47917953,0.4135385,0.56451285,0.65312827,0.6432821,0.65641034,0.9747693,1.4276924,1.4834872,1.204513,0.9485129,1.3784616,1.8642052,1.7723079,1.4539489,1.1716924,1.0994873,1.4802053,1.5556924,1.3850257,1.204513,1.4375386,1.8313848,1.6147693,1.2471796,1.086359,1.4145643,2.281026,3.6594875,4.388103,3.9122055,2.3105643,1.5524104,1.4244103,1.9692309,2.8324106,3.2787695,2.868513,2.228513,1.5622566,1.0535386,0.84348726,0.7417436,1.079795,1.9561027,3.318154,4.95918,5.651693,5.989744,5.6418467,4.8804107,4.5817437,5.100308,6.6527185,9.035488,11.398565,12.225642,10.962052,9.961026,9.93477,10.896411,12.156719,11.897437,9.511385,6.567385,4.204308,3.131077,3.8498464,5.346462,7.250052,9.429334,11.989334,13.66318,13.08554,11.920411,11.562668,13.13477,16.656412,19.203283,20.775387,22.075079,24.523489,28.248617,32.11159,35.9319,39.36821,41.928207,39.151592,33.319386,26.74872,21.034668,17.03713,14.299898,12.422565,10.571488,8.448001,6.314667,4.8344617,4.1878977,3.9647183,3.8662567,3.6857438,3.1442053,2.8980515,3.2295387,3.8859491,4.086154,2.9407182,2.0906668,1.5195899,1.1848207,1.0108719,0.9124103,1.0010257,1.6508719,3.0260515,5.097026,5.651693,5.612308,5.425231,5.3005133,5.221744,4.273231,3.4658465,3.2065644,4.138667,7.1548724,9.892103,10.020103,7.788308,4.4242053,2.1398976,1.4441026,1.1158975,0.95835906,0.8598975,0.79425645,0.48246157,0.38728207,0.44964105,0.56123084,0.5349744,0.4660513,0.33476925,0.19364104,0.0951795,0.0951795,0.08205129,0.08205129,0.09189744,0.1148718,0.16082053,0.16738462,0.13128206,0.08861539,0.059076928,0.04594872,0.049230773,0.06564103,0.098461546,0.128,0.14769232,0.128,0.11158975,0.09189744,0.07876924,0.08205129,0.07876924,0.07876924,0.07876924,0.07876924,0.08861539,0.15097436,0.21333335,0.27241027,0.32164106,0.36430773,0.36430773,0.36430773,0.3511795,0.3249231,0.30851284,0.3511795,0.45292312,0.71548724,1.0765129,1.3128207,1.4408206,1.4933335,1.5327181,1.6311796,1.913436,2.5206156,2.7142565,2.5271797,2.0742567,1.5392822,1.2898463,1.1520001,1.0436924,0.9353847,0.8598975,0.86646163,0.955077,1.1716924,1.5458462,2.0742567,2.605949,2.9801028,3.245949,3.4724104,3.7218463,3.7907696,3.9122055,4.0008206,4.0336413,4.059898,10.975181,11.37559,11.175385,10.358154,9.321027,8.884514,8.293744,8.12636,8.674462,9.665642,10.262975,10.348309,10.656821,10.453334,9.668923,8.907488,9.019077,8.408616,7.5388722,6.8299494,6.678975,6.3934364,6.11118,6.265436,6.875898,7.5487185,7.962257,8.4283085,8.986258,9.511385,9.728001,9.586872,9.7903595,10.039796,10.322052,10.919386,10.998155,11.0375395,10.939077,10.912822,11.441232,11.329642,10.71918,9.872411,9.02236,8.36595,8.260923,8.4972315,8.681026,8.592411,8.178872,7.456821,6.5411286,5.7435904,5.330052,5.5269747,5.8223596,6.2194877,6.7150774,7.200821,7.460103,8.100103,8.513641,8.710565,8.707283,8.507077,8.086975,7.3321033,7.1220517,7.6176414,8.264206,8.700719,8.835282,8.641642,7.9524107,6.4656415,5.330052,4.601436,4.0008206,3.6463592,4.076308,5.3234878,7.466667,9.783795,11.621744,12.412719,12.186257,12.544001,13.042872,13.4170265,13.548308,13.042872,12.675283,12.09436,11.349334,10.909539,10.6469755,10.404103,9.833026,9.133949,9.078155,9.330873,7.24677,5.35959,4.604718,4.3290257,3.3476925,3.0490258,3.259077,3.7710772,4.3618464,4.0303593,4.06318,4.4373336,4.955898,5.2447186,5.2676926,5.4941545,5.8092313,6.163693,6.557539,6.2162056,5.077334,3.692308,2.3860514,1.273436,1.5589745,1.273436,0.76800007,0.3446154,0.27569234,0.35446155,0.49230772,0.67610264,0.85005134,0.90256417,0.9419488,1.0075898,1.2274873,1.6278975,2.1431797,2.989949,3.4560003,3.8498464,4.279795,4.6572313,5.2512827,5.917539,6.675693,7.6898465,9.26195,8.94359,7.515898,5.421949,3.501949,3.0227695,3.5774362,4.3716927,5.658257,7.312411,8.809027,8.746667,8.802463,9.426052,11.004719,13.866668,14.506668,13.15118,9.498257,5.0838976,3.2853336,2.3663592,1.8313848,1.463795,1.1191796,0.7187693,0.33805132,0.43323082,0.6268718,0.73517954,0.76800007,0.8992821,0.92553854,0.8763078,0.9288206,1.4276924,1.2964103,0.9288206,0.42338464,0.0,0.0,0.0,0.7089231,1.148718,1.0994873,1.083077,1.0962052,1.2603078,1.401436,1.4244103,1.3029745,0.98461545,0.69907695,0.446359,0.3052308,0.39712822,0.46276927,0.47589746,0.38728207,0.24943592,0.24943592,0.33476925,0.38728207,0.40697438,0.39712822,0.36758977,0.35446155,0.31507695,0.2855385,0.2986667,0.3708718,0.34133336,0.29210258,0.21989745,0.15753847,0.15097436,0.190359,0.25928208,0.2986667,0.29538465,0.29210258,0.24287182,0.09189744,0.0,0.0,0.0,0.0,0.0,0.009846155,0.02297436,0.0,0.04266667,0.08861539,0.06564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.01969231,0.032820515,0.029538464,0.016410258,0.016410258,0.04266667,0.108307704,0.13456412,0.15097436,0.28882053,0.40369233,0.5152821,0.7844103,1.1191796,1.2012309,0.8598975,0.9944616,1.4309745,1.8215386,1.6311796,1.2209232,1.1618463,1.3226668,1.4933335,1.3817437,1.5556924,2.1202054,2.802872,3.2164104,2.858667,2.2908719,1.6443079,1.2504616,1.1946667,1.2898463,1.3751796,1.2635899,1.394872,1.7887181,2.0709746,2.034872,1.5163078,0.8533334,0.35446155,0.3117949,0.39056414,0.56123084,0.7975385,1.0436924,1.2012309,1.3029745,1.585231,2.0611284,2.681436,3.3509746,3.8038976,3.7743592,3.4133337,2.8488207,2.1891284,1.9954873,2.103795,2.3466668,2.4188719,1.8674873,1.4998976,1.847795,2.809436,4.082872,5.1626673,3.3444104,1.8051283,0.76800007,0.29538465,0.2986667,0.256,0.40697438,0.7187693,1.2307693,2.048,1.9298463,2.0676925,2.5895386,3.255795,3.4264617,3.1048207,2.300718,1.4703591,0.9288206,0.8369231,1.0075898,1.1093334,1.2832822,1.4506668,1.2898463,0.9517949,1.083077,1.6672822,2.2580514,1.9987694,1.2012309,0.8205129,0.6432821,0.58092314,0.67282057,0.7975385,0.9485129,1.3718976,2.0020514,2.4484105,2.4484105,2.228513,2.044718,2.028308,2.176,2.2186668,2.038154,1.6344616,1.1848207,1.0371283,0.9682052,0.8795898,0.74830776,0.61374366,0.57764107,0.57764107,0.6071795,0.636718,0.65312827,0.6662565,0.47261542,0.34133336,0.25928208,0.2231795,0.2231795,0.36758977,0.574359,0.73517954,0.8566154,1.0765129,1.394872,1.024,0.51856416,0.2100513,0.23302566,0.37743592,0.41025645,0.41682056,0.43651286,0.45620516,0.39712822,0.38728207,0.36430773,0.36430773,0.51856416,0.7384616,0.8730257,0.88615394,0.78769237,0.6301539,0.6104616,0.64000005,0.5973334,0.51856416,0.57764107,0.76800007,0.7450257,0.6104616,0.60389745,1.0994873,1.6738462,1.7394873,1.4145643,0.98133343,0.8467693,1.332513,1.5097437,1.3587693,1.1126155,1.2668719,1.5097437,1.2504616,0.85005134,0.6170257,0.83035904,1.8609232,3.698872,5.5302567,6.1538467,4.0008206,1.8674873,1.6902566,2.4352822,3.2787695,3.6069746,3.2229745,2.425436,1.5753847,0.9682052,0.83035904,1.2077949,2.1891284,3.6824617,5.142975,5.5696416,5.044513,4.8049235,4.772103,4.903385,5.2020516,5.687795,6.9021544,8.756514,10.709334,11.749744,11.638155,11.136001,10.929232,11.204924,11.644719,10.299078,7.4830775,5.1298466,3.9975388,3.6627696,4.378257,5.8880005,7.8539495,9.961026,11.9171295,13.206975,12.99036,12.173129,11.720206,12.658873,14.854566,17.864206,20.804924,23.299284,25.475285,28.337233,30.84472,33.53272,36.529232,39.53559,39.141747,34.87508,28.977234,23.168001,18.619078,15.796514,13.656616,11.431385,8.969847,6.73477,5.605744,5.0576415,4.7425647,4.397949,3.8498464,3.186872,2.930872,3.6824617,5.1232824,6.0225644,4.59159,3.2164104,2.100513,1.4080001,1.2603078,1.401436,1.8182565,2.4910772,3.3805132,4.4307694,4.2535386,4.0533338,4.2272825,4.7983594,5.405539,5.2578464,4.516103,3.69559,3.5478978,5.0642056,7.525744,7.8441033,6.764308,4.955898,2.986667,1.6180514,1.1355898,1.0896411,1.1552821,1.1290257,0.6859488,0.47589746,0.446359,0.51856416,0.5940513,0.571077,0.47917953,0.42994875,0.46933338,0.5940513,0.42994875,0.23958977,0.11158975,0.07876924,0.0951795,0.098461546,0.08533334,0.072205134,0.055794876,0.02297436,0.029538464,0.049230773,0.072205134,0.09189744,0.108307704,0.07876924,0.055794876,0.036102567,0.026256412,0.026256412,0.036102567,0.049230773,0.052512825,0.052512825,0.059076928,0.10502565,0.14769232,0.18707694,0.22646156,0.27241027,0.3249231,0.34133336,0.32164106,0.28225642,0.23630771,0.24287182,0.33805132,0.5316923,0.8041026,1.1224617,1.3620514,1.5031796,1.4342566,1.2570257,1.2964103,1.6836925,1.9232821,1.9626669,1.8806155,1.8674873,1.5491283,1.3751796,1.2537436,1.1257436,0.94523084,0.88615394,0.9288206,1.079795,1.3489232,1.7690258,2.349949,2.7667694,3.0916924,3.3969233,3.764513,3.8498464,3.892513,3.82359,3.6758976,3.6135387,7.076103,8.162462,8.769642,8.63836,8.083693,8.01477,7.834257,7.8112826,8.2215395,8.845129,8.976411,9.554052,10.555078,10.79795,10.194052,9.728001,10.194052,9.399796,8.103385,6.8627696,6.012718,5.2578464,4.906667,4.8311796,5.0838976,5.8978467,6.117744,6.452513,6.685539,6.5378466,5.664821,5.395693,5.7698464,6.245744,6.491898,6.370462,5.937231,5.789539,6.2194877,7.2960005,8.864821,9.29477,9.088,8.644924,8.116513,7.387898,7.0498466,7.3386674,7.5946674,7.506052,7.138462,6.485334,5.651693,5.349744,5.7534366,6.5083084,6.4557953,6.672411,7.1909747,7.7981544,8.018052,8.595693,9.035488,9.07159,8.615385,7.75877,6.741334,5.8880005,5.8420515,6.5870776,7.4469748,7.778462,7.9294367,7.936001,7.716103,7.066257,6.242462,6.0324106,6.2227697,6.8496413,8.192,9.488411,11.040821,12.885334,14.385232,14.247386,13.026463,12.517745,12.4685135,12.694975,13.069129,13.08554,14.237539,15.297642,15.455181,14.329437,12.675283,11.37559,10.496001,9.69518,8.2215395,6.810257,5.5991797,5.028103,4.9099493,4.457026,3.4789746,3.0162053,3.1934361,4.0369234,5.4580517,5.2053337,5.907693,7.171283,8.628513,9.954462,8.996103,7.3682055,5.8092313,4.916513,5.1298466,5.1265645,4.2436924,2.9801028,1.7263591,0.7844103,1.6475899,1.4408206,0.86974365,0.4660513,0.58092314,0.50543594,0.57764107,0.8008206,1.0535386,1.0962052,1.1290257,1.2176411,1.7558975,2.7044106,3.570872,4.2207184,3.8498464,3.4691284,3.5938463,4.210872,4.903385,5.7501545,6.616616,7.463385,8.329846,8.201847,7.5979495,6.3376417,4.926359,4.5554876,5.3103595,6.9842057,8.923898,10.742155,12.343796,13.686155,13.413745,12.84595,12.796719,13.571283,13.748514,12.324103,9.209436,5.353026,2.7503593,1.5688206,1.276718,1.2242053,1.086359,0.8960001,0.71548724,0.88287187,1.0272821,0.9911796,0.827077,0.5907693,0.5546667,0.60389745,0.71548724,0.9517949,1.3587693,1.529436,1.0765129,0.32820517,0.3314872,0.3249231,1.214359,1.6213335,1.3292309,1.276718,1.847795,1.7165129,1.4080001,1.211077,1.1651284,0.9517949,0.7253334,0.49887183,0.3511795,0.4135385,0.36758977,0.24943592,0.15425642,0.14769232,0.26256412,0.4004103,0.3117949,0.21333335,0.18707694,0.2100513,0.22646156,0.256,0.28882053,0.3052308,0.28225642,0.26584616,0.24287182,0.18707694,0.12143591,0.098461546,0.13784617,0.2231795,0.31507695,0.38400003,0.4135385,0.3708718,0.14441027,0.0,0.0,0.0,0.0,0.0,0.01969231,0.036102567,0.0,0.0,0.04266667,0.04266667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.01969231,0.01969231,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.04266667,0.055794876,0.052512825,0.032820515,0.013128206,0.08205129,0.19364104,0.26912823,0.2986667,0.36430773,0.49230772,0.5874872,0.7778462,1.0732309,1.3653334,1.3751796,1.7296412,2.0742567,2.1891284,2.0118976,1.6147693,1.339077,1.3456411,1.5655385,1.6935385,2.176,2.3860514,2.284308,1.9659488,1.6705642,1.142154,0.7515898,0.5481026,0.51856416,0.6104616,0.61374366,0.8205129,1.086359,1.270154,1.2176411,0.764718,0.37415388,0.26256412,0.39384618,0.45620516,0.3708718,0.39056414,0.54482055,0.8041026,1.0666667,1.2077949,1.6836925,2.3630772,3.1343591,3.8990772,4.204308,4.194462,3.8859491,3.3378465,2.6486156,2.2514873,2.1333334,2.0709746,1.9068719,1.5524104,1.3423591,2.0578463,3.8465643,6.1997952,7.939283,4.3618464,2.28759,1.1618463,0.69579494,0.86974365,0.8533334,0.5021539,0.22646156,0.2231795,0.47261542,1.0666667,1.522872,1.585231,1.2504616,0.7811283,0.7220513,0.63343596,0.53825647,0.49887183,0.60061544,0.86974365,1.4342566,2.2186668,2.8258464,2.540308,2.0676925,2.412308,3.4527183,4.4274874,3.948308,2.2383592,1.4998976,1.2635899,1.2504616,1.3751796,1.3653334,1.522872,1.6410258,1.6705642,1.7099489,2.0151796,2.1300514,2.1891284,2.4516926,3.2853336,5.152821,4.850872,3.4724104,2.1333334,1.9922053,1.8871796,1.657436,1.3587693,1.0962052,1.0371283,0.94523084,0.85005134,0.77128214,0.7253334,0.7417436,0.6892308,0.5907693,0.47261542,0.36758977,0.28225642,0.4955898,0.7450257,0.85005134,0.88943595,1.211077,2.0873847,1.8412309,1.1651284,0.56451285,0.36430773,0.24943592,0.19692309,0.16410258,0.14441027,0.14112821,0.24943592,0.37743592,0.47261542,0.5481026,0.67282057,0.83035904,0.9616411,1.0404103,1.0338463,0.9124103,0.85005134,0.9124103,0.8041026,0.5218462,0.3314872,0.57764107,0.77128214,0.67938465,0.5316923,1.014154,1.4441026,1.3817437,1.1224617,0.8795898,0.78769237,0.9353847,1.0075898,0.9747693,0.85005134,0.6859488,0.79425645,0.8467693,0.7384616,0.57764107,0.6826667,1.4244103,2.7306669,5.21518,7.4141545,5.789539,2.5731285,2.284308,3.0424619,3.7448208,4.0303593,3.751385,2.5435898,1.4769232,1.0765129,1.3259488,2.4057438,3.9187696,5.4383593,6.160411,4.903385,3.5478978,2.9571285,3.3542566,4.535795,5.874872,6.3934364,7.026872,8.185436,9.711591,10.883283,11.572514,12.153437,12.304411,11.956513,11.303386,8.87795,6.744616,5.3694363,4.788513,4.598154,5.4843082,7.213949,9.357129,11.35918,12.540719,13.069129,12.199386,11.766154,12.373334,13.400617,14.749539,17.368616,21.129848,25.091284,27.529848,29.830566,31.271387,33.017437,35.669334,39.27303,40.772926,38.006157,32.958363,27.19508,21.861746,18.661745,16.269129,13.725539,10.81436,8.096821,7.003898,6.2818465,5.7468724,5.1856413,4.342154,3.4560003,3.0326157,3.7973337,5.533539,7.072821,6.547693,4.8640003,3.1245131,2.0020514,1.7657437,2.2514873,3.0949745,3.876103,4.161641,3.5216413,2.356513,1.6344616,1.7985642,2.8553848,4.3716927,5.293949,4.7425647,3.6857438,2.937436,3.170462,5.504,6.705231,6.695385,5.4941545,3.2032824,2.353231,2.0709746,1.9561027,1.785436,1.5097437,0.9944616,0.69579494,0.5481026,0.48574364,0.47589746,0.5152821,0.574359,0.7581539,1.0338463,1.2209232,0.7975385,0.37415388,0.11158975,0.036102567,0.032820515,0.07548718,0.1148718,0.12143591,0.09189744,0.03938462,0.036102567,0.052512825,0.06564103,0.08861539,0.15097436,0.2100513,0.15425642,0.068923086,0.013128206,0.0,0.0,0.0,0.0032820515,0.013128206,0.02297436,0.04266667,0.072205134,0.0951795,0.118153855,0.17723078,0.29538465,0.3446154,0.33476925,0.28225642,0.19692309,0.15425642,0.24943592,0.3708718,0.5021539,0.74830776,0.96492314,1.3489232,1.3751796,1.0699488,1.0108719,1.1618463,1.3620514,1.6508719,2.0053334,2.3466668,2.097231,1.8445129,1.6180514,1.3981539,1.1257436,0.99774367,1.0108719,1.1355898,1.3423591,1.6082052,2.038154,2.412308,2.7437952,3.0490258,3.3641028,3.5446157,3.6463592,3.6890259,3.7448208,3.9351797,5.477744,5.733744,6.889026,7.515898,7.328821,7.171283,7.50277,7.6110773,7.8736415,8.500513,9.537642,10.328616,10.886565,11.113027,11.0605135,10.925949,11.500309,12.356924,12.130463,10.673231,9.065026,7.4896417,7.453539,7.9786673,8.461129,8.681026,7.975385,7.4404106,6.921847,6.1997952,5.0051284,5.028103,5.4843082,6.2588725,6.99077,7.066257,6.6133337,5.786257,5.737026,6.633026,7.643898,8.132924,7.1187696,6.009436,5.677949,6.485334,6.058667,5.5204105,4.9821544,4.647385,4.8082056,4.2338467,3.0818465,3.4921029,5.349744,6.301539,6.229334,6.4754877,7.269744,8.553026,9.993847,9.176616,8.3593855,7.584821,6.806975,5.8912826,5.2545643,4.8049235,4.6211286,4.6276927,4.578462,4.578462,4.7327185,4.768821,4.6966157,4.8082056,5.5269747,7.1089234,9.18318,11.500309,13.932309,14.736411,15.195899,15.133539,14.723283,14.480412,14.076719,13.5089245,13.174155,13.069129,12.786873,12.530872,15.543797,18.569847,19.98113,19.77436,15.894976,13.239796,11.382154,9.846154,8.086975,6.9382567,6.1407185,5.8092313,5.7009234,5.1889234,4.457026,3.7218463,3.5938463,4.197744,5.1889234,6.419693,8.881231,11.628308,14.057027,15.898257,13.164309,9.91836,6.5444107,3.6890259,2.2744617,1.5655385,1.4244103,1.3522053,1.1257436,0.80738467,0.29538465,0.2855385,0.60389745,1.1290257,1.8018463,0.9944616,0.58420515,0.47261542,0.508718,0.47261542,0.69251287,1.1782565,2.2416413,3.764513,5.218462,6.0849237,5.5236926,4.388103,3.2722054,2.5042052,3.3312824,4.850872,6.498462,7.817847,8.454565,8.73354,9.133949,9.7673855,10.194052,9.412924,9.964309,12.150155,14.27036,15.51754,16.006565,15.432206,13.505642,11.575796,10.325335,9.750975,9.957745,9.15036,7.460103,5.093744,2.3335385,1.0666667,0.6301539,0.76800007,1.214359,1.6771283,2.0939488,2.225231,1.8937438,1.1552821,0.28882053,0.13128206,0.9419488,1.8510771,1.8904617,0.0,0.26912823,0.6104616,1.1290257,1.6377437,1.6640002,1.6278975,1.6804104,1.7657437,1.8018463,1.6771283,1.276718,0.8172308,0.446359,0.23958977,0.21333335,0.8598975,1.020718,0.74830776,0.4397949,0.8533334,0.7581539,0.39384618,0.14441027,0.10502565,0.09189744,0.09189744,0.036102567,0.0,0.026256412,0.13784617,0.25928208,0.35446155,0.39712822,0.35446155,0.18379489,0.15753847,0.16082053,0.16082053,0.12143591,0.0,0.0,0.23958977,0.35446155,0.27897438,0.2297436,0.31507695,0.13456412,0.0,0.0,0.0,0.0,0.0,0.09189744,0.18379489,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.04266667,0.10502565,0.09189744,0.01969231,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.15425642,0.25271797,0.21661541,0.108307704,0.21661541,0.30851284,0.45620516,0.72861546,1.204513,1.6082052,1.782154,1.6344616,1.3751796,1.5097437,1.6705642,1.5360001,1.4244103,1.595077,2.2416413,3.2918978,2.4188719,1.273436,0.65641034,0.5349744,0.28882053,0.14769232,0.072205134,0.06235898,0.12143591,0.34133336,0.571077,0.67938465,0.6301539,0.47261542,0.26584616,0.16738462,0.25271797,0.4660513,0.6268718,0.3446154,0.30194873,0.4004103,0.57764107,0.80738467,1.3226668,2.0086155,2.8914874,3.826872,4.4865646,4.6802053,4.417641,3.9318976,3.3312824,2.6256413,1.7591796,1.2668719,0.9321026,0.6498462,0.44307697,0.6498462,0.85005134,1.0633847,1.3817437,1.9692309,2.0676925,1.9265642,1.7591796,1.8707694,2.6387694,3.190154,2.034872,0.88287187,0.44964105,0.47261542,1.6804104,2.5435898,2.9210258,2.6256413,1.404718,1.1093334,0.9911796,0.7187693,0.30851284,0.13784617,0.5021539,1.2898463,2.9440002,4.969026,5.920821,4.8344617,4.97559,5.1889234,4.890257,4.059898,2.6912823,1.9298463,1.8182565,2.3269746,3.3411283,3.7316926,3.6726158,2.8488207,1.6738462,1.2832822,1.5392822,1.4276924,1.782154,3.249231,6.301539,15.05477,13.617231,7.3485136,1.5786668,1.6016412,2.0545642,2.359795,2.2482052,1.9298463,2.0742567,2.1956925,2.1267693,1.8773335,1.5360001,1.2668719,1.401436,1.3981539,1.2570257,0.97805136,0.56451285,0.9911796,1.1257436,0.9353847,0.7844103,1.4178462,2.1891284,2.281026,1.9987694,1.5721027,1.1454359,0.5349744,0.318359,0.23958977,0.16410258,0.09189744,0.23958977,0.3117949,0.32820517,0.32820517,0.36758977,0.4266667,0.50543594,0.58092314,0.67938465,0.8992821,1.4736412,2.5796926,2.5600002,1.2964103,0.19692309,0.40697438,0.55794877,0.636718,0.6235898,0.48902568,0.5481026,0.51856416,0.39056414,0.23958977,0.21333335,0.22646156,0.24615386,0.27897438,0.32164106,0.380718,0.47917953,0.99774367,1.3587693,1.3915899,1.3423591,2.9538465,4.2371287,4.9788723,4.8377438,3.31159,2.5665643,2.4155898,3.045744,4.1156926,4.775385,4.066462,2.28759,1.3259488,1.7624617,2.8980515,4.1550775,5.4416413,6.0816417,5.4908724,3.1573336,2.2908719,2.166154,2.733949,3.9581542,5.8125134,6.413129,6.0750775,6.7117953,8.329846,9.065026,8.710565,9.409642,10.112,10.30236,10.010257,9.363693,8.293744,7.1089234,6.186667,5.9667697,6.9809237,8.661334,10.948924,12.78359,12.100924,10.256411,9.7673855,10.725744,12.593232,14.204719,14.204719,17.135592,21.205336,25.051899,27.726772,30.825027,33.184822,34.54031,35.92862,39.686565,41.970875,41.88226,38.610054,33.043694,27.769438,23.584822,20.256823,17.02072,13.564719,10.023385,8.805744,7.939283,7.3714876,6.806975,5.720616,4.414359,3.5938463,4.0533338,6.012718,9.124104,11.040821,8.664616,5.691077,3.8531284,2.9144619,3.18359,3.5052311,3.6463592,3.4002054,2.5928206,1.9954873,1.6278975,1.4736412,1.9692309,3.9811285,4.4832826,3.1540515,1.8215386,1.339077,1.5721027,2.6945643,4.082872,4.5522056,3.570872,1.2504616,3.3017437,4.1911798,3.9581542,2.937436,1.7558975,1.020718,0.51856416,0.32820517,0.40369233,0.5481026,0.69579494,0.7220513,0.764718,0.83035904,0.79425645,0.37743592,0.15425642,0.04594872,0.009846155,0.04594872,0.20348719,0.318359,0.28225642,0.13784617,0.07548718,0.06564103,0.06235898,0.08533334,0.17723078,0.39712822,0.78769237,0.56451285,0.21661541,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.02297436,0.04266667,0.09189744,0.14112821,0.18051283,0.2100513,0.21989745,0.18379489,0.12143591,0.12471796,0.16082053,0.23630771,0.380718,0.5415385,0.90912825,1.020718,0.8763078,0.9616411,1.1323078,1.2931283,1.7099489,2.359795,2.9440002,3.2623591,2.9013336,2.3466668,1.8576412,1.4802053,1.2242053,1.1782565,1.2635899,1.4375386,1.6935385,1.8412309,1.9331284,2.1464617,2.484513,2.7766156,3.0096412,3.1573336,3.5610259,4.2863593,5.142975,3.8531284,3.1934361,3.370667,4.092718,5.1298466,6.3277955,6.961231,7.1483083,7.240206,7.532308,8.267488,9.275078,10.213744,10.70277,10.551796,9.754257,7.3583593,7.460103,8.454565,8.992821,7.9786673,7.6931286,7.6701546,7.466667,7.1647186,7.3649235,7.4174366,7.1680007,7.020308,7.020308,6.8594875,6.5247183,6.7544622,7.13518,7.253334,6.7117953,6.3573337,6.0160003,5.8847184,5.914257,5.8125134,5.6385646,5.1626673,5.730462,7.3091288,8.474257,8.185436,7.9228725,7.565129,7.0925136,6.5772314,6.6560006,6.3868723,6.124308,6.0652313,6.265436,6.193231,6.11118,6.117744,6.1997952,6.235898,5.8092313,5.3792825,5.356308,5.805949,6.452513,5.72718,5.034667,4.466872,4.197744,4.493129,5.3136415,6.3179493,7.2664623,7.890052,7.8834877,8.464411,11.001437,13.833847,16.009848,17.27672,14.995693,13.899488,13.3251295,12.813129,12.100924,11.579078,11.497026,12.09436,13.000206,13.226667,13.124924,13.446565,14.736411,16.295385,16.17395,12.576821,11.618463,11.208206,10.161232,8.198565,7.4010262,6.7610264,6.311385,5.9569235,5.4941545,4.8771286,4.197744,3.82359,4.059898,5.1265645,7.0531287,9.882257,11.697231,11.733335,10.394258,7.9819493,6.7938466,6.363898,6.2818465,6.2030773,5.533539,4.788513,4.07959,3.3969233,2.5895386,1.7460514,1.0305642,0.6892308,0.7220513,0.88615394,0.71548724,0.702359,0.8041026,0.97805136,1.204513,1.2406155,1.6935385,2.8291285,4.4734364,6.0225644,6.626462,5.970052,4.9854364,4.2601027,4.027077,4.788513,6.6560006,8.241231,8.763078,8.050873,8.165744,9.051898,10.7158985,12.901745,15.090873,16.928822,18.596104,18.848822,17.650873,16.177233,14.588719,14.024206,13.4170265,12.337232,10.971898,9.636104,7.4075904,4.7261543,2.3236926,1.2373334,0.9714873,1.3357949,2.665026,4.0303593,3.2525132,1.9593848,1.522872,1.4572309,1.4178462,1.204513,0.53825647,0.43323082,0.5284103,0.48574364,0.0,0.052512825,0.12143591,0.7778462,1.657436,1.4572309,1.214359,1.1093334,0.79425645,0.36102566,0.33476925,1.2012309,0.636718,0.08861539,0.07548718,0.17723078,0.3249231,0.34789747,0.2297436,0.08861539,0.17066668,0.15097436,0.3052308,0.4266667,0.42994875,0.34789747,0.2100513,0.13784617,0.118153855,0.15097436,0.2100513,0.20676924,0.20348719,0.19692309,0.18707694,0.18379489,0.16738462,0.17394873,0.23630771,0.29538465,0.18379489,0.036102567,0.049230773,0.072205134,0.06564103,0.0951795,0.072205134,0.026256412,0.0,0.0,0.0,0.0,0.0,0.01969231,0.036102567,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.03938462,0.1148718,0.072205134,0.02297436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.29210258,0.36102566,0.30851284,0.2100513,0.118153855,0.2297436,0.446359,0.8008206,1.2242053,1.5360001,1.7033848,1.7165129,1.4966155,1.204513,1.2406155,1.4605129,1.2964103,1.332513,1.8379488,2.7667694,2.353231,1.5458462,0.7318975,0.21333335,0.21661541,0.18707694,0.14769232,0.098461546,0.07548718,0.14769232,0.30851284,0.4135385,0.43323082,0.3708718,0.23958977,0.15097436,0.10502565,0.11158975,0.16410258,0.23630771,0.21661541,0.26912823,0.4266667,0.67282057,0.955077,1.3981539,2.048,2.9013336,3.7907696,4.352,3.95159,3.387077,2.8849232,2.6190772,2.7208207,2.5698464,2.2186668,1.5524104,0.76800007,0.40697438,0.37743592,0.56123084,0.9124103,1.3226668,1.6147693,1.5064616,1.270154,1.1979488,1.4506668,2.0545642,2.300718,1.9790771,1.332513,0.69907695,0.49887183,0.955077,1.4441026,1.5721027,1.5163078,2.0151796,4.056616,10.735591,13.561437,9.780514,2.3827693,1.1290257,0.764718,1.0896411,1.657436,1.7690258,1.9922053,2.7076926,3.9680004,5.031385,4.388103,3.2361028,3.1048207,3.4297438,3.9023592,4.4767184,4.9854364,4.598154,3.636513,2.4681027,1.4998976,1.5031796,1.4539489,1.463795,1.7493335,2.6518977,4.7360005,4.8607183,3.4888208,1.8149745,1.7624617,2.484513,3.446154,3.9712822,3.7874875,3.0260515,2.9636924,3.446154,4.3585644,4.962462,3.9023592,2.8750772,1.8215386,1.2635899,1.2176411,1.1749744,1.2603078,0.9944616,0.6826667,0.7778462,1.8838975,6.813539,7.328821,5.5007186,3.4231799,3.2328207,2.3958976,1.6246156,1.0305642,0.64000005,0.4201026,0.3446154,0.31507695,0.40369233,0.62030774,0.93866676,1.4309745,1.4572309,1.2964103,1.1454359,1.1323078,0.8960001,0.8369231,0.6892308,0.40697438,0.19692309,0.24943592,0.25928208,0.29210258,0.33805132,0.34133336,0.3446154,0.3511795,0.33805132,0.32164106,0.33476925,0.318359,0.28882053,0.26912823,0.28225642,0.3446154,0.48246157,0.761436,1.1060513,1.5655385,2.3072822,3.8006158,5.720616,7.515898,8.746667,9.084719,5.536821,5.0838976,6.4689236,7.9130263,7.1089234,4.630975,2.412308,1.7526156,2.930872,5.169231,6.5345645,5.6943593,4.2601027,2.92759,1.4736412,1.2307693,1.585231,2.3729234,3.4691284,4.788513,5.044513,5.868308,7.968821,10.492719,11.027693,10.55836,9.954462,10.459898,11.943385,12.891898,12.632616,10.512411,8.329846,7.062975,6.882462,7.5421543,9.429334,12.337232,14.116103,10.660104,9.07159,9.435898,10.771693,12.130463,12.619488,12.619488,15.307488,19.295181,23.588104,27.592207,30.280207,32.40698,34.248207,36.63426,40.92062,42.79467,42.184208,38.275284,32.118156,26.660105,22.728207,20.447182,18.166155,15.399385,12.796719,11.808822,11.142565,10.633847,10.003693,8.858257,6.87918,5.648411,5.579488,6.5870776,8.100103,8.326565,6.810257,5.1265645,3.9220517,2.9144619,2.0217438,1.9003079,2.0118976,2.0644104,2.0217438,2.359795,2.5042052,2.409026,2.2350771,2.3335385,1.9954873,1.2603078,0.67610264,0.49230772,0.65641034,1.086359,1.4080001,1.4834872,1.2537436,0.7515898,1.2307693,1.5327181,1.5327181,1.2504616,0.8763078,0.56451285,0.33476925,0.31507695,0.49887183,0.7450257,0.8533334,0.6432821,0.44964105,0.37743592,0.28225642,0.128,0.052512825,0.026256412,0.03938462,0.0951795,0.23302566,0.2986667,0.23302566,0.09189744,0.03938462,0.036102567,0.029538464,0.03938462,0.07876924,0.15097436,0.27897438,0.2100513,0.08861539,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.01969231,0.029538464,0.059076928,0.118153855,0.190359,0.256,0.26912823,0.14769232,0.108307704,0.12143591,0.16082053,0.19692309,0.41682056,0.7253334,0.90912825,0.86317956,0.6071795,0.6235898,0.67282057,0.86646163,1.214359,1.6147693,2.038154,2.3368206,2.5271797,2.5993848,2.5042052,1.9462565,1.6278975,1.591795,1.7460514,1.8773335,1.9856411,2.0512822,2.231795,2.5632823,2.9735386,3.4789746,3.7776413,3.8432825,3.6693337,3.2754874,4.4373336,4.007385,3.6102567,3.5347695,3.9253337,4.781949,5.9963083,6.5903597,6.8430777,7.1023593,7.77518,8.375795,8.828718,9.051898,8.982975,8.582564,7.0400004,7.125334,7.529026,7.3485136,6.0849237,6.245744,6.452513,6.426257,6.2490263,6.3573337,6.0652313,5.8256416,5.989744,6.426257,6.547693,6.3967185,6.3474874,6.3507695,6.304821,6.0652313,5.989744,6.1538467,6.3540516,6.422975,6.242462,5.805949,5.5663595,6.262154,7.529026,7.899898,7.6143594,7.387898,7.0465646,6.633026,6.3868723,6.705231,7.076103,7.1614366,6.9054365,6.521436,6.0324106,5.796103,5.786257,5.924103,6.0816417,6.1046157,6.11118,6.6100516,7.4043083,7.571693,6.5050263,5.5729237,5.2578464,5.802667,7.197539,7.315693,7.7423596,8.457847,9.051898,8.717129,8.297027,9.110975,12.212514,16.571077,19.055592,19.27877,19.882668,19.032618,16.331488,12.852514,12.580104,11.949949,11.365745,10.8996935,10.289231,9.370257,8.5661545,8.743385,9.672206,10.026668,9.035488,9.304616,9.67877,9.504821,8.618668,7.748924,6.9776416,6.413129,6.170257,6.38359,6.229334,5.9602056,5.737026,5.737026,6.1538467,6.8562055,7.8473854,8.41518,8.155898,6.994052,5.3891287,4.7261543,4.778667,5.287385,5.9602056,6.0192823,5.756718,5.2742567,4.768821,4.529231,3.9876926,2.9965131,2.169436,1.6869745,1.3062565,0.9419488,0.92553854,1.079795,1.3161026,1.654154,2.3302567,3.2951798,4.70318,6.636308,9.081436,8.989539,7.2927184,5.536821,4.59159,4.6834874,5.8978467,8.149334,10.095591,10.994873,10.7158985,8.861539,8.569437,9.5606165,11.585642,14.404924,16.843489,18.658463,18.625643,16.873028,14.8939495,13.138052,12.882052,12.694975,11.904001,10.59118,8.408616,5.7698464,3.117949,1.1158975,0.6498462,1.6049232,2.4615386,2.8291285,2.678154,2.3466668,1.7624617,1.1782565,0.90912825,0.93866676,0.9124103,0.35446155,0.47261542,0.6892308,0.6170257,0.06564103,0.48902568,0.92553854,1.6246156,2.172718,1.4769232,1.0896411,1.1618463,0.9124103,0.318359,0.09189744,0.49230772,0.23630771,0.0,0.013128206,0.06564103,0.07548718,0.072205134,0.03938462,0.0,0.0,0.0,0.38400003,0.6170257,0.55794877,0.42994875,0.25271797,0.18707694,0.17066668,0.17066668,0.17394873,0.26256412,0.24943592,0.15753847,0.059076928,0.072205134,0.068923086,0.072205134,0.101743594,0.13456412,0.09189744,0.068923086,0.026256412,0.0,0.0032820515,0.02297436,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016410258,0.08533334,0.04266667,0.013128206,0.0,0.0032820515,0.01969231,0.01969231,0.006564103,0.0,0.009846155,0.055794876,0.06235898,0.026256412,0.0,0.049230773,0.24615386,0.58420515,0.7253334,0.7122052,0.6235898,0.5973334,0.7089231,0.88943595,1.1913847,1.5261539,1.6640002,1.467077,1.2406155,1.086359,1.0994873,1.3686155,1.4309745,1.3620514,1.404718,1.6147693,1.8543591,1.339077,0.8041026,0.41682056,0.24943592,0.30194873,0.34133336,0.28225642,0.190359,0.11158975,0.098461546,0.2231795,0.28882053,0.3052308,0.26256412,0.14769232,0.09189744,0.0951795,0.15097436,0.2297436,0.256,0.2231795,0.24943592,0.36102566,0.56451285,0.827077,1.3259488,1.9790771,2.7011285,3.308308,3.4855387,2.9440002,2.484513,2.353231,2.5961027,3.0752823,3.2918978,3.1113849,2.3762052,1.3259488,0.6170257,0.4201026,0.8205129,1.6016412,2.5173335,3.3017437,3.0030773,2.5074873,1.847795,1.401436,1.8904617,2.162872,2.0578463,1.5524104,0.8763078,0.5316923,0.7253334,1.2865642,1.7001027,1.8904617,2.1956925,3.0096412,6.0619493,7.3714876,5.7665644,2.8980515,2.8882053,4.391385,4.6276927,3.1048207,1.6377437,1.0010257,1.142154,1.9068719,2.7602053,2.7766156,2.2350771,2.353231,2.7175386,3.006359,2.993231,3.5314875,3.7251284,3.495385,2.917744,2.225231,1.9232821,2.2350771,2.3991797,2.2186668,2.041436,2.7044106,2.8488207,2.5206156,2.2613335,3.117949,3.2229745,3.0260515,2.8422565,2.6584618,2.1398976,2.2055387,2.733949,3.3476925,3.5872824,2.9243078,2.300718,1.6607181,1.3226668,1.3653334,1.6475899,2.556718,2.3236926,1.5458462,0.9911796,1.595077,4.9788723,6.701949,7.6931286,8.178872,7.6996927,3.761231,2.3335385,1.9659488,1.7427694,1.2832822,1.0305642,0.85005134,0.77456415,0.84348726,1.1093334,1.3653334,1.3686155,1.2209232,1.020718,0.8598975,0.65641034,0.44964105,0.36758977,0.4594872,0.69251287,0.69907695,0.6104616,0.4660513,0.33476925,0.34133336,0.35774362,0.41025645,0.508718,0.61374366,0.6301539,0.5546667,0.54482055,0.58092314,0.65312827,0.764718,0.81066674,0.86646163,0.98461545,1.2570257,1.8149745,2.8192823,4.204308,5.4875903,6.226052,6.042257,4.4012313,4.9460516,6.6461544,8.257642,8.329846,5.362872,3.7382567,3.8432825,5.0051284,5.5007186,4.972308,3.6529233,2.353231,1.4769232,1.0075898,1.1126155,1.4473847,2.048,2.8192823,3.5347695,3.8662567,5.4383593,7.8670774,10.059488,10.210463,10.075898,10.44677,11.746463,13.328411,13.472821,12.143591,10.121847,8.605539,8.080411,8.320001,8.694155,9.324308,10.213744,10.515693,8.533334,8.838565,9.655796,10.686359,11.536411,11.736616,12.074668,14.020925,17.335796,21.520412,25.846155,29.400618,32.384003,34.845543,37.014977,39.28944,39.939285,38.79713,35.44944,30.559181,25.898668,23.56513,22.54113,21.297232,19.242668,16.722052,14.020925,13.003489,12.632616,12.225642,11.474052,9.31118,7.6668725,6.7314878,6.7183595,7.8441033,7.9786673,7.026872,5.6385646,4.263385,3.1442053,2.1136413,1.6213335,1.4703591,1.4933335,1.5655385,1.7591796,1.8674873,1.8149745,1.6049232,1.3259488,1.3128207,1.2898463,1.0436924,0.69579494,0.702359,0.9353847,0.9419488,0.77456415,0.56123084,0.50543594,0.636718,0.7515898,0.8402052,0.9124103,1.0043077,0.71548724,0.48902568,0.45292312,0.5513847,0.56451285,0.49230772,0.3249231,0.2100513,0.17723078,0.12471796,0.07548718,0.06235898,0.11158975,0.24615386,0.48246157,0.37415388,0.3117949,0.22646156,0.118153855,0.03938462,0.06235898,0.09189744,0.108307704,0.1148718,0.13784617,0.15425642,0.101743594,0.03938462,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.016410258,0.026256412,0.049230773,0.08861539,0.12471796,0.14441027,0.08861539,0.11158975,0.16082053,0.18379489,0.14441027,0.24287182,0.42338464,0.6892308,0.83035904,0.43651286,0.39712822,0.38728207,0.5415385,0.8467693,1.1355898,1.5491283,2.0676925,2.5698464,2.934154,3.0194874,2.5731285,2.1530259,1.8937438,1.8674873,2.0676925,2.1891284,2.1989746,2.2908719,2.5173335,2.802872,3.2000003,3.5741541,3.7284105,3.5478978,3.0096412,4.5423594,4.453744,4.1222568,3.6463592,3.2886157,3.501949,4.673641,5.664821,6.3507695,6.8430777,7.4830775,7.430565,7.026872,6.629744,6.5837955,7.213949,7.53559,8.214975,8.234667,7.4207187,6.445949,6.518154,6.314667,5.930667,5.504,5.1856413,4.9920006,4.97559,5.2676926,5.723898,5.917539,6.1505647,6.232616,6.2162056,6.1472826,6.052103,6.052103,6.442667,6.8594875,7.1089234,7.1483083,7.1187696,6.892308,6.948103,7.273026,7.3452315,7.1220517,6.941539,6.7774363,6.6461544,6.5837955,6.5870776,6.409847,6.294975,6.2162056,5.8880005,5.4449234,5.3202057,5.477744,5.8978467,6.5706673,6.8693337,6.9382567,7.171283,7.532308,7.5421543,6.9776416,6.5870776,6.8430777,7.9228725,9.714872,10.000411,10.597744,11.250873,11.319796,9.777231,9.504821,9.682052,11.82195,15.113848,16.406975,17.293129,18.277744,17.880617,15.707899,12.455385,11.979488,10.873437,9.475283,8.024616,6.6560006,6.3277955,6.1440005,6.2720003,6.633026,6.8955903,7.2960005,7.748924,8.283898,8.707283,8.582564,7.7325134,6.8266673,6.2194877,6.1472826,6.738052,7.194257,7.3747697,7.2992826,7.1023593,7.0400004,6.875898,6.5805135,6.442667,6.3442054,5.737026,4.8082056,4.7327185,4.716308,4.4964104,4.325744,4.890257,4.9985647,4.6966157,4.2830772,4.2962055,4.0500517,3.436308,2.9407182,2.6945643,2.4582565,2.1924105,2.028308,1.910154,1.8313848,1.8379488,2.484513,3.9253337,6.0816417,9.091283,13.305437,13.02318,10.774975,7.837539,5.5269747,5.1856413,6.2227697,7.9885135,9.580308,10.499283,10.640411,8.369231,7.6668725,8.119796,9.462154,11.572514,13.699283,15.287796,15.363283,14.057027,12.609642,11.54954,11.641437,11.690667,11.0605135,9.6754875,6.5345645,4.023795,2.0775387,0.8598975,0.75487185,1.7033848,2.3204105,2.028308,1.2307693,1.3161026,1.4276924,1.0962052,0.81394875,0.73517954,0.65641034,0.16082053,0.51856416,0.96492314,1.0994873,0.86974365,1.3292309,1.6607181,1.8116925,1.7099489,1.2570257,0.9485129,0.892718,0.7220513,0.39056414,0.17723078,0.10502565,0.032820515,0.0,0.02297436,0.108307704,0.02297436,0.0,0.0,0.029538464,0.14112821,0.16082053,0.4004103,0.48574364,0.35446155,0.26584616,0.2100513,0.18707694,0.16410258,0.13128206,0.08205129,0.24287182,0.26256412,0.17723078,0.052512825,0.0,0.0,0.0,0.0,0.0,0.0,0.052512825,0.026256412,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.06564103,0.03938462,0.013128206,0.006564103,0.01969231,0.01969231,0.01969231,0.013128206,0.01969231,0.036102567,0.055794876,0.18051283,0.16738462,0.12143591,0.18707694,0.56451285,0.7778462,0.82379496,0.79425645,0.761436,0.7450257,0.7975385,1.0305642,1.2996924,1.4867693,1.5097437,1.0732309,0.90912825,1.1257436,1.5819489,1.8970258,1.6377437,1.4145643,1.3817437,1.404718,1.0666667,0.67282057,0.39384618,0.29538465,0.33476925,0.38728207,0.40369233,0.30851284,0.19364104,0.108307704,0.072205134,0.13784617,0.17394873,0.18707694,0.17066668,0.108307704,0.0951795,0.10502565,0.17723078,0.27897438,0.3052308,0.2100513,0.190359,0.24615386,0.3708718,0.571077,1.1454359,1.7887181,2.3958976,2.7667694,2.6190772,2.2022567,2.1103592,2.425436,3.0326157,3.6069746,3.6890259,3.4198978,2.733949,1.8149745,1.1060513,0.827077,1.1520001,1.972513,3.0785644,4.1550775,4.089436,3.5282054,2.8160002,2.3696413,2.681436,2.4385643,2.1530259,1.6804104,1.0896411,0.67282057,1.1388719,2.034872,2.7470772,2.9604106,2.6518977,2.0939488,1.4539489,1.142154,1.3981539,2.284308,2.9604106,4.716308,5.182359,4.1156926,3.4133337,1.8543591,1.1618463,1.0338463,1.270154,1.7526156,1.8018463,1.719795,1.7657437,1.9265642,1.9495386,2.605949,3.2065644,3.4034874,3.131077,2.6026669,2.1136413,2.4418464,2.7503593,2.6584618,2.2383592,2.8816411,3.0654361,3.121231,3.436308,4.450462,4.017231,2.6289232,1.6049232,1.3128207,1.1684103,1.204513,1.4342566,1.522872,1.3915899,1.214359,1.1355898,1.0502565,1.017436,1.1290257,1.5130258,2.5435898,2.553436,2.0053334,1.4933335,1.7427694,3.1967182,4.896821,7.0859494,9.508103,11.385437,9.409642,10.220308,9.682052,7.0400004,4.919795,3.9581542,2.868513,2.9702566,4.273231,5.4908724,3.4756925,2.3302567,1.5819489,1.0338463,0.7515898,0.6826667,0.64000005,0.6695385,0.827077,1.1815386,1.4309745,1.3751796,1.0929232,0.75487185,0.6170257,0.571077,0.63343596,0.75487185,0.8566154,0.8336411,0.9517949,1.3686155,1.9068719,2.3302567,2.3401027,2.0086155,1.7427694,1.8182565,2.2711797,2.9078977,3.2196925,3.7448208,4.2371287,4.325744,3.5282054,4.089436,5.58277,6.9021544,7.571693,7.7390776,6.0291286,5.218462,5.481026,5.986462,4.8836927,2.9833848,1.9364104,1.3883078,1.1979488,1.4112822,1.7296412,2.03159,2.4713848,3.0293336,3.5347695,3.7973337,4.9887185,6.872616,8.730257,9.380103,9.435898,10.410667,11.848206,13.046155,13.065847,11.680821,10.125129,9.199591,9.117539,9.501539,9.701744,9.852718,9.396514,8.3823595,7.460103,8.52677,9.728001,10.827488,11.608616,11.884309,12.5374365,14.024206,16.551386,19.830154,23.056412,27.188515,31.855593,36.102566,39.13518,40.31344,39.926155,37.586056,33.988926,29.902771,26.154669,25.281643,24.530054,23.250053,21.238155,18.73395,16.039387,14.890668,14.391796,13.978257,13.413745,11.487181,9.412924,7.748924,7.0104623,7.6668725,7.9852314,7.3616414,6.1013336,4.644103,3.5774362,2.9604106,2.4615386,2.1070771,1.8937438,1.7920002,1.5885129,1.4769232,1.3456411,1.1585642,0.9321026,1.0469744,1.2242053,1.1290257,0.8172308,0.7318975,0.90256417,0.8992821,0.7318975,0.5284103,0.5316923,0.8992821,1.6672822,2.3630772,2.6322052,2.2350771,1.5097437,0.8763078,0.574359,0.69579494,1.1881026,1.3357949,1.1946667,1.0108719,0.8730257,0.69907695,0.3314872,0.19692309,0.27897438,0.55794877,0.9878975,1.0075898,0.88943595,0.64000005,0.52512825,1.0601027,1.1749744,0.8041026,0.4201026,0.22646156,0.16082053,0.13128206,0.07548718,0.029538464,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.016410258,0.04594872,0.059076928,0.059076928,0.04594872,0.032820515,0.032820515,0.08205129,0.13456412,0.16082053,0.13128206,0.13456412,0.21333335,0.43651286,0.6432821,0.42994875,0.4201026,0.42994875,0.574359,0.8533334,1.1355898,1.4342566,1.8445129,2.359795,2.8947694,3.2918978,3.186872,2.8356924,2.428718,2.1431797,2.1792822,2.2482052,2.2153847,2.2121027,2.294154,2.4484105,2.7241027,3.1081028,3.3444104,3.318154,3.0523078,3.892513,3.8564105,3.8629746,3.5478978,3.0391798,2.9440002,3.4034874,4.348718,5.3136415,6.055385,6.564103,6.121026,5.225026,4.381539,4.20759,5.4153852,6.764308,8.1066675,8.635077,8.470975,8.648206,8.388924,7.397744,6.196513,5.149539,4.4307694,4.8771286,5.1987696,5.4383593,5.6418467,5.865026,6.2523084,6.705231,6.997334,7.059693,6.961231,6.8365135,7.000616,7.138462,7.197539,7.3714876,8.041026,7.9425645,7.512616,7.213949,7.522462,7.3091288,7.128616,7.13518,7.2237954,7.02359,6.6133337,5.5105643,4.818052,4.844308,5.100308,5.3103595,5.586052,6.012718,6.701949,7.75877,8.149334,8.100103,7.7325134,7.4010262,7.702975,8.2904625,9.015796,9.829744,10.683078,11.510155,12.3306675,13.348104,14.01436,13.636924,11.362462,12.553847,13.522053,13.892924,13.426873,11.989334,10.489437,9.688616,9.80677,10.348309,10.112,9.209436,8.165744,7.1548724,6.163693,4.95918,6.0258465,7.1614366,7.9425645,8.103385,7.5421543,7.3386674,7.138462,7.2631803,7.6012316,7.6110773,7.2270775,6.6100516,6.0717955,5.8912826,6.304821,7.712821,8.448001,8.579283,8.326565,8.077128,8.0377445,7.6931286,7.256616,6.8004107,6.2588725,5.786257,6.3310776,6.1407185,4.7360005,2.9210258,3.3476925,3.3509746,3.0129232,2.5435898,2.284308,2.3204105,2.5829747,3.0523078,3.5380516,3.6529233,3.7054362,3.4724104,3.0523078,2.550154,2.0611284,1.9003079,3.2984617,6.0324106,10.125129,15.845745,16.577642,15.113848,11.569232,7.525744,6.0291286,5.910975,6.2752824,6.747898,7.0957956,7.2369237,6.705231,6.948103,7.6964107,8.776206,10.108719,10.998155,11.497026,11.23118,10.43036,9.941334,9.941334,10.59118,10.86359,10.180923,8.4053335,4.414359,2.3696413,1.3817437,0.9944616,1.1749744,1.2077949,1.1749744,1.2832822,1.4211283,1.1520001,1.0502565,1.079795,0.99774367,0.7811283,0.63343596,0.51856416,0.86317956,1.2931283,1.7099489,2.300718,2.1858463,1.8346668,1.1913847,0.57764107,0.6826667,0.60389745,0.27569234,0.0951795,0.14112821,0.17066668,0.17066668,0.068923086,0.0,0.04266667,0.21989745,0.04266667,0.0,0.029538464,0.13128206,0.36758977,0.38728207,0.28882053,0.13128206,0.0,0.0,0.128,0.17066668,0.16410258,0.12471796,0.04266667,0.12471796,0.16082053,0.15753847,0.108307704,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.01969231,0.016410258,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.0032820515,0.0,0.0,0.0032820515,0.01969231,0.029538464,0.032820515,0.02297436,0.013128206,0.06235898,0.06235898,0.02297436,0.013128206,0.029538464,0.0,0.0032820515,0.026256412,0.049230773,0.052512825,0.013128206,0.28882053,0.39056414,0.36102566,0.38728207,0.7975385,0.892718,0.7089231,0.6268718,0.71548724,0.7515898,0.7318975,1.0436924,1.2832822,1.2537436,0.9878975,0.5973334,0.8041026,1.5491283,2.3860514,2.4648206,1.8543591,1.2603078,1.0666667,1.1224617,0.76800007,0.37743592,0.25271797,0.24287182,0.26584616,0.29538465,0.26584616,0.18707694,0.12143591,0.098461546,0.108307704,0.09189744,0.07548718,0.068923086,0.07548718,0.09189744,0.13784617,0.128,0.14112821,0.18707694,0.22646156,0.190359,0.21661541,0.2231795,0.2231795,0.318359,0.827077,1.3718976,1.8838975,2.1989746,2.041436,1.8281027,2.0611284,2.6190772,3.3444104,4.0434875,3.9089234,3.508513,2.9440002,2.359795,1.9396925,1.6311796,1.585231,1.9331284,2.6026669,3.3214362,3.623385,3.3378465,3.3214362,3.7415388,4.073026,2.9965131,2.3040001,1.7362052,1.2242053,0.8795898,1.7723079,2.9768207,3.7251284,3.7185643,3.0982566,2.3466668,1.6738462,1.3784616,1.5097437,1.8543591,1.7723079,1.5819489,1.910154,2.930872,4.3716927,3.0523078,2.1989746,1.6377437,1.4112822,1.7558975,2.0841026,1.7624617,1.5195899,1.6738462,2.1530259,2.878359,3.3050258,3.2787695,2.861949,2.3401027,1.9626669,1.972513,2.162872,2.28759,2.0644104,2.4549747,3.045744,3.7743592,4.414359,4.585026,4.0303593,2.4615386,1.2898463,0.9517949,0.90912825,0.7253334,0.5677949,0.44307697,0.36102566,0.3314872,0.39056414,0.512,0.6629744,0.85005134,1.1158975,1.3686155,1.5753847,1.8281027,2.225231,2.8914874,3.9286156,4.3585644,4.768821,6.301539,10.676514,13.863386,17.61477,16.705643,11.533129,8.093539,6.629744,4.9920006,5.5269747,8.093539,10.066052,6.482052,5.225026,3.9056413,2.0512822,1.0896411,0.955077,0.98133343,1.0404103,1.1454359,1.4506668,1.9659488,2.0151796,1.7558975,1.3653334,1.0469744,0.8795898,0.9124103,0.96492314,0.9616411,0.9189744,1.339077,2.2777438,3.4494362,4.4242053,4.6080003,3.9286156,3.508513,3.9351797,5.0576415,5.9536414,5.8256416,5.717334,5.543385,5.146257,4.2896414,5.159385,6.9021544,7.709539,7.171283,6.2752824,6.363898,6.49518,7.066257,7.240206,4.955898,2.8389745,2.1169233,2.0676925,2.294154,2.737231,3.1606157,3.4691284,3.82359,4.2994876,4.890257,4.896821,5.100308,6.12759,7.817847,9.225847,9.170052,9.659078,10.44677,11.34277,12.199386,11.844924,10.768411,10.066052,10.121847,10.624001,10.620719,11.175385,10.8996935,9.531077,7.962257,8.303591,9.737847,11.378873,12.57354,12.898462,13.289026,14.418053,16.196924,18.340103,20.33231,24.192001,30.286772,36.883694,42.2039,44.438976,43.74975,40.323284,35.633232,30.946465,27.32636,26.53867,24.979694,22.89231,20.617847,18.586258,17.624617,16.672821,15.894976,15.317334,14.831591,13.449847,11.300103,9.3078985,8.0377445,7.6635904,7.7390776,7.1515903,6.170257,5.1626673,4.6112823,4.7491283,4.325744,3.5577438,2.7700515,2.3926156,1.9692309,1.6672822,1.394872,1.1257436,0.88615394,0.6859488,0.61374366,0.6071795,0.5973334,0.5152821,0.5940513,0.6104616,0.574359,0.55794877,0.6892308,1.3915899,2.934154,4.1780515,4.3651285,3.1245131,1.9954873,1.0338463,0.7187693,1.3259488,2.9505644,3.436308,3.2754874,2.8816411,2.3794873,1.585231,0.75487185,0.46276927,0.6465641,1.1913847,1.910154,2.2580514,1.847795,1.2964103,1.3161026,2.7273848,2.8521028,1.8609232,0.8369231,0.2855385,0.13128206,0.07876924,0.049230773,0.029538464,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.01969231,0.08533334,0.14112821,0.17066668,0.16082053,0.09189744,0.04594872,0.032820515,0.049230773,0.07876924,0.1148718,0.13456412,0.18379489,0.28225642,0.42338464,0.56451285,0.636718,0.7056411,0.81394875,1.0010257,1.3128207,1.4572309,1.6344616,1.9987694,2.5895386,3.3214362,3.6496413,3.5282054,3.1409233,2.678154,2.3302567,2.2547693,2.162872,2.0742567,2.0250258,2.097231,2.3105643,2.6289232,2.8291285,2.8750772,2.930872,4.6244106,4.598154,4.2272825,3.7087183,3.249231,3.0654361,2.9210258,2.8553848,3.1606157,3.7087183,3.95159,4.0369234,3.9778464,3.7152824,3.3050258,2.9144619,3.5971284,4.6834874,5.9667697,7.3419495,8.818872,8.257642,7.466667,6.5772314,5.858462,5.737026,6.0192823,6.114462,6.2063594,6.3179493,6.3179493,6.1472826,6.3868723,6.9054365,7.6077952,8.438154,8.402052,7.824411,6.9382567,6.2227697,6.3934364,7.017026,7.77518,8.067283,7.778462,7.27959,6.6067696,6.0192823,5.5105643,5.156103,5.080616,5.179077,5.330052,5.6352825,6.1374364,6.820103,7.686565,8.598975,9.819899,11.313231,12.740924,13.216822,13.673027,13.856822,13.525334,12.452104,13.341539,14.54277,15.593027,15.855591,14.5263605,12.816411,11.319796,10.581334,10.752001,11.58236,13.889642,13.988104,13.39077,13.174155,13.991385,12.051693,10.210463,9.068309,8.67118,8.500513,8.2445135,7.6307697,7.397744,7.6307697,7.765334,7.4371285,8.333129,9.31118,9.419488,7.9195905,7.1023593,6.4032826,5.609026,5.034667,5.5236926,6.242462,6.892308,6.547693,5.5958977,5.7074876,8.989539,10.84718,11.736616,11.848206,11.093334,11.142565,10.614155,9.137232,7.529026,7.7981544,7.968821,7.525744,6.0356927,3.8728209,2.2121027,1.9068719,1.8215386,1.7920002,1.719795,1.5885129,2.5632823,3.6594875,4.6966157,5.142975,4.1058464,3.446154,3.3903592,3.3969233,3.2196925,2.9144619,2.4615386,2.9078977,4.4898467,7.460103,12.084514,15.504412,16.439796,14.273643,10.253129,7.506052,5.687795,4.57518,4.201026,4.46359,5.113436,6.370462,7.634052,9.081436,10.804514,12.816411,11.756309,10.381129,8.802463,7.5585647,7.643898,8.096821,8.749949,8.841846,7.965539,6.0717955,2.5829747,1.4080001,1.1323078,1.017436,0.9911796,1.2471796,1.2209232,1.8674873,2.6420515,1.4966155,0.88615394,0.82379496,0.5316923,0.0,0.0,1.9528207,2.6322052,2.9013336,3.1803079,3.4494362,2.5337439,1.8182565,1.3423591,0.88943595,0.0,0.0,0.2100513,0.2100513,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.14769232,0.37743592,0.4266667,0.34133336,0.128,0.0,0.0,0.0,0.108307704,0.21989745,0.2855385,0.2855385,0.21333335,0.04266667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01969231,0.09189744,0.07876924,0.029538464,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.06235898,0.013128206,0.0,0.0,0.01969231,0.09189744,0.14112821,0.17066668,0.108307704,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02297436,0.059076928,0.04594872,0.013128206,0.06235898,0.26912823,0.5218462,0.5940513,0.56451285,0.80738467,1.0404103,0.9419488,1.017436,1.3850257,1.8018463,1.847795,1.8806155,1.7690258,1.270154,0.0,0.0,0.5316923,1.5261539,2.4549747,2.3204105,1.5491283,0.80738467,0.32164106,0.13456412,0.12143591,0.072205134,0.06235898,0.06564103,0.07548718,0.07548718,0.06564103,0.07876924,0.14769232,0.21661541,0.16738462,0.0951795,0.049230773,0.036102567,0.055794876,0.09189744,0.17723078,0.17066668,0.128,0.09189744,0.09189744,0.36102566,0.5907693,0.5316923,0.256,0.18379489,0.29210258,0.5316923,0.8730257,1.2603078,1.6016412,1.467077,1.5458462,1.8609232,2.5665643,3.9220517,4.4701543,4.644103,4.338872,3.7218463,3.2361028,2.8553848,2.6617439,2.4484105,2.172718,1.9528207,1.8084104,2.044718,2.674872,3.6332312,4.8049235,3.9023592,2.7076926,1.6082052,0.93866676,0.97805136,1.6344616,2.7076926,3.2131286,2.9013336,2.2416413,1.719795,1.7624617,2.0906668,2.6617439,3.6627696,3.0030773,2.1431797,1.5064616,1.2340513,1.1585642,1.5983591,2.2383592,2.2777438,1.6705642,1.1454359,1.2800001,1.5327181,1.7755898,1.9692309,2.1530259,2.4681027,2.4188719,1.9856411,1.5097437,1.6935385,1.9003079,1.9364104,1.7887181,1.5491283,1.404718,1.8937438,2.3991797,2.7634873,2.8258464,2.412308,1.8379488,1.4276924,1.2406155,1.214359,1.1913847,1.0075898,0.7318975,0.54482055,0.49230772,0.5021539,0.6498462,0.9616411,1.2800001,1.5064616,1.6180514,1.654154,1.7263591,2.0578463,2.989949,5.0051284,5.5893335,5.5007186,4.394667,2.678154,1.4966155,1.3751796,1.3456411,1.4244103,1.6475899,2.0742567,2.3794873,3.4921029,3.9909747,3.4002054,2.166154,4.571898,9.731283,10.023385,5.080616,1.785436,1.5031796,1.3686155,1.2964103,1.3161026,1.5721027,1.657436,1.6968206,1.6672822,1.5360001,1.2668719,1.1093334,1.0765129,1.0601027,1.0404103,1.1126155,1.3587693,1.9593848,2.917744,4.240411,5.9503593,5.730462,5.9503593,7.171283,8.713847,8.651488,9.078155,8.809027,7.6012316,5.8289237,4.4865646,3.8038976,5.142975,6.669129,7.2631803,6.5312824,6.042257,7.906462,11.497026,13.512206,7.9950776,5.5663595,4.7294364,4.7655387,5.1298466,5.4482055,5.7534366,5.7107697,5.7468724,6.0028725,6.3310776,6.3573337,6.7117953,7.450257,8.237949,8.346257,8.162462,8.2904625,9.035488,10.112,10.650257,10.039796,9.531077,9.849437,11.113027,12.832822,12.2847185,12.11077,11.913847,11.1983595,9.353847,9.547488,10.548513,12.3306675,14.070155,14.145642,12.924719,12.675283,13.548308,15.707899,19.334566,22.50831,27.867899,35.13764,42.584618,47.028515,46.85785,44.708107,40.001644,33.746056,28.534157,25.481848,23.033438,21.11672,19.70872,18.82913,17.69354,16.741745,16.068924,15.819489,16.17395,15.514257,14.378668,12.5374365,10.33518,8.713847,8.018052,7.0104623,6.294975,6.2588725,7.066257,8.346257,7.24677,5.0149746,2.9046156,2.1956925,1.7329233,1.3784616,1.0994873,0.8730257,0.702359,0.58092314,0.55794877,0.60061544,0.636718,0.56451285,0.56451285,0.508718,0.42994875,0.43323082,0.702359,1.4703591,2.028308,1.9495386,1.3062565,0.67282057,0.24287182,0.15425642,1.1126155,3.0982566,5.356308,5.1954875,5.2020516,4.9296412,3.892513,1.5721027,0.9353847,0.86974365,1.4802053,2.6551797,4.059898,3.9975388,2.297436,1.4605129,2.1792822,3.3280003,3.0227695,2.0742567,0.9353847,0.08205129,0.04594872,0.032820515,0.02297436,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.029538464,0.07876924,0.20020515,0.40369233,0.5546667,0.39712822,0.16410258,0.068923086,0.04594872,0.055794876,0.09189744,0.23958977,0.30194873,0.380718,0.5415385,0.80738467,0.9682052,1.0535386,1.1323078,1.2504616,1.4342566,1.5195899,1.6246156,1.8182565,2.1858463,2.806154,3.626667,3.8301542,3.6758976,3.3312824,2.868513,2.5764105,2.3368206,2.1530259,2.0217438,1.9364104,1.9364104,2.0841026,2.3236926,2.6256413,2.989949,4.7327185,4.923077,4.5390773,3.7710772,2.8947694,2.2613335,2.3105643,2.359795,2.481231,2.6551797,2.793026,3.1015387,3.3247182,3.3214362,3.1770258,3.1967182,3.4297438,3.626667,4.309334,5.3891287,6.183385,5.0642056,4.457026,4.128821,3.9417439,3.8695388,3.8006158,3.8301542,4.161641,4.6572313,4.850872,5.1889234,6.121026,7.509334,9.137232,10.709334,11.529847,10.692924,9.051898,7.3419495,6.186667,6.242462,6.6034875,6.9743595,7.2927184,7.7292314,7.9097443,7.450257,7.2960005,7.7423596,8.4512825,8.996103,9.577026,10.226872,11.001437,11.946668,12.668719,13.184001,13.371078,13.4400015,13.961847,14.418053,14.578873,14.116103,13.088821,11.926975,12.386462,13.042872,13.774771,14.477129,15.051488,14.834873,14.480412,14.283488,14.713437,16.403694,18.340103,17.952822,16.728617,15.402668,13.955283,10.41395,8.129642,6.889026,6.5739493,7.1548724,6.9382567,6.482052,6.3540516,6.5444107,6.4722056,6.3474874,7.128616,7.578257,7.177847,6.124308,5.796103,5.3792825,4.9920006,4.9854364,5.9634876,6.058667,5.756718,5.080616,4.585026,5.3760004,7.5388722,9.275078,10.541949,11.30995,11.569232,10.817642,9.6065645,8.03118,6.557539,6.0160003,5.1331286,4.1189747,3.4133337,2.9604106,2.1891284,1.4539489,1.1716924,1.1355898,1.2209232,1.3784616,1.719795,3.3608208,5.717334,7.4404106,6.413129,6.124308,6.1308722,5.4941545,4.4340515,4.3552823,4.9493337,4.7524104,5.2447186,7.020308,9.7903595,10.729027,11.805539,12.524308,11.785847,7.88677,6.1538467,5.7435904,6.744616,8.237949,8.297027,7.181129,7.1581545,7.5552826,8.024616,8.546462,7.90318,7.315693,6.7938466,6.5083084,6.7774363,7.7948723,9.110975,9.222565,7.7292314,5.3398976,2.0545642,0.892718,0.56123084,0.39056414,0.35774362,0.6826667,0.47261542,0.40369233,0.64000005,0.8598975,0.9156924,0.85005134,0.5677949,0.4135385,1.1946667,3.3247182,3.8432825,3.5413337,2.8192823,1.6902566,1.0108719,0.574359,0.32820517,0.23302566,0.28225642,0.4266667,0.5349744,0.47589746,0.29210258,0.19692309,0.20348719,0.14112821,0.059076928,0.0,0.0,0.08861539,0.22646156,0.446359,0.6268718,0.49887183,0.40369233,0.32164106,0.22646156,0.13456412,0.08533334,0.118153855,0.15753847,0.17066668,0.13456412,0.04266667,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.01969231,0.016410258,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.06235898,0.052512825,0.01969231,0.0,0.03938462,0.19692309,0.17723078,0.17723078,0.25271797,0.33476925,0.24943592,0.15097436,0.118153855,0.06564103,0.0,0.0,0.049230773,0.06235898,0.055794876,0.03938462,0.0,0.0032820515,0.03938462,0.03938462,0.0032820515,0.013128206,0.052512825,0.7122052,0.9944616,0.69579494,0.39384618,0.4594872,0.9288206,1.5721027,2.1070771,2.1924105,1.6344616,1.0896411,0.90584624,0.9911796,0.8041026,0.8041026,0.8402052,1.7887181,3.4133337,4.332308,1.8445129,0.636718,0.20676924,0.18707694,0.34133336,0.25271797,0.108307704,0.01969231,0.016410258,0.016410258,0.013128206,0.016410258,0.032820515,0.059076928,0.059076928,0.04266667,0.032820515,0.04266667,0.07876924,0.16410258,0.16082053,0.118153855,0.072205134,0.04594872,0.055794876,0.21661541,0.54482055,0.761436,0.79097444,0.7581539,0.61374366,0.5152821,0.5415385,0.81066674,1.5031796,1.4375386,1.2471796,1.1815386,1.5425643,2.6518977,3.8859491,4.8607183,5.077334,4.4898467,3.501949,2.4910772,2.2744617,2.481231,2.7109745,2.550154,2.0053334,1.6016412,1.9035898,2.8356924,3.69559,3.767795,2.6847181,1.7099489,1.4244103,1.7460514,2.9604106,3.636513,3.761231,3.4822567,3.0982566,2.7667694,2.6683078,3.1245131,3.9614363,4.493129,4.273231,3.6102567,2.9111798,2.3893335,2.0644104,2.5993848,2.8553848,2.7798977,2.5271797,2.4516926,2.4681027,2.5829747,3.1474874,3.9318976,4.1058464,3.7185643,2.733949,1.7952822,1.273436,1.2406155,1.8116925,2.4549747,3.0884104,3.43959,3.0391798,2.9702566,3.0227695,3.190154,3.2689233,2.8750772,2.162872,1.8970258,1.9265642,2.1234872,2.3630772,1.3686155,0.81066674,0.636718,0.7253334,0.892718,1.148718,1.4506668,1.6311796,1.6410258,1.5556924,1.3981539,1.3718976,1.4276924,1.5819489,1.9167181,2.1234872,2.1924105,2.044718,1.6869745,1.2274873,1.2012309,1.3292309,1.6902566,2.1924105,2.550154,2.806154,4.8377438,5.7698464,4.384821,1.079795,1.591795,3.4888208,5.10359,5.3103595,3.5183592,2.740513,2.2678976,1.7985642,1.3686155,1.3522053,1.7394873,1.972513,1.9823592,1.7296412,1.2176411,1.1191796,1.079795,1.0699488,1.1224617,1.3226668,1.6147693,2.0020514,2.7208207,3.5478978,3.8038976,2.7437952,4.128821,6.5083084,8.94359,11.021129,9.816616,8.385642,6.741334,5.940513,8.073847,8.434873,7.5388722,5.8912826,4.1124105,2.930872,3.1737437,3.889231,5.100308,6.232616,6.114462,7.5913854,8.707283,9.222565,9.163487,8.815591,9.317744,10.551796,11.034257,10.627283,10.555078,11.08677,10.65354,10.020103,9.537642,9.140513,7.4929237,6.6822567,6.9842057,7.8441033,7.90318,8.162462,9.005949,9.93477,11.017847,12.895181,15.684924,14.132514,11.83836,10.8996935,11.9171295,13.528616,14.605129,14.916924,14.470565,13.5089245,12.62277,12.320822,12.872206,14.329437,16.538258,19.429745,24.359386,30.5559,37.284107,43.86462,44.320824,43.11303,40.139492,35.285336,28.422565,23.263182,20.309336,18.648617,17.680412,17.132309,16.994463,17.293129,17.70995,18.038155,18.189129,16.787693,15.274668,13.778052,12.393026,11.191795,10.036513,8.585847,7.899898,8.113232,8.418462,8.011488,6.1997952,4.0336413,2.3696413,1.8674873,1.5392822,1.2438976,0.93866676,0.67938465,0.6170257,0.62030774,0.6695385,0.9616411,1.4112822,1.6508719,1.2209232,1.0601027,0.98461545,0.8763078,0.67610264,0.9189744,1.1257436,1.1191796,0.88943595,0.5874872,0.38400003,0.35774362,0.5874872,1.0765129,1.7427694,2.3663592,2.28759,1.8773335,1.394872,0.99774367,0.9485129,0.90256417,0.7811283,0.69579494,0.95835906,1.0338463,0.8172308,0.7253334,0.86646163,1.0568206,0.955077,0.7122052,0.41682056,0.16738462,0.08205129,0.03938462,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.029538464,0.055794876,0.055794876,0.055794876,0.08205129,0.11158975,0.07876924,0.032820515,0.013128206,0.01969231,0.03938462,0.06564103,0.16410258,0.3117949,0.512,0.74830776,0.9682052,1.0075898,0.98461545,0.9911796,1.0633847,1.1782565,1.3029745,1.6869745,1.9889232,2.166154,2.4648206,3.0982566,3.4100516,3.5216413,3.498667,3.3575387,2.937436,2.4910772,2.225231,2.1464617,2.0611284,1.9922053,2.03159,2.3138463,2.8389745,3.4789746,3.8071797,4.397949,4.585026,4.4307694,4.0041027,3.370667,3.131077,2.9702566,2.7700515,2.546872,2.4746668,2.7109745,3.0752823,3.4067695,3.6857438,4.0434875,4.1058464,4.073026,4.2863593,4.7917953,5.349744,4.7655387,4.0434875,3.6332312,3.6135387,3.6693337,3.7743592,3.9712822,4.3552823,4.9526157,5.6943593,6.9776416,8.267488,9.449026,10.8537445,13.226667,14.54277,13.236514,11.096616,9.275078,8.277334,9.888822,10.880001,11.54954,12.07795,12.521027,12.803283,12.560411,12.0549755,11.759591,12.3306675,13.019898,13.213539,13.4400015,13.899488,14.473847,15.304206,15.225437,14.454155,13.4400015,12.875488,12.662155,12.360206,11.949949,11.290257,10.128411,9.429334,9.777231,10.276103,10.57477,10.860309,11.004719,10.811078,10.420513,10.384411,11.657847,13.50236,14.326155,13.971693,12.471796,10.04636,6.3540516,4.7983594,4.535795,5.097026,6.4000006,6.045539,6.2785645,7.145026,8.2904625,8.960001,9.091283,9.245539,9.097847,8.51036,7.53559,6.675693,5.83877,5.225026,5.0543594,5.549949,5.8945646,5.7698464,5.293949,4.7294364,4.5062566,5.3037953,6.6461544,7.5520005,7.722667,7.5421543,6.449231,5.533539,4.604718,3.7120004,3.1343591,2.6223593,2.3630772,2.6617439,3.0916924,2.4746668,1.6705642,1.2012309,1.079795,1.2406155,1.5458462,1.9790771,2.9833848,4.46359,5.989744,6.7872825,6.738052,6.7183595,6.36718,5.8092313,5.6320004,5.9634876,6.157129,6.75118,7.8802056,9.271795,9.485129,10.673231,12.012309,12.09436,8.933744,7.7357955,7.3616414,7.650462,8.155898,8.113232,7.394462,6.921847,6.6625648,6.5936418,6.7249236,7.213949,7.1614366,6.987488,7.2960005,8.89436,9.842873,10.33518,9.298052,7.0498466,5.3136415,3.69559,2.3072822,1.2537436,0.5513847,0.13456412,0.2986667,0.42994875,0.702359,1.1027694,1.4441026,1.1946667,0.78769237,1.0338463,1.8445129,2.228513,2.3926156,2.425436,2.28759,1.9331284,1.3062565,0.82379496,0.44307697,0.190359,0.08533334,0.14112821,0.21333335,0.30851284,0.446359,0.571077,0.53825647,0.33805132,0.20020515,0.101743594,0.036102567,0.0,0.12471796,0.24287182,0.36102566,0.46933338,0.51856416,0.47261542,0.3446154,0.190359,0.06564103,0.04266667,0.049230773,0.055794876,0.055794876,0.03938462,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.04594872,0.059076928,0.06564103,0.06564103,0.06235898,0.055794876,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02297436,0.12143591,0.108307704,0.098461546,0.1148718,0.17723078,0.30194873,0.3052308,0.27569234,0.2231795,0.16410258,0.1148718,0.16410258,0.09189744,0.02297436,0.0,0.0,0.02297436,0.029538464,0.07876924,0.14441027,0.108307704,0.13128206,0.21333335,0.21333335,0.12143591,0.06564103,0.07876924,0.46933338,0.78769237,0.9485129,1.2340513,1.148718,1.3456411,1.7132308,1.9626669,1.6377437,1.1224617,0.74830776,0.65312827,0.761436,0.7975385,0.827077,1.4375386,2.4976413,3.370667,2.9407182,1.2176411,0.39056414,0.098461546,0.08205129,0.15753847,0.118153855,0.068923086,0.036102567,0.02297436,0.0,0.0,0.0,0.0032820515,0.009846155,0.029538464,0.029538464,0.026256412,0.036102567,0.06564103,0.09189744,0.06564103,0.049230773,0.036102567,0.03938462,0.072205134,0.14112821,0.40369233,0.6892308,0.9321026,1.1552821,0.9419488,0.65641034,0.5349744,0.7417436,1.3620514,1.6771283,1.4342566,1.142154,1.142154,1.585231,2.806154,4.0336413,4.8771286,4.916513,3.6890259,2.7963078,2.481231,2.5895386,2.7634873,2.4352822,1.591795,1.1027694,1.3292309,2.2022567,3.2164104,3.6004105,2.934154,1.8707694,1.2931283,2.3236926,3.508513,4.197744,4.31918,4.027077,3.69559,3.1967182,3.2328207,3.7710772,4.525949,4.955898,4.414359,3.8367183,3.498667,3.5446157,3.9811285,4.1911798,3.7349746,3.0687182,2.5042052,2.2186668,2.2219489,2.6715899,3.3050258,3.7120004,3.3575387,2.7437952,1.9823592,1.4605129,1.4080001,1.9068719,3.1737437,4.667077,5.5926156,5.691077,5.2414365,4.916513,4.647385,4.535795,4.535795,4.4373336,3.7284105,3.3476925,3.2722054,3.3247182,3.1770258,2.5895386,2.231795,2.0250258,1.8904617,1.7624617,1.7427694,1.7558975,1.7296412,1.6869745,1.7526156,1.6968206,1.7165129,1.9003079,2.2383592,2.6354873,3.0162053,2.937436,2.7503593,2.5961027,2.4057438,2.484513,2.5337439,2.7208207,3.0687182,3.43959,3.0096412,3.876103,6.229334,8.178872,5.7435904,2.9078977,2.1169233,3.9089234,7.5881033,11.247591,10.433641,8.329846,5.182359,2.6256413,3.6693337,3.8695388,3.387077,2.858667,2.5107694,2.156308,2.2186668,2.231795,2.0808206,1.7755898,1.4736412,1.7427694,2.0873847,2.422154,2.6912823,2.8914874,3.0326157,4.637539,6.6100516,8.333129,9.672206,8.441437,7.062975,6.2687182,6.7117953,8.953437,9.921641,9.120821,7.174565,5.2315903,4.9788723,5.280821,5.609026,5.87159,6.038975,6.166975,7.02359,8.3593855,9.386667,9.777231,9.659078,10.289231,11.08677,11.54954,11.684103,11.995898,12.412719,12.27159,12.022155,11.936821,12.084514,11.644719,10.266257,8.940309,8.03118,7.253334,7.824411,8.874667,10.092308,11.421539,13.082257,14.313026,12.868924,11.378873,11.162257,12.228924,13.709129,15.169642,15.894976,15.458463,13.718975,12.888617,12.688411,12.980514,13.725539,14.985847,17.161848,21.008411,26.65354,33.618053,40.815594,42.003696,41.603287,39.584824,35.649643,29.239798,24.480822,21.540104,19.59713,18.248207,17.513027,17.493334,18.248207,19.111385,19.623386,19.551182,17.77559,16.331488,15.31077,14.539488,13.594257,12.347078,10.916103,9.816616,9.117539,8.464411,7.269744,5.3891287,3.629949,2.4943593,2.1530259,1.7985642,1.4408206,1.0896411,0.8467693,0.8960001,0.9911796,1.1191796,1.2077949,1.2504616,1.3193847,1.2931283,1.4900514,1.5392822,1.2438976,0.5874872,0.5677949,0.61374366,0.64000005,0.6498462,0.7384616,0.69579494,0.5677949,0.7384616,1.332513,2.2383592,3.498667,3.1540515,2.428718,2.1530259,2.7503593,2.1956925,1.3883078,0.7253334,0.6826667,1.8313848,2.6223593,2.156308,1.4145643,0.86974365,0.50543594,0.47917953,0.42338464,0.34133336,0.23958977,0.128,0.06564103,0.026256412,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.02297436,0.01969231,0.006564103,0.0,0.0,0.0,0.0,0.006564103,0.016410258,0.03938462,0.068923086,0.15425642,0.26256412,0.40369233,0.571077,0.7417436,0.85005134,0.9419488,1.020718,1.086359,1.1323078,1.1946667,1.4966155,1.8707694,2.2022567,2.4451284,2.802872,3.0424619,3.2361028,3.4297438,3.626667,3.4297438,3.05559,2.7273848,2.5140514,2.356513,2.2350771,2.2449234,2.481231,2.9636924,3.6660516,3.5938463,3.876103,4.1222568,4.309334,4.3684106,4.194462,4.1485133,4.086154,3.820308,3.3444104,2.8422565,2.6551797,2.7864618,3.2820516,4.007385,4.647385,4.7983594,4.9099493,5.0182567,5.1626673,5.362872,5.533539,5.284103,5.0543594,4.9362054,4.6802053,4.7360005,5.280821,5.7764106,6.186667,6.957949,8.631796,9.83959,10.541949,11.313231,13.331694,14.313026,13.318565,11.894155,10.880001,10.387693,12.27159,13.686155,14.690463,15.363283,15.82277,16.23631,16.15754,15.55036,14.880821,15.133539,15.225437,14.838155,14.598565,14.6182575,14.500104,14.605129,14.158771,13.213539,11.995898,10.886565,10.496001,10.203898,10.098872,9.970873,9.31118,8.146052,7.8539495,7.8473854,7.778462,7.5585647,7.5421543,7.4404106,7.030154,6.521436,6.554257,7.9458466,9.242257,9.580308,8.740103,7.13518,4.818052,3.8104618,3.8662567,4.6572313,5.7632823,5.333334,6.2785645,7.9294367,9.593436,10.55836,10.486155,10.026668,9.429334,8.779488,8.018052,7.056411,6.121026,5.5007186,5.277539,5.356308,5.5597954,5.5630774,5.3037953,4.70318,3.6660516,3.3969233,3.8695388,4.197744,4.0008206,3.4100516,2.4582565,2.0742567,1.8412309,1.5786668,1.3456411,1.2471796,1.4375386,1.9823592,2.481231,2.097231,1.585231,1.2438976,1.2209232,1.4834872,1.8281027,2.3466668,2.8980515,3.5216413,4.352,5.602462,6.51159,7.0793853,7.3353853,7.174565,6.380308,6.160411,6.5903597,7.3616414,8.2904625,9.32759,10.220308,10.935796,11.188514,10.410667,7.7357955,7.515898,7.4174366,7.138462,6.8955903,7.4240007,7.7292314,7.3682055,6.810257,6.426257,6.49518,7.9195905,8.408616,8.5202055,8.92718,10.433641,10.489437,9.826463,8.057437,5.7107697,4.2502565,3.383795,2.2646155,1.3095386,0.6859488,0.318359,0.41025645,0.5874872,0.8598975,1.148718,1.2865642,1.2307693,1.1355898,1.5261539,2.2022567,2.2416413,1.6738462,1.5097437,1.4080001,1.2012309,0.8730257,0.6859488,0.4955898,0.3511795,0.24943592,0.10502565,0.16082053,0.3511795,0.5284103,0.6071795,0.54482055,0.2986667,0.190359,0.14112821,0.10502565,0.06564103,0.0951795,0.128,0.16738462,0.23302566,0.35446155,0.34133336,0.21333335,0.07548718,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.04594872,0.08533334,0.07548718,0.06564103,0.06235898,0.055794876,0.009846155,0.0,0.0,0.0,0.0,0.0,0.02297436,0.06564103,0.12143591,0.16410258,0.11158975,0.08533334,0.07876924,0.0951795,0.15753847,0.15753847,0.18051283,0.23302566,0.2986667,0.33805132,0.34133336,0.29538465,0.18051283,0.059076928,0.049230773,0.16738462,0.12143591,0.07548718,0.06235898,0.0,0.0,0.059076928,0.15425642,0.23302566,0.21989745,0.26584616,0.38728207,0.39712822,0.27241027,0.13128206,0.30851284,0.55794877,0.892718,1.2668719,1.591795,1.5622566,1.8215386,1.8674873,1.5130258,0.88287187,0.6268718,0.56123084,0.58092314,0.6235898,0.67938465,1.5885129,2.8488207,3.5511796,3.1737437,1.6049232,0.65312827,0.19364104,0.026256412,0.0,0.0,0.029538464,0.036102567,0.032820515,0.026256412,0.02297436,0.0032820515,0.0,0.0,0.0032820515,0.01969231,0.02297436,0.016410258,0.01969231,0.032820515,0.01969231,0.0032820515,0.006564103,0.02297436,0.049230773,0.072205134,0.12143591,0.26912823,0.53825647,0.88943595,1.2176411,1.1257436,0.9124103,0.827077,0.9878975,1.3915899,1.9298463,1.7165129,1.2471796,0.8763078,0.80738467,1.6935385,2.8258464,3.8629746,4.3060517,3.4888208,2.9078977,2.6486156,2.681436,2.7700515,2.477949,1.6738462,1.3029745,1.4539489,2.0742567,2.9965131,3.2131286,2.7536411,1.785436,1.079795,2.0118976,3.1113849,4.0041027,4.2896414,3.9680004,3.446154,3.0424619,3.1540515,3.6036925,4.1222568,4.345436,3.761231,3.511795,3.6660516,4.2141542,5.0871797,5.0674877,4.128821,2.92759,2.0184617,1.8707694,2.169436,2.7142565,3.0030773,2.8160002,2.2219489,1.8149745,1.6246156,1.7920002,2.3696413,3.3280003,4.781949,6.23918,7.0432825,7.145026,7.1154876,6.7872825,6.1505647,5.353026,4.7655387,4.9854364,4.9329233,4.5456414,4.1550775,3.7743592,3.1048207,3.3509746,3.4494362,3.2032824,2.7536411,2.5665643,2.5895386,2.7766156,2.8389745,2.7831798,2.934154,3.1606157,3.314872,3.6890259,4.3684106,5.2545643,5.3858466,5.1265645,4.824616,4.818052,5.4186673,5.8912826,5.536821,4.9526157,4.466872,4.1517954,3.2262566,2.802872,4.519385,7.0367184,6.0356927,3.4888208,2.5107694,3.367385,6.055385,10.28595,11.175385,11.21477,9.042052,6.373744,8.001641,8.283898,7.1548724,5.868308,5.034667,4.6244106,4.854154,5.3037953,4.5390773,2.7273848,1.6213335,1.8937438,2.1858463,2.169436,1.972513,2.176,3.4198978,4.8147697,6.0291286,6.8955903,7.4075904,6.4590774,5.4875903,5.9995904,8.060719,10.295795,10.84718,10.121847,8.536616,6.9809237,6.813539,7.141744,7.6603084,7.9950776,7.9491286,7.509334,7.3353853,7.939283,8.907488,9.8592825,10.410667,11.0145645,10.886565,10.850462,11.362462,12.484924,12.829539,13.092104,13.499078,13.974976,14.155488,14.401642,13.650052,11.85477,9.593436,8.021334,8.375795,9.081436,10.315488,11.772718,12.668719,13.331694,13.620514,13.607386,13.410462,13.167591,12.800001,13.522053,14.276924,14.358975,13.3940525,13.249642,13.315283,13.433437,13.810873,14.998976,17.184822,20.617847,25.422771,31.074465,36.4078,37.993027,38.419697,37.231594,34.208824,29.348104,25.508104,23.076105,21.362873,20.01395,19.016207,18.806156,19.295181,19.905643,20.243694,20.059898,18.530462,17.408,16.725334,16.265848,15.553642,14.214565,12.859077,11.58236,10.417232,9.357129,7.9097443,5.865026,4.0402055,2.8717952,2.409026,2.1398976,1.9331284,1.7558975,1.6902566,1.9396925,1.9396925,1.7526156,1.3718976,0.9353847,0.7187693,1.0732309,1.9954873,2.481231,2.0611284,0.81394875,0.48574364,0.4397949,0.58420515,0.8205129,1.0502565,0.9878975,0.75487185,1.1979488,2.5009232,4.1878977,5.093744,4.420923,3.5249233,3.2820516,4.0992823,3.314872,1.9167181,0.9485129,1.0010257,2.1924105,2.986667,2.3696413,1.4178462,0.7253334,0.38400003,0.41682056,0.42338464,0.38728207,0.30851284,0.20020515,0.12471796,0.06564103,0.029538464,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.016410258,0.026256412,0.052512825,0.13128206,0.21989745,0.33805132,0.48574364,0.6301539,0.78769237,0.955077,1.0601027,1.0732309,1.024,1.0305642,1.2931283,1.7296412,2.2022567,2.487795,2.6322052,2.7995899,3.0424619,3.3575387,3.7054362,3.8038976,3.6332312,3.3280003,3.006359,2.7831798,2.6256413,2.5895386,2.7536411,3.1803079,3.9154875,4.3552823,3.9089234,3.7185643,3.761231,3.9712822,4.273231,4.6867695,4.9296412,4.841026,4.3716927,3.564308,3.05559,2.8356924,3.186872,3.9975388,4.7524104,5.1626673,5.540103,5.8092313,5.8945646,5.7042055,6.2785645,6.9120007,7.273026,7.1515903,6.491898,5.986462,6.5050263,7.0859494,7.4174366,7.821129,9.068309,9.944616,10.361437,10.57477,11.201642,11.113027,11.027693,11.142565,11.336206,11.158976,11.493745,12.42913,13.361232,14.040616,14.565744,15.002257,15.209026,15.169642,15.035078,15.117129,14.496821,13.896206,13.51877,13.269335,12.714667,11.736616,11.191795,10.686359,10.006975,9.120821,9.107693,9.229129,9.357129,9.412924,9.363693,8.55959,7.6176414,7.0957956,6.994052,6.7544622,6.564103,6.6494365,6.550975,6.042257,5.146257,5.661539,6.170257,6.413129,6.3573337,6.2063594,5.730462,4.841026,4.4012313,4.644103,5.1856413,5.2512827,6.47877,8.090257,9.4916935,10.249847,9.494975,8.661334,7.88677,7.282872,6.9382567,6.554257,6.1341543,5.9634876,6.0192823,5.9503593,5.356308,5.0642056,4.7425647,4.1025643,2.9013336,2.1825643,1.723077,1.585231,1.5622566,1.1782565,0.7220513,0.6892308,0.78769237,0.88287187,0.9714873,0.9124103,0.98461545,1.1355898,1.2504616,1.1454359,1.0929232,1.1520001,1.404718,1.7985642,2.1530259,2.6223593,3.387077,3.9187696,4.0533338,3.9975388,5.917539,7.4075904,8.28718,8.224821,6.7577443,6.245744,6.432821,6.9677954,7.8047185,9.206155,11.185231,10.660104,9.07159,7.0859494,4.594872,5.3202057,5.7698464,5.7403083,5.7632823,7.1187696,7.9524107,7.939283,7.397744,6.806975,6.7971287,8.356103,9.163487,9.478565,9.494975,9.330873,8.12636,6.7577443,5.280821,3.7448208,2.2022567,1.0305642,0.5907693,0.54482055,0.65969235,0.7844103,0.75487185,0.5907693,0.39384618,0.27241027,0.3708718,1.1158975,1.8116925,1.8346668,1.3981539,1.522872,1.8707694,1.723077,1.3128207,0.79097444,0.21661541,0.33805132,0.4266667,0.48902568,0.47917953,0.3052308,0.42338464,0.67610264,0.6859488,0.43651286,0.26584616,0.16410258,0.15097436,0.15425642,0.14769232,0.13456412,0.026256412,0.0,0.029538464,0.07548718,0.08533334,0.07548718,0.029538464,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.01969231,0.016410258,0.013128206,0.052512825,0.02297436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.04266667,0.13128206,0.24287182,0.34133336,0.26256412,0.23958977,0.25271797,0.26256412,0.20348719,0.18379489,0.20676924,0.26584616,0.3314872,0.32820517,0.3249231,0.27569234,0.20348719,0.13784617,0.12143591,0.16082053,0.17723078,0.17394873,0.128,0.0,0.0,0.128,0.2855385,0.4135385,0.49230772,0.37743592,0.44307697,0.48246157,0.4004103,0.20020515,0.60389745,1.024,1.3489232,1.4572309,1.1979488,1.3292309,1.8642052,1.7887181,1.0108719,0.380718,0.3314872,0.4397949,0.6235898,0.9321026,1.5327181,3.5807183,4.821334,4.516103,2.9111798,1.2537436,0.42994875,0.11158975,0.03938462,0.029538464,0.0,0.059076928,0.029538464,0.0,0.009846155,0.049230773,0.009846155,0.0,0.0,0.0,0.0,0.009846155,0.0032820515,0.0,0.0,0.0,0.009846155,0.009846155,0.02297436,0.052512825,0.06235898,0.14112821,0.21989745,0.45292312,0.81394875,1.083077,1.2603078,1.3161026,1.3620514,1.4506668,1.6082052,1.9232821,1.6935385,1.1355898,0.56451285,0.4004103,0.9189744,1.7985642,2.5961027,3.0490258,3.0949745,2.8324106,2.8422565,2.9997952,3.1376412,3.05559,2.6223593,2.3991797,2.3991797,2.6157951,3.0260515,2.917744,2.3991797,1.7165129,1.1848207,1.1749744,2.2908719,3.3476925,3.820308,3.56759,2.8324106,2.6847181,2.6322052,2.8225644,3.114667,3.058872,2.793026,3.006359,3.5249233,4.204308,4.9296412,4.699898,3.5807183,2.231795,1.3817437,1.8379488,2.6322052,3.006359,2.8127182,2.225231,1.7099489,1.8116925,2.1136413,2.7536411,3.6594875,4.5456414,5.4580517,6.0652313,6.76759,7.5979495,8.241231,7.716103,6.7544622,5.3760004,4.161641,4.273231,4.854154,4.598154,4.0402055,3.4198978,2.6880002,3.4133337,3.761231,3.5183592,3.0194874,3.1409233,3.190154,3.639795,3.9154875,4.027077,4.5554876,5.4974365,6.0258465,6.235898,6.4590774,7.273026,7.1122055,7.276308,7.3321033,7.5191803,8.730257,9.796924,9.137232,7.8112826,6.3376417,4.706462,3.564308,2.6157951,2.1530259,2.0512822,1.7591796,2.3762052,3.6036925,3.820308,2.9997952,2.7044106,5.152821,8.63836,9.974154,9.547488,11.34277,12.379898,11.756309,10.184206,8.392206,7.138462,6.954667,7.5585647,6.2162056,3.1770258,1.6771283,1.9068719,2.0512822,1.8609232,1.4703591,1.4145643,2.6584618,3.761231,4.562052,5.0674877,5.4580517,4.588308,4.322462,5.9470773,9.019077,11.372309,10.9686165,9.865847,8.618668,7.5454364,6.7314878,7.24677,8.155898,8.828718,8.969847,8.602257,8.2445135,8.004924,8.4512825,9.504821,10.456616,11.313231,11.411694,11.221334,11.365745,12.655591,13.033027,13.380924,13.952001,14.503386,14.283488,14.148924,14.720001,13.991385,11.825232,9.95118,9.728001,10.000411,10.801231,11.680821,11.69395,13.797745,15.812924,16.498873,15.730873,14.523078,12.058257,11.204924,11.204924,11.700514,12.754052,13.814155,14.536206,15.041642,15.760411,17.404718,20.240412,23.798155,27.313232,30.276926,32.42667,33.64103,34.20554,33.375183,31.077745,27.923695,24.966566,23.446976,22.629745,21.96349,21.07077,20.680206,20.496412,20.41436,20.289642,19.928617,19.003078,18.310566,17.920002,17.667284,17.161848,15.579899,14.070155,12.803283,11.792411,10.857026,9.304616,6.987488,4.7655387,3.18359,2.4582565,2.3335385,2.359795,2.4155898,2.537026,2.9243078,2.8192823,2.2055387,1.4867693,0.90584624,0.54482055,0.9517949,2.4320002,3.5314875,3.370667,1.654154,0.7844103,0.5415385,0.7515898,1.1323078,1.2603078,1.0535386,0.9911796,1.9561027,4.013949,6.413129,6.3343596,5.2020516,4.020513,3.4100516,3.6036925,3.1442053,1.8970258,1.0338463,0.8795898,0.92553854,1.0075898,0.8205129,0.47261542,0.16410258,0.17066668,0.25271797,0.33476925,0.37415388,0.3511795,0.2855385,0.20676924,0.128,0.068923086,0.029538464,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.006564103,0.0032820515,0.02297436,0.10502565,0.24287182,0.44307697,0.65969235,0.80738467,0.9124103,1.0108719,1.0404103,0.98133343,0.8598975,0.90912825,1.2635899,1.7493335,2.2088206,2.5009232,2.550154,2.7142565,3.0096412,3.4002054,3.7973337,4.0992823,4.1452312,3.9384618,3.5938463,3.3476925,3.1770258,3.0654361,3.2065644,3.6660516,4.4012313,4.8672824,4.7327185,4.7556925,4.8836927,4.9920006,4.8836927,4.6145644,4.5390773,4.4701543,4.332308,4.1517954,4.332308,4.397949,4.2830772,4.201026,4.6539493,5.3366156,5.8912826,6.1505647,6.180103,6.301539,6.633026,7.3452315,8.113232,8.651488,8.713847,7.322257,6.377026,6.629744,7.785026,8.530052,8.992821,9.787078,10.256411,10.200616,9.856001,8.5891285,8.690872,9.442462,10.148104,10.148104,9.475283,8.841846,8.592411,8.635077,8.438154,7.7292314,8.815591,9.944616,10.377847,10.390975,10.624001,10.673231,10.505847,10.295795,10.407386,10.016821,9.330873,8.809027,8.572719,8.438154,8.316719,8.467693,8.546462,8.349539,7.8112826,7.020308,6.629744,6.488616,6.3868723,6.058667,6.0816417,5.8781543,5.8223596,6.0225644,6.3179493,6.0717955,5.930667,5.720616,5.2676926,4.3651285,3.9745643,3.6660516,3.3247182,3.4166157,4.9887185,6.931693,7.6077952,8.254359,9.360411,10.666668,9.225847,8.178872,7.5552826,7.27959,7.1548724,7.1089234,7.3321033,7.7292314,7.9524107,7.4141545,6.0619493,5.474462,4.7425647,3.4625645,1.7558975,1.2800001,0.86646163,0.51856416,0.3249231,0.45620516,0.5677949,0.5940513,0.5415385,0.45620516,0.45620516,0.65312827,1.0962052,1.4375386,1.401436,0.7778462,0.9616411,1.2996924,1.7263591,2.1924105,2.6551797,3.373949,4.634257,5.1232824,4.594872,3.876103,4.6802053,6.12759,7.6898465,8.513641,7.4141545,7.0137444,6.9842057,6.997334,7.27959,8.621949,10.453334,8.090257,5.228308,3.6069746,3.0227695,3.7054362,4.1222568,4.31918,4.716308,6.117744,6.8627696,7.076103,6.820103,6.4065647,6.3934364,6.9677954,7.1483083,6.8955903,6.193231,5.0215387,3.2984617,2.0709746,1.5491283,1.4473847,1.0075898,0.6170257,0.32820517,0.49887183,1.017436,1.2964103,0.5152821,0.23958977,0.21989745,0.3446154,0.6268718,1.529436,2.1300514,1.9396925,1.3259488,1.5097437,1.8773335,1.1979488,0.54482055,0.3511795,0.4135385,0.5349744,0.56451285,0.5284103,0.47589746,0.48902568,0.48902568,0.46933338,0.4266667,0.36430773,0.28882053,0.18051283,0.13456412,0.10502565,0.06235898,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.06564103,0.101743594,0.08533334,0.06235898,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.06235898,0.19692309,0.32820517,0.47589746,0.54482055,0.3511795,0.20348719,0.11158975,0.15097436,0.28225642,0.36758977,0.39056414,0.3052308,0.190359,0.108307704,0.12143591,0.17066668,0.18379489,0.108307704,0.0,0.0,0.0,0.055794876,0.40369233,0.9682052,1.3587693,0.5513847,0.3314872,0.4135385,0.50543594,0.33476925,0.7384616,1.1881026,1.3029745,1.1520001,1.2373334,1.2471796,0.8763078,0.5415385,0.39384618,0.32164106,0.25928208,0.48246157,1.0929232,2.3729234,4.7917953,6.242462,6.3310776,4.604718,1.8904617,0.28882053,0.118153855,0.15097436,0.19364104,0.14769232,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.049230773,0.04266667,0.02297436,0.036102567,0.12143591,0.18379489,0.30851284,0.49887183,0.7778462,1.204513,1.6935385,1.9626669,2.0545642,1.9987694,1.8149745,1.3883078,0.9419488,0.571077,0.36430773,0.4135385,0.75487185,1.4080001,2.0709746,2.6420515,3.2032824,3.4592824,3.826872,4.1452312,4.263385,4.0434875,4.07959,4.023795,3.9220517,3.7973337,3.6627696,3.501949,3.0982566,2.5238976,1.8707694,1.2373334,2.2744617,3.2000003,3.8071797,3.9187696,3.4166157,2.8192823,2.3401027,2.2547693,2.484513,2.5928206,2.1530259,2.3729234,2.9111798,3.5971284,4.4406157,3.3411283,1.9396925,0.9517949,0.78769237,1.5556924,2.605949,3.2262566,3.121231,2.3926156,1.5261539,2.2350771,2.9144619,3.4560003,3.8137438,3.9975388,4.059898,4.2568207,5.661539,7.8014364,8.667898,6.921847,6.009436,5.5072823,4.969026,3.9056413,3.245949,2.9538465,2.9735386,3.2131286,3.5544617,3.6168208,3.3280003,3.1638978,3.31159,3.6758976,2.3696413,1.6968206,1.6344616,2.4681027,4.775385,7.53559,9.028924,8.218257,6.0750775,5.5991797,6.8562055,9.02236,10.082462,9.632821,8.864821,10.282667,10.341744,9.714872,8.392206,5.7074876,4.010667,3.117949,3.0030773,3.1606157,2.6256413,2.6847181,6.3901544,9.015796,8.881231,7.3550773,6.170257,4.3552823,3.5511796,4.7261543,8.195283,10.696206,12.914873,12.566976,9.603283,6.2096415,3.9286156,2.7634873,2.176,1.8018463,1.4342566,1.3128207,1.2373334,1.1323078,1.0469744,1.1454359,1.4605129,2.356513,3.259077,3.7349746,3.4789746,2.7470772,4.2305646,6.3179493,7.7325134,7.5388722,7.1844106,6.774154,6.688821,6.9382567,7.171283,7.7948723,8.736821,8.907488,8.103385,7.003898,5.6976414,5.435077,5.677949,6.012718,6.1341543,8.464411,11.995898,13.643488,12.924719,11.946668,11.936821,12.1238985,12.35036,12.672001,13.367796,13.866668,14.641232,14.936617,14.418053,13.197129,12.379898,12.452104,11.936821,10.912822,10.985026,12.658873,12.993642,12.901745,12.875488,12.983796,11.300103,10.026668,9.924924,11.21477,13.594257,15.291079,17.473642,19.843283,22.019283,23.545437,26.351591,28.947695,31.218874,32.964924,33.90359,33.575386,32.00985,29.686155,27.129438,24.933746,23.72595,23.368206,23.384617,23.476515,23.512617,22.977642,22.291695,21.615591,20.880411,19.80718,19.035898,18.7799,19.06872,19.446156,18.983387,17.076513,15.0088215,13.154463,11.638155,10.345026,8.392206,6.419693,4.588308,3.1803079,2.5928206,2.300718,2.044718,1.8379488,1.7263591,1.8018463,2.1070771,1.9167181,1.5688206,1.2504616,1.0075898,1.4342566,2.3269746,3.7448208,4.7294364,3.3247182,1.6180514,0.8336411,0.67282057,0.8205129,0.9321026,0.67282057,1.4342566,3.3312824,6.1308722,9.232411,9.097847,7.076103,4.6769233,2.678154,1.1126155,0.7122052,0.56451285,0.49230772,0.4004103,0.28882053,0.21661541,0.18051283,0.15425642,0.13456412,0.12143591,0.13456412,0.20020515,0.26912823,0.3117949,0.33476925,0.27569234,0.19692309,0.1148718,0.049230773,0.0,0.0,0.009846155,0.009846155,0.0032820515,0.016410258,0.016410258,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.04594872,0.16738462,0.39056414,0.67610264,0.955077,1.1126155,1.1027694,1.0535386,1.0043077,0.9714873,0.94523084,1.1913847,1.5721027,2.0217438,2.412308,2.546872,2.609231,2.7634873,3.0654361,3.564308,4.273231,4.663795,4.8344617,4.699898,4.3618464,4.1058464,3.9351797,3.8071797,4.0402055,4.594872,5.097026,5.4547696,4.529231,3.8334363,3.4067695,3.3903592,4.0041027,4.6834874,5.297231,5.3234878,4.9427695,5.041231,5.733744,6.619898,7.0892315,6.87918,6.0816417,5.8289237,5.901129,6.2555904,6.7085133,6.948103,7.003898,6.9120007,6.99077,7.200821,7.125334,6.114462,6.0652313,6.6100516,7.3091288,7.6635904,8.1755905,8.805744,9.373539,9.55077,8.854975,8.192,9.685334,11.099898,11.441232,10.952206,10.125129,9.370257,8.779488,8.556309,9.02236,9.206155,9.537642,10.594462,11.818667,11.539693,9.53436,8.474257,7.9885135,7.939283,8.4283085,7.7948723,7.1876926,6.7216415,6.265436,5.4482055,5.366154,6.340924,6.9021544,6.692103,6.4590774,7.138462,6.692103,5.976616,5.8223596,7.0465646,6.445949,5.543385,5.5072823,6.311385,6.7183595,6.738052,6.6822567,6.8562055,7.2927184,7.7456417,6.3573337,5.142975,4.066462,3.3575387,3.4756925,3.9417439,4.315898,4.4406157,4.453744,4.781949,4.9821544,4.97559,4.818052,4.5128207,4.020513,5.356308,5.835488,4.926359,3.3575387,3.0818465,2.9078977,2.8160002,2.4352822,1.7033848,0.86317956,0.60389745,0.40369233,0.256,0.2100513,0.3708718,0.46276927,0.5152821,0.5973334,0.73517954,0.90912825,1.0962052,1.2209232,1.273436,1.2406155,1.0962052,1.4834872,1.8970258,2.3269746,2.8225644,3.4724104,3.56759,3.3247182,3.2229745,3.4330258,3.826872,4.8672824,6.488616,8.241231,9.777231,10.84718,9.905231,9.869129,11.536411,12.941129,9.340718,5.7534366,3.948308,3.2098465,3.0654361,3.2886157,3.8564105,4.414359,4.97559,5.6320004,6.557539,7.1647186,7.387898,6.6560006,5.435077,5.2447186,5.937231,5.7074876,4.972308,3.9680004,2.737231,2.2744617,2.176,2.4615386,2.5862565,1.4342566,1.014154,1.273436,1.273436,0.827077,0.5021539,0.41682056,0.5907693,0.7417436,0.6465641,0.12471796,0.6268718,0.9682052,0.92553854,0.636718,0.5940513,0.571077,0.446359,0.3446154,0.3249231,0.38728207,0.65641034,0.6432821,0.46933338,0.29210258,0.29210258,0.3314872,0.37415388,0.4004103,0.39056414,0.3249231,0.21661541,0.09189744,0.01969231,0.029538464,0.08533334,0.016410258,0.0,0.02297436,0.049230773,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.055794876,0.28225642,0.055794876,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.01969231,0.016410258,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.03938462,0.06564103,0.26584616,0.51856416,0.4135385,0.20676924,0.16738462,0.256,0.42994875,0.6235898,0.6170257,0.48902568,0.27897438,0.0951795,0.098461546,0.08861539,0.055794876,0.08533334,0.2297436,0.512,1.0010257,1.1552821,1.2307693,1.3456411,1.4933335,0.9321026,0.54482055,0.37415388,0.3052308,0.06564103,0.14769232,1.1388719,1.7165129,1.5195899,1.1257436,0.65969235,0.33476925,0.15097436,0.07876924,0.06564103,0.052512825,0.46933338,1.5097437,3.495385,6.87918,10.246565,8.746667,5.658257,2.809436,0.5940513,0.5316923,0.44964105,0.3249231,0.16738462,0.0,0.0,0.036102567,0.036102567,0.0,0.0,0.0,0.013128206,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.009846155,0.0032820515,0.006564103,0.02297436,0.12471796,0.25271797,0.42994875,0.6892308,1.0601027,1.2931283,1.4112822,1.3653334,1.1848207,0.9747693,0.7122052,0.5218462,0.40369233,0.36102566,0.4004103,0.63343596,0.94523084,1.2832822,1.7690258,2.6912823,3.495385,4.2240005,4.2994876,3.7120004,3.0424619,2.553436,2.4516926,2.5632823,2.7766156,3.0523078,2.6289232,2.2153847,2.0512822,2.097231,2.028308,2.3236926,2.7536411,3.1409233,3.3805132,3.4166157,2.9965131,2.6256413,2.3762052,2.2514873,2.2153847,2.0676925,2.0906668,2.353231,2.6420515,2.4516926,1.332513,0.761436,0.6071795,0.827077,1.4572309,1.9331284,2.1530259,2.1070771,1.9790771,2.1497438,2.806154,3.5413337,3.7185643,3.3608208,3.1442053,3.7809234,4.2240005,4.8377438,5.622154,6.226052,4.6276927,3.3772311,3.31159,4.086154,4.1747694,4.06318,4.1189747,4.535795,5.412103,6.7282057,7.765334,7.1154876,5.651693,4.6112823,5.5926156,5.2644105,4.562052,3.69559,3.0654361,3.2623591,4.263385,7.752206,9.7903595,8.461129,3.8531284,5.356308,7.0104623,7.6307697,7.1483083,6.5837955,6.9152827,7.5618467,9.258667,11.208206,11.090053,5.7796926,3.9187696,3.754667,3.9909747,3.7973337,3.1343591,3.1803079,3.2328207,3.1967182,3.5938463,4.384821,5.395693,5.7698464,5.2676926,4.2994876,5.2315903,7.145026,9.143796,9.764103,6.9677954,4.841026,3.4297438,2.8521028,2.8750772,2.8980515,2.7963078,2.2055387,1.6278975,1.2668719,1.020718,1.4080001,2.231795,3.3805132,4.0992823,3.0030773,2.2514873,3.05559,4.6211286,6.1341543,6.76759,5.9963083,7.062975,8.667898,9.350565,7.50277,7.578257,8.12636,7.7325134,6.226052,4.709744,3.6660516,3.9680004,4.8311796,5.8518977,6.987488,7.1515903,8.897642,11.556104,13.397334,11.631591,10.729027,10.607591,10.200616,9.537642,9.7673855,11.329642,12.964104,13.955283,13.781334,12.114052,12.662155,12.875488,11.762873,10.112,10.499283,11.71036,12.393026,12.750771,12.842668,12.583385,11.2672825,10.807796,11.050668,11.920411,13.413745,16.935387,20.978874,23.860516,25.350567,26.679796,28.639181,30.628105,33.348927,36.88698,40.717133,40.15262,37.750156,33.906876,30.211285,29.449848,30.25067,31.812925,31.497849,29.295591,27.798977,27.46749,26.04308,24.431591,23.171284,22.416412,20.778667,19.544617,19.06872,19.26236,19.580719,19.081848,17.312822,15.192616,13.177437,11.247591,9.130668,7.387898,5.937231,4.7425647,3.8137438,3.1606157,2.5796926,2.034872,1.5819489,1.3718976,1.3062565,1.2898463,1.214359,1.0338463,0.7515898,0.9616411,1.270154,1.6705642,1.8543591,1.2012309,0.6268718,0.380718,0.39384618,0.5513847,0.7122052,0.9321026,1.9528207,3.6890259,6.1538467,9.452309,9.442462,8.297027,6.5083084,4.4045134,2.1398976,0.7220513,0.32164106,0.256,0.19364104,0.14441027,0.21661541,0.2986667,0.33476925,0.29538465,0.14769232,0.098461546,0.0951795,0.118153855,0.17066668,0.26256412,0.37743592,0.28225642,0.15097436,0.059076928,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.029538464,0.108307704,0.26912823,0.574359,0.9485129,1.3128207,1.5885129,1.4506668,1.3029745,1.1815386,1.1257436,1.1782565,1.401436,1.719795,2.0611284,2.3466668,2.5009232,2.6387694,3.2295387,3.945026,4.6080003,5.1889234,5.3234878,5.431795,5.5138464,5.467898,5.106872,4.7491283,4.453744,4.630975,5.2414365,5.792821,7.532308,7.463385,6.294975,4.821334,3.626667,3.0785644,3.95159,4.46359,4.522667,4.394667,4.6966157,5.3169236,6.0356927,6.567385,6.6625648,6.1013336,5.5171285,5.2578464,5.3694363,5.7468724,6.1407185,5.586052,5.1364107,5.0051284,5.159385,5.330052,5.1298466,5.3366156,5.8978467,6.626462,7.1909747,7.6701546,8.516924,9.468719,10.151385,10.089026,9.816616,10.394258,10.742155,10.538668,10.220308,9.852718,9.42277,9.02236,8.79918,8.940309,8.779488,8.963283,9.82318,10.893129,10.883283,9.527796,8.339693,8.0377445,8.51036,8.795898,7.6964107,7.2664623,7.030154,6.5378466,5.395693,5.858462,6.688821,6.7971287,6.2752824,6.4032826,7.204103,7.2960005,6.9710774,6.6560006,6.928411,6.6822567,6.2555904,6.186667,6.47877,6.619898,6.8430777,7.1187696,7.030154,6.6527185,6.567385,5.83877,5.1659493,4.772103,4.8607183,5.6320004,5.504,5.5007186,5.4941545,5.533539,5.8486156,6.157129,5.917539,5.0084105,3.5971284,2.1530259,2.7470772,2.8717952,2.2678976,1.401436,1.4506668,1.4473847,1.3522053,1.1979488,0.98133343,0.65969235,0.39384618,0.256,0.2231795,0.2855385,0.46933338,0.5415385,0.5907693,0.6465641,0.7417436,0.892718,1.0108719,1.0469744,1.1815386,1.4703591,1.8346668,2.4713848,2.9111798,3.2754874,3.6726158,4.20759,4.013949,3.626667,3.754667,4.601436,5.865026,7.351795,8.474257,9.4457445,10.384411,11.290257,11.805539,12.383181,13.46954,13.384206,8.323282,5.100308,4.7261543,5.139693,5.3760004,5.5532312,5.5926156,5.910975,6.1768208,6.1505647,5.6976414,6.1997952,6.6592827,6.5903597,5.901129,4.886975,4.2371287,4.0500517,3.5807183,2.5993848,1.3981539,1.1913847,1.2012309,1.4441026,1.847795,2.2383592,1.9790771,1.5327181,1.142154,0.92553854,0.8730257,1.1782565,1.6016412,2.0020514,2.1989746,1.9692309,1.7985642,1.4276924,0.97805136,0.574359,0.33805132,0.23958977,0.30851284,0.446359,0.56123084,0.5546667,0.5021539,0.44307697,0.39384618,0.39712822,0.5284103,0.512,0.43651286,0.38400003,0.35774362,0.28225642,0.18707694,0.098461546,0.049230773,0.03938462,0.04266667,0.009846155,0.0,0.013128206,0.02297436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.029538464,0.14112821,0.029538464,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08533334,0.20348719,0.17066668,0.23630771,0.30194873,0.38400003,0.47261542,0.5316923,0.47589746,0.37415388,0.24615386,0.13456412,0.09189744,0.03938462,0.18051283,0.4004103,0.6432821,0.92553854,1.0305642,1.0272821,1.0601027,1.148718,1.204513,0.8598975,0.40369233,0.14769232,0.101743594,0.0,0.101743594,0.9747693,1.5786668,1.4375386,0.6301539,0.30851284,0.190359,0.21661541,0.318359,0.4135385,0.48574364,0.7450257,1.467077,2.8422565,4.965744,7.3682055,6.626462,4.7524104,2.8160002,0.94523084,0.55794877,0.39384618,0.24287182,0.068923086,0.0,0.0,0.052512825,0.07548718,0.052512825,0.0,0.0,0.006564103,0.006564103,0.0032820515,0.009846155,0.009846155,0.0032820515,0.0,0.0032820515,0.009846155,0.0032820515,0.0,0.0,0.0032820515,0.01969231,0.128,0.26256412,0.40697438,0.55794877,0.72861546,0.67282057,0.64000005,0.5907693,0.52512825,0.48902568,0.42994875,0.40369233,0.39712822,0.41682056,0.4594872,0.5874872,0.761436,1.0404103,1.4933335,2.1956925,2.8291285,3.058872,2.8160002,2.28759,1.8871796,2.0250258,2.4582565,2.9768207,3.2853336,2.9801028,2.103795,1.7263591,1.8313848,2.284308,2.806154,2.8553848,2.8356924,2.7109745,2.7437952,3.508513,3.5544617,3.259077,2.9440002,2.7109745,2.4320002,1.9692309,1.8806155,1.9429746,1.8806155,1.3489232,0.6071795,0.3052308,0.33476925,0.7778462,1.910154,2.612513,2.1070771,1.4736412,1.2865642,1.5819489,2.6453335,3.314872,3.3936412,3.0358977,2.7470772,3.117949,3.43959,4.276513,5.3727183,5.661539,4.0336413,2.8849232,2.5600002,2.8488207,3.0162053,3.5511796,4.4274874,5.8453336,8.136206,11.769437,13.702565,12.747488,10.016821,7.0990777,6.045539,8.5891285,9.170052,8.772923,8.786052,11.0145645,8.579283,6.442667,6.1538467,6.62318,4.141949,4.378257,6.5444107,8.119796,8.254359,7.768616,6.7249236,6.314667,6.7971287,7.9786673,9.212719,6.941539,5.3727183,4.9362054,5.284103,5.3070774,4.273231,3.6036925,3.3411283,3.6102567,4.604718,4.6276927,4.8836927,5.097026,4.8804107,3.764513,4.3749747,7.8736415,11.096616,12.045129,9.892103,8.129642,6.9152827,6.294975,6.308103,7.0104623,6.7216415,5.668103,4.6211286,3.9351797,3.5446157,4.1550775,3.6660516,3.058872,2.6387694,2.0512822,2.1497438,3.1048207,4.6112823,5.976616,6.1013336,5.3891287,6.055385,6.8693337,6.87918,5.395693,5.4514875,5.832206,5.7435904,4.9329233,3.7054362,3.4822567,4.161641,5.0871797,6.1997952,8.054154,9.527796,10.226872,11.040821,11.477334,9.665642,9.179898,9.199591,9.012513,8.549745,8.388924,8.953437,9.465437,9.55077,9.078155,8.152616,10.059488,11.126155,11.08677,10.427077,10.384411,11.18195,11.733335,11.37559,10.440206,10.246565,10.791386,11.835078,12.924719,13.866668,14.739694,17.634462,20.804924,23.289438,24.789335,25.652515,27.75631,30.887386,35.10154,39.85395,44.01231,43.703796,40.74667,36.62113,33.250465,32.994465,33.847797,35.11795,36.102566,36.434055,36.082874,35.538055,33.913437,32.006565,30.240824,28.681849,25.655796,23.322258,21.842052,21.31036,21.769848,21.448206,19.990976,17.742771,15.094155,12.461949,9.833026,8.198565,6.99077,5.87159,4.6966157,4.1485133,3.5971284,2.8849232,2.1792822,1.9790771,1.9035898,1.7985642,1.6672822,1.4834872,1.1913847,0.7844103,0.63343596,0.64000005,0.6826667,0.5973334,0.48246157,0.39712822,0.4266667,0.65312827,1.1684103,2.2219489,3.43959,4.772103,6.2720003,8.077128,7.3419495,6.0783596,4.5587697,2.9702566,1.4539489,0.60061544,0.38728207,0.380718,0.42338464,0.6301539,1.4933335,1.6377437,1.3193847,0.7975385,0.3446154,0.15097436,0.055794876,0.032820515,0.055794876,0.108307704,0.17723078,0.14441027,0.09189744,0.055794876,0.04594872,0.029538464,0.02297436,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.036102567,0.12143591,0.32164106,0.7122052,1.1290257,1.4834872,1.7362052,1.6082052,1.5031796,1.4342566,1.4178462,1.4933335,1.6672822,1.9200002,2.1070771,2.1858463,2.2121027,2.2908719,3.0030773,3.8728209,4.601436,5.077334,5.225026,5.5762057,5.9569235,6.1538467,5.924103,5.549949,5.208616,5.290667,5.8190775,6.432821,7.7390776,8.4972315,7.755488,5.979898,3.9023592,2.5107694,2.7831798,2.9210258,3.0194874,3.18359,3.5249233,3.9253337,4.2896414,4.6145644,4.827898,4.781949,4.4767184,4.315898,4.276513,4.3618464,4.601436,4.066462,3.8400004,3.8662567,4.066462,4.3290257,4.6605134,4.9854364,5.533539,6.3212314,7.1581545,7.7390776,8.664616,9.540924,10.092308,10.174359,9.777231,9.458873,9.117539,8.786052,8.608821,8.612103,8.579283,8.530052,8.4283085,8.172308,7.4699492,7.6603084,8.3823595,9.235693,9.796924,9.350565,8.743385,8.891078,9.5606165,9.393231,8.464411,8.516924,8.776206,8.828718,8.605539,9.770667,9.708308,8.644924,7.453539,7.653744,8.021334,8.293744,8.375795,8.188719,7.6603084,7.2631803,6.8627696,6.491898,6.180103,5.940513,5.986462,6.186667,5.9470773,5.2447186,4.650667,4.5095387,4.6145644,5.037949,5.805949,6.9021544,6.3474874,5.802667,5.356308,5.0871797,5.0543594,5.1298466,4.8804107,3.9909747,2.6322052,1.4572309,1.467077,1.3226668,1.1552821,1.0568206,1.0896411,1.2537436,1.2832822,1.270154,1.2242053,1.0929232,0.7417436,0.44964105,0.32164106,0.35774362,0.47589746,0.5284103,0.5874872,0.636718,0.7089231,0.88287187,1.083077,1.2635899,1.7066668,2.4385643,3.2065644,3.9844105,4.135385,4.141949,4.263385,4.5456414,4.4964104,4.31918,4.3290257,4.8311796,6.0849237,7.5979495,8.704,9.737847,10.752001,11.546257,12.028719,12.153437,11.894155,10.505847,6.550975,5.0084105,5.2315903,5.72718,5.8814363,5.9503593,5.9470773,6.3868723,6.8693337,7.138462,7.062975,6.954667,6.941539,6.8299494,6.160411,4.201026,2.5271797,2.2219489,2.0053334,1.3784616,0.6235898,0.52512825,0.5349744,0.6432821,0.95835906,1.7066668,1.7099489,1.2603078,0.92225647,0.94523084,1.2635899,1.910154,2.3827693,2.7142565,2.7700515,2.2383592,1.9331284,1.3489232,0.82379496,0.47261542,0.19364104,0.14112821,0.28882053,0.45620516,0.53825647,0.5021539,0.39384618,0.35774362,0.37743592,0.44307697,0.54482055,0.5152821,0.42994875,0.37415388,0.3446154,0.24943592,0.1148718,0.08205129,0.07876924,0.06235898,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01969231,0.009846155,0.0,0.013128206,0.06235898,0.4004103,0.57764107,0.6301539,0.571077,0.39056414,0.26256412,0.2100513,0.18707694,0.17066668,0.16410258,0.23958977,0.49230772,0.77128214,1.0010257,1.1979488,1.0075898,0.8763078,0.8533334,0.9124103,0.9485129,0.7450257,0.35774362,0.12143591,0.10502565,0.10502565,0.16738462,0.5677949,0.88943595,0.8467693,0.28225642,0.26584616,0.34789747,0.47589746,0.5874872,0.62030774,0.571077,0.8041026,1.3128207,2.0512822,2.937436,3.7776413,3.6890259,2.989949,1.972513,0.90256417,0.44307697,0.2986667,0.20676924,0.08861539,0.055794876,0.055794876,0.08533334,0.1148718,0.10502565,0.0,0.0,0.0,0.0032820515,0.006564103,0.016410258,0.009846155,0.0032820515,0.0,0.0032820515,0.009846155,0.016410258,0.01969231,0.009846155,0.0032820515,0.01969231,0.08861539,0.18379489,0.26912823,0.3314872,0.37415388,0.22646156,0.14769232,0.128,0.15425642,0.21989745,0.27897438,0.35446155,0.4201026,0.47261542,0.5284103,0.5677949,0.6826667,0.9616411,1.4539489,2.1497438,2.665026,2.6387694,2.103795,1.3981539,1.1848207,1.7591796,2.793026,3.6660516,3.9286156,3.2918978,2.166154,1.6902566,1.7690258,2.3204105,3.2820516,3.43959,3.1934361,2.7306669,2.4943593,3.1803079,3.56759,3.501949,3.31159,3.0752823,2.5895386,2.041436,1.9200002,1.9331284,1.7690258,1.0994873,0.46933338,0.19364104,0.17394873,0.49887183,1.4211283,2.2121027,1.8313848,1.3653334,1.4112822,2.0578463,3.0096412,2.9801028,2.6683078,2.425436,2.294154,2.4024618,2.5993848,3.511795,4.8049235,5.1922054,3.826872,3.2886157,3.2295387,3.3345644,3.3017437,3.7940516,4.857436,6.626462,9.370257,13.505642,14.191591,12.773745,10.420513,8.333129,7.748924,10.692924,12.048411,11.477334,10.614155,13.039591,12.694975,7.9950776,5.0477953,5.7042055,7.5454364,5.717334,5.85518,6.6560006,7.5979495,8.966565,9.626257,8.605539,7.351795,6.820103,7.4797955,6.806975,5.7796926,5.691077,6.7314878,7.9917955,7.509334,6.5903597,6.0192823,6.1341543,6.803693,6.2884107,5.8518977,5.730462,5.658257,4.841026,5.0215387,7.8047185,10.463181,11.500309,10.633847,9.83959,10.089026,10.614155,11.0605135,11.490462,13.748514,13.413745,11.539693,9.344001,8.214975,7.5979495,5.4514875,3.3444104,2.0939488,1.7690258,2.100513,3.1015387,4.5489235,5.835488,5.989744,5.9930263,6.38359,6.678975,6.669129,6.439385,6.196513,5.802667,5.4875903,5.2447186,4.821334,5.1265645,5.5729237,6.124308,6.882462,8.103385,10.469745,11.621744,11.884309,11.424822,10.243283,9.754257,9.301334,8.707283,8.050873,7.6701546,7.3780518,7.4436927,7.936001,8.425026,7.9983597,8.0377445,7.9458466,8.36595,9.104411,9.140513,9.186462,9.554052,9.061745,7.9885135,8.070564,9.6525135,11.339488,12.724514,13.715693,14.5263605,16.659693,18.855387,20.87713,22.521437,23.591387,26.335182,30.25395,34.59939,38.623184,41.58359,41.58359,39.45354,36.644104,34.44513,33.952824,34.563286,35.843285,38.035694,40.31344,40.789337,39.45026,37.569645,35.797337,34.287594,32.699078,29.866669,27.552822,25.862566,24.894361,24.74995,23.689848,21.779694,19.055592,15.858873,12.849232,10.197334,8.940309,8.132924,7.1515903,5.7107697,5.0543594,4.585026,4.0402055,3.4560003,3.1573336,2.92759,2.5665643,2.1858463,1.8018463,1.3489232,0.7187693,0.43651286,0.3708718,0.4135385,0.48902568,0.46933338,0.46276927,0.55794877,0.92225647,1.8084104,3.43959,4.1911798,4.414359,4.450462,4.640821,3.8990772,3.0654361,2.2088206,1.4309745,0.8533334,0.74830776,0.8369231,1.014154,1.3456411,2.0676925,3.383795,3.5741541,2.8192823,1.5885129,0.6268718,0.21333335,0.049230773,0.006564103,0.006564103,0.016410258,0.032820515,0.08861539,0.13128206,0.14112821,0.12471796,0.12143591,0.10502565,0.072205134,0.029538464,0.01969231,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.02297436,0.072205134,0.17723078,0.4201026,0.8566154,1.3095386,1.6640002,1.8937438,1.8740515,1.8510771,1.8116925,1.7723079,1.7723079,1.847795,1.975795,2.0217438,1.9561027,1.8510771,1.910154,2.5895386,3.5052311,4.3651285,4.962462,5.3858466,5.9536414,6.4623594,6.7314878,6.5870776,6.3212314,5.9963083,5.927385,6.229334,6.7938466,5.3070774,6.0947695,6.294975,5.277539,3.4560003,2.2678976,1.8149745,1.7263591,1.8215386,2.0020514,2.225231,2.4943593,2.7109745,2.8389745,2.92759,3.1343591,3.4297438,3.6529233,3.6660516,3.5314875,3.501949,3.629949,3.9351797,4.309334,4.6605134,4.906667,5.3234878,5.7009234,6.170257,6.820103,7.6964107,8.297027,8.868103,9.110975,8.946873,8.507077,7.722667,7.2960005,7.1647186,7.174565,7.072821,6.9710774,7.0498466,7.1548724,7.1154876,6.7150774,5.943795,6.173539,6.8299494,7.6274877,8.530052,8.28718,8.704,9.488411,10.079181,9.642668,9.662359,10.35159,11.234463,12.2387705,13.676309,15.382976,14.139078,11.690667,9.563898,9.058462,8.868103,8.664616,8.553026,8.434873,7.9786673,6.961231,6.1046157,5.533539,5.211898,4.9362054,4.640821,4.4274874,4.279795,4.0992823,3.7054362,3.6036925,4.0500517,4.673641,5.221744,5.5926156,4.7392826,3.8071797,2.8324106,1.910154,1.1946667,1.1979488,1.3850257,1.4309745,1.3259488,1.3883078,1.5556924,1.4309745,1.3095386,1.270154,1.1454359,1.7099489,2.048,2.100513,1.9626669,1.8838975,1.4539489,0.86646163,0.4955898,0.4135385,0.40369233,0.41682056,0.508718,0.65312827,0.8795898,1.2668719,1.6344616,2.0217438,2.7011285,3.6627696,4.598154,5.35959,5.211898,4.919795,4.8311796,4.8705645,4.7655387,4.585026,4.201026,3.9122055,4.4274874,5.61559,7.3485136,9.265231,10.985026,12.117334,11.057232,9.813334,8.408616,6.7610264,4.6933336,4.194462,4.263385,4.5554876,4.8311796,4.9460516,5.159385,5.756718,6.5936418,7.6274877,8.917334,8.152616,7.240206,6.2030773,4.844308,2.740513,1.2471796,0.73517954,0.574359,0.4594872,0.40369233,0.58092314,0.79425645,0.9682052,0.9517949,0.5415385,0.6432821,0.88287187,0.86317956,0.7811283,1.4408206,2.5600002,2.6715899,2.425436,1.9561027,0.8566154,0.764718,0.4660513,0.25271797,0.190359,0.12143591,0.14769232,0.2855385,0.3446154,0.29210258,0.26256412,0.38400003,0.40697438,0.380718,0.3314872,0.256,0.26584616,0.29210258,0.318359,0.3052308,0.20676924,0.04266667,0.036102567,0.07548718,0.07876924,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.01969231,0.02297436,0.052512825,0.032820515,0.032820515,0.108307704,0.3052308,0.67282057,0.8566154,0.84348726,0.65312827,0.318359,0.12143591,0.128,0.17066668,0.2100513,0.32164106,0.69907695,0.94523084,1.1027694,1.1618463,1.0633847,0.955077,0.9616411,0.9714873,0.9714873,1.0371283,0.8960001,0.6662565,0.48574364,0.39056414,0.30194873,0.190359,0.13128206,0.118153855,0.14441027,0.21989745,0.35446155,0.508718,0.5907693,0.56123084,0.43323082,0.17394873,0.49230772,1.1027694,1.7493335,2.1792822,2.0873847,1.7887181,1.3161026,0.8041026,0.47261542,0.2986667,0.26584616,0.25271797,0.19692309,0.1148718,0.12143591,0.12143591,0.13128206,0.12471796,0.009846155,0.0032820515,0.0032820515,0.006564103,0.016410258,0.016410258,0.0032820515,0.0032820515,0.0032820515,0.0032820515,0.006564103,0.03938462,0.052512825,0.03938462,0.013128206,0.006564103,0.01969231,0.049230773,0.08205129,0.118153855,0.15425642,0.0951795,0.049230773,0.032820515,0.049230773,0.07876924,0.14441027,0.29538465,0.446359,0.5546667,0.6301539,0.6301539,0.69251287,0.88615394,1.339077,2.2350771,2.8553848,3.0260515,2.3893335,1.3292309,1.0010257,1.4933335,2.806154,3.8662567,4.1452312,3.6529233,2.6387694,2.0841026,2.038154,2.5304618,3.564308,3.9318976,3.761231,3.3608208,2.9965131,2.858667,3.2098465,3.3476925,3.2656412,2.9472823,2.3696413,2.0742567,1.9922053,2.034872,1.9331284,1.2307693,0.49887183,0.23958977,0.21661541,0.2855385,0.37415388,0.92553854,1.4572309,2.028308,2.806154,4.0500517,4.128821,3.05559,2.0709746,1.6869745,1.6902566,1.8773335,2.1497438,2.6157951,3.2262566,3.764513,3.0490258,3.190154,3.7809234,4.3684106,4.453744,4.6867695,5.622154,7.3452315,9.603283,11.812103,9.810052,7.5913854,6.6527185,7.509334,9.718155,10.253129,11.418258,10.607591,8.316719,8.162462,12.442257,10.217027,6.7577443,5.8814363,9.947898,7.3386674,5.2742567,5.0642056,7.1154876,10.94236,13.5318985,12.228924,10.121847,8.736821,8.064001,6.2555904,5.32677,5.5762057,7.0498466,9.531077,10.371283,9.252103,8.185436,8.027898,8.480822,8.569437,8.562873,8.293744,7.5388722,6.0258465,5.21518,5.3825645,6.6461544,8.195283,8.28718,8.237949,9.984001,12.11077,13.453129,13.075693,18.487797,20.027079,18.12677,14.614976,12.73436,10.459898,7.387898,4.7392826,3.121231,2.5271797,2.9636924,4.312616,5.7468724,6.8594875,7.686565,8.556309,9.097847,9.540924,10.006975,10.522257,9.593436,7.936001,6.685539,6.340924,6.7807183,7.282872,7.5618467,7.9819493,8.375795,8.04759,9.6754875,11.766154,13.144616,13.512206,13.479385,12.2847185,10.397539,8.592411,7.3780518,6.987488,6.669129,7.145026,8.644924,10.213744,9.728001,7.02359,5.61559,5.687795,6.5345645,6.5772314,6.2555904,6.885744,7.1680007,6.885744,6.928411,8.277334,9.537642,10.482873,11.21477,12.160001,13.98154,15.973744,17.893745,19.728413,21.684515,24.963284,28.55713,31.520823,33.555695,34.993233,35.11795,34.770054,34.195694,33.490055,32.597336,33.201233,35.058876,37.454773,39.427284,39.762054,37.763287,35.7678,34.29744,33.3719,32.502155,31.087593,29.781336,28.767181,27.969643,27.03754,25.212719,22.426258,19.098257,15.691488,12.704822,10.59118,9.796924,9.547488,9.074872,7.637334,6.416411,5.7764106,5.346462,4.8804107,4.240411,3.5905645,2.8947694,2.2547693,1.6836925,1.1093334,0.7975385,0.69251287,0.67938465,0.6662565,0.5677949,0.47589746,0.5152821,0.7056411,1.1913847,2.2416413,4.128821,4.33559,3.3476925,1.8970258,0.95835906,0.8795898,0.99774367,1.0765129,1.0568206,1.024,1.3292309,1.7985642,2.3335385,2.9538465,3.817026,4.568616,4.4406157,3.4198978,1.9068719,0.71548724,0.2100513,0.04266667,0.013128206,0.016410258,0.01969231,0.059076928,0.18707694,0.27569234,0.27569234,0.20676924,0.2297436,0.21661541,0.15753847,0.07548718,0.04266667,0.01969231,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.02297436,0.072205134,0.16410258,0.3117949,0.5973334,1.017436,1.4736412,1.8674873,2.1300514,2.2482052,2.294154,2.2383592,2.1070771,1.975795,1.913436,1.8642052,1.7952822,1.6869745,1.5425643,1.6640002,2.2383592,3.1540515,4.2141542,5.1298466,5.858462,6.4032826,6.774154,6.9710774,6.9809237,6.921847,6.705231,6.547693,6.62318,7.069539,2.0611284,2.231795,2.4746668,2.6518977,2.546872,1.8773335,1.9626669,2.0939488,1.9954873,1.7493335,1.785436,2.0545642,2.3236926,2.5665643,2.806154,3.0982566,3.7448208,4.06318,4.135385,4.161641,4.457026,4.9427695,5.4416413,6.0947695,6.885744,7.6307697,8.057437,8.054154,8.077128,8.379078,9.002667,8.930462,8.635077,8.241231,7.788308,7.2631803,6.6527185,6.114462,5.9995904,6.340924,6.8660517,6.11118,5.664821,5.395693,5.113436,4.578462,4.5423594,4.9821544,5.543385,5.989744,6.2096415,6.173539,7.785026,9.504821,10.473026,10.499283,11.670976,12.668719,13.892924,15.520822,17.48677,19.282053,17.266872,14.007796,10.925949,8.300308,7.506052,6.51159,5.3037953,4.1091285,3.387077,2.8521028,2.6256413,2.8980515,3.5544617,4.164923,4.1550775,3.9680004,3.6693337,3.387077,3.3280003,3.498667,3.751385,3.6824617,3.2722054,2.868513,2.4648206,2.0250258,1.5753847,1.1191796,0.65641034,0.58420515,0.62030774,0.7975385,0.99774367,0.9616411,0.9124103,0.8008206,0.79425645,0.9747693,1.3259488,2.0118976,2.3204105,2.3630772,2.3335385,2.5173335,2.028308,1.2307693,0.7187693,0.6104616,0.5481026,0.47589746,0.5940513,0.9321026,1.5097437,2.3663592,2.6453335,2.9440002,3.318154,3.8301542,4.562052,5.1987696,5.6385646,6.0356927,6.3343596,6.2851286,4.5423594,4.023795,4.2601027,4.6966157,4.6834874,5.979898,8.1066675,9.898667,10.873437,11.21477,10.545232,9.002667,7.128616,5.169231,3.0818465,3.5577438,4.6112823,6.1078978,7.4010262,7.3386674,6.692103,6.11118,5.481026,4.8147697,4.2436924,4.2305646,3.5052311,2.1792822,0.8730257,0.702359,0.60389745,0.5874872,0.6695385,0.84348726,1.0994873,1.4998976,1.8313848,2.0808206,2.1530259,1.847795,1.4309745,1.079795,0.63343596,0.5874872,2.0742567,3.9187696,2.8324106,1.5130258,1.1881026,1.6016412,0.892718,0.40697438,0.118153855,0.12143591,0.6104616,0.7450257,0.5874872,0.43323082,0.38400003,0.33476925,0.26256412,0.24287182,0.23958977,0.20676924,0.12143591,0.12143591,0.13128206,0.108307704,0.049230773,0.0,0.0,0.036102567,0.06235898,0.049230773,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.036102567,0.0951795,0.108307704,0.068923086,0.068923086,0.16738462,0.4266667,0.9156924,0.90256417,0.8008206,0.6170257,0.40369233,0.24287182,0.049230773,0.128,0.24943592,0.3446154,0.5021539,1.2242053,1.5031796,1.4867693,1.086359,0.0,0.0,0.60389745,1.1716924,1.463795,1.6475899,1.5261539,1.404718,1.214359,0.9124103,0.47261542,0.30194873,0.2231795,0.19692309,0.19692309,0.18379489,0.17066668,0.15097436,0.12471796,0.10502565,0.09189744,0.01969231,0.0,0.6235898,1.5556924,1.5556924,1.3489232,0.9321026,0.54482055,0.28882053,0.108307704,0.108307704,0.17066668,0.17066668,0.09189744,0.029538464,0.055794876,0.08861539,0.101743594,0.08205129,0.04594872,0.02297436,0.016410258,0.016410258,0.016410258,0.016410258,0.0032820515,0.009846155,0.016410258,0.01969231,0.029538464,0.055794876,0.07876924,0.08533334,0.06564103,0.029538464,0.04266667,0.072205134,0.12143591,0.18051283,0.2297436,0.16738462,0.07876924,0.02297436,0.01969231,0.029538464,0.06564103,0.3052308,0.5677949,0.764718,0.8992821,0.9485129,0.9353847,0.8533334,0.892718,1.404718,1.9167181,2.0250258,1.7329233,1.2209232,0.8533334,1.4539489,2.425436,3.5380516,4.2141542,3.5544617,2.9210258,2.7700515,3.0818465,3.6627696,4.1517954,4.4800005,4.663795,4.699898,4.5062566,3.9220517,3.7743592,3.5446157,3.0326157,2.3204105,1.7690258,1.4769232,1.4572309,1.404718,1.1815386,0.8402052,0.55794877,0.4594872,0.5940513,0.86317956,1.020718,1.585231,2.5107694,3.8367183,5.280821,6.2720003,5.1954875,3.8301542,2.5009232,1.5327181,1.2504616,1.6902566,2.2777438,2.1956925,1.4933335,1.0535386,1.1027694,1.0601027,1.1323078,1.522872,2.425436,3.9384618,6.1768208,9.199591,11.825232,11.641437,8.94359,5.4416413,4.135385,5.4580517,7.2631803,6.2752824,7.207385,9.130668,10.469745,9.019077,7.273026,5.8486156,4.1025643,2.3794873,2.0151796,3.370667,7.2336416,11.890873,16.019693,18.707693,14.362258,10.748719,8.454565,7.6110773,7.90318,7.709539,6.0750775,4.568616,4.0008206,4.4406157,6.491898,6.885744,6.994052,7.785026,9.810052,10.505847,10.535385,9.813334,8.323282,6.088206,4.1714873,4.818052,6.4065647,7.213949,5.431795,3.8104618,3.8071797,5.2709746,7.1581545,7.522462,9.475283,12.885334,14.434463,13.676309,13.016617,12.2847185,10.28595,7.197539,4.2830772,3.9056413,6.8233852,10.538668,12.570257,12.754052,13.22995,13.961847,13.676309,12.980514,12.291283,11.841642,10.423796,8.103385,6.235898,5.5597954,6.196513,7.3419495,9.314463,11.067078,11.795693,10.939077,11.661129,12.425847,13.154463,14.004514,15.396104,13.955283,10.052924,7.384616,6.87918,6.6822567,6.304821,5.733744,4.5062566,3.0752823,2.809436,4.417641,7.9425645,8.759795,6.2588725,3.8301542,5.3431797,7.269744,8.136206,7.6110773,6.5017443,7.7325134,8.664616,9.091283,9.179898,9.462154,10.279386,11.930258,14.116103,16.594053,19.18031,22.209642,24.923899,27.103182,28.645746,29.571285,29.607388,30.037336,30.880823,31.59631,31.081028,31.327183,32.377438,33.860924,35.331284,36.26995,35.367386,34.36308,33.014156,31.425644,30.06031,28.46195,27.648003,27.342772,27.136002,26.489437,25.317745,22.672413,19.557745,16.551386,13.778052,12.045129,11.024411,11.241027,12.032001,11.58236,9.531077,8.139488,6.820103,5.4514875,4.3651285,3.2525132,2.2514873,1.591795,1.3062565,1.2209232,1.270154,1.3915899,1.4769232,1.4473847,1.2504616,0.9944616,0.86646163,0.9353847,1.3161026,2.1825643,4.4767184,5.8190775,5.2020516,3.0326157,1.1290257,0.6892308,0.7089231,0.9944616,1.3423591,1.5261539,2.2580514,3.4297438,4.5095387,4.965744,4.2568207,3.0851285,1.5392822,0.56123084,0.3117949,0.15425642,0.07876924,0.02297436,0.006564103,0.01969231,0.029538464,0.14112821,0.26912823,0.3249231,0.29210258,0.24287182,0.256,0.23958977,0.18707694,0.10502565,0.029538464,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02297436,0.07548718,0.17394873,0.3249231,0.51856416,0.82379496,1.148718,1.5130258,1.8970258,2.228513,2.4352822,2.5238976,2.487795,2.3401027,2.1202054,1.9626669,1.7591796,1.5556924,1.4080001,1.3587693,1.529436,1.9462565,2.7963078,3.9811285,5.142975,5.7042055,5.8978467,5.924103,6.091488,6.8365135,7.066257,7.1909747,7.256616,7.4141545,7.890052,2.2416413,2.3860514,2.3072822,2.048,1.7394873,1.595077,1.8379488,2.1267693,2.3204105,2.425436,2.5796926,3.0818465,3.6135387,4.132103,4.785231,5.930667,7.4174366,8.3593855,8.605539,8.274052,7.77518,7.4732313,6.944821,6.2785645,5.83877,6.2490263,6.3245134,5.904411,5.540103,5.464616,5.609026,5.8486156,6.1407185,6.4065647,6.419693,5.799385,5.293949,4.9460516,4.7294364,4.59159,4.460308,4.1550775,3.9680004,3.9909747,4.2568207,4.7228723,4.6867695,4.673641,4.6178465,4.5554876,4.598154,4.601436,4.5587697,5.0838976,6.2555904,7.6176414,7.9885135,8.448001,9.042052,9.639385,9.944616,10.400822,10.174359,9.048616,7.4371285,6.38359,6.5280004,5.6943593,4.5390773,3.5938463,3.2525132,2.9111798,2.6683078,2.678154,2.793026,2.553436,1.975795,1.4802053,1.4441026,2.03159,3.1934361,2.8455386,2.6387694,2.5042052,2.3630772,2.1366155,1.8904617,1.6869745,1.654154,1.7723079,1.8642052,2.0939488,2.281026,2.3401027,2.1333334,1.4605129,1.3456411,1.4408206,1.4736412,1.4080001,1.4506668,1.723077,1.6443079,1.5458462,1.6278975,1.9692309,1.3522053,0.7844103,0.571077,0.72861546,1.0010257,1.2800001,1.4998976,2.0644104,3.0654361,4.2830772,3.8990772,4.588308,6.0816417,7.525744,7.466667,7.427283,7.4010262,7.318975,6.961231,5.943795,3.4756925,3.442872,4.397949,5.35959,5.805949,6.5247183,7.269744,7.522462,7.2664623,6.99077,6.62318,6.432821,6.262154,6.058667,5.865026,7.824411,9.462154,10.748719,11.195078,9.865847,8.027898,6.114462,4.210872,2.540308,1.4605129,2.8521028,3.3050258,3.0687182,2.3105643,1.1060513,0.6859488,0.6170257,0.8598975,1.1881026,1.2209232,1.2832822,1.270154,1.2898463,1.3620514,1.4178462,0.8763078,0.52512825,0.5218462,0.9911796,2.0020514,2.809436,1.9692309,1.0436924,0.67610264,0.60061544,0.39056414,0.3511795,0.46276927,0.6235898,0.63343596,0.63343596,0.6301539,0.54482055,0.39384618,0.2855385,0.28225642,0.28225642,0.26584616,0.21333335,0.108307704,0.072205134,0.03938462,0.02297436,0.009846155,0.0,0.0,0.006564103,0.013128206,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.029538464,0.049230773,0.03938462,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.032820515,0.07876924,0.049230773,0.009846155,0.0,0.006564103,0.01969231,0.02297436,0.013128206,0.013128206,0.052512825,0.13784617,0.24287182,0.23302566,0.18051283,0.41025645,0.84348726,0.9878975,0.45292312,0.3446154,0.5152821,0.8533334,1.2832822,1.467077,1.4900514,1.4506668,1.3161026,0.90256417,0.6104616,0.61374366,0.7811283,1.0601027,1.4769232,1.6377437,1.6443079,1.4703591,1.1126155,0.5940513,0.25928208,0.16738462,0.17066668,0.18707694,0.19692309,0.17394873,0.15097436,0.0951795,0.06564103,0.20020515,0.49887183,0.88287187,1.083077,1.0272821,0.81066674,0.6235898,0.39384618,0.21333335,0.12471796,0.118153855,0.08861539,0.06564103,0.04266667,0.01969231,0.006564103,0.009846155,0.026256412,0.032820515,0.029538464,0.02297436,0.006564103,0.009846155,0.009846155,0.0032820515,0.0032820515,0.0,0.009846155,0.009846155,0.0032820515,0.006564103,0.01969231,0.04266667,0.059076928,0.06564103,0.07876924,0.14112821,0.20348719,0.23302566,0.22646156,0.21661541,0.19364104,0.15097436,0.108307704,0.068923086,0.04266667,0.029538464,0.13128206,0.3314872,0.61374366,0.9747693,1.2570257,1.3817437,1.4867693,1.6640002,1.9528207,1.8609232,1.8182565,1.7755898,1.5983591,1.086359,1.1684103,1.5261539,1.9790771,2.3368206,2.4188719,2.665026,3.2984617,3.8137438,3.9089234,3.4789746,3.5347695,3.6430771,3.8695388,4.056616,3.8104618,3.4198978,3.2984617,3.0884104,2.6551797,2.0873847,1.7362052,1.4605129,1.2209232,1.024,0.9353847,0.73517954,0.4660513,0.5021539,0.84348726,1.1191796,1.4080001,2.0906668,2.9571285,3.754667,4.197744,4.089436,3.7842054,3.0490258,2.1792822,1.9954873,2.4155898,2.5206156,2.353231,2.0086155,1.6278975,1.5491283,1.6935385,2.3236926,3.370667,4.4406157,6.0028725,7.9294367,10.066052,11.651283,11.300103,6.7085133,4.4012313,4.338872,6.2096415,9.42277,9.508103,7.8637953,6.7577443,6.7150774,6.491898,4.8640003,3.9581542,3.564308,3.5314875,3.761231,4.4406157,5.661539,6.2752824,6.3606157,7.2205133,7.200821,6.8594875,7.282872,8.65477,10.246565,7.0531287,5.654975,6.3179493,7.6603084,6.626462,6.340924,5.3398976,6.8496413,11.053949,15.07118,13.764924,11.585642,9.288206,7.4371285,6.4065647,7.3682055,8.832001,10.072617,10.200616,8.152616,4.644103,3.4625645,3.9548721,5.5269747,7.634052,10.502565,13.197129,13.784616,12.481642,11.634872,12.662155,14.355694,13.735386,10.706052,8.093539,9.5835905,10.988309,11.720206,11.277129,9.212719,8.851693,9.9282055,10.604308,10.496001,10.66995,10.873437,8.664616,6.2851286,5.182359,6.012718,7.1483083,8.182155,8.5661545,7.9983597,6.413129,6.3310776,8.03118,10.020103,11.69395,13.35795,12.931283,10.571488,7.578257,5.464616,5.9634876,5.8781543,5.034667,4.3716927,4.2371287,4.4077954,5.0018463,5.7764106,5.87159,5.159385,4.2338467,4.778667,5.425231,5.7140517,5.61559,5.5105643,6.196513,7.584821,8.720411,9.107693,8.717129,9.435898,10.571488,11.828514,13.430155,16.105026,19.026052,21.507284,23.512617,25.051899,26.2039,26.738874,27.349335,27.953234,28.425848,28.616207,29.669746,31.17949,32.541542,33.493336,34.110363,34.20226,33.870773,33.05026,31.727592,29.94872,28.048412,26.53867,25.501541,24.854977,24.352823,23.93272,22.646156,20.818052,18.592821,15.937642,13.161027,11.303386,10.509129,10.476309,10.433641,9.330873,7.788308,6.23918,4.890257,3.7054362,2.8291285,2.2744617,2.162872,2.4418464,2.8914874,2.7470772,2.3794873,2.1792822,2.28759,2.6289232,3.1638978,3.8367183,4.2207184,3.9942567,2.937436,3.367385,3.748103,3.6036925,2.937436,2.2022567,2.028308,2.2350771,2.7076926,3.3017437,3.8465643,3.9909747,4.3716927,4.6802053,4.417641,2.878359,2.487795,2.5042052,2.2055387,1.4375386,0.60389745,0.15097436,0.013128206,0.006564103,0.016410258,0.01969231,0.098461546,0.16082053,0.16082053,0.128,0.15753847,0.20020515,0.2231795,0.20020515,0.13784617,0.055794876,0.029538464,0.016410258,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.032820515,0.12471796,0.26584616,0.45620516,0.702359,0.9485129,1.1913847,1.4703591,1.782154,2.0939488,2.3696413,2.5632823,2.6486156,2.6256413,2.5238976,2.3171284,2.0841026,1.8379488,1.6475899,1.6377437,1.8970258,2.4549747,3.318154,4.3060517,5.044513,4.854154,4.4964104,4.240411,4.391385,5.2742567,6.363898,7.515898,8.602257,9.386667,9.511385,4.5587697,5.674667,6.124308,6.042257,5.4547696,4.273231,3.2787695,2.3696413,2.097231,2.4713848,2.9702566,3.7874875,4.31918,4.7491283,5.3103595,6.2720003,7.968821,9.38995,9.856001,9.4457445,8.989539,8.664616,8.001641,7.1220517,6.2490263,5.720616,5.3792825,4.97559,4.778667,4.8377438,4.972308,5.2676926,5.6976414,6.0652313,6.189949,5.917539,5.47118,5.1364107,4.8607183,4.604718,4.3651285,4.2207184,4.161641,4.450462,5.106872,5.8781543,6.3179493,5.609026,4.568616,3.82359,3.8301542,3.5282054,2.9669745,2.674872,2.937436,3.7842054,4.2994876,4.778667,5.2348723,5.602462,5.7403083,6.2720003,6.6100516,6.311385,5.5893335,5.3202057,5.543385,5.349744,5.10359,5.041231,5.2512827,5.297231,4.8311796,4.076308,3.1934361,2.28759,1.6213335,1.2635899,1.1323078,1.2340513,1.6672822,1.4178462,1.3522053,1.3620514,1.332513,1.1191796,1.4834872,2.1103592,3.1606157,4.312616,4.7491283,4.650667,4.263385,3.620103,2.7109745,1.4867693,1.1749744,1.0633847,1.0010257,1.0108719,1.2603078,1.4375386,1.142154,0.8533334,0.7975385,0.9419488,0.83035904,0.72861546,0.77128214,1.1355898,2.048,2.3335385,2.166154,2.7798977,4.332308,5.8945646,6.560821,8.723693,10.965334,11.733335,9.337437,9.18318,9.199591,8.267488,6.692103,6.226052,5.9995904,5.32677,4.7360005,4.3716927,4.010667,4.9296412,5.6385646,5.970052,5.8092313,5.10359,4.342154,3.748103,3.9056413,4.896821,6.304821,8.914052,10.06277,10.194052,9.810052,9.472001,7.351795,4.1747694,2.3236926,2.1891284,2.172718,2.9669745,3.367385,3.2918978,2.5632823,0.88615394,1.5425643,2.4549747,2.6584618,2.1103592,1.6804104,1.4441026,1.529436,1.5031796,1.1651284,0.5349744,0.3249231,0.56451285,1.3883078,2.0250258,0.79425645,1.014154,1.2570257,1.1749744,0.7450257,0.2855385,0.3708718,0.4660513,0.5973334,0.71548724,0.6859488,0.6071795,0.512,0.43651286,0.39384618,0.37415388,0.41682056,0.37743592,0.3052308,0.22646156,0.15097436,0.14112821,0.12471796,0.072205134,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.02297436,0.01969231,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.04266667,0.06235898,0.03938462,0.02297436,0.049230773,0.02297436,0.0,0.0,0.0,0.029538464,0.04266667,0.055794876,0.07548718,0.10502565,0.12143591,0.049230773,0.14441027,0.380718,0.46933338,0.21989745,0.15753847,0.3511795,0.6892308,0.8763078,0.955077,1.1093334,1.1585642,1.0338463,0.7811283,0.3708718,0.24615386,0.37743592,0.69579494,1.1060513,1.2406155,1.2077949,0.90584624,0.4660513,0.24943592,0.12143591,0.11158975,0.12471796,0.13456412,0.15097436,0.13456412,0.101743594,0.06235898,0.08861539,0.3117949,0.61374366,0.69907695,0.5973334,0.40369233,0.29538465,0.25928208,0.20020515,0.14112821,0.108307704,0.13128206,0.118153855,0.055794876,0.009846155,0.0,0.0,0.0,0.0032820515,0.006564103,0.006564103,0.016410258,0.009846155,0.013128206,0.009846155,0.0,0.0,0.0,0.013128206,0.02297436,0.01969231,0.01969231,0.016410258,0.016410258,0.029538464,0.04594872,0.06564103,0.101743594,0.13784617,0.15425642,0.15097436,0.14112821,0.15753847,0.15097436,0.118153855,0.07548718,0.04594872,0.029538464,0.068923086,0.25928208,0.60389745,1.0108719,1.3653334,1.585231,1.7460514,1.8773335,1.9364104,1.5721027,1.1848207,1.0075898,1.0043077,0.84348726,0.9189744,1.0732309,1.2471796,1.401436,1.5327181,1.9462565,2.4976413,2.9046156,2.9833848,2.6617439,2.5304618,2.5140514,2.7766156,3.2722054,3.7185643,3.2984617,3.05559,2.8389745,2.540308,2.1202054,1.7985642,1.4998976,1.1651284,0.82379496,0.5874872,0.5415385,0.39712822,0.37415388,0.5546667,0.8960001,1.3226668,1.9462565,2.4057438,2.6026669,2.7175386,2.8356924,3.045744,2.9833848,2.6289232,2.300718,2.5042052,2.5107694,2.3302567,2.0217438,1.7066668,1.5589745,1.6705642,2.28759,3.4100516,4.8049235,8.408616,10.092308,9.7903595,8.43159,7.9097443,5.6352825,4.604718,4.571898,5.3169236,6.6395903,6.373744,5.3366156,4.598154,4.352,3.9089234,2.8521028,2.1956925,2.0709746,2.353231,2.6683078,3.1081028,3.8662567,4.312616,4.4898467,5.1265645,5.398975,5.8518977,7.532308,9.83959,10.541949,8.04759,6.4032826,6.6034875,8.149334,9.028924,6.9842057,5.5696416,6.2588725,8.605539,10.236719,9.878975,9.833026,9.222565,8.119796,7.5552826,8.815591,8.914052,8.421744,8.018052,8.503796,6.6067696,5.0838976,4.9788723,6.2227697,7.640616,8.999385,11.1983595,12.363488,11.897437,10.496001,13.98154,17.076513,16.708925,13.955283,14.04718,16.626873,17.178257,15.862155,12.839386,8.274052,8.267488,8.881231,9.130668,8.996103,9.416205,9.357129,7.5421543,5.786257,5.074052,5.5630774,6.954667,7.3058467,6.941539,6.308103,5.9667697,5.8847184,6.5936418,7.90318,9.42277,10.5780525,10.59118,9.012513,7.2992826,6.8299494,8.914052,9.114257,8.592411,7.8703594,7.4469748,7.8080006,8.260923,7.8802056,7.8080006,8.411898,9.268514,8.152616,6.738052,4.95918,3.570872,4.1189747,5.146257,6.803693,8.316719,9.26195,9.573745,9.882257,10.663385,11.621744,12.711386,14.162052,15.819489,17.381744,19.078566,20.962463,22.889027,24.805746,25.659079,26.056208,26.318771,26.479591,27.897438,29.48595,30.84472,31.721027,31.993439,32.000004,31.8359,31.284515,30.28349,28.914873,27.815386,26.791388,25.911797,25.370258,25.48513,26.548515,28.15672,27.966362,25.432617,21.83549,16.876308,13.794462,11.976206,10.909539,10.194052,9.363693,8.303591,6.9087186,5.3694363,4.1517954,3.3805132,3.6463592,4.276513,4.8705645,5.280821,3.9942567,2.678154,1.8084104,1.5425643,1.7132308,2.0841026,2.4549747,2.733949,2.7995899,2.4681027,2.8717952,3.3378465,3.7185643,4.073026,4.6867695,4.7622566,4.338872,4.056616,4.1485133,4.414359,4.781949,4.266667,3.3312824,2.300718,1.3620514,2.294154,3.7152824,3.7349746,2.2580514,1.0010257,0.21661541,0.013128206,0.006564103,0.006564103,0.006564103,0.06564103,0.101743594,0.09189744,0.06564103,0.101743594,0.15753847,0.20676924,0.2231795,0.20020515,0.14441027,0.07548718,0.032820515,0.009846155,0.0032820515,0.009846155,0.009846155,0.0032820515,0.0,0.0032820515,0.01969231,0.08533334,0.2100513,0.3708718,0.56451285,0.7844103,1.0305642,1.2898463,1.5786668,1.8871796,2.169436,2.4188719,2.5993848,2.7076926,2.740513,2.6978464,2.5961027,2.4484105,2.2350771,2.0086155,1.8838975,1.9528207,2.3138463,2.8914874,3.5478978,4.086154,3.7874875,3.5314875,3.4297438,3.6758976,4.516103,5.786257,7.3485136,8.677744,9.4457445,9.53436,5.2381544,6.6461544,7.50277,8.060719,8.237949,7.604513,6.1407185,4.9329233,4.493129,4.7392826,4.9887185,5.5138464,5.7501545,5.7140517,5.664821,6.11118,7.9228725,8.641642,8.369231,7.8441033,8.4283085,8.684308,8.530052,8.113232,7.5618467,6.9677954,6.7872825,6.6428723,6.5903597,6.6133337,6.6067696,6.554257,6.6002054,6.626462,6.5378466,6.242462,5.648411,5.21518,4.841026,4.4800005,4.1452312,3.9286156,3.7874875,3.9581542,4.4045134,4.827898,5.2676926,4.7228723,3.8006158,3.0358977,2.9013336,2.477949,1.9528207,1.4309745,1.1684103,1.5556924,2.3630772,3.1442053,3.6758976,3.9581542,4.1911798,4.7524104,5.041231,4.9526157,4.630975,4.4832826,4.7458467,5.1232824,5.5138464,5.8125134,5.8814363,5.6320004,5.0609236,4.1780515,3.1245131,2.1530259,1.7362052,1.6246156,1.5392822,1.3784616,1.2340513,1.2471796,1.4998976,1.6475899,1.5360001,1.1815386,1.5753847,2.2219489,3.2262566,4.332308,4.9329233,4.972308,4.6900516,4.0402055,3.0654361,1.8838975,1.1684103,0.7844103,0.6235898,0.64000005,0.8402052,0.955077,0.75487185,0.64000005,0.7122052,0.7844103,0.88287187,1.0043077,1.1749744,1.5655385,2.5107694,3.2656412,3.5478978,4.332308,5.979898,8.228104,10.230155,11.644719,12.895181,13.61395,12.632616,10.505847,9.15036,7.650462,6.12759,5.756718,6.4623594,6.0816417,5.4449234,4.9099493,4.3651285,4.1058464,4.1780515,4.4012313,4.460308,3.9056413,3.1638978,2.3696413,2.7273848,4.4800005,6.87918,10.029949,10.7158985,9.941334,8.661334,7.781744,6.1046157,3.6463592,2.6912823,3.5314875,4.466872,5.2315903,5.3398976,5.074052,4.466872,3.2886157,3.058872,3.0884104,2.6518977,1.8904617,1.8281027,1.9823592,2.2055387,2.0053334,1.2209232,0.009846155,0.40697438,0.97805136,1.7952822,2.103795,0.318359,0.16082053,0.6498462,0.9189744,0.7056411,0.38400003,0.5152821,0.5513847,0.5546667,0.58420515,0.6859488,0.5874872,0.39384618,0.34133336,0.43651286,0.49230772,0.49230772,0.39712822,0.27569234,0.17394873,0.108307704,0.118153855,0.118153855,0.08205129,0.029538464,0.02297436,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.032820515,0.036102567,0.026256412,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.04266667,0.04266667,0.0,0.0,0.04266667,0.02297436,0.0,0.0,0.0,0.029538464,0.04266667,0.04594872,0.052512825,0.072205134,0.1148718,0.049230773,0.0,0.0,0.0,0.0,0.14769232,0.34133336,0.47261542,0.42338464,0.46276927,0.761436,0.9156924,0.76800007,0.41025645,0.08205129,0.0,0.11158975,0.3446154,0.60389745,0.6662565,0.56451285,0.29210258,0.0,0.0,0.02297436,0.049230773,0.068923086,0.07876924,0.07876924,0.07548718,0.059076928,0.052512825,0.101743594,0.24943592,0.37743592,0.27569234,0.13128206,0.04594872,0.04594872,0.08205129,0.098461546,0.101743594,0.108307704,0.118153855,0.0951795,0.049230773,0.01969231,0.013128206,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.013128206,0.016410258,0.013128206,0.0032820515,0.0,0.0032820515,0.01969231,0.029538464,0.026256412,0.029538464,0.01969231,0.009846155,0.013128206,0.026256412,0.03938462,0.052512825,0.059076928,0.06235898,0.06564103,0.07876924,0.1148718,0.128,0.1148718,0.08861539,0.08205129,0.08533334,0.128,0.28882053,0.55794877,0.8402052,1.0601027,1.1979488,1.3292309,1.4539489,1.4966155,1.2996924,0.86646163,0.574359,0.53825647,0.5874872,0.764718,0.90584624,0.98133343,0.99774367,0.9944616,1.2176411,1.5031796,1.7723079,1.9626669,2.03159,1.975795,2.0217438,2.294154,2.7667694,3.249231,2.9702566,2.7602053,2.5337439,2.2580514,1.9561027,1.7132308,1.591795,1.4703591,1.1946667,0.5874872,0.40369233,0.27897438,0.2297436,0.34789747,0.79425645,1.5491283,1.9265642,1.9035898,1.6607181,1.5819489,1.8084104,2.1956925,2.3827693,2.284308,2.0676925,2.300718,2.2613335,2.0512822,1.7887181,1.6147693,1.4769232,1.5688206,2.034872,3.045744,4.8114877,8.592411,9.724719,8.553026,6.482052,5.9634876,5.4514875,5.280821,5.4843082,6.048821,6.928411,6.439385,5.398975,4.594872,4.1189747,3.3608208,2.8882053,2.7142565,2.934154,3.436308,3.9253337,3.8104618,3.6660516,3.7185643,3.9975388,4.2962055,4.2568207,4.854154,6.925129,9.96759,12.150155,11.234463,9.540924,8.096821,7.6996927,8.907488,7.53559,6.7872825,6.2194877,5.4974365,4.381539,4.7983594,6.189949,7.269744,7.387898,6.5378466,6.7577443,6.196513,5.720616,6.23918,8.700719,8.274052,7.197539,6.8627696,7.4010262,7.6668725,7.125334,7.578257,8.231385,8.582564,8.43159,13.367796,16.659693,16.75159,14.943181,15.382976,17.631182,18.034874,16.370872,12.993642,8.828718,8.556309,9.6754875,10.522257,10.364718,9.419488,8.342975,6.770872,5.474462,4.8049235,4.6900516,5.6287184,5.901129,5.7731285,5.6352825,6.0160003,6.3606157,6.380308,6.7216415,7.6176414,8.868103,8.713847,7.059693,6.038975,6.62318,8.621949,9.426052,9.987283,10.079181,9.862565,9.865847,9.718155,8.776206,8.234667,8.539898,9.403078,8.034462,6.452513,4.6112823,3.2262566,3.761231,4.854154,6.3540516,8.024616,9.567181,10.630565,11.083488,11.707078,12.435693,13.157744,13.692719,13.889642,14.339283,15.458463,17.306257,19.600412,21.888002,23.105642,23.722668,24.050873,24.241232,25.636105,26.935797,27.9959,28.586668,28.432413,28.117336,27.871181,27.536413,27.083488,26.62072,26.532104,26.25313,25.862566,25.603285,25.888823,27.050669,29.128208,29.787899,28.114054,24.595694,19.131079,15.881847,14.020925,12.973949,12.412719,10.84718,9.206155,7.397744,5.6451287,4.4898467,3.7940516,3.9778464,4.3027697,4.397949,4.266667,3.0129232,1.8970258,1.1716924,0.92225647,1.0699488,1.2340513,1.1355898,1.1323078,1.3620514,1.7624617,2.162872,2.6880002,3.4330258,4.7556925,7.276308,7.768616,6.564103,5.077334,4.0500517,3.5380516,3.6102567,2.7831798,1.6705642,0.79425645,0.5874872,1.5786668,2.8258464,2.934154,1.8609232,0.9156924,0.20348719,0.02297436,0.013128206,0.0,0.0,0.052512825,0.07876924,0.06564103,0.03938462,0.059076928,0.10502565,0.15097436,0.18707694,0.20348719,0.18707694,0.09189744,0.036102567,0.009846155,0.0032820515,0.009846155,0.009846155,0.0032820515,0.006564103,0.029538464,0.072205134,0.17394873,0.32820517,0.50543594,0.6826667,0.8467693,1.083077,1.3718976,1.6968206,2.0184617,2.2744617,2.4549747,2.5829747,2.681436,2.7634873,2.8258464,2.8980515,2.9013336,2.789744,2.5796926,2.353231,2.2153847,2.3171284,2.5731285,2.917744,3.2853336,3.1245131,3.0326157,3.0326157,3.239385,3.889231,4.8738465,6.114462,7.174565,7.837539,8.113232,4.6834874,5.5105643,6.340924,7.5191803,8.969847,10.203898,9.642668,9.524513,9.662359,9.819899,9.682052,8.891078,8.136206,7.1122055,6.2588725,6.75118,8.618668,7.8145647,6.186667,5.346462,6.675693,7.5191803,8.14277,8.612103,8.982975,9.288206,9.796924,10.148104,10.164514,9.892103,9.596719,9.202872,8.5891285,7.9228725,7.2336416,6.413129,5.612308,5.0838976,4.6112823,4.082872,3.511795,3.0260515,2.740513,2.609231,2.553436,2.4681027,2.5600002,2.865231,2.9472823,2.7011285,2.3302567,2.048,1.8379488,1.6705642,1.6902566,2.2055387,2.9046156,3.767795,4.31918,4.4800005,4.6080003,4.788513,4.8607183,4.772103,4.532513,4.194462,4.279795,4.588308,4.841026,4.8049235,4.2863593,3.387077,2.8882053,2.5895386,2.3401027,2.048,2.2449234,2.4549747,2.6847181,2.9210258,3.1245131,3.3772311,3.7940516,3.9154875,3.6135387,3.0916924,2.8816411,2.5764105,2.2908719,2.2219489,2.6584618,3.1442053,3.498667,3.4724104,3.0260515,2.3433847,1.2635899,0.80738467,0.67282057,0.65969235,0.6301539,0.7975385,1.0108719,1.401436,1.8215386,1.8116925,1.585231,1.7132308,2.1989746,2.993231,3.9975388,5.287385,6.2096415,6.675693,7.4896417,10.31877,12.859077,12.153437,11.634872,12.836103,15.392821,10.929232,7.837539,6.38359,5.937231,4.965744,4.634257,5.2676926,5.989744,6.3606157,6.36718,4.57518,3.4330258,2.878359,2.7864618,2.9505644,2.868513,2.7011285,3.3772311,5.1331286,7.496206,10.650257,10.965334,9.95118,8.3593855,6.196513,5.668103,5.5007186,5.504,5.786257,6.7544622,8.165744,8.165744,7.7325134,7.328821,6.925129,4.6145644,2.5862565,1.2340513,0.83035904,1.5458462,2.349949,2.5829747,2.1858463,1.2800001,0.17394873,1.0502565,1.4276924,1.401436,1.1093334,0.7450257,0.43323082,0.28882053,0.32820517,0.47917953,0.5940513,0.5677949,0.48902568,0.40697438,0.40369233,0.6104616,0.5415385,0.3708718,0.34789747,0.47917953,0.5218462,0.4397949,0.3249231,0.20676924,0.10502565,0.01969231,0.013128206,0.006564103,0.026256412,0.059076928,0.049230773,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02297436,0.06564103,0.08861539,0.068923086,0.026256412,0.0,0.0,0.0,0.013128206,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03938462,0.01969231,0.0,0.0,0.0,0.0,0.32820517,0.49230772,0.39056414,0.3117949,0.26584616,0.51856416,0.702359,0.6104616,0.17723078,0.049230773,0.013128206,0.029538464,0.07548718,0.15097436,0.18707694,0.07876924,0.0,0.0032820515,0.0,0.0,0.0,0.01969231,0.04266667,0.013128206,0.036102567,0.03938462,0.052512825,0.072205134,0.06235898,0.02297436,0.036102567,0.036102567,0.013128206,0.016410258,0.006564103,0.0032820515,0.029538464,0.068923086,0.072205134,0.032820515,0.032820515,0.03938462,0.032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.013128206,0.013128206,0.016410258,0.016410258,0.02297436,0.026256412,0.02297436,0.016410258,0.026256412,0.016410258,0.013128206,0.013128206,0.016410258,0.026256412,0.04266667,0.049230773,0.052512825,0.059076928,0.09189744,0.108307704,0.13456412,0.14769232,0.14769232,0.15097436,0.15425642,0.20348719,0.28882053,0.39384618,0.48246157,0.4955898,0.49887183,0.5907693,0.7811283,0.9747693,1.1093334,0.9288206,0.6859488,0.5349744,0.5349744,0.7220513,0.8795898,0.92225647,0.8566154,0.78769237,0.7811283,0.95835906,1.2176411,1.5097437,1.8445129,2.0053334,2.1825643,2.3762052,2.5107694,2.428718,2.4549747,2.5206156,2.4320002,2.1398976,1.7362052,1.5130258,1.5327181,1.6968206,1.6705642,0.8992821,0.44964105,0.21333335,0.17723078,0.37415388,0.8992821,1.7952822,1.8215386,1.4506668,1.0469744,0.8960001,1.2012309,1.4933335,1.5097437,1.3489232,1.4769232,1.9889232,1.9889232,1.8215386,1.6935385,1.6869745,1.6311796,1.6705642,1.9232821,2.6847181,4.417641,6.5017443,7.1122055,6.921847,6.51159,6.3606157,5.989744,6.262154,6.8988724,7.958975,9.810052,10.115283,8.208411,6.2227697,5.0477953,4.3290257,4.20759,4.667077,5.3792825,6.117744,6.76759,6.242462,4.8049235,3.4855387,2.733949,2.3926156,2.9735386,3.8071797,5.4908724,8.438154,12.885334,12.727796,11.592206,9.412924,7.197539,7.062975,7.8145647,7.7981544,6.3179493,3.879385,2.1825643,2.3072822,2.8717952,3.9712822,4.7655387,3.501949,2.865231,2.9833848,3.9745643,5.76,8.050873,7.9786673,8.050873,8.090257,7.9885135,7.712821,6.173539,4.4340515,3.5314875,4.132103,6.5312824,11.178667,14.017642,15.031796,14.36554,12.320822,12.445539,12.803283,12.544001,11.503591,10.220308,8.749949,10.673231,12.626052,12.688411,10.397539,8.910769,7.256616,5.691077,4.466872,3.817026,3.7120004,4.2174363,4.8804107,5.3792825,5.5302567,6.2851286,6.426257,6.2490263,6.449231,8.1066675,8.057437,6.3376417,4.9821544,4.7294364,5.0018463,6.2227697,7.7456417,8.999385,9.55077,9.120821,8.3364105,7.0531287,5.799385,4.97559,4.850872,4.709744,4.844308,4.9099493,4.821334,4.7425647,5.2020516,6.160411,7.7948723,9.770667,11.241027,12.235488,12.826258,13.4170265,14.112822,14.6871805,14.076719,13.640206,13.945437,15.130258,16.922258,18.021746,19.209848,20.279797,21.14954,21.85518,23.030155,23.945848,24.497232,24.582565,24.109951,23.70954,23.417439,23.361643,23.545437,23.857233,24.175592,24.30031,24.346258,24.38236,24.44472,24.388926,24.4119,24.726976,24.65149,22.613335,19.177027,17.106052,16.036104,15.658668,15.734155,13.197129,10.272821,7.6570263,5.7468724,4.630975,4.013949,3.3017437,2.4943593,1.6672822,0.9747693,0.9321026,1.079795,1.3029745,1.5064616,1.6180514,1.6311796,1.2832822,1.0338463,1.0732309,1.3193847,1.2471796,1.4539489,2.176,3.9187696,7.463385,8.408616,7.138462,5.100308,3.249231,2.048,1.394872,0.8795898,0.5874872,0.5218462,0.5940513,0.6892308,0.84348726,1.0732309,1.211077,0.8992821,0.30851284,0.0951795,0.032820515,0.006564103,0.0032820515,0.068923086,0.12143591,0.14769232,0.14112821,0.0951795,0.07548718,0.128,0.19692309,0.25271797,0.27569234,0.14769232,0.06235898,0.016410258,0.0032820515,0.0,0.0032820515,0.0032820515,0.02297436,0.068923086,0.15097436,0.2855385,0.47917953,0.67938465,0.8566154,0.9682052,1.1585642,1.4276924,1.7493335,2.0676925,2.300718,2.4385643,2.537026,2.6322052,2.7602053,2.9407182,3.1573336,3.2984617,3.31159,3.190154,2.9636924,2.7569232,2.665026,2.6912823,2.8258464,3.0293336,3.0949745,3.1113849,3.0884104,3.114667,3.3575387,3.754667,4.2469745,4.8804107,5.58277,6.173539,7.4929237,8.152616,8.874667,9.833026,10.889847,11.595488,12.3536415,13.449847,14.736411,16.02954,17.106052,13.820719,10.584617,7.817847,6.629744,8.789334,10.217027,8.805744,6.892308,5.540103,4.562052,4.9788723,6.1538467,7.824411,9.485129,10.374565,11.352616,12.612924,13.082257,12.73436,12.586668,12.819694,11.871181,10.197334,8.375795,7.0957956,6.4590774,6.0258465,5.612308,5.074052,4.31918,3.4034874,3.2656412,3.436308,3.639795,3.8006158,4.397949,4.821334,4.8771286,4.578462,4.1517954,3.9056413,4.312616,4.8672824,5.330052,5.720616,5.5991797,5.61559,5.8420515,6.170257,6.3179493,6.439385,6.377026,6.2129235,5.986462,5.7074876,4.240411,3.242667,2.7011285,2.4648206,2.2580514,1.8674873,1.4211283,1.4145643,1.9987694,2.9768207,4.3552823,5.2020516,5.796103,6.409847,7.325539,7.860513,8.041026,7.890052,7.499488,7.0334363,6.521436,5.35959,4.1025643,3.1573336,2.793026,2.6322052,2.4385643,2.231795,1.9396925,1.404718,0.5973334,0.40697438,0.57764107,0.9485129,1.4506668,2.231795,3.0194874,3.7907696,4.1452312,3.3247182,2.678154,3.1113849,4.827898,7.6242056,10.893129,11.1983595,10.305642,8.444718,7.145026,9.232411,10.758565,11.579078,11.792411,11.585642,11.23118,9.472001,8.300308,7.499488,6.8463597,6.088206,5.7107697,5.5958977,5.110154,4.3027697,3.9384618,4.460308,3.5216413,2.3696413,1.9626669,2.9768207,3.5380516,4.1517954,4.4898467,4.713026,5.4941545,6.518154,5.5762057,4.630975,4.706462,5.8912826,7.3550773,8.306872,8.251078,7.6209235,7.765334,8.132924,8.077128,7.6635904,6.8988724,5.7534366,5.093744,4.086154,2.6157951,1.2504616,1.2504616,1.4703591,1.654154,1.5458462,1.1749744,0.86974365,1.4933335,1.4572309,0.9485129,0.4135385,0.5481026,0.5481026,0.48574364,0.5021539,0.5940513,0.5940513,0.31507695,0.25271797,0.27897438,0.34133336,0.48902568,0.48902568,0.44307697,0.40697438,0.38728207,0.3511795,0.28882053,0.26584616,0.23958977,0.190359,0.09189744,0.06564103,0.032820515,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016410258,0.07548718,0.07548718,0.029538464,0.0,0.0,0.0,0.06235898,0.029538464,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02297436,0.049230773,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.18379489,0.26912823,0.20020515,0.15097436,0.128,0.15097436,0.19692309,0.21333335,0.09189744,0.09189744,0.072205134,0.049230773,0.026256412,0.016410258,0.0032820515,0.0,0.006564103,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.072205134,0.036102567,0.006564103,0.013128206,0.0,0.013128206,0.016410258,0.032820515,0.06564103,0.07548718,0.026256412,0.02297436,0.029538464,0.02297436,0.0,0.036102567,0.06564103,0.059076928,0.02297436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.03938462,0.07548718,0.06564103,0.032820515,0.009846155,0.0032820515,0.016410258,0.016410258,0.006564103,0.0,0.0032820515,0.016410258,0.03938462,0.06564103,0.12471796,0.20020515,0.21333335,0.15097436,0.20020515,0.26912823,0.28225642,0.19692309,0.12471796,0.08861539,0.08205129,0.10502565,0.15097436,0.21333335,0.37415388,0.5513847,0.7187693,0.8992821,0.88943595,0.77456415,0.63343596,0.55794877,0.65641034,0.764718,0.8763078,0.9124103,0.8598975,0.761436,0.78769237,1.020718,1.4080001,1.8543591,2.2580514,2.3926156,2.297436,2.0709746,1.8313848,1.7099489,2.2219489,2.6157951,2.7864618,2.553436,1.6640002,1.2373334,0.88287187,0.7187693,0.7056411,0.65641034,0.508718,0.4004103,0.40697438,0.58420515,0.9616411,1.2307693,1.3522053,1.2898463,1.142154,1.1290257,1.0436924,0.892718,0.8041026,0.83035904,0.97805136,1.5753847,2.1267693,2.3335385,2.2482052,2.2744617,2.3335385,1.9561027,1.6640002,1.7460514,2.2580514,4.6145644,5.7632823,5.865026,5.651693,6.409847,7.200821,7.968821,7.8145647,6.882462,6.3310776,8.628513,8.303591,6.485334,4.460308,3.692308,3.6332312,4.201026,4.5554876,4.4996924,4.4865646,5.330052,4.962462,3.8695388,2.8192823,2.868513,4.650667,5.4613338,5.5532312,5.2545643,4.97559,4.1813335,4.378257,5.0904617,6.183385,7.8441033,8.342975,6.994052,4.71959,2.9997952,3.889231,4.023795,3.4002054,2.733949,2.2711797,1.7690258,2.2449234,2.7602053,2.9111798,2.789744,2.9604106,3.767795,5.6352825,7.1220517,7.686565,7.6767187,6.5772314,5.277539,4.4964104,5.10359,8.116513,10.998155,12.770463,13.252924,12.675283,11.674257,11.08677,11.07036,11.592206,12.343796,12.711386,10.587898,9.462154,9.179898,9.567181,10.420513,10.752001,8.772923,6.373744,4.6605134,3.95159,3.4264617,3.5347695,4.332308,5.4449234,6.042257,6.6527185,6.521436,6.1013336,5.8486156,6.226052,8.3364105,8.408616,7.003898,5.2447186,4.8049235,4.903385,5.3398976,5.549949,5.5204105,5.8125134,6.521436,5.362872,4.1550775,4.059898,5.586052,6.196513,7.2270775,7.6110773,7.0990777,6.2555904,5.671385,6.045539,7.4075904,9.4457445,11.52,12.251899,12.78359,13.896206,15.530668,16.800821,16.774565,16.009848,15.497848,15.602873,16.068924,15.212309,14.880821,15.862155,17.900309,19.669334,20.768822,21.691078,22.150566,22.130873,21.910976,21.717335,21.730463,22.06195,22.501745,22.537848,21.940514,21.83549,22.06195,22.465643,22.918566,22.59036,21.819078,20.880411,20.036924,19.561028,19.561028,19.186872,18.422155,17.296412,15.868719,14.01436,11.516719,9.015796,6.961231,5.6320004,5.044513,4.082872,3.0227695,2.1464617,1.7558975,1.9856411,2.6945643,3.495385,3.754667,2.5928206,1.8248206,1.276718,1.0305642,1.0502565,1.1585642,0.9517949,0.8533334,0.892718,1.1060513,1.5556924,2.5074873,2.9472823,2.7470772,2.0611284,1.3259488,0.98461545,0.79097444,0.65641034,0.571077,0.5940513,1.2537436,2.1136413,2.878359,3.1573336,2.487795,0.98461545,0.3249231,0.0951795,0.026256412,0.016410258,0.101743594,0.29538465,0.5284103,0.6301539,0.3511795,0.15425642,0.318359,0.52512825,0.64000005,0.702359,0.41025645,0.17066668,0.04266667,0.013128206,0.0,0.013128206,0.016410258,0.032820515,0.08861539,0.19692309,0.39384618,0.6432821,0.8992821,1.1126155,1.2373334,1.3587693,1.5163078,1.7296412,1.9823592,2.228513,2.4352822,2.5698464,2.678154,2.7963078,2.930872,3.1245131,3.2853336,3.3805132,3.3903592,3.2820516,3.170462,2.9801028,2.8488207,2.8717952,3.0654361,3.5446157,3.945026,4.1485133,4.0402055,3.5413337,3.1376412,3.2098465,3.6857438,4.46359,5.4153852,5.674667,7.7390776,9.714872,11.497026,13.02318,14.27036,14.539488,14.9398985,16.052513,17.266872,16.787693,13.88636,12.068104,10.748719,9.803488,9.570462,8.743385,7.4436927,6.232616,5.5762057,5.8190775,6.957949,8.064001,9.110975,9.974154,10.423796,10.94236,11.766154,12.632616,13.075693,12.442257,11.559385,10.686359,9.6754875,8.595693,7.6931286,7.499488,7.204103,6.7610264,6.2030773,5.661539,5.2644105,5.175795,5.290667,5.5302567,5.8256416,6.6002054,7.2960005,7.8047185,7.955693,7.5191803,7.4010262,7.574975,7.827693,8.080411,8.3823595,8.818872,8.621949,8.109949,7.512616,6.9776416,7.177847,7.4929237,7.3058467,6.488616,5.425231,4.0500517,2.9636924,2.1366155,1.5031796,0.96492314,0.827077,0.8763078,1.2438976,1.9561027,2.9636924,4.4012313,5.835488,6.7544622,6.9842057,6.688821,6.0750775,5.4908724,5.0609236,4.7228723,4.240411,3.5807183,2.425436,1.5425643,1.2373334,1.339077,1.142154,1.0338463,1.020718,1.2537436,2.0250258,2.4713848,2.993231,3.2000003,3.058872,2.9144619,3.0326157,4.4110775,6.5280004,8.740103,10.282667,11.2672825,12.064821,12.475078,12.4685135,12.176412,10.499283,9.931488,9.869129,10.128411,10.916103,11.825232,13.065847,12.99036,11.707078,11.0605135,10.962052,9.40636,7.578257,6.2162056,5.6352825,4.8377438,4.0434875,3.6857438,3.6332312,3.1671798,2.861949,2.989949,2.9604106,2.5435898,1.8773335,2.156308,2.553436,3.2656412,4.532513,6.6527185,8.694155,8.904206,8.507077,7.9425645,6.892308,7.3583593,7.9163084,8.579283,8.815591,7.5454364,7.8637953,10.55836,12.018872,11.073642,8.999385,5.605744,3.748103,3.0030773,2.3696413,0.24943592,0.29538465,1.1585642,1.6771283,1.5425643,1.2832822,1.017436,0.7811283,0.5874872,0.5677949,0.97805136,1.014154,0.955077,0.9682052,1.0272821,0.8992821,0.45292312,0.2855385,0.2297436,0.20348719,0.18379489,0.2231795,0.26584616,0.27897438,0.26256412,0.26584616,0.27241027,0.23630771,0.18379489,0.1148718,0.01969231,0.02297436,0.026256412,0.016410258,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016410258,0.08861539,0.13784617,0.14112821,0.12471796,0.101743594,0.072205134,0.026256412,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03938462,0.055794876,0.036102567,0.0,0.0,0.0,0.0951795,0.17066668,0.17066668,0.10502565,0.098461546,0.0951795,0.0951795,0.11158975,0.16410258,0.08533334,0.032820515,0.009846155,0.006564103,0.0032820515,0.0,0.0,0.0,0.0032820515,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.016410258,0.006564103,0.0,0.0032820515,0.0,0.013128206,0.029538464,0.072205134,0.118153855,0.101743594,0.02297436,0.04266667,0.049230773,0.029538464,0.072205134,0.16738462,0.101743594,0.026256412,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.026256412,0.026256412,0.013128206,0.0032820515,0.0,0.0032820515,0.0032820515,0.0,0.0032820515,0.009846155,0.0032820515,0.016410258,0.03938462,0.07548718,0.12143591,0.15097436,0.11158975,0.12143591,0.18379489,0.24287182,0.18707694,0.08205129,0.055794876,0.059076928,0.072205134,0.09189744,0.1148718,0.19364104,0.29538465,0.38728207,0.42338464,0.42338464,0.40697438,0.43323082,0.5152821,0.6301539,0.7220513,0.79097444,0.80738467,0.76800007,0.6892308,0.8008206,1.1158975,1.4769232,1.7690258,1.9167181,1.9922053,1.9987694,1.9265642,1.7263591,1.3292309,1.4441026,1.6410258,1.9298463,2.1136413,1.7985642,1.2242053,0.9124103,0.7778462,0.7089231,0.58420515,0.43651286,0.39384618,0.50543594,0.81066674,1.3161026,1.9167181,2.1136413,1.9659488,1.5819489,1.1290257,0.94523084,0.764718,0.5940513,0.5481026,0.83035904,1.5163078,2.6256413,3.2820516,3.2131286,2.7503593,2.5271797,2.3630772,2.162872,2.0808206,2.5140514,3.7185643,4.585026,5.3431797,6.1768208,7.2270775,8.12636,7.90318,6.7774363,5.7731285,6.698667,7.8703594,7.3485136,6.3868723,5.6320004,5.106872,4.850872,4.906667,4.844308,4.5423594,4.1682053,4.9526157,5.2447186,4.381539,3.006359,3.0752823,4.525949,4.384821,3.9023592,4.092718,5.7074876,5.3825645,5.211898,5.5138464,6.157129,6.547693,5.8092313,4.8082056,3.9253337,3.3214362,2.9636924,2.806154,2.4713848,2.4615386,2.681436,2.4648206,2.1891284,2.1267693,2.1136413,2.100513,2.1530259,2.7733335,3.6726158,4.138667,4.073026,4.013949,3.7251284,3.515077,4.096,5.668103,7.9228725,9.5146675,10.167795,9.941334,9.4457445,9.842873,10.427077,10.315488,10.463181,10.850462,10.463181,9.268514,9.078155,9.393231,10.095591,11.447796,9.403078,6.5903597,4.7458467,4.128821,3.5478978,2.9669745,3.006359,3.7021542,4.9952826,6.7249236,6.701949,6.2490263,5.989744,6.2063594,6.8496413,8.178872,9.130668,9.216001,8.234667,6.2720003,5.5302567,5.1856413,5.172513,5.346462,5.47118,5.349744,5.2578464,4.886975,4.315898,3.9844105,4.4012313,4.775385,4.97559,4.955898,4.778667,4.5456414,4.6112823,5.113436,6.055385,7.322257,8.306872,9.42277,11.10318,13.525334,16.580925,17.8839,17.808413,16.689232,15.218873,14.431181,14.592001,14.7790785,15.350155,16.41354,17.801847,18.244925,18.441847,18.379488,18.192411,18.189129,18.550156,19.121233,19.734976,20.178053,20.194464,19.662771,19.334566,19.259079,19.446156,19.879387,20.30277,20.378258,20.489847,20.804924,21.293951,21.001848,20.115694,18.970259,17.723078,16.331488,14.634667,12.527591,10.240001,8.057437,6.3277955,5.5072823,4.588308,3.5511796,2.5665643,1.9987694,2.4155898,3.7349746,4.9526157,5.4514875,4.9854364,3.3772311,3.0129232,3.5347695,4.3060517,4.4077954,4.5029745,4.4077954,4.092718,3.6693337,3.387077,3.6660516,4.2502565,4.6178465,4.4964104,3.889231,2.9636924,1.9462565,1.3653334,1.339077,1.6082052,2.28759,3.05559,3.748103,4.1452312,4.0008206,2.7831798,1.585231,0.6695385,0.15097436,0.0032820515,0.049230773,0.21989745,0.37415388,0.4135385,0.27897438,0.4135385,0.6301539,0.78769237,0.83035904,0.761436,0.49887183,0.23958977,0.072205134,0.013128206,0.013128206,0.013128206,0.02297436,0.04594872,0.101743594,0.2100513,0.41682056,0.67610264,0.9321026,1.142154,1.273436,1.394872,1.522872,1.6836925,1.8871796,2.1431797,2.3794873,2.556718,2.6880002,2.7864618,2.8914874,3.058872,3.2853336,3.5282054,3.7316926,3.817026,3.7087183,3.4855387,3.2295387,3.062154,3.1409233,3.626667,4.2207184,4.6867695,4.854154,4.6276927,4.2240005,4.092718,4.3716927,5.0642056,6.0258465,3.2951798,4.5554876,5.9470773,7.312411,8.5891285,9.793642,10.614155,10.985026,11.464206,11.959796,11.71036,11.201642,11.464206,11.611898,11.254155,10.499283,8.79918,7.571693,6.633026,5.976616,5.7501545,6.547693,7.4043083,8.146052,8.743385,9.275078,9.964309,10.985026,12.015591,12.672001,12.524308,11.730052,10.932513,10.085744,9.202872,8.346257,7.837539,8.054154,8.303591,8.241231,7.8637953,8.123077,8.470975,8.851693,9.104411,8.950154,8.891078,9.074872,9.344001,9.521232,9.432616,9.15036,8.973129,8.805744,8.641642,8.572719,8.576,7.9786673,7.0334363,5.986462,5.07077,5.723898,6.3310776,6.6067696,6.2785645,5.110154,4.0992823,3.4921029,3.0162053,2.5862565,2.3171284,3.0424619,3.629949,4.164923,4.713026,5.330052,6.3967185,7.6668725,8.904206,9.737847,9.642668,7.6635904,5.5630774,3.6168208,2.1924105,1.7558975,1.7394873,1.785436,1.8281027,1.913436,2.176,2.409026,2.6880002,3.0490258,3.5840003,4.4340515,4.33559,4.096,4.023795,4.1682053,4.325744,4.5456414,6.1440005,8.402052,10.761847,12.839386,14.5952835,15.91795,16.452925,15.927796,14.135796,11.1294365,11.23118,12.599796,14.247386,16.052513,15.415796,14.578873,12.750771,10.35159,8.992821,8.372514,7.0334363,5.717334,4.850872,4.535795,4.604718,4.1025643,3.1474874,2.3466668,2.7733335,3.0293336,2.5895386,2.166154,2.0151796,1.9396925,3.1737437,3.4789746,3.0654361,2.9571285,5.0018463,6.51159,6.987488,7.1187696,7.131898,6.803693,7.9228725,8.920616,9.90195,10.213744,8.444718,8.310155,10.121847,10.81436,9.596719,7.936001,6.2096415,4.900103,4.017231,3.2361028,1.9035898,1.404718,1.2077949,0.96492314,0.65312827,0.5546667,1.0272821,1.0338463,0.9288206,0.9747693,1.3489232,1.148718,0.81066674,0.69579494,0.7811283,0.67282057,0.318359,0.2100513,0.21661541,0.256,0.2986667,0.29538465,0.2855385,0.24615386,0.190359,0.15097436,0.118153855,0.09189744,0.06564103,0.03938462,0.0,0.0032820515,0.009846155,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.032820515,0.16410258,0.128,0.049230773,0.0,0.0,0.0,0.0,0.08861539,0.16738462,0.18379489,0.108307704,0.06564103,0.02297436,0.0,0.006564103,0.036102567,0.11158975,0.09189744,0.06235898,0.052512825,0.036102567,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01969231,0.04266667,0.036102567,0.026256412,0.029538464,0.01969231,0.0,0.0,0.006564103,0.03938462,0.068923086,0.08205129,0.08205129,0.08205129,0.07876924,0.059076928,0.04266667,0.08205129,0.036102567,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.04594872,0.08861539,0.098461546,0.06235898,0.01969231,0.02297436,0.01969231,0.013128206,0.036102567,0.08205129,0.04266667,0.006564103,0.0,0.0,0.006564103,0.0032820515,0.0032820515,0.009846155,0.009846155,0.0032820515,0.0,0.0,0.0,0.006564103,0.006564103,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0,0.013128206,0.02297436,0.03938462,0.101743594,0.29210258,0.3511795,0.33805132,0.2855385,0.21333335,0.118153855,0.11158975,0.1148718,0.118153855,0.118153855,0.12143591,0.14112821,0.18379489,0.23958977,0.29210258,0.3052308,0.29210258,0.318359,0.39712822,0.51856416,0.6629744,0.7122052,0.7253334,0.73517954,0.7515898,0.7811283,0.90912825,1.3292309,1.7755898,2.038154,1.9692309,1.7887181,1.6114873,1.5721027,1.6082052,1.4736412,1.4802053,1.7132308,1.9987694,2.1431797,1.9593848,1.4080001,1.0075898,0.7844103,0.7089231,0.69251287,0.7089231,0.6498462,0.80738467,1.3029745,2.0808206,1.9003079,1.5983591,1.2406155,0.88943595,0.6071795,0.5021539,0.43323082,0.39056414,0.42994875,0.67282057,1.6246156,2.4943593,2.861949,2.6453335,2.0808206,2.1825643,3.0916924,3.3772311,2.8291285,2.422154,3.5938463,4.850872,5.976616,6.633026,6.3507695,6.738052,7.0892315,6.695385,5.8289237,5.737026,5.3234878,4.6080003,4.082872,4.0008206,4.3716927,4.8672824,5.549949,5.7632823,5.297231,4.4012313,3.2229745,2.789744,2.3663592,2.041436,2.7536411,3.9647183,4.3585644,4.138667,3.8400004,4.325744,3.8301542,4.420923,5.346462,5.933949,5.5663595,4.069744,2.8816411,2.8849232,3.6430771,3.3805132,2.6223593,2.789744,3.6496413,4.9132314,6.23918,5.730462,5.0182567,4.2141542,3.5905645,3.564308,3.948308,3.9089234,3.4592824,2.793026,2.2646155,2.8324106,3.8728209,5.789539,8.018052,9.025641,8.92718,7.8145647,7.0531287,7.3747697,8.881231,10.492719,10.827488,10.384411,9.452309,8.109949,7.3419495,7.6964107,8.149334,8.388924,8.818872,7.765334,6.2096415,4.886975,4.092718,3.7054362,3.2525132,3.121231,3.6726158,4.8311796,6.0816417,5.5532312,5.037949,4.850872,5.280821,6.5837955,7.9819493,9.4457445,10.44677,10.44677,8.881231,6.2523084,5.152821,4.9493337,4.9887185,4.6276927,4.1222568,4.027077,4.1025643,4.1517954,4.017231,4.132103,4.276513,4.4307694,4.594872,4.7589746,4.46359,4.315898,4.919795,6.1440005,7.1056414,7.466667,7.939283,8.772923,10.112,12.002462,13.200411,13.5548725,13.042872,12.212514,12.182976,12.95754,13.551591,14.027489,14.450873,14.916924,14.634667,14.506668,14.631386,15.081027,15.911386,16.918976,17.975796,18.638771,18.753643,18.44513,17.874052,17.70995,17.992207,18.569847,19.091694,19.534771,19.846565,20.22072,20.630976,20.850874,19.692308,18.231796,16.715488,15.510976,15.113848,14.112822,12.425847,10.453334,8.513641,6.8562055,5.8978467,5.0642056,4.2469745,3.4166157,2.6354873,2.5140514,2.9833848,3.5347695,3.8367183,3.7349746,2.9111798,2.8717952,3.373949,4.06318,4.466872,4.893539,5.1954875,5.4613338,5.786257,6.2523084,7.0137444,6.3343596,5.21518,4.269949,3.7251284,2.8291285,1.8806155,1.2504616,1.0666667,1.2209232,1.6640002,2.0906668,2.3893335,2.4582565,2.2186668,1.5556924,0.8763078,0.38400003,0.13784617,0.06564103,0.07876924,0.17723078,0.25271797,0.25928208,0.21333335,0.31507695,0.39384618,0.41682056,0.380718,0.32164106,0.21661541,0.118153855,0.04594872,0.016410258,0.016410258,0.02297436,0.04594872,0.07876924,0.14441027,0.26912823,0.46276927,0.71548724,0.955077,1.142154,1.2635899,1.3423591,1.4539489,1.6049232,1.8149745,2.0939488,2.3433847,2.556718,2.7011285,2.7864618,2.8914874,3.0884104,3.4002054,3.7776413,4.1583595,4.44718,4.460308,4.31918,3.9844105,3.56759,3.3247182,3.446154,3.9318976,4.519385,5.0182567,5.32677,5.4908724,5.720616,6.088206,6.5444107,6.921847,3.1442053,3.1442053,3.5249233,4.1714873,4.95918,5.7468724,6.6002054,6.8529234,6.8299494,6.803693,6.997334,8.264206,9.760821,10.919386,11.401847,11.10318,9.924924,9.035488,7.9524107,6.6625648,5.6320004,6.377026,6.9382567,7.256616,7.4174366,7.6570263,8.51036,9.93477,11.260718,12.182976,12.750771,12.747488,12.297847,11.654565,11.008,10.482873,9.7903595,9.803488,9.938052,9.882257,9.567181,9.888822,10.774975,11.720206,12.186257,11.618463,10.952206,10.492719,9.787078,8.904206,8.421744,8.0377445,7.7423596,7.4699492,7.204103,6.9382567,6.665847,6.1374364,5.398975,4.57518,3.8498464,4.384821,4.962462,5.5105643,5.786257,5.366154,4.6276927,4.3290257,4.532513,5.113436,5.7764106,7.0498466,6.918565,6.3212314,5.7501545,5.2709746,6.173539,7.3091288,8.621949,9.593436,9.216001,6.7774363,4.5489235,2.7175386,1.6640002,1.9495386,2.8488207,3.8498464,4.4898467,4.588308,4.2568207,4.0041027,4.1025643,4.7524104,5.9602056,7.522462,6.669129,5.7764106,5.35959,5.6976414,6.813539,7.8769236,9.347282,10.893129,12.3536415,13.74195,15.330462,17.05354,18.596104,19.429745,18.835693,16.49559,15.307488,14.903796,15.028514,15.540514,13.925745,12.071385,9.980719,8.214975,7.890052,7.6964107,7.3682055,6.564103,5.435077,4.6145644,5.402257,5.044513,3.6496413,2.3138463,3.114667,3.3542566,2.2153847,1.4408206,1.6180514,2.172718,3.4592824,3.5511796,2.6584618,1.9035898,3.31159,4.089436,4.493129,5.169231,6.229334,7.240206,8.812308,9.708308,10.345026,10.742155,10.525539,10.47959,10.820924,9.885539,7.6701546,5.8420515,5.100308,4.1485133,3.1474874,2.3401027,2.0709746,1.6443079,1.1027694,0.5874872,0.24287182,0.23302566,0.9485129,1.0305642,0.9156924,0.88287187,1.0633847,0.8960001,0.6301539,0.5973334,0.764718,0.7056411,0.4397949,0.58420515,0.7515898,0.7253334,0.45620516,0.27569234,0.19692309,0.14769232,0.098461546,0.055794876,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.02297436,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.026256412,0.06235898,0.098461546,0.128,0.13784617,0.10502565,0.049230773,0.032820515,0.16410258,0.128,0.06235898,0.098461546,0.24943592,0.39056414,0.512,0.53825647,0.47261542,0.34133336,0.21333335,0.12471796,0.04266667,0.0,0.0,0.0,0.07548718,0.03938462,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.02297436,0.0032820515,0.0,0.029538464,0.07548718,0.072205134,0.03938462,0.03938462,0.036102567,0.026256412,0.029538464,0.03938462,0.03938462,0.026256412,0.016410258,0.04594872,0.04594872,0.04594872,0.029538464,0.009846155,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.006564103,0.006564103,0.03938462,0.06235898,0.059076928,0.029538464,0.01969231,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.0032820515,0.0032820515,0.009846155,0.009846155,0.0032820515,0.0,0.0,0.0,0.006564103,0.006564103,0.0032820515,0.0,0.0,0.0,0.0032820515,0.006564103,0.006564103,0.0032820515,0.0,0.032820515,0.059076928,0.06564103,0.098461546,0.26912823,0.34789747,0.34789747,0.29538465,0.2297436,0.20348719,0.2986667,0.37743592,0.39712822,0.380718,0.39056414,0.45292312,0.49887183,0.512,0.48574364,0.40369233,0.34789747,0.3511795,0.42994875,0.56123084,0.67282057,0.6826667,0.6695385,0.65969235,0.67938465,0.7318975,0.8598975,1.2898463,1.9003079,2.3663592,2.1530259,1.595077,1.3062565,1.3226668,1.5491283,1.7657437,2.0939488,2.4910772,2.6387694,2.4451284,2.044718,1.4473847,1.0469744,0.8598975,0.8730257,1.0338463,1.2832822,1.4605129,1.8510771,2.349949,2.4648206,1.463795,0.85005134,0.49230772,0.31507695,0.29538465,0.3511795,0.40369233,0.4397949,0.60061544,1.1552821,2.2580514,2.8849232,2.9078977,2.4188719,1.7591796,2.8127182,4.2141542,4.637539,4.020513,3.5511796,4.4110775,5.149539,5.5729237,5.4908724,4.709744,5.208616,6.121026,6.5345645,6.0324106,4.706462,3.6594875,3.4330258,3.4855387,3.629949,4.020513,3.882667,4.706462,5.58277,5.6418467,4.0336413,2.038154,1.2800001,1.2406155,1.657436,2.5435898,3.4133337,4.1189747,4.2338467,3.7021542,2.8291285,2.3171284,3.259077,4.082872,4.076308,3.387077,2.2514873,1.4145643,1.6869745,2.7503593,3.1442053,3.3345644,4.6605134,5.796103,6.5444107,7.824411,7.755488,6.73477,5.5762057,5.1167183,6.2194877,6.0160003,4.893539,3.6004105,2.612513,2.1234872,3.0654361,4.6802053,6.8397956,8.805744,9.229129,7.8769236,5.835488,4.8016415,5.356308,6.944821,8.763078,8.953437,8.14277,6.9776416,6.1078978,6.0783596,6.6527185,6.9743595,6.8299494,6.688821,6.820103,6.925129,6.688821,6.229334,6.0849237,4.827898,3.9581542,4.082872,4.8607183,4.9887185,4.027077,3.5807183,3.6496413,4.3651285,5.979898,7.2664623,8.707283,10.036513,10.656821,9.655796,6.8660517,5.6352825,5.2644105,5.074052,4.417641,3.8564105,3.5478978,3.5314875,3.7743592,4.161641,4.309334,4.397949,4.4865646,4.630975,4.8672824,4.7392826,4.6572313,5.2381544,6.38359,7.269744,7.4075904,7.5881033,8.024616,8.769642,9.718155,10.404103,10.909539,11.162257,11.300103,11.680821,12.1238985,12.304411,12.389745,12.455385,12.488206,12.458668,12.875488,13.751796,14.989129,16.393847,17.46708,18.277744,18.46154,18.034874,17.375181,16.823795,16.8599,17.394873,18.14318,18.6519,18.763489,18.822565,19.157335,19.587284,19.423182,17.667284,15.931078,14.309745,13.164309,13.092104,12.544001,11.378873,9.885539,8.392206,7.2369237,6.672411,5.930667,5.1954875,4.568616,4.076308,3.623385,3.3509746,3.3050258,3.3575387,3.2098465,2.7864618,2.868513,3.3017437,4.013949,5.0116925,4.841026,4.4832826,4.3749747,4.706462,5.4186673,6.3934364,5.609026,4.2994876,3.2164104,2.6289232,2.0118976,1.4703591,1.1552821,1.0404103,0.9156924,0.8402052,0.90584624,0.92553854,0.8041026,0.54482055,0.318359,0.18051283,0.18707694,0.34133336,0.5940513,0.81066674,0.702359,0.5546667,0.512,0.5677949,0.72861546,0.7318975,0.5513847,0.27569234,0.11158975,0.029538464,0.013128206,0.013128206,0.009846155,0.016410258,0.02297436,0.052512825,0.098461546,0.17723078,0.3117949,0.508718,0.77128214,1.024,1.2274873,1.3686155,1.3915899,1.463795,1.5819489,1.7591796,2.03159,2.2777438,2.4910772,2.6289232,2.7044106,2.7963078,2.9997952,3.3312824,3.7448208,4.201026,4.6539493,4.906667,5.0182567,4.824616,4.3716927,3.895795,3.5413337,3.6594875,4.056616,4.601436,5.225026,5.8289237,6.432821,6.961231,7.3058467,7.3353853,4.9296412,4.263385,3.9942567,4.132103,4.5489235,4.972308,5.0051284,4.8311796,4.5817437,4.4307694,4.578462,5.914257,7.50277,9.025641,10.131693,10.427077,10.305642,9.931488,8.809027,7.2303596,6.2818465,7.3616414,7.712821,7.581539,7.1876926,6.75118,7.3583593,8.841846,10.44677,11.759591,12.688411,13.653335,14.191591,14.326155,14.244103,14.290052,13.6237955,12.839386,12.156719,11.644719,11.227899,10.9456415,11.867898,12.973949,13.4629755,12.744206,12.320822,11.608616,9.970873,7.7259493,6.163693,5.5729237,5.1987696,5.0576415,5.0477953,4.923077,4.850872,4.827898,4.7491283,4.588308,4.414359,4.397949,4.7392826,5.2644105,5.8518977,6.416411,5.7107697,5.1987696,5.5893335,6.8463597,8.192,9.176616,7.7948723,5.7435904,3.9056413,2.356513,3.1606157,4.1550775,5.146257,5.602462,4.667077,3.170462,2.481231,2.4320002,2.986667,4.240411,5.8781543,7.282872,8.264206,8.411898,7.1089234,5.6451287,4.8377438,5.3792825,7.2631803,9.80677,9.002667,8.375795,8.057437,8.503796,10.518975,12.511181,13.824001,14.519796,14.844719,15.209026,16.20677,17.959387,20.279797,22.62318,24.096823,23.128616,19.380514,15.320617,12.045129,9.268514,7.8637953,6.987488,6.445949,6.5805135,8.251078,9.216001,9.639385,8.631796,6.550975,5.0084105,5.8912826,5.3398976,4.076308,3.05559,3.4658465,3.006359,1.913436,1.3620514,1.6082052,1.9922053,2.3466668,2.28759,2.0545642,2.028308,2.7273848,3.4658465,4.066462,5.1626673,6.7872825,8.3593855,9.649232,9.878975,9.875693,10.410667,12.2387705,12.944411,12.905026,11.053949,7.778462,4.896821,2.733949,1.6049232,0.94523084,0.5316923,0.47589746,0.5973334,0.72861546,0.7122052,0.5874872,0.574359,0.6826667,0.67282057,0.6104616,0.53825647,0.46933338,0.5513847,0.64000005,0.8402052,1.0929232,1.1716924,1.0929232,1.4276924,1.6016412,1.2964103,0.45620516,0.09189744,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01969231,0.052512825,0.06235898,0.068923086,0.07548718,0.072205134,0.055794876,0.049230773,0.016410258,0.01969231,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.016410258,0.059076928,0.12471796,0.21333335,0.3314872,0.4135385,0.34133336,0.16738462,0.0032820515,0.016410258,0.06564103,0.19364104,0.44964105,0.79097444,1.083077,1.2209232,1.020718,0.67282057,0.34789747,0.20676924,0.118153855,0.03938462,0.0032820515,0.013128206,0.01969231,0.052512825,0.02297436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.049230773,0.009846155,0.0,0.029538464,0.07548718,0.08205129,0.07876924,0.098461546,0.098461546,0.07876924,0.07548718,0.068923086,0.072205134,0.04266667,0.0,0.0,0.009846155,0.006564103,0.0032820515,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.013128206,0.013128206,0.013128206,0.016410258,0.02297436,0.02297436,0.013128206,0.006564103,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.013128206,0.0032820515,0.0,0.0032820515,0.006564103,0.013128206,0.016410258,0.016410258,0.013128206,0.006564103,0.059076928,0.1148718,0.12471796,0.098461546,0.08533334,0.0951795,0.128,0.18051283,0.256,0.3708718,0.5021539,0.64000005,0.69579494,0.6892308,0.72861546,0.8402052,0.892718,0.8763078,0.77128214,0.5481026,0.44964105,0.4135385,0.47589746,0.58420515,0.60061544,0.571077,0.5481026,0.53825647,0.5415385,0.55794877,0.6859488,1.0010257,1.6836925,2.3958976,2.2744617,1.5524104,1.3620514,1.4998976,1.8313848,2.284308,2.9997952,3.4166157,3.3247182,2.789744,2.1333334,1.6180514,1.401436,1.3620514,1.4408206,1.657436,2.038154,2.5665643,3.1442053,3.2984617,2.1792822,0.9353847,0.40369233,0.24287182,0.25928208,0.38728207,0.57764107,0.65969235,0.6695385,0.88943595,1.8412309,3.0523078,3.8629746,3.9811285,3.4560003,2.6518977,4.2962055,5.211898,5.3037953,5.0018463,5.2447186,5.2742567,4.71959,3.9384618,3.3476925,3.446154,4.571898,5.330052,5.786257,5.6254363,4.1583595,3.4822567,4.059898,4.7655387,4.900103,4.1911798,2.553436,2.789744,3.9811285,4.670359,2.8291285,1.7657437,1.5064616,1.6968206,2.0906668,2.5271797,2.9505644,3.3280003,3.564308,3.367385,2.231795,1.8838975,2.3827693,2.3171284,1.4473847,0.7122052,0.571077,0.53825647,0.6662565,1.0601027,1.8904617,3.6791797,5.8814363,6.6527185,6.0258465,5.8912826,6.3868723,5.546667,4.71959,5.0084105,7.243488,6.547693,4.857436,3.2689233,2.422154,2.5206156,3.4625645,4.972308,6.413129,7.3452315,7.522462,5.737026,4.073026,3.2098465,3.3345644,4.161641,5.349744,5.0871797,4.457026,4.1682053,4.562052,5.2611284,5.792821,5.9602056,5.8781543,5.98318,6.4590774,7.581539,8.4053335,8.556309,8.231385,5.8781543,4.4077954,4.1583595,4.4898467,3.764513,2.7798977,2.605949,3.1015387,4.0992823,5.395693,6.1538467,7.3353853,8.694155,9.554052,8.786052,7.4075904,6.36718,5.720616,5.3136415,4.7622566,4.397949,4.1189747,3.7842054,3.5577438,3.9089234,4.391385,4.667077,4.7983594,4.8836927,5.0510774,5.362872,5.477744,5.5269747,5.7107697,6.304821,6.892308,7.568411,8.444718,9.501539,10.594462,11.0605135,11.602052,12.2847185,12.885334,12.895181,12.544001,11.963078,11.569232,11.536411,11.805539,12.708103,13.991385,15.537232,17.122463,18.418873,18.97354,18.960411,18.422155,17.572104,16.820515,16.459488,16.57436,16.984617,17.476925,17.811693,17.56554,17.211079,17.411283,17.962667,17.785437,16.219898,14.742975,13.436719,12.425847,11.894155,11.346052,10.614155,9.580308,8.441437,7.7259493,7.6209235,6.954667,6.2096415,5.7468724,5.792821,5.5302567,5.1987696,5.0051284,4.854154,4.3716927,3.5478978,3.4133337,3.7940516,4.6539493,6.0980515,5.208616,3.7448208,2.425436,1.6738462,1.6016412,2.1333334,2.481231,2.5764105,2.3663592,1.8346668,1.4276924,1.1716924,1.1881026,1.3161026,1.0732309,0.6465641,0.45292312,0.35446155,0.28225642,0.23630771,0.18707694,0.190359,0.31507695,0.63343596,1.2373334,1.6968206,1.3883078,1.0305642,0.9747693,1.1848207,1.5655385,1.6344616,1.3161026,0.764718,0.35446155,0.101743594,0.01969231,0.006564103,0.009846155,0.02297436,0.01969231,0.04266667,0.09189744,0.17394873,0.30851284,0.52512825,0.8172308,1.1257436,1.394872,1.5885129,1.5688206,1.5786668,1.6246156,1.7362052,1.972513,2.2055387,2.3926156,2.5107694,2.5764105,2.6322052,2.806154,3.0785644,3.4231799,3.8432825,4.3585644,4.8377438,5.2512827,5.3924108,5.211898,4.821334,4.197744,3.876103,3.82359,4.0336413,4.5456414,5.175795,5.868308,6.491898,6.931693,7.1023593,5.293949,4.893539,4.460308,4.4012313,4.824616,5.5696416,4.8114877,4.2207184,3.761231,3.4166157,3.1737437,3.3575387,4.7655387,6.11118,6.813539,7.0334363,6.76759,6.5903597,6.5903597,6.9677954,8.041026,8.687591,9.051898,9.094564,8.802463,8.178872,7.9458466,8.503796,9.7214365,11.067078,11.565949,13.115078,15.75713,17.77559,18.58954,18.720821,17.526155,16.705643,16.246155,15.891693,15.120412,14.145642,13.673027,13.177437,12.475078,11.720206,12.3766165,12.232206,11.260718,9.593436,7.506052,5.87159,4.7589746,4.378257,4.568616,4.775385,4.850872,5.0674877,5.3792825,5.661539,5.720616,5.930667,6.311385,6.9645133,7.712821,8.103385,7.24677,6.055385,4.8082056,3.895795,3.7842054,3.5413337,3.0949745,2.3302567,1.3686155,0.5481026,0.36758977,0.38400003,0.574359,0.9321026,1.4802053,2.1989746,3.1573336,3.7448208,4.096,5.097026,6.928411,8.996103,11.090053,12.258463,10.817642,9.170052,7.322257,6.99077,8.234667,9.429334,9.892103,10.522257,11.510155,12.898462,14.572309,16.328207,18.06113,18.835693,18.75036,18.921026,20.04349,21.211899,22.416412,23.364925,23.499489,20.667078,16.810667,12.672001,8.914052,6.117744,5.8880005,6.2687182,6.76759,7.312411,8.241231,7.496206,6.1013336,4.3060517,2.6880002,2.1530259,3.006359,2.6420515,2.038154,1.7690258,2.0151796,1.9528207,1.8838975,1.6213335,1.273436,1.2373334,1.6377437,2.097231,2.4943593,2.740513,2.7766156,4.6080003,6.3376417,7.4141545,7.968821,8.835282,9.908514,10.243283,10.28595,10.308924,10.407386,11.835078,12.796719,12.150155,9.69518,6.180103,1.7985642,0.8763078,1.0272821,1.014154,0.7318975,0.6104616,0.52512825,0.49887183,0.52512825,0.5481026,0.6104616,0.94523084,1.1946667,1.1782565,0.88615394,0.7515898,0.7253334,0.82379496,1.0994873,1.6475899,2.281026,2.231795,1.8051283,1.1520001,0.27569234,0.055794876,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.098461546,0.256,0.3052308,0.34133336,0.37743592,0.35446155,0.23302566,0.0,0.036102567,0.09189744,0.072205134,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.06235898,0.08533334,0.036102567,0.0,0.07548718,0.380718,0.6859488,0.6629744,0.35774362,0.016410258,0.07548718,0.3314872,0.827077,1.2471796,1.4605129,1.5097437,0.9747693,0.58420515,0.3314872,0.17066668,0.0,0.0,0.0,0.02297436,0.06564103,0.09189744,0.01969231,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02297436,0.059076928,0.04594872,0.08205129,0.108307704,0.13456412,0.13784617,0.07548718,0.03938462,0.049230773,0.036102567,0.0,0.0,0.049230773,0.032820515,0.016410258,0.016410258,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.016410258,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.01969231,0.029538464,0.01969231,0.016410258,0.016410258,0.01969231,0.029538464,0.055794876,0.08861539,0.118153855,0.13456412,0.12143591,0.12143591,0.12143591,0.14112821,0.18707694,0.25928208,0.3446154,0.40369233,0.46276927,0.54482055,0.65641034,0.72861546,0.7581539,0.7450257,0.6826667,0.5481026,0.4397949,0.47589746,0.51856416,0.49230772,0.380718,0.27241027,0.24287182,0.318359,0.4594872,0.5940513,0.69251287,0.8533334,1.1979488,1.7001027,2.2121027,2.1136413,2.1530259,2.4352822,2.9440002,3.5544617,3.8596926,3.7251284,3.370667,2.937436,2.487795,2.793026,2.9407182,2.8882053,2.7076926,2.609231,2.7569232,3.1671798,3.1803079,2.5435898,1.4342566,0.67610264,0.3052308,0.19692309,0.27897438,0.5349744,0.7056411,0.6662565,0.6662565,0.8402052,1.204513,2.92759,4.381539,5.395693,5.717334,5.0215387,4.886975,4.962462,4.772103,4.4274874,4.6244106,4.2207184,3.4527183,2.8849232,2.9440002,3.9220517,4.7261543,4.781949,4.4701543,4.1124105,3.95159,3.3542566,3.5971284,4.31918,4.532513,2.6387694,1.9790771,2.0644104,2.0250258,1.6705642,1.4506668,1.2176411,1.3620514,1.7099489,2.0644104,2.1956925,2.3204105,2.605949,2.9111798,2.9997952,2.546872,1.8412309,1.847795,1.7362052,1.1979488,0.44307697,0.32164106,0.30851284,0.40697438,0.6071795,0.8992821,1.2537436,1.7263591,2.2219489,2.6683078,3.0227695,2.9735386,2.6683078,2.3269746,2.0545642,1.847795,1.9331284,1.7066668,1.3751796,1.2274873,1.6180514,2.9111798,4.5062566,5.605744,5.605744,4.1058464,2.6026669,2.1103592,2.103795,2.294154,2.6256413,2.989949,3.6857438,3.9811285,3.69559,3.2196925,3.1967182,3.4724104,3.7973337,4.076308,4.394667,5.467898,6.5706673,6.636308,5.435077,3.5544617,2.2482052,2.1891284,2.5042052,2.605949,2.166154,2.3138463,2.8521028,3.6529233,4.4800005,5.0051284,5.3727183,6.8004107,8.52677,9.750975,9.6295395,8.152616,6.426257,5.1331286,4.5029745,4.332308,4.417641,4.450462,4.315898,4.0303593,3.7382567,4.397949,5.477744,6.180103,6.3573337,6.514872,7.003898,6.941539,6.2818465,5.3398976,4.7917953,5.7665644,7.020308,8.057437,8.825437,9.705027,10.620719,11.424822,12.274873,13.056001,13.397334,13.298873,13.302155,13.328411,13.466257,13.991385,14.834873,15.760411,16.748308,17.664001,18.248207,18.323694,17.893745,17.270155,16.699078,16.357744,16.406975,16.528412,16.699078,16.869745,16.968206,16.626873,16.239592,16.114874,16.246155,16.295385,15.894976,15.343591,14.788924,14.296617,13.869949,13.236514,12.455385,11.378873,10.082462,8.848411,7.8736415,7.253334,6.8332314,6.5247183,6.3179493,6.4754877,6.3245134,6.0225644,5.5663595,4.7622566,3.9187696,3.2951798,3.0260515,3.2656412,4.1813335,5.0116925,4.640821,3.4198978,1.9331284,0.9911796,1.0535386,1.3522053,1.7001027,1.9561027,2.028308,1.467077,1.017436,0.74830776,0.7187693,0.97805136,1.2832822,0.955077,0.56451285,0.380718,0.380718,0.380718,0.318359,0.27569234,0.39384618,0.86974365,1.0272821,0.88615394,0.78769237,0.9288206,1.3423591,1.782154,1.9823592,1.8379488,1.3686155,0.7318975,0.3052308,0.098461546,0.029538464,0.032820515,0.04594872,0.032820515,0.03938462,0.06564103,0.12471796,0.25928208,0.4660513,0.79425645,1.1782565,1.5425643,1.785436,1.723077,1.6804104,1.6869745,1.7755898,1.9823592,2.228513,2.4155898,2.5271797,2.5731285,2.609231,2.7306669,2.92759,3.1967182,3.5282054,3.9056413,4.3585644,4.8016415,5.2348723,5.5893335,5.737026,5.4449234,4.9493337,4.4373336,4.1091285,4.1813335,4.4865646,4.9821544,5.58277,6.173539,6.636308,5.1364107,4.9296412,4.598154,4.1124105,3.6332312,3.5183592,3.698872,4.007385,4.0336413,3.626667,2.8914874,2.550154,2.809436,3.7940516,5.149539,6.0324106,6.340924,6.7544622,6.987488,6.9809237,6.8955903,7.2369237,7.5191803,7.634052,7.7325134,8.201847,9.212719,9.754257,10.105436,10.35159,10.381129,10.801231,11.72677,13.147899,14.674052,15.560206,15.360002,15.432206,15.589745,15.77354,16.049232,14.234258,12.42913,11.132719,10.305642,9.363693,9.242257,10.085744,10.896411,11.080206,10.436924,7.512616,5.0215387,3.9023592,4.1058464,4.6178465,5.110154,5.1200004,5.139693,5.4153852,5.9667697,6.7872825,7.529026,7.9885135,8.008205,7.4929237,6.3245134,4.6572313,3.0949745,2.0250258,1.6114873,1.463795,1.3357949,1.1585642,1.1355898,1.7329233,2.5764105,4.138667,5.8847184,7.5585647,9.18318,9.6295395,9.895386,9.655796,9.235693,9.613129,10.732308,12.432411,13.801026,14.280207,13.650052,12.314258,10.71918,9.143796,7.955693,7.5979495,7.6734366,9.45559,11.972924,14.726565,17.696821,16.866463,16.229744,15.760411,15.228719,14.198155,12.340514,12.566976,13.6008215,14.575591,15.051488,13.459693,11.569232,9.622975,7.939283,6.8988724,6.6592827,6.3573337,5.7534366,4.775385,3.515077,2.917744,2.4385643,2.1136413,1.9987694,2.162872,2.7142565,2.7536411,2.5206156,2.1956925,1.8904617,1.910154,2.0644104,2.4910772,2.9604106,2.8849232,2.4188719,2.3072822,2.6157951,3.3509746,4.460308,5.5991797,6.7971287,8.086975,9.222565,9.688616,9.93477,9.93477,9.67877,9.186462,8.503796,9.872411,10.33518,9.078155,6.4032826,3.7382567,1.1815386,0.5546667,0.5513847,0.512,0.4266667,0.77456415,0.92225647,0.8008206,0.60389745,0.79425645,1.2537436,2.1825643,2.7864618,2.7306669,2.1070771,1.7558975,1.4506668,1.2471796,1.1749744,1.2438976,1.3128207,1.1191796,0.81394875,0.4660513,0.055794876,0.009846155,0.0,0.0,0.0,0.0,0.098461546,0.049230773,0.0,0.0,0.0,0.108307704,0.14112821,0.108307704,0.052512825,0.06235898,0.068923086,0.07548718,0.072205134,0.04594872,0.0,0.006564103,0.01969231,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.06235898,0.10502565,0.10502565,0.08205129,0.06564103,0.07548718,0.13784617,0.13128206,0.17723078,0.38400003,0.8467693,1.2570257,1.3456411,1.2668719,1.1224617,0.9353847,0.60389745,0.3446154,0.17394873,0.072205134,0.0,0.0,0.036102567,0.06564103,0.06235898,0.01969231,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.029538464,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.02297436,0.01969231,0.02297436,0.026256412,0.026256412,0.016410258,0.006564103,0.009846155,0.013128206,0.009846155,0.0,0.01969231,0.013128206,0.0032820515,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0032820515,0.013128206,0.013128206,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.02297436,0.032820515,0.029538464,0.016410258,0.006564103,0.01969231,0.026256412,0.026256412,0.026256412,0.026256412,0.01969231,0.02297436,0.036102567,0.059076928,0.08861539,0.13456412,0.18379489,0.20348719,0.21989745,0.24943592,0.28225642,0.34133336,0.38400003,0.41025645,0.42994875,0.4594872,0.4955898,0.49887183,0.49230772,0.47917953,0.45292312,0.46933338,0.49230772,0.50543594,0.47589746,0.35774362,0.29538465,0.39056414,0.53825647,0.65312827,0.67938465,1.2176411,1.972513,2.7208207,3.2295387,3.2754874,3.0982566,2.8849232,2.8324106,3.0096412,3.3345644,3.9253337,3.8006158,3.31159,2.92759,3.2689233,3.6529233,3.95159,4.0041027,3.7809234,3.3903592,2.609231,1.9922053,1.4572309,0.9682052,0.5316923,0.30194873,0.2231795,0.30194873,0.50543594,0.7417436,0.7253334,0.6695385,0.7056411,0.9616411,1.5721027,3.0687182,4.7392826,5.6385646,5.622154,5.32677,6.1078978,5.9602056,5.1331286,4.007385,3.1113849,2.540308,2.1464617,1.9954873,2.1792822,2.8356924,3.4264617,3.4198978,3.1442053,2.8553848,2.7569232,2.5665643,2.6945643,3.1409233,3.5971284,3.4330258,2.793026,2.4910772,2.0512822,1.4506668,1.1454359,1.0502565,1.0371283,1.4441026,2.15959,2.6256413,1.9659488,1.5655385,1.3193847,1.204513,1.2800001,1.2832822,1.276718,1.0765129,0.6892308,0.3314872,0.26912823,0.30851284,0.4266667,0.57764107,0.7056411,0.79425645,0.9156924,1.0075898,1.0535386,1.1060513,1.2209232,1.1552821,1.024,0.90256417,0.8336411,0.8598975,0.88943595,0.9124103,0.9485129,1.0568206,1.7558975,2.3893335,2.6683078,2.477949,1.8937438,1.3784616,1.1093334,1.0010257,0.99774367,1.0732309,1.2537436,1.5392822,1.7296412,1.7460514,1.6213335,1.7624617,2.0676925,2.4155898,2.7667694,3.1606157,4.381539,6.1440005,7.571693,7.7948723,5.924103,4.0303593,3.0490258,2.8127182,2.9801028,3.0096412,3.7021542,4.2535386,4.647385,4.8738465,4.9329233,5.1626673,6.180103,7.322257,8.044309,7.9327188,6.9809237,5.8945646,5.0018463,4.420923,4.066462,4.1714873,4.5128207,4.6080003,4.4307694,4.420923,7.1909747,9.757539,11.290257,11.040821,8.3593855,7.2172313,6.5805135,5.612308,4.5128207,4.5095387,6.23918,7.0990777,7.282872,7.506052,9.02236,10.171078,10.860309,11.523283,12.258463,12.836103,13.2562065,13.476104,13.489232,13.4170265,13.492514,13.689437,14.020925,14.473847,14.943181,15.248411,15.212309,14.887385,14.480412,14.247386,14.503386,14.697027,14.513232,14.043899,13.495796,13.184001,12.852514,12.422565,12.179693,12.248616,12.609642,13.213539,13.74195,14.007796,13.932309,13.551591,12.95754,12.2157955,11.286975,10.203898,9.068309,8.231385,7.4830775,6.770872,6.121026,5.671385,5.1265645,5.172513,5.428513,5.5926156,5.431795,4.532513,3.5216413,2.5961027,1.9987694,1.9954873,2.484513,2.044718,1.332513,0.7515898,0.4660513,0.5284103,0.8205129,1.1520001,1.3981539,1.4802053,1.142154,0.9156924,0.92225647,1.1224617,1.3292309,1.3226668,1.1093334,0.7384616,0.37415388,0.29538465,0.23630771,0.14441027,0.08205129,0.09189744,0.19692309,0.43651286,0.67610264,0.8730257,1.024,1.1946667,1.2635899,1.2635899,1.1355898,0.8730257,0.49887183,0.2297436,0.08205129,0.029538464,0.036102567,0.059076928,0.055794876,0.04266667,0.055794876,0.1148718,0.2100513,0.41682056,0.72861546,1.1060513,1.463795,1.6869745,1.6836925,1.657436,1.6836925,1.7920002,1.9593848,2.1530259,2.359795,2.550154,2.7011285,2.806154,2.917744,3.1015387,3.3509746,3.639795,3.9318976,4.2272825,4.453744,4.6769233,4.9296412,5.211898,5.4482055,5.481026,5.395693,5.2611284,5.110154,4.9854364,4.8114877,4.7261543,4.8672824,5.3792825,5.280821,4.9362054,4.5029745,3.945026,3.3805132,3.0785644,3.1442053,3.2361028,3.318154,3.2886157,3.006359,2.7569232,2.8356924,3.3542566,4.240411,5.21518,5.835488,6.5312824,7.2861543,8.004924,8.5202055,9.074872,9.173334,9.012513,8.684308,8.192,8.467693,8.832001,9.18318,9.452309,9.609847,9.6065645,9.5835905,9.760821,9.997129,9.780514,9.662359,10.06277,10.870154,11.851488,12.675283,11.746463,10.686359,9.803488,9.360411,9.590155,9.682052,9.954462,10.381129,10.676514,10.308924,7.5881033,5.3694363,4.069744,4.017231,5.4383593,6.2916927,6.370462,6.091488,5.789539,5.6976414,5.940513,6.521436,7.181129,7.509334,6.954667,6.377026,5.648411,5.106872,4.850872,4.71959,4.276513,4.7458467,5.691077,6.7249236,7.522462,8.848411,11.053949,12.76718,13.650052,14.385232,16.354464,16.498873,15.251694,13.994668,15.07118,16.22318,17.391592,18.07754,18.01518,17.168411,14.483693,12.593232,11.277129,10.213744,8.999385,8.937026,10.571488,12.757335,14.79877,16.456207,14.683899,13.679591,13.282462,13.564719,14.818462,14.41477,13.6008215,12.947693,12.609642,12.297847,11.733335,10.676514,9.186462,7.702975,7.076103,6.0061545,4.1714873,2.6584618,1.7788719,1.0699488,1.1191796,1.273436,1.5786668,1.9889232,2.3696413,2.6453335,2.7109745,2.7733335,2.878359,2.9144619,2.0873847,1.6902566,1.8018463,2.3762052,3.249231,3.3641028,2.8947694,2.9702566,3.948308,5.3858466,6.0652313,6.921847,8.021334,8.946873,8.776206,8.402052,7.965539,7.4469748,6.8365135,6.1407185,5.868308,5.284103,4.086154,2.5731285,1.6278975,0.8369231,0.5415385,0.47589746,0.4955898,0.56123084,0.7318975,0.761436,0.5415385,0.3249231,0.7253334,1.1848207,1.8379488,2.2186668,2.1464617,1.723077,1.276718,0.9124103,0.65312827,0.508718,0.4660513,0.42994875,0.34133336,0.23630771,0.12471796,0.0,0.052512825,0.059076928,0.032820515,0.0,0.0,0.049230773,0.06235898,0.08205129,0.1148718,0.13784617,0.14769232,0.12471796,0.06564103,0.0032820515,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.02297436,0.04266667,0.12471796,0.17723078,0.14112821,0.0,0.2986667,0.6268718,1.0699488,1.5491283,1.8248206,1.8215386,1.3850257,0.8992821,0.56123084,0.380718,0.32164106,0.25928208,0.14769232,0.01969231,0.0,0.0,0.01969231,0.029538464,0.02297436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.068923086,0.06564103,0.036102567,0.009846155,0.009846155,0.009846155,0.0032820515,0.0,0.0,0.0,0.013128206,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.0032820515,0.0032820515,0.006564103,0.006564103,0.013128206,0.013128206,0.006564103,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.02297436,0.026256412,0.01969231,0.006564103,0.0,0.006564103,0.01969231,0.016410258,0.013128206,0.009846155,0.006564103,0.013128206,0.02297436,0.03938462,0.059076928,0.09189744,0.13128206,0.15425642,0.18707694,0.23958977,0.30851284,0.35774362,0.39056414,0.39056414,0.3708718,0.38400003,0.41025645,0.41682056,0.42338464,0.4397949,0.49230772,0.5481026,0.571077,0.6465641,0.76800007,0.8369231,0.7417436,0.8960001,1.1618463,1.4309745,1.6082052,2.481231,3.5807183,3.9417439,3.4789746,2.9801028,2.989949,2.868513,2.7208207,2.5698464,2.356513,2.5600002,2.6256413,2.740513,3.0194874,3.4921029,3.7021542,4.164923,4.5554876,4.516103,3.639795,2.4451284,1.2931283,0.61374366,0.43323082,0.3708718,0.3446154,0.3446154,0.41682056,0.58092314,0.8467693,0.82379496,0.69579494,0.892718,1.5688206,2.6157951,3.879385,5.028103,5.5171285,5.1856413,4.266667,4.634257,4.916513,4.532513,3.4855387,2.3663592,1.595077,1.2832822,1.3161026,1.7493335,2.7831798,3.6069746,4.023795,3.7907696,3.1343591,2.7503593,2.7602053,2.7602053,2.806154,2.917744,3.0818465,2.5074873,1.7132308,1.1191796,0.8566154,0.77456415,0.71548724,0.69579494,0.8992821,1.3259488,1.7788719,1.5097437,1.2340513,0.92553854,0.65641034,0.57764107,0.6859488,0.65969235,0.5152821,0.3446154,0.31507695,0.36102566,0.44307697,0.58092314,0.75487185,0.8763078,0.86317956,0.8041026,0.69579494,0.57764107,0.56123084,0.6465641,0.67610264,0.63343596,0.54482055,0.47917953,0.49230772,0.51856416,0.55794877,0.67282057,1.017436,1.719795,2.3105643,2.550154,2.3860514,1.975795,1.2800001,0.90584624,0.75487185,0.69579494,0.5677949,0.57764107,0.6892308,0.8992821,1.1520001,1.3128207,1.2406155,1.3817437,1.6640002,1.9954873,2.284308,3.2722054,5.139693,7.02359,8.080411,7.4863596,4.8672824,3.4100516,3.114667,3.4756925,3.4658465,4.3618464,5.5893335,5.8157954,4.841026,3.5872824,3.6791797,4.4898467,5.612308,6.416411,6.052103,5.349744,4.788513,4.3290257,3.9844105,3.82359,4.394667,4.6966157,4.634257,4.4996924,4.9394875,6.7938466,8.146052,8.766359,8.441437,6.987488,6.3540516,6.055385,5.8781543,5.7009234,5.474462,5.4514875,5.139693,5.1856413,5.973334,7.634052,8.15918,8.720411,9.521232,10.525539,11.460924,12.1468725,12.419283,12.340514,12.041847,11.72677,11.618463,11.61518,11.746463,11.926975,11.969642,12.009027,12.068104,11.98277,11.798975,11.739899,11.766154,11.529847,11.1064625,10.66995,10.489437,10.371283,10.177642,10.134975,10.371283,10.929232,12.084514,13.013334,13.5089245,13.423591,12.678565,11.723488,10.807796,9.908514,9.042052,8.2445135,7.6077952,7.076103,6.5706673,6.183385,6.1768208,5.9634876,5.4843082,5.0871797,4.8705645,4.6933336,3.9548721,3.05559,2.1924105,1.5688206,1.394872,1.6377437,1.4244103,1.1158975,0.95835906,1.086359,1.1618463,1.2635899,1.3029745,1.270154,1.2242053,1.0535386,0.92553854,0.92553854,1.0272821,1.0994873,0.86646163,0.6498462,0.42994875,0.24287182,0.18379489,0.118153855,0.055794876,0.02297436,0.01969231,0.029538464,0.21333335,0.42994875,0.6071795,0.7253334,0.81066674,0.82379496,0.8795898,0.8533334,0.6826667,0.3708718,0.17394873,0.06235898,0.02297436,0.02297436,0.032820515,0.026256412,0.016410258,0.032820515,0.08205129,0.15097436,0.3446154,0.6235898,0.9714873,1.3226668,1.5360001,1.591795,1.5885129,1.6082052,1.6869745,1.8149745,1.9987694,2.1924105,2.4057438,2.6190772,2.806154,2.9768207,3.1803079,3.4166157,3.6824617,3.9647183,4.1485133,4.269949,4.352,4.457026,4.6867695,4.9788723,5.2315903,5.467898,5.684513,5.835488,5.5729237,5.1856413,4.824616,4.7360005,5.277539,5.927385,5.9930263,6.0356927,5.677949,4.9394875,4.2436924,3.761231,3.4067695,3.2984617,3.3805132,3.4330258,3.442872,3.6890259,4.086154,4.6211286,5.349744,5.3792825,5.8092313,6.705231,7.8834877,8.910769,9.67877,9.95118,9.757539,9.101129,7.958975,7.5585647,7.824411,8.4972315,9.137232,9.120821,8.848411,8.530052,8.090257,7.463385,6.619898,6.422975,6.695385,7.4174366,8.392206,9.248821,9.396514,9.419488,9.409642,9.67877,10.735591,11.766154,12.074668,12.045129,11.670976,10.535385,8.195283,6.5444107,5.504,5.356308,6.7314878,7.2894363,7.1876926,6.5378466,5.6352825,4.9821544,4.6605134,4.906667,5.4875903,6.009436,5.930667,5.654975,5.6385646,6.1472826,7.2894363,9.02236,10.673231,12.924719,14.92677,15.954053,15.412514,15.602873,16.594053,17.601643,18.22195,18.46154,20.358566,21.001848,20.565334,20.09272,21.504002,21.461334,21.152822,21.074053,20.906668,19.524925,15.9573345,13.10195,11.372309,10.735591,10.732308,11.447796,12.84595,13.856822,13.935591,13.062565,10.102155,9.189744,9.557334,11.277129,15.271386,16.479181,15.704617,14.36554,13.108514,11.792411,10.584617,9.238976,7.581539,5.858462,4.7261543,3.7743592,2.4320002,1.4145643,0.9485129,0.80738467,0.8795898,1.0765129,1.3915899,1.7788719,2.166154,2.5632823,2.9571285,3.117949,3.1967182,3.751385,4.378257,4.2174363,3.7776413,3.495385,3.751385,4.2305646,4.4242053,4.637539,5.074052,5.8125134,6.2096415,6.7314878,7.3419495,7.6077952,6.701949,5.914257,5.277539,4.6244106,3.9581542,3.436308,3.0687182,2.5140514,1.8510771,1.211077,0.7844103,0.5874872,0.4594872,0.42994875,0.48574364,0.5874872,0.60061544,0.571077,0.42338464,0.29538465,0.51856416,0.72861546,0.9944616,1.1158975,1.0404103,0.85005134,0.54482055,0.31507695,0.15425642,0.059076928,0.026256412,0.009846155,0.006564103,0.009846155,0.009846155,0.006564103,0.055794876,0.06564103,0.036102567,0.0,0.0,0.0,0.068923086,0.12471796,0.14112821,0.13784617,0.09189744,0.055794876,0.02297436,0.0032820515,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.029538464,0.006564103,0.0,0.0,0.0,0.0,0.0,0.07548718,0.13456412,0.20020515,0.4135385,0.82379496,1.2209232,1.6443079,1.9528207,1.8510771,1.3718976,0.8795898,0.50543594,0.32164106,0.3314872,0.30194873,0.2100513,0.09189744,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.036102567,0.052512825,0.02297436,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.068923086,0.06564103,0.036102567,0.009846155,0.009846155,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.009846155,0.02297436,0.02297436,0.009846155,0.0,0.0,0.0,0.006564103,0.009846155,0.006564103,0.0,0.0,0.0032820515,0.006564103,0.0032820515,0.0032820515,0.009846155,0.009846155,0.006564103,0.0032820515,0.0,0.0,0.006564103,0.0032820515,0.0,0.0,0.0,0.013128206,0.02297436,0.032820515,0.04266667,0.049230773,0.06235898,0.08205129,0.118153855,0.17394873,0.23958977,0.28882053,0.3314872,0.34789747,0.35446155,0.39056414,0.40369233,0.41025645,0.42338464,0.44964105,0.49887183,0.5152821,0.5415385,0.827077,1.5097437,2.6420515,2.2121027,1.7526156,1.7952822,2.3040001,2.6945643,3.442872,4.138667,4.020513,3.1376412,2.3401027,2.2908719,2.2022567,1.9987694,1.7329233,1.591795,2.0611284,2.5731285,3.2000003,3.817026,4.076308,4.07959,4.33559,4.59159,4.453744,3.383795,1.8904617,0.7975385,0.30194873,0.30194873,0.39384618,0.43323082,0.44964105,0.5513847,0.7450257,0.93866676,0.72861546,0.64000005,0.99774367,1.9528207,3.4822567,4.7917953,5.792821,5.9536414,5.211898,3.9548721,3.748103,3.8596926,3.570872,2.7208207,1.719795,1.020718,0.8008206,0.9321026,1.404718,2.3138463,2.8816411,3.2295387,3.0129232,2.5304618,2.7306669,2.9702566,2.7963078,2.4057438,1.9954873,1.7690258,1.4178462,0.79097444,0.45620516,0.5218462,0.6465641,0.61374366,0.5415385,0.508718,0.58420515,0.8041026,0.8795898,0.8369231,0.69251287,0.49230772,0.3249231,0.36758977,0.35774362,0.30851284,0.27569234,0.33805132,0.4135385,0.47589746,0.5677949,0.6892308,0.8041026,0.8008206,0.73517954,0.6465641,0.5907693,0.6235898,0.6301539,0.64000005,0.5940513,0.48574364,0.37415388,0.34789747,0.33476925,0.40697438,0.6662565,1.2373334,1.6935385,2.156308,2.4681027,2.4681027,1.9790771,1.142154,0.85005134,0.78769237,0.7253334,0.52512825,0.47261542,0.5218462,0.702359,0.9616411,1.1782565,1.0568206,1.0765129,1.2209232,1.4276924,1.595077,2.284308,3.8432825,5.973334,7.9524107,8.664616,6.9349747,5.156103,4.378257,4.785231,5.7009234,5.72718,6.0947695,5.796103,4.571898,2.9078977,2.3171284,2.9702566,4.1058464,4.9493337,4.7327185,3.9187696,3.245949,2.809436,2.6584618,2.7864618,3.6102567,3.7382567,3.5872824,3.639795,4.420923,5.8453336,6.9382567,7.2369237,6.9743595,7.0793853,7.6176414,7.131898,6.5017443,5.970052,5.113436,3.7907696,2.7109745,2.7306669,3.826872,5.0642056,5.218462,5.684513,6.4722056,7.529026,8.730257,9.537642,9.947898,10.052924,9.944616,9.714872,9.511385,9.255385,9.03877,8.874667,8.690872,8.746667,8.976411,9.147078,9.163487,9.055181,9.019077,8.858257,8.635077,8.470975,8.553026,8.704,8.838565,9.078155,9.508103,10.171078,11.497026,12.675283,13.5548725,13.810873,12.921437,11.841642,10.791386,9.645949,8.461129,7.4699492,7.0531287,6.6494365,6.2129235,5.8157954,5.6287184,5.431795,4.785231,4.2863593,4.132103,4.1091285,3.3247182,2.5206156,1.7985642,1.3062565,1.2307693,1.3784616,1.4900514,1.595077,1.7558975,2.0873847,1.9922053,1.8084104,1.5261539,1.2668719,1.2832822,1.273436,1.1552821,1.0371283,0.9517949,0.8730257,0.5481026,0.3249231,0.22646156,0.20676924,0.16410258,0.10502565,0.068923086,0.059076928,0.06564103,0.07876924,0.18379489,0.26584616,0.3117949,0.33476925,0.38400003,0.45620516,0.67938465,0.7975385,0.6892308,0.37415388,0.190359,0.06564103,0.013128206,0.009846155,0.009846155,0.0032820515,0.0,0.016410258,0.055794876,0.1148718,0.28882053,0.5284103,0.84348726,1.1749744,1.3751796,1.4867693,1.5261539,1.5589745,1.6180514,1.7132308,1.8609232,2.0217438,2.2121027,2.4418464,2.6978464,2.9440002,3.1540515,3.3509746,3.5511796,3.751385,3.945026,4.1222568,4.279795,4.4242053,4.588308,4.7360005,4.9493337,5.21518,5.5007186,5.7731285,5.5991797,5.349744,5.1331286,5.159385,5.733744,7.453539,7.860513,8.267488,7.88677,6.698667,5.4613338,4.647385,4.4110775,4.4077954,4.4274874,4.4045134,4.460308,4.778667,5.35959,6.0258465,6.439385,5.618872,5.4580517,5.9470773,6.8430777,7.6898465,8.241231,8.717129,8.736821,8.260923,7.5881033,7.2336416,7.3353853,8.011488,8.786052,8.572719,8.241231,8.162462,8.119796,7.955693,7.571693,7.2992826,6.99077,6.806975,6.882462,7.3091288,7.762052,8.152616,8.713847,9.524513,10.505847,12.278154,13.292309,13.426873,12.635899,10.94236,9.189744,8.136206,7.568411,7.387898,7.6110773,7.315693,6.744616,5.7796926,4.670359,4.0467696,3.82359,4.023795,4.3749747,4.827898,5.579488,6.045539,6.816821,8.264206,10.5780525,13.745232,17.762463,21.234873,23.250053,23.273027,21.152822,19.62995,18.678156,18.868515,19.938463,20.78195,21.175797,22.298258,23.282873,23.811283,24.103386,22.170258,20.33559,19.712002,19.75795,18.281027,15.510976,12.409437,9.997129,9.18318,10.774975,12.491488,13.702565,13.525334,11.835078,9.229129,5.4843082,4.4996924,5.287385,7.6307697,12.087796,13.403898,13.659899,13.266052,12.406155,11.017847,8.749949,6.6395903,4.71959,2.9636924,1.2635899,1.3784616,2.0775387,2.422154,2.162872,1.7362052,1.1749744,1.0305642,1.079795,1.2176411,1.4703591,2.4648206,3.56759,3.7907696,3.5183592,4.4964104,7.9294367,8.5202055,7.719385,6.488616,5.3103595,5.3431797,6.2523084,6.6067696,6.121026,5.674667,5.6451287,5.664821,5.651693,5.3431797,4.263385,3.4691284,2.986667,2.5074873,2.0020514,1.7066668,2.5600002,2.930872,2.9111798,2.4516926,1.3522053,0.7220513,0.508718,0.47261542,0.48246157,0.49887183,0.55794877,0.5907693,0.6071795,0.56123084,0.36430773,0.29210258,0.35774362,0.38728207,0.32164106,0.21989745,0.15097436,0.11158975,0.08205129,0.055794876,0.036102567,0.016410258,0.0032820515,0.0032820515,0.009846155,0.013128206,0.013128206,0.01969231,0.013128206,0.0,0.0,0.0,0.06235898,0.08861539,0.055794876,0.009846155,0.013128206,0.009846155,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016410258,0.08205129,0.026256412,0.0032820515,0.0,0.0,0.0,0.0,0.006564103,0.013128206,0.190359,0.86317956,1.083077,1.2274873,1.2931283,1.2307693,0.93866676,0.4135385,0.27241027,0.28225642,0.35446155,0.5513847,0.38400003,0.13784617,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.072205134,0.101743594,0.04266667,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.01969231,0.049230773,0.029538464,0.009846155,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.02297436,0.029538464,0.02297436,0.009846155,0.0032820515,0.0032820515,0.0032820515,0.009846155,0.009846155,0.0,0.0,0.0032820515,0.0032820515,0.0032820515,0.0,0.0,0.009846155,0.026256412,0.03938462,0.055794876,0.06564103,0.06564103,0.072205134,0.08861539,0.11158975,0.128,0.16410258,0.21333335,0.26256412,0.318359,0.38728207,0.4004103,0.40369233,0.43323082,0.47917953,0.49887183,0.47917953,0.512,0.9156924,2.0053334,4.092718,3.4756925,2.4320002,2.156308,2.737231,3.170462,3.387077,3.2525132,2.917744,2.4418464,1.7920002,1.5753847,1.4605129,1.3029745,1.270154,1.847795,3.249231,4.352,5.1364107,5.5597954,5.579488,5.4613338,5.149539,4.6867695,3.9975388,2.8816411,1.2438976,0.5152821,0.2986667,0.3249231,0.43651286,0.44964105,0.44307697,0.5940513,0.8467693,0.9353847,0.54482055,0.6071795,1.1749744,2.3269746,4.1747694,5.674667,6.6067696,6.262154,5.028103,4.4045134,4.082872,3.4297438,2.7241027,2.0611284,1.3620514,0.9189744,0.78769237,0.892718,1.1290257,1.3817437,1.3357949,1.1946667,1.0043077,1.1224617,2.2088206,2.5042052,2.162872,1.5491283,0.8992821,0.318359,0.24943592,0.26256412,0.36102566,0.51856416,0.69251287,0.7122052,0.5513847,0.39384618,0.31507695,0.28882053,0.30194873,0.30851284,0.318359,0.32820517,0.318359,0.34789747,0.39712822,0.43651286,0.4594872,0.4594872,0.47917953,0.46933338,0.44964105,0.43323082,0.44964105,0.48574364,0.4955898,0.5316923,0.6071795,0.67938465,0.6465641,0.61374366,0.5513847,0.44964105,0.3249231,0.24615386,0.25928208,0.5349744,1.0601027,1.657436,1.6082052,1.5458462,1.6180514,1.6672822,1.2373334,0.7318975,0.72861546,0.7975385,0.7417436,0.5907693,0.571077,0.62030774,0.71548724,0.8041026,0.8402052,0.8598975,0.85005134,0.88615394,0.9878975,1.1355898,1.6016412,2.8291285,5.159385,7.8047185,8.835282,8.720411,6.921847,5.6418467,6.052103,8.300308,7.7390776,6.488616,5.402257,4.601436,3.4560003,2.1956925,2.7503593,3.6627696,4.1780515,4.2436924,3.0162053,1.8051283,1.0699488,0.94523084,1.2340513,1.8609232,1.8806155,1.8281027,2.0775387,2.8291285,4.8377438,6.8332314,7.706257,7.6898465,8.349539,9.619693,8.651488,6.957949,5.4843082,4.6178465,3.511795,2.3860514,1.9396925,2.169436,2.3827693,2.4057438,2.7044106,3.1967182,3.9089234,4.97559,5.7107697,6.2720003,6.7216415,7.072821,7.2992826,7.2205133,6.9054365,6.47877,6.0685134,5.7665644,5.7009234,5.7796926,6.0192823,6.3573337,6.6494365,6.7774363,6.7610264,6.705231,6.741334,7.026872,7.427283,7.8703594,8.362667,8.94359,9.6984625,10.971898,12.389745,13.771488,14.5952835,13.988104,13.203693,12.268309,11.126155,9.800206,8.392206,7.5946674,6.7610264,5.8847184,4.969026,4.017231,3.3608208,3.0227695,3.1113849,3.495385,3.8006158,2.9046156,2.1169233,1.4506668,1.0108719,0.98133343,1.0896411,1.3456411,1.6869745,2.0644104,2.4320002,2.2646155,2.1891284,2.1825643,2.15959,2.0053334,1.8281027,1.5655385,1.3029745,1.083077,0.8992821,0.56451285,0.35774362,0.2855385,0.3052308,0.3052308,0.3249231,0.4201026,0.47917953,0.4594872,0.37743592,0.3249231,0.24943592,0.15425642,0.072205134,0.07548718,0.18379489,0.51856416,0.75487185,0.7417436,0.50543594,0.2855385,0.1148718,0.02297436,0.0032820515,0.0,0.0,0.0032820515,0.016410258,0.049230773,0.11158975,0.26912823,0.47917953,0.761436,1.0666667,1.2832822,1.4572309,1.5556924,1.6213335,1.6935385,1.7788719,1.8806155,1.9987694,2.1530259,2.3630772,2.6551797,2.9702566,3.170462,3.3050258,3.3969233,3.4166157,3.6562054,3.95159,4.309334,4.663795,4.8771286,4.9427695,4.9952826,5.024821,5.037949,5.0510774,5.031385,5.0576415,5.2414365,5.6418467,6.301539,10.407386,8.979693,7.4765134,5.933949,4.532513,3.6168208,3.3608208,4.532513,5.832206,6.5280004,6.4557953,6.052103,6.088206,6.619898,7.3682055,7.719385,7.719385,7.3649235,7.210667,7.496206,8.116513,7.640616,7.276308,7.1581545,7.269744,7.4141545,7.171283,6.4689236,6.091488,6.413129,7.4010262,7.890052,8.441437,9.350565,10.305642,10.390975,9.609847,8.178872,6.8529234,6.0160003,5.661539,5.293949,4.97559,4.9920006,5.3924108,5.9667697,6.7117953,7.0432825,7.2336416,7.453539,7.781744,8.198565,8.592411,8.385642,7.5881033,6.806975,5.914257,4.9952826,4.1222568,3.4592824,3.2656412,3.9122055,4.9526157,5.8453336,6.8004107,8.789334,13.08554,16.94195,20.279797,22.288412,21.421951,21.044514,20.775387,20.404514,19.761232,18.724104,18.100513,17.650873,17.161848,17.11918,18.707693,19.892515,20.14195,18.743795,15.996719,13.213539,11.749744,10.8996935,10.660104,10.712616,10.407386,10.420513,10.696206,10.299078,9.140513,7.9819493,8.897642,9.032206,8.306872,7.0793853,6.163693,5.2611284,4.322462,3.7415388,3.639795,3.8596926,4.7294364,5.6320004,6.5772314,7.525744,8.392206,8.625232,6.567385,4.204308,2.5074873,1.4342566,1.8116925,2.2547693,2.5665643,2.5435898,1.9692309,1.1618463,1.017436,1.0108719,0.8960001,0.702359,2.5928206,4.2568207,4.965744,5.2020516,6.669129,9.147078,8.89436,8.011488,7.716103,8.362667,7.5913854,6.5312824,5.7796926,5.330052,4.562052,3.4034874,2.5731285,2.0545642,1.9429746,2.4582565,2.4943593,2.3926156,2.6354873,3.18359,3.4625645,3.2918978,3.4789746,3.6791797,3.5380516,2.6715899,2.0118976,1.4539489,1.1093334,0.96492314,0.8533334,0.84348726,0.79425645,0.7253334,0.6301539,0.47261542,0.36430773,0.27241027,0.2231795,0.20676924,0.18379489,0.036102567,0.0,0.0,0.0,0.0,0.0,0.0,0.01969231,0.036102567,0.0,0.013128206,0.04266667,0.036102567,0.0,0.0,0.0,0.01969231,0.029538464,0.032820515,0.04594872,0.059076928,0.052512825,0.026256412,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02297436,0.108307704,0.068923086,0.02297436,0.0,0.0,0.0,0.0,0.026256412,0.068923086,0.118153855,0.16738462,0.19364104,0.20676924,0.19692309,0.19692309,0.3052308,0.5973334,0.5152821,0.24615386,0.016410258,0.07548718,0.06564103,0.02297436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02297436,0.108307704,0.108307704,0.052512825,0.016410258,0.016410258,0.016410258,0.016410258,0.016410258,0.009846155,0.0,0.0,0.013128206,0.016410258,0.009846155,0.0,0.0,0.0,0.026256412,0.08205129,0.15097436,0.21333335,0.21333335,0.20348719,0.18707694,0.16410258,0.15097436,0.14112821,0.14769232,0.15753847,0.18051283,0.2297436,0.28882053,0.3511795,0.44307697,0.571077,0.7187693,0.81394875,0.8467693,0.76800007,0.7122052,0.9911796,1.4802053,1.8773335,2.103795,2.169436,2.1825643,1.9495386,1.6738462,1.3915899,1.1946667,1.204513,1.4998976,1.7001027,2.0053334,2.6157951,3.7382567,5.47118,7.003898,7.893334,8.14277,8.178872,8.080411,7.2336416,5.943795,4.394667,2.6256413,1.4769232,0.71548724,0.4955898,0.65641034,0.7187693,0.5349744,0.37743592,0.29210258,0.33805132,0.5940513,0.72861546,0.90912825,1.9659488,3.8334363,5.5532312,6.8496413,6.0816417,4.1124105,2.5009232,3.5249233,3.6332312,2.8849232,2.353231,2.3368206,2.349949,1.847795,1.4769232,1.2077949,1.1126155,1.3587693,1.5163078,1.6016412,1.585231,1.4900514,1.404718,0.9288206,0.5513847,0.3446154,0.26912823,0.18379489,0.13456412,0.13128206,0.19692309,0.3249231,0.47261542,0.5218462,0.47917953,0.3708718,0.26584616,0.28882053,0.30194873,0.27897438,0.25271797,0.24287182,0.24287182,0.34133336,0.4660513,0.60061544,0.72861546,0.8402052,0.8402052,0.764718,0.65641034,0.5218462,0.3511795,0.33805132,0.33476925,0.32820517,0.31507695,0.28882053,0.26584616,0.3249231,0.3708718,0.3708718,0.33476925,0.2855385,0.4135385,0.97805136,1.8412309,2.425436,2.425436,1.847795,1.1848207,0.761436,0.74830776,0.77128214,0.761436,0.73517954,0.702359,0.64000005,0.6301539,0.761436,0.88615394,0.8763078,0.65641034,0.508718,0.446359,0.574359,0.86646163,1.1585642,1.4408206,2.9571285,5.093744,6.747898,6.3310776,5.024821,4.096,4.017231,4.857436,6.2884107,8.851693,8.950154,7.6077952,5.786257,4.394667,4.161641,4.818052,5.3005133,5.1232824,4.378257,2.6322052,1.401436,0.65641034,0.37743592,0.5481026,0.7089231,0.86646163,0.90256417,0.86317956,0.9616411,2.1103592,2.9440002,3.5610259,4.2601027,5.5532312,6.38359,6.5378466,6.7577443,7.499488,8.92718,8.717129,7.75877,5.8912826,3.639795,2.2121027,1.1979488,1.020718,1.1355898,1.2635899,1.3751796,1.6804104,2.0020514,2.3433847,2.7241027,3.1737437,3.564308,3.7809234,3.8596926,3.8137438,3.6332312,3.4002054,3.2689233,3.3411283,3.6102567,3.95159,4.2929235,4.5062566,4.7392826,5.074052,5.540103,6.160411,6.8660517,7.5913854,8.369231,9.3078985,10.551796,11.963078,13.13477,13.75836,13.610668,13.292309,12.895181,13.216822,13.860104,13.213539,10.259693,7.9097443,5.970052,4.4438977,3.5413337,2.9407182,2.5829747,2.4484105,2.4582565,2.4582565,2.0906668,1.6246156,1.2274873,0.95835906,0.761436,0.6170257,0.46933338,0.4201026,0.5284103,0.80738467,1.4309745,2.7503593,4.6112823,5.802667,4.0434875,2.674872,1.9692309,1.5589745,1.2668719,1.083077,0.67938465,0.43323082,0.34789747,0.4135385,0.6104616,0.9517949,1.5589745,1.8838975,1.7329233,1.2832822,0.76800007,0.37415388,0.13784617,0.03938462,0.016410258,0.06564103,0.25928208,0.48574364,0.65312827,0.702359,0.43323082,0.21989745,0.08533334,0.02297436,0.0,0.0,0.009846155,0.026256412,0.06564103,0.13784617,0.28225642,0.48574364,0.74830776,1.0502565,1.3423591,1.6344616,1.7920002,1.8904617,1.9856411,2.1202054,2.231795,2.3302567,2.4648206,2.6683078,2.9604106,3.314872,3.5314875,3.629949,3.6135387,3.4789746,3.5511796,3.754667,4.125539,4.6080003,5.034667,5.366154,5.3366156,5.1232824,4.8311796,4.5029745,4.453744,4.604718,5.0674877,5.8125134,6.669129,6.5739493,5.976616,5.802667,5.7665644,5.5597954,4.84759,4.210872,4.5128207,5.21518,5.933949,6.416411,6.7085133,6.954667,7.1056414,6.928411,6.012718,6.186667,6.5837955,6.9349747,7.1089234,7.1154876,6.688821,7.4699492,8.464411,8.982975,8.661334,7.8014364,6.931693,6.9677954,7.9458466,9.02236,9.813334,9.908514,9.655796,9.291488,8.92718,8.1066675,6.738052,5.6254363,4.97559,4.417641,3.620103,3.2951798,3.249231,3.255795,3.0490258,3.314872,4.0041027,4.8344617,5.6254363,6.3179493,6.770872,7.1056414,7.1515903,7.000616,7.000616,6.987488,6.918565,7.0859494,7.6110773,8.441437,9.291488,10.164514,10.988309,12.137027,14.427898,17.729643,20.824617,23.256617,24.497232,23.962257,20.099283,17.273438,15.954053,15.845745,15.891693,15.698052,13.922462,12.051693,11.063796,11.421539,12.320822,12.911591,12.626052,11.697231,11.139283,11.441232,11.874462,12.09436,11.792411,10.686359,10.04636,9.45559,8.89436,8.395488,8.067283,8.237949,8.044309,7.5421543,6.8693337,6.23918,5.149539,3.7809234,3.0851285,3.117949,3.05559,2.3991797,2.546872,3.2000003,4.056616,4.8147697,4.900103,3.9581542,3.0687182,2.6945643,2.6551797,2.858667,3.255795,3.7874875,4.086154,3.495385,2.9997952,3.5544617,4.31918,4.8607183,5.1331286,4.699898,5.0510774,5.9930263,7.125334,7.827693,8.536616,7.955693,6.7577443,5.3694363,3.9548721,3.3312824,2.7241027,2.349949,2.2121027,2.097231,1.9626669,2.0906668,2.3729234,2.7963078,3.446154,3.8531284,4.007385,3.9220517,3.6758976,3.3903592,2.92759,3.0982566,3.2886157,3.0720003,2.2055387,1.8707694,1.6902566,1.4834872,1.2012309,0.96492314,0.7975385,0.7220513,0.67610264,0.56451285,0.28882053,0.16082053,0.108307704,0.098461546,0.101743594,0.098461546,0.01969231,0.0,0.0,0.0,0.0,0.0,0.006564103,0.009846155,0.009846155,0.013128206,0.0032820515,0.009846155,0.006564103,0.0,0.0,0.0,0.0032820515,0.006564103,0.006564103,0.009846155,0.013128206,0.009846155,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.02297436,0.068923086,0.108307704,0.16738462,0.24943592,0.17723078,0.0,0.0,0.0,0.006564103,0.013128206,0.098461546,0.4004103,0.47261542,0.43323082,0.45620516,0.55794877,0.5973334,0.22646156,0.101743594,0.049230773,0.0032820515,0.016410258,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.013128206,0.013128206,0.013128206,0.013128206,0.013128206,0.0032820515,0.0,0.006564103,0.032820515,0.052512825,0.04594872,0.036102567,0.026256412,0.026256412,0.016410258,0.016410258,0.013128206,0.013128206,0.013128206,0.02297436,0.026256412,0.029538464,0.036102567,0.036102567,0.036102567,0.04266667,0.098461546,0.19364104,0.27569234,0.36102566,0.4201026,0.4266667,0.40697438,0.43323082,0.39056414,0.26584616,0.2297436,0.31507695,0.4135385,0.35446155,0.37415388,0.4594872,0.60389745,0.79097444,0.9353847,0.9517949,0.90912825,0.88943595,1.0043077,1.1224617,1.214359,1.276718,1.2800001,1.1454359,0.9517949,0.80738467,0.8205129,1.0469744,1.4998976,1.9003079,2.4484105,3.6004105,5.3070774,7.0465646,8.536616,9.685334,10.295795,10.33518,9.911796,9.07159,7.75877,5.989744,3.9975388,2.2449234,1.1191796,0.67610264,0.5513847,0.52512825,0.49887183,0.51856416,0.53825647,0.53825647,0.5546667,0.69251287,0.8763078,1.1716924,1.8510771,2.9669745,4.345436,4.6539493,4.086154,3.3772311,3.0424619,3.4133337,3.2820516,2.8422565,2.3860514,2.169436,2.4352822,2.8914874,3.4330258,3.8334363,4.066462,4.2994876,4.020513,3.446154,2.7569232,2.2088206,2.1234872,1.785436,1.1585642,0.63343596,0.36758977,0.29210258,0.2231795,0.16410258,0.16410258,0.2297436,0.3249231,0.37415388,0.34133336,0.28225642,0.24615386,0.23958977,0.3314872,0.4135385,0.4594872,0.45620516,0.4266667,0.36758977,0.38728207,0.48902568,0.65312827,0.85005134,0.81394875,0.67938465,0.5349744,0.43651286,0.4135385,0.4201026,0.40697438,0.39712822,0.38728207,0.36430773,0.33805132,0.31507695,0.29538465,0.27569234,0.23958977,0.27569234,0.702359,1.2996924,1.785436,1.8051283,1.6771283,1.3817437,1.0338463,0.77128214,0.761436,0.79425645,0.7187693,0.6071795,0.52512825,0.5316923,0.65641034,0.88943595,1.0765129,1.1191796,0.99774367,0.8402052,0.7318975,0.7089231,0.8566154,1.3062565,2.3958976,3.882667,4.926359,5.034667,4.06318,3.56759,3.6890259,4.3027697,5.146257,5.8223596,6.442667,6.5280004,6.1013336,5.733744,6.5312824,6.0258465,5.21518,4.6178465,4.1583595,3.1573336,1.9495386,1.0633847,0.508718,0.28225642,0.36758977,0.4660513,0.5513847,0.7089231,0.8795898,0.8402052,1.273436,2.028308,2.609231,2.9407182,3.3575387,3.4756925,3.3608208,3.511795,4.007385,4.5062566,4.535795,4.197744,4.069744,4.5128207,5.691077,6.0849237,6.2129235,5.277539,3.5807183,2.5074873,1.972513,1.654154,1.4309745,1.2635899,1.1979488,1.2931283,1.4375386,1.6246156,1.8149745,1.9364104,1.8674873,1.8248206,1.8806155,2.1267693,2.6322052,3.121231,3.4100516,3.629949,3.9187696,4.4045134,5.533539,6.8266673,8.116513,9.245539,10.089026,11.011283,12.2617445,13.24636,13.6008215,13.170873,12.347078,11.769437,11.798975,12.265027,12.458668,10.683078,8.2215395,5.83877,3.9876926,2.7700515,2.2711797,1.9856411,1.8379488,1.7263591,1.5425643,1.3226668,1.0535386,0.9517949,1.0666667,1.2504616,0.9189744,0.6170257,0.50543594,0.62030774,0.88287187,1.6114873,3.170462,5.280821,7.0859494,7.145026,4.926359,3.0096412,1.8445129,1.394872,1.1323078,0.8763078,0.6662565,0.52512825,0.47261542,0.49887183,0.7450257,1.1290257,1.4080001,1.3981539,0.97805136,0.60061544,0.35774362,0.19364104,0.07876924,0.016410258,0.026256412,0.16082053,0.41025645,0.6892308,0.8369231,0.5481026,0.2855385,0.108307704,0.02297436,0.0,0.009846155,0.049230773,0.08861539,0.10502565,0.101743594,0.19692309,0.37415388,0.6268718,0.93866676,1.270154,1.5721027,1.7952822,1.975795,2.1464617,2.3401027,2.4713848,2.5600002,2.6847181,2.878359,3.1442053,3.4888208,3.820308,4.056616,4.1550775,4.089436,3.9975388,4.023795,4.279795,4.7425647,5.2676926,5.7435904,5.8256416,5.5204105,4.965744,4.4406157,4.352,4.670359,5.280821,6.0980515,7.059693,5.139693,5.0642056,5.0543594,5.1889234,5.408821,5.4974365,5.546667,5.3760004,5.3891287,5.979898,7.515898,7.8112826,7.4108725,6.6560006,5.7632823,4.8147697,5.028103,5.3825645,5.7435904,6.124308,6.665847,6.7249236,6.7216415,7.204103,8.080411,8.615385,7.6077952,7.00718,7.171283,8.1755905,9.787078,10.522257,9.796924,8.963283,8.582564,8.421744,7.00718,5.4547696,4.204308,3.4133337,2.9505644,2.422154,2.1989746,2.1956925,2.3171284,2.4484105,3.4592824,4.7425647,6.0258465,7.00718,7.3714876,7.24677,7.77518,8.421744,8.910769,9.245539,9.403078,9.521232,9.905231,10.594462,11.372309,12.09436,13.190565,14.500104,16.059078,18.12677,20.54236,23.000618,24.871386,25.767387,25.550772,22.308104,19.078566,16.30195,14.536206,14.460719,13.965129,12.2847185,10.919386,10.640411,11.503591,14.742975,16.341335,16.187078,14.946463,14.080001,13.689437,13.755078,13.696001,13.2562065,12.4685135,11.59877,10.601027,9.554052,8.536616,7.637334,6.7314878,5.9634876,5.5565133,5.5762057,5.907693,6.163693,6.226052,6.045539,5.586052,4.821334,3.498667,2.605949,2.1398976,2.1103592,2.556718,3.18359,3.6627696,3.882667,3.9154875,4.0402055,4.076308,5.32677,7.0432825,8.04759,6.7314878,5.7665644,5.5565133,5.467898,5.2611284,5.0871797,5.0838976,5.346462,5.8945646,6.2752824,5.5729237,5.080616,4.568616,3.9384618,3.170462,2.3302567,2.3171284,2.1136413,1.8084104,1.6049232,1.8281027,2.162872,2.7011285,3.2000003,3.5905645,3.9680004,4.3716927,4.493129,4.2371287,3.7251284,3.2886157,2.868513,2.9472823,3.0358977,2.8553848,2.3204105,2.2449234,2.2055387,1.9626669,1.5097437,1.0732309,0.65312827,0.45620516,0.35446155,0.27897438,0.20676924,0.13784617,0.08533334,0.049230773,0.029538464,0.029538464,0.006564103,0.0,0.013128206,0.029538464,0.0,0.0,0.0032820515,0.0032820515,0.0,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.03938462,0.08861539,0.118153855,0.108307704,0.14769232,0.2231795,0.2100513,0.13784617,0.17394873,0.18051283,0.17723078,0.10502565,0.036102567,0.18379489,0.21661541,0.19692309,0.2100513,0.25928208,0.26912823,0.09189744,0.04594872,0.026256412,0.0,0.0,0.006564103,0.009846155,0.009846155,0.009846155,0.009846155,0.0032820515,0.0,0.0,0.0032820515,0.009846155,0.016410258,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.006564103,0.006564103,0.006564103,0.013128206,0.006564103,0.0032820515,0.009846155,0.016410258,0.026256412,0.026256412,0.026256412,0.02297436,0.02297436,0.02297436,0.01969231,0.01969231,0.02297436,0.02297436,0.052512825,0.07548718,0.0951795,0.118153855,0.14769232,0.17723078,0.16082053,0.17066668,0.23958977,0.35446155,0.64000005,0.8598975,0.83035904,0.60061544,0.47589746,0.43323082,0.32164106,0.27241027,0.33805132,0.48574364,0.44307697,0.4266667,0.5513847,0.78769237,0.98133343,1.0601027,1.0535386,0.9878975,0.88615394,0.76800007,0.8598975,1.083077,1.1323078,0.95835906,0.7581539,0.77128214,0.90256417,1.079795,1.3226668,1.7460514,2.612513,4.1124105,6.048821,8.090257,9.777231,10.450052,10.886565,10.988309,10.656821,9.80677,8.536616,6.921847,5.1298466,3.3509746,1.8051283,1.1060513,0.79425645,0.6465641,0.56123084,0.5349744,0.5940513,0.6432821,0.69251287,0.77456415,0.9353847,1.270154,1.6968206,2.172718,2.7142565,3.383795,3.754667,3.754667,3.515077,3.1245131,2.6354873,2.3696413,2.2153847,2.028308,1.8149745,1.7427694,1.8609232,2.1333334,2.4549747,2.9046156,3.7448208,3.4330258,2.6715899,2.0086155,1.6738462,1.5885129,1.723077,1.3259488,0.7384616,0.28225642,0.23958977,0.19364104,0.14441027,0.13456412,0.17066668,0.22646156,0.24615386,0.23630771,0.2297436,0.25928208,0.35774362,0.5021539,0.6170257,0.63343596,0.5546667,0.43651286,0.35446155,0.34133336,0.38728207,0.48246157,0.5973334,0.57764107,0.5021539,0.43651286,0.4135385,0.41682056,0.41682056,0.4135385,0.39056414,0.3446154,0.2986667,0.27569234,0.24287182,0.21989745,0.21333335,0.20348719,0.7844103,1.8871796,2.858667,3.2262566,2.7011285,1.6836925,1.1782565,0.92225647,0.8008206,0.8172308,0.8041026,0.7056411,0.636718,0.62030774,0.5874872,0.5677949,0.72861546,0.9419488,1.079795,1.020718,0.8960001,0.8336411,0.827077,0.9288206,1.2340513,2.0873847,2.9440002,3.4658465,3.4691284,2.8980515,2.861949,3.501949,4.342154,4.9788723,5.093744,4.7655387,4.460308,4.1682053,4.2338467,5.3792825,5.4941545,4.7261543,4.020513,3.5282054,2.605949,1.6049232,0.8336411,0.38400003,0.23302566,0.26584616,0.32164106,0.380718,0.48574364,0.58092314,0.5152821,0.6268718,1.014154,1.4933335,1.9298463,2.2580514,2.4549747,2.6354873,3.0687182,3.629949,3.7874875,3.6102567,3.495385,3.4133337,3.4198978,3.6758976,4.056616,4.3552823,4.210872,3.7087183,3.387077,3.5216413,3.570872,3.1934361,2.4582565,1.8379488,1.5819489,1.4736412,1.4834872,1.522872,1.4473847,1.2832822,1.2242053,1.3029745,1.5458462,1.9561027,2.1431797,2.2482052,2.3630772,2.5764105,2.9768207,3.9680004,5.6418467,7.273026,8.516924,9.3768215,10.453334,11.67754,12.645744,13.010053,12.458668,11.264001,10.197334,9.416205,8.966565,8.753231,7.7357955,6.3540516,4.9394875,3.7087183,2.7536411,2.1431797,1.7591796,1.4900514,1.270154,1.083077,1.0108719,0.955077,1.0108719,1.1979488,1.463795,1.5983591,1.3784616,1.0601027,0.8336411,0.8172308,1.3620514,2.6912823,4.3552823,5.8518977,6.629744,5.76,4.709744,3.4724104,2.2777438,1.6016412,1.339077,1.3686155,1.463795,1.4867693,1.3784616,1.1454359,1.0962052,1.0994873,1.0010257,0.6432821,0.4201026,0.27569234,0.16738462,0.07548718,0.016410258,0.016410258,0.12471796,0.38728207,0.71548724,0.8795898,0.65969235,0.40369233,0.190359,0.06564103,0.01969231,0.06564103,0.12471796,0.14441027,0.12471796,0.09189744,0.13456412,0.25271797,0.43323082,0.67282057,0.97805136,1.2438976,1.4769232,1.6738462,1.8609232,2.0841026,2.3138463,2.4648206,2.5862565,2.733949,2.9702566,3.31159,3.698872,4.0533338,4.315898,4.4340515,4.3585644,4.3290257,4.4274874,4.6966157,5.142975,5.5532312,5.737026,5.602462,5.218462,4.7917953,4.699898,4.886975,5.3070774,5.9963083,7.072821,4.571898,4.667077,4.670359,4.788513,5.093744,5.5138464,5.937231,5.861744,5.687795,5.904411,7.076103,6.99077,6.298257,5.362872,4.4996924,3.9614363,4.066462,4.342154,4.6834874,5.10359,5.723898,5.933949,5.720616,6.2588725,7.506052,8.182155,7.200821,6.6002054,6.5050263,7.072821,8.500513,9.081436,8.513641,8.008205,8.011488,8.2215395,7.3780518,5.920821,4.5062566,3.6036925,3.511795,3.1967182,2.861949,2.737231,2.9210258,3.373949,4.7655387,6.49518,8.27077,9.636104,9.980719,10.112,11.067078,12.107488,12.855796,13.298873,13.4170265,13.46954,13.617231,13.850258,14.011078,14.290052,15.2155905,16.666258,18.491077,20.512821,22.340925,23.968822,24.868105,24.822155,23.906464,21.572926,19.429745,17.109335,15.00554,14.263796,12.987078,11.464206,10.9226675,11.825232,13.892924,18.51077,20.834463,21.024822,19.403488,16.449642,14.677335,13.778052,13.315283,13.000206,12.701539,12.143591,11.286975,10.200616,8.973129,7.748924,6.160411,4.5554876,3.8498464,4.1878977,4.9427695,5.533539,6.3868723,6.9809237,6.9349747,5.9995904,4.594872,2.878359,1.5360001,0.9189744,1.0732309,1.7887181,2.7076926,3.383795,3.9351797,5.0609236,6.3343596,8.083693,10.013539,11.349334,10.807796,9.458873,8.178872,6.738052,5.353026,4.70318,5.402257,5.4843082,5.3234878,4.9394875,3.9909747,3.186872,2.7044106,2.3860514,2.176,2.1300514,2.612513,2.6157951,2.300718,2.0151796,2.2744617,2.6289232,3.0851285,3.442872,3.626667,3.7054362,3.8071797,3.751385,3.4691284,3.0293336,2.6486156,2.3105643,2.1825643,2.2055387,2.3171284,2.4582565,2.665026,2.6551797,2.2153847,1.4703591,0.892718,0.38400003,0.19364104,0.1148718,0.072205134,0.108307704,0.0951795,0.059076928,0.02297436,0.0,0.0,0.0,0.0,0.013128206,0.029538464,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.08205129,0.16410258,0.22646156,0.24615386,0.2100513,0.3511795,0.6465641,1.0010257,1.3357949,1.6082052,1.394872,1.1290257,0.761436,0.380718,0.19364104,0.098461546,0.101743594,0.13784617,0.17066668,0.19364104,0.14769232,0.08861539,0.03938462,0.013128206,0.013128206,0.013128206,0.013128206,0.009846155,0.009846155,0.009846155,0.0032820515,0.0032820515,0.006564103,0.006564103,0.016410258,0.026256412,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.0032820515,0.0032820515,0.009846155,0.016410258,0.029538464,0.04594872,0.04594872,0.036102567,0.016410258,0.026256412,0.029538464,0.03938462,0.06564103,0.1148718,0.14769232,0.14441027,0.15425642,0.19692309,0.256,0.26584616,0.2297436,0.190359,0.21333335,0.3708718,0.702359,0.9517949,0.9124103,0.6235898,0.3708718,0.36102566,0.3117949,0.27241027,0.28882053,0.4004103,0.42338464,0.47261542,0.6498462,0.9189744,1.1355898,1.3883078,1.5688206,1.4473847,1.0699488,0.7581539,0.827077,1.0108719,1.0568206,1.0404103,1.3357949,1.7657437,2.2153847,2.5304618,2.7864618,3.2820516,4.604718,6.442667,8.379078,10.04636,11.139283,11.208206,10.994873,10.509129,9.737847,8.621949,7.1876926,5.5696416,3.9876926,2.605949,1.522872,1.1126155,0.892718,0.8598975,0.9911796,1.2176411,1.0108719,0.8730257,0.892718,1.1520001,1.7132308,2.4188719,2.6880002,2.7175386,2.6190772,2.425436,3.308308,4.07959,4.089436,3.4002054,2.7963078,2.9505644,2.6026669,2.0676925,1.5753847,1.2668719,1.3456411,1.7493335,1.7952822,1.5655385,1.913436,1.7296412,1.3522053,1.1848207,1.2570257,1.204513,1.4145643,1.204513,0.75487185,0.3117949,0.19692309,0.18051283,0.15753847,0.13784617,0.14441027,0.19692309,0.24943592,0.318359,0.36430773,0.38728207,0.43651286,0.4955898,0.5349744,0.508718,0.41682056,0.31507695,0.27897438,0.2855385,0.30851284,0.33805132,0.3708718,0.41682056,0.44964105,0.47589746,0.48246157,0.45620516,0.40369233,0.40697438,0.4004103,0.3511795,0.256,0.2231795,0.21333335,0.2231795,0.23958977,0.23958977,0.76800007,1.8838975,2.930872,3.31159,2.487795,1.339077,0.8533334,0.6826667,0.6301539,0.65312827,0.71548724,0.7515898,0.83035904,0.90584624,0.81066674,0.65312827,0.64000005,0.7450257,0.88615394,0.9288206,0.8992821,0.92553854,0.9911796,1.1684103,1.6114873,2.3630772,2.740513,2.9407182,2.9768207,2.6617439,2.868513,3.564308,4.2272825,4.568616,4.5029745,3.9975388,3.370667,2.8356924,2.6486156,3.114667,3.6791797,3.7743592,3.6594875,3.367385,2.678154,1.5130258,0.7450257,0.35774362,0.24943592,0.24615386,0.256,0.27569234,0.3052308,0.3249231,0.30851284,0.3314872,0.48246157,0.8336411,1.273436,1.5327181,1.7657437,1.9922053,2.3794873,2.8389745,3.0293336,3.0490258,3.2065644,3.1507695,2.858667,2.6223593,3.0030773,3.6726158,4.2502565,4.4438977,4.0467696,4.394667,4.6244106,4.4964104,4.1025643,3.889231,4.0500517,3.817026,3.3903592,2.7864618,1.8379488,1.3029745,1.0666667,1.0502565,1.1716924,1.3522053,1.3193847,1.339077,1.4145643,1.5688206,1.8281027,2.4057438,3.620103,4.8738465,5.917539,6.8332314,8.392206,9.4457445,9.898667,9.796924,9.314463,8.490667,7.781744,7.056411,6.3310776,5.756718,5.2709746,4.844308,4.4045134,3.9023592,3.3247182,2.6978464,2.0808206,1.5556924,1.1716924,0.9485129,0.9878975,1.0601027,1.0732309,1.079795,1.2570257,1.6804104,1.6836925,1.4506668,1.1355898,0.8730257,1.0994873,1.8182565,2.7995899,3.8432825,4.778667,5.3169236,5.72718,5.5532312,4.5817437,2.8717952,1.9823592,1.8740515,2.156308,2.484513,2.556718,2.0184617,1.6410258,1.3554872,1.0601027,0.60061544,0.32820517,0.19692309,0.118153855,0.055794876,0.016410258,0.009846155,0.101743594,0.34789747,0.6892308,0.94523084,0.9714873,0.7318975,0.44307697,0.2231795,0.098461546,0.098461546,0.1148718,0.11158975,0.09189744,0.072205134,0.09189744,0.16738462,0.2855385,0.45292312,0.6892308,0.92553854,1.1585642,1.3751796,1.585231,1.8149745,2.0709746,2.2350771,2.3302567,2.4188719,2.5796926,2.868513,3.245949,3.6857438,4.135385,4.519385,4.647385,4.709744,4.7228723,4.7524104,4.893539,5.0477953,5.2414365,5.366154,5.398975,5.402257,5.3202057,5.3169236,5.435077,5.8256416,6.7249236,4.027077,4.0500517,4.2240005,4.5522056,4.9526157,5.2742567,5.543385,5.7698464,5.677949,5.297231,4.97559,4.568616,4.3290257,4.1189747,3.9023592,3.7415388,3.629949,3.8367183,4.0533338,4.1780515,4.325744,4.5062566,5.0182567,6.2129235,7.568411,7.686565,6.774154,5.796103,5.21518,5.2348723,5.8157954,6.4557953,6.921847,7.243488,7.4863596,7.765334,8.224821,7.3616414,6.157129,5.3858466,5.5893335,5.362872,4.97559,4.821334,5.044513,5.5269747,6.626462,8.470975,10.597744,12.442257,13.321847,14.381949,15.668514,16.715488,17.355488,17.742771,17.792002,17.831387,17.686975,17.253744,16.502155,16.111591,16.269129,17.234053,18.947283,20.998566,22.531284,23.312412,23.19754,22.216208,20.578463,18.491077,17.634462,17.10277,16.36431,15.254975,13.682873,12.360206,12.274873,13.620514,15.812924,19.078566,20.955898,21.507284,20.178053,15.786668,13.515489,12.071385,11.378873,11.188514,11.076924,11.057232,10.758565,10.148104,9.235693,8.054154,6.180103,3.8531284,2.7306669,3.0326157,3.5544617,3.4592824,3.9220517,4.8804107,5.648411,4.9394875,3.8334363,2.103795,0.7975385,0.30851284,0.4004103,0.88615394,1.394872,1.9954873,3.0490258,5.225026,8.011488,9.701744,10.774975,11.595488,12.389745,11.208206,9.728001,8.0377445,6.5772314,6.12759,6.8562055,6.5050263,5.8092313,5.228308,4.97559,4.5423594,4.020513,3.5314875,3.2229745,3.2722054,4.0402055,3.7842054,3.1540515,2.665026,2.7208207,2.917744,3.1376412,3.186872,3.0358977,2.8160002,2.481231,2.2350771,2.028308,1.8346668,1.6508719,1.3850257,1.0502565,1.014154,1.3883078,2.034872,2.3958976,2.4155898,1.910154,1.0896411,0.5481026,0.16410258,0.06235898,0.052512825,0.029538464,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.21989745,0.35774362,0.45620516,0.6859488,1.3456411,1.9561027,2.3335385,2.7011285,3.0916924,3.3280003,2.7208207,2.0775387,1.4473847,0.88615394,0.48246157,0.23302566,0.22646156,0.29538465,0.35774362,0.41025645,0.24287182,0.10502565,0.03938462,0.03938462,0.032820515,0.016410258,0.006564103,0.0032820515,0.0,0.0032820515,0.0,0.006564103,0.013128206,0.013128206,0.013128206,0.02297436,0.016410258,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.006564103,0.016410258,0.04594872,0.07548718,0.08205129,0.06235898,0.026256412,0.036102567,0.04266667,0.072205134,0.13128206,0.23630771,0.24615386,0.18707694,0.17066668,0.22646156,0.29538465,0.256,0.2100513,0.16082053,0.17394873,0.36102566,0.5874872,0.7122052,0.6892308,0.51856416,0.27241027,0.27897438,0.2855385,0.27241027,0.25928208,0.28882053,0.380718,0.56123084,0.78769237,1.0436924,1.3554872,1.9396925,2.3138463,2.103795,1.4539489,1.017436,0.9714873,0.90912825,1.0108719,1.4703591,2.4648206,3.2229745,3.9286156,4.4800005,4.9920006,5.805949,7.1581545,8.385642,9.419488,10.134975,10.374565,10.358154,9.921641,9.186462,8.182155,6.8529234,5.3858466,4.017231,2.7995899,1.8510771,1.3489232,1.086359,1.024,1.2077949,1.6311796,2.2416413,1.8806155,1.3751796,1.204513,1.6311796,2.733949,3.7842054,3.7874875,3.1770258,2.3893335,1.8576412,3.4855387,4.388103,4.132103,3.2328207,3.1638978,3.9614363,3.4002054,2.3991797,1.5885129,1.3128207,1.719795,2.5665643,2.4484105,1.3226668,0.49887183,0.43651286,0.62030774,0.9353847,1.211077,1.2012309,1.1257436,0.9878975,0.8172308,0.6301539,0.4201026,0.4201026,0.40697438,0.35774362,0.29538465,0.30194873,0.39384618,0.512,0.5677949,0.5284103,0.40369233,0.2986667,0.2297436,0.190359,0.16738462,0.17066668,0.19692309,0.2297436,0.256,0.26584616,0.2855385,0.38728207,0.5874872,0.764718,0.8205129,0.67938465,0.512,0.4397949,0.42338464,0.39712822,0.27897438,0.22646156,0.23302566,0.26912823,0.29538465,0.28225642,0.22646156,0.65641034,1.2964103,1.6344616,0.9353847,0.54482055,0.4135385,0.36102566,0.32164106,0.33476925,0.54482055,0.764718,0.98461545,1.142154,1.1027694,0.9517949,0.8041026,0.7417436,0.78769237,0.90584624,0.9616411,1.083077,1.2307693,1.4933335,2.1103592,3.006359,3.3608208,3.383795,3.170462,2.7175386,3.0424619,3.6660516,4.2436924,4.588308,4.673641,4.2994876,3.4133337,2.5074873,1.8576412,1.4998976,1.8543591,2.6256413,3.190154,3.239385,2.7798977,1.4506668,0.73517954,0.4135385,0.30194873,0.26912823,0.23958977,0.21661541,0.21989745,0.24943592,0.28225642,0.29210258,0.41025645,0.62030774,0.82379496,0.85005134,0.88943595,0.83035904,0.8533334,1.0436924,1.3817437,1.8740515,2.28759,2.5829747,2.868513,3.373949,3.9712822,4.827898,5.287385,4.965744,3.751385,3.7087183,3.7382567,3.9286156,4.338872,5.0018463,5.8912826,5.832206,5.182359,4.06318,2.3696413,1.5688206,1.1716924,1.0108719,0.97805136,1.020718,1.0896411,1.2373334,1.4080001,1.5688206,1.719795,1.782154,1.8510771,2.162872,2.7864618,3.629949,5.428513,6.0750775,5.756718,5.037949,4.8705645,4.9493337,5.2545643,5.395693,5.2315903,4.84759,4.644103,4.450462,4.263385,4.0369234,3.6890259,3.2065644,2.4746668,1.7887181,1.2964103,0.9944616,1.0305642,1.086359,0.9911796,0.8566154,1.079795,1.585231,1.7591796,1.7788719,1.7132308,1.5031796,1.4703591,1.4966155,1.7591796,2.3401027,3.2229745,4.6244106,6.1374364,7.397744,7.466667,4.84759,3.062154,2.3040001,2.5042052,3.242667,3.751385,3.190154,2.5731285,1.9265642,1.2865642,0.69251287,0.30194873,0.14441027,0.07876924,0.036102567,0.016410258,0.006564103,0.068923086,0.24615386,0.5513847,0.97805136,1.3653334,1.2274873,0.90256417,0.574359,0.26912823,0.12143591,0.04594872,0.02297436,0.032820515,0.04266667,0.068923086,0.128,0.2231795,0.35774362,0.53825647,0.77128214,1.0404103,1.3095386,1.5655385,1.8051283,1.9954873,2.1169233,2.1792822,2.1956925,2.2088206,2.359795,2.6486156,3.0916924,3.6529233,4.2338467,4.6539493,4.9329233,5.0543594,5.0215387,4.8640003,4.7556925,4.857436,5.1265645,5.5236926,6.0192823,5.9503593,5.8157954,5.684513,5.720616,6.186667,3.3575387,3.3214362,3.4198978,3.8596926,4.637539,5.5532312,6.114462,5.9634876,5.1331286,4.069744,3.6332312,3.5577438,4.0992823,4.634257,4.890257,4.9132314,4.5456414,4.023795,3.3969233,3.0194874,3.5544617,4.667077,5.034667,5.3398976,5.940513,6.882462,6.124308,4.8640003,3.9975388,3.8629746,4.2436924,5.4875903,6.3376417,6.8627696,7.0104623,6.6067696,6.5083084,6.6034875,6.5017443,6.163693,5.920821,6.2490263,6.7610264,7.456821,8.274052,9.078155,10.19077,11.858052,13.610668,15.212309,16.676104,17.591797,18.500925,19.331284,19.91549,19.987694,19.794052,20.066463,20.004105,19.111385,17.19795,16.036104,15.2155905,15.412514,16.544823,17.77559,19.094976,19.728413,20.027079,20.322464,20.919796,20.345438,19.075283,18.080822,17.673847,17.503181,17.795284,18.06113,18.261335,18.048002,16.754873,15.986873,15.455181,14.772514,13.820719,12.770463,12.245335,11.621744,10.896411,10.246565,10.039796,10.026668,10.31877,10.112,8.969847,6.820103,4.3290257,2.1530259,1.3226668,1.785436,2.3958976,3.1277952,3.4133337,3.3378465,2.806154,1.5097437,0.9485129,0.69907695,0.6071795,0.69251287,1.1454359,2.4976413,3.314872,3.820308,4.1025643,4.089436,4.9821544,6.9152827,7.8014364,7.069539,5.677949,5.287385,5.674667,6.918565,8.54318,9.521232,10.180923,10.180923,9.764103,9.091283,8.224821,8.103385,7.8802056,7.4108725,6.9087186,6.957949,8.165744,6.820103,4.854154,3.4921029,3.2361028,3.5282054,3.948308,3.7120004,2.793026,1.9364104,1.2800001,0.9682052,0.86317956,0.9189744,1.1749744,1.1618463,0.8763078,0.62030774,0.49887183,0.4135385,0.44964105,0.5481026,0.71548724,0.8172308,0.6104616,0.39056414,0.13456412,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.26912823,0.53825647,0.78769237,1.8215386,5.2644105,6.997334,6.2030773,4.7261543,3.4527183,2.3040001,1.4506668,0.8795898,0.65312827,0.6301539,0.45620516,0.190359,0.10502565,0.08533334,0.07876924,0.09189744,0.09189744,0.08205129,0.08205129,0.08205129,0.04594872,0.009846155,0.009846155,0.009846155,0.0032820515,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.02297436,0.026256412,0.016410258,0.016410258,0.016410258,0.026256412,0.052512825,0.07548718,0.06564103,0.06235898,0.10502565,0.17394873,0.19692309,0.15097436,0.128,0.128,0.15097436,0.19692309,0.19692309,0.190359,0.21989745,0.3117949,0.45620516,0.71548724,0.761436,0.65641034,0.49230772,0.380718,0.32164106,0.3314872,0.3708718,0.4135385,0.47261542,0.6301539,0.8369231,1.086359,1.4408206,2.0151796,2.550154,2.5009232,2.15959,1.7001027,1.1749744,1.0535386,1.086359,1.5327181,2.3072822,2.989949,3.3575387,4.161641,5.182359,6.2720003,7.3714876,7.8703594,8.096821,7.8080006,7.177847,6.774154,7.030154,7.131898,7.1122055,6.5870776,4.7294364,3.1540515,2.0676925,1.4244103,1.1158975,0.94523084,1.2406155,1.4867693,1.6443079,1.8904617,2.609231,3.1343591,2.2678976,1.6443079,1.9790771,3.0523078,3.8071797,4.06318,3.1343591,1.8838975,2.7011285,5.47118,4.315898,2.1234872,0.6859488,0.6859488,1.1979488,1.7755898,2.0217438,1.847795,1.4966155,1.142154,0.9714873,0.8730257,0.7811283,0.67282057,0.6465641,0.6859488,0.7056411,0.67610264,0.64000005,0.7515898,0.9156924,1.1093334,1.2635899,1.2504616,1.2373334,1.2176411,1.1126155,0.9124103,0.65641034,0.58420515,0.51856416,0.46276927,0.40369233,0.3052308,0.21989745,0.18051283,0.16738462,0.17066668,0.18379489,0.20676924,0.21333335,0.21333335,0.22646156,0.27569234,0.33476925,0.827077,1.4244103,1.7427694,1.3259488,0.92553854,0.55794877,0.3511795,0.30194873,0.28882053,0.2297436,0.20348719,0.20348719,0.2100513,0.19692309,0.19692309,0.23630771,0.25928208,0.25271797,0.2297436,0.2297436,0.2297436,0.2100513,0.20020515,0.27569234,0.38400003,0.5218462,0.7056411,0.9419488,1.2373334,1.273436,1.2438976,1.1946667,1.1520001,1.1126155,1.0896411,1.3029745,1.5458462,1.6311796,1.3883078,1.7296412,2.3926156,2.6420515,2.353231,1.9987694,2.3401027,3.387077,4.8640003,6.186667,6.4557953,5.805949,4.2830772,2.9636924,2.2580514,1.8904617,1.463795,1.404718,1.7591796,2.1464617,1.7558975,1.0601027,0.6662565,0.446359,0.318359,0.24287182,0.24287182,0.24287182,0.26256412,0.28225642,0.24287182,0.14769232,0.15753847,0.20020515,0.23958977,0.28882053,0.33805132,0.2855385,0.35446155,0.5874872,0.86974365,1.0404103,1.0929232,1.0633847,1.0404103,1.1749744,1.1388719,0.9288206,0.78769237,0.8205129,0.9911796,1.6147693,1.8609232,1.8084104,1.6443079,1.6935385,1.8904617,2.3302567,2.5698464,2.409026,1.9068719,1.7001027,1.585231,1.5425643,1.6180514,1.9232821,2.3729234,2.7700515,3.1081028,3.3805132,3.6004105,3.0260515,2.1956925,1.8248206,2.0545642,2.4582565,3.249231,3.373949,3.1737437,3.0654361,3.5413337,4.027077,4.4800005,4.827898,5.044513,5.142975,4.70318,4.135385,3.43959,2.7634873,2.3958976,2.0775387,1.7985642,1.5458462,1.3128207,1.0666667,0.8598975,0.7450257,0.77456415,1.1060513,1.9823592,3.1442053,3.1507695,2.9111798,2.9440002,3.370667,3.3476925,3.1113849,2.5764105,2.1858463,2.930872,5.5893335,7.427283,8.5202055,8.582564,6.957949,5.175795,3.56759,3.318154,4.2994876,5.080616,4.4340515,3.3378465,1.8871796,0.571077,0.28882053,0.19364104,0.12143591,0.06564103,0.026256412,0.016410258,0.016410258,0.016410258,0.03938462,0.2100513,0.74830776,1.4080001,1.6443079,1.5589745,1.1946667,0.5481026,0.256,0.09189744,0.029538464,0.029538464,0.029538464,0.06564103,0.12143591,0.20676924,0.34133336,0.5481026,0.84348726,1.1979488,1.5458462,1.8510771,2.1202054,2.2908719,2.4155898,2.477949,2.428718,2.1956925,2.1103592,2.2186668,2.487795,2.878359,3.3411283,3.9384618,4.5095387,5.041231,5.4383593,5.5236926,5.474462,5.435077,5.533539,5.8223596,6.2851286,6.23918,6.052103,5.805949,5.648411,5.7829747,4.5423594,3.9286156,3.4592824,3.308308,3.501949,3.9318976,4.3651285,4.640821,4.706462,4.571898,4.325744,3.7284105,3.3214362,3.0293336,2.7864618,2.556718,2.2514873,1.9200002,1.7493335,2.100513,3.5052311,4.07959,4.007385,4.263385,5.077334,5.930667,5.835488,5.395693,4.8738465,4.460308,4.240411,4.4340515,4.926359,5.612308,6.3376417,6.9120007,6.738052,6.6002054,6.4754877,6.4754877,6.8365135,7.5454364,8.323282,9.061745,9.685334,10.128411,11.424822,13.029744,14.634667,15.90154,16.459488,16.006565,16.351181,17.05354,17.80513,18.41559,18.921026,19.400208,19.045746,17.78872,16.292105,15.31077,15.061335,15.616001,16.94195,18.888206,20.762259,21.986464,22.265438,21.67795,20.676924,20.23713,19.771078,19.767796,19.971283,19.370668,18.304,17.900309,17.591797,16.918976,15.547078,14.483693,13.768207,13.594257,13.63036,13.039591,11.234463,9.6984625,8.346257,7.450257,7.6242056,8.342975,9.6525135,9.878975,8.553026,6.3934364,3.9712822,2.4681027,1.9659488,2.028308,1.7132308,1.6836925,1.9659488,2.3335385,2.6223593,2.7569232,2.537026,2.3433847,2.166154,2.0709746,2.1825643,2.5600002,2.2219489,1.7132308,1.4342566,1.6344616,2.1858463,3.0523078,4.417641,5.8190775,6.1768208,4.8672824,4.46359,4.7294364,5.395693,6.12759,7.000616,8.0377445,9.101129,10.098872,10.971898,10.975181,10.587898,9.770667,8.572719,7.1154876,5.602462,4.269949,3.367385,3.0851285,3.5413337,3.3050258,2.92759,2.1924105,1.2537436,0.6432821,0.43323082,0.3511795,0.34133336,0.3511795,0.3446154,0.34133336,0.32820517,0.29210258,0.24615386,0.2297436,0.24615386,0.27569234,0.33805132,0.3708718,0.23302566,0.108307704,0.032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.06235898,0.17394873,0.5481026,1.1520001,2.0611284,3.4822567,4.1911798,3.6824617,2.809436,1.9954873,1.2176411,0.7450257,0.48246157,0.46933338,0.58092314,0.50543594,0.26584616,0.18051283,0.15425642,0.13128206,0.10502565,0.13456412,0.18379489,0.13456412,0.016410258,0.009846155,0.013128206,0.013128206,0.08205129,0.14769232,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.009846155,0.0032820515,0.0,0.0,0.0,0.009846155,0.013128206,0.02297436,0.029538464,0.026256412,0.016410258,0.016410258,0.016410258,0.026256412,0.03938462,0.036102567,0.04266667,0.06235898,0.08205129,0.08861539,0.118153855,0.14441027,0.15097436,0.14112821,0.15097436,0.14112821,0.14441027,0.16738462,0.21333335,0.26256412,0.41025645,0.4955898,0.4397949,0.29210258,0.2231795,0.26912823,0.380718,0.52512825,0.63343596,0.6071795,0.6892308,0.8795898,1.0962052,1.3062565,1.5392822,1.8609232,1.8740515,1.6804104,1.3883078,1.1257436,0.96492314,0.75487185,0.9944616,1.8313848,3.0523078,4.1517954,5.3792825,6.4065647,7.1614366,7.857231,8.379078,7.3780518,5.9536414,4.9394875,4.906667,4.919795,4.8114877,4.824616,4.8082056,4.240411,2.5796926,1.6672822,1.2898463,1.211077,1.1651284,1.4309745,1.8740515,2.5796926,3.56759,4.7950773,3.190154,1.8871796,1.3620514,1.8084104,3.1376412,4.342154,3.4330258,1.8904617,0.81066674,0.90584624,2.2711797,2.2416413,1.4178462,0.5415385,0.49230772,0.6432821,0.79097444,0.85005134,0.79097444,0.65312827,0.62030774,0.6629744,0.77456415,0.88287187,0.84348726,0.65312827,0.6268718,0.67938465,0.761436,0.8598975,0.8336411,0.8336411,1.014154,1.3259488,1.5064616,1.2800001,1.0896411,0.8960001,0.79425645,0.98461545,1.3620514,1.079795,0.6432821,0.33805132,0.23302566,0.2231795,0.21333335,0.19364104,0.18051283,0.18379489,0.19692309,0.24615386,0.2986667,0.32164106,0.26256412,0.31507695,0.4594872,0.574359,0.6104616,0.5940513,1.1093334,1.1651284,0.84348726,0.39384618,0.21661541,0.16410258,0.20348719,0.256,0.2855385,0.28225642,0.3708718,0.45292312,0.45292312,0.39384618,0.4004103,0.42994875,0.40697438,0.3511795,0.29538465,0.2986667,0.36102566,0.44964105,0.5284103,0.6268718,0.8205129,1.1520001,1.4539489,1.6771283,1.7427694,1.529436,1.339077,1.4211283,1.5163078,1.4900514,1.3653334,1.4802053,1.719795,1.9528207,2.0611284,1.9626669,2.1103592,2.5271797,3.117949,3.7054362,4.06318,4.1780515,3.9253337,3.387077,2.7602053,2.356513,2.0151796,1.7362052,1.5524104,1.4178462,1.1946667,0.90912825,0.6662565,0.56451285,0.58092314,0.5874872,0.380718,0.27897438,0.23958977,0.23302566,0.24287182,0.21333335,0.20020515,0.20020515,0.20348719,0.19364104,0.24943592,0.25928208,0.28225642,0.33805132,0.39384618,0.50543594,0.6170257,0.77128214,1.083077,1.7362052,2.2088206,2.100513,1.7624617,1.5064616,1.6377437,2.0086155,2.353231,2.5173335,2.5271797,2.5961027,2.7634873,2.9702566,3.190154,3.2196925,2.7011285,1.8084104,1.4933335,1.6278975,1.9396925,2.0217438,1.9823592,1.9429746,1.9823592,2.1497438,2.4648206,2.6453335,2.3236926,1.9823592,1.8313848,1.8346668,1.8281027,1.6771283,1.7755898,2.3171284,3.3214362,3.9351797,4.1780515,4.007385,3.495385,2.8225644,2.4024618,2.1989746,2.1136413,2.048,1.9068719,1.7558975,1.6180514,1.4802053,1.3259488,1.1290257,0.90256417,0.86317956,1.083077,1.5392822,2.1070771,2.4746668,2.5009232,2.6026669,3.0752823,4.128821,5.169231,5.799385,5.618872,4.699898,3.5872824,3.495385,4.066462,4.4767184,4.325744,3.636513,2.861949,2.477949,2.8521028,3.754667,4.3618464,3.6758976,2.546872,1.3357949,0.4135385,0.19364104,0.14441027,0.09189744,0.052512825,0.026256412,0.016410258,0.006564103,0.0032820515,0.016410258,0.08205129,0.24615386,0.61374366,0.98461545,1.1323078,0.9747693,0.56123084,0.26912823,0.10502565,0.032820515,0.01969231,0.029538464,0.06564103,0.128,0.23302566,0.39712822,0.6235898,0.96492314,1.3784616,1.7887181,2.1431797,2.4024618,2.5042052,2.5829747,2.5961027,2.5074873,2.294154,2.100513,2.041436,2.1070771,2.2744617,2.5238976,2.9078977,3.3575387,3.8662567,4.384821,4.841026,5.1922054,5.5597954,5.937231,6.298257,6.616616,6.4590774,6.0258465,5.605744,5.3891287,5.464616,4.8016415,4.138667,3.6332312,3.3280003,3.2262566,3.3050258,3.318154,3.3312824,3.4625645,3.639795,3.6036925,3.0851285,2.5238976,1.9954873,1.5589745,1.273436,1.0469744,0.8730257,0.9714873,1.5064616,2.5895386,3.2623591,3.515077,3.8071797,4.3060517,4.893539,5.1889234,5.477744,5.609026,5.5138464,5.211898,5.0871797,5.2742567,5.6418467,6.1407185,6.806975,7.282872,7.53559,7.716103,7.9852314,8.51036,9.009232,9.416205,9.8363085,10.305642,10.811078,11.897437,13.37436,15.051488,16.387283,16.512001,15.80636,15.340309,15.461744,16.213335,17.362053,18.556719,19.528206,19.777643,19.373951,18.934155,18.563284,18.198977,18.310566,19.2,20.995283,22.790565,24.329847,24.42831,23.184412,21.979898,21.714052,21.704206,21.927387,22.071796,21.54995,19.794052,17.322668,16.978052,19.094976,21.497438,23.151592,22.357334,18.60595,13.423591,10.371283,7.8080006,6.7544622,6.232616,5.8978467,6.048821,6.416411,7.138462,7.702975,7.860513,7.604513,7.059693,5.9930263,4.8738465,3.9318976,3.170462,2.8258464,2.865231,3.0162053,3.1376412,3.2229745,2.7602053,2.4188719,2.2088206,2.4582565,3.8137438,4.9362054,5.07077,5.464616,6.770872,9.042052,10.912822,12.76718,14.424617,15.100719,13.397334,9.353847,6.6034875,4.7294364,3.7120004,3.9056413,4.5489235,5.622154,6.7610264,7.6996927,8.280616,7.817847,7.003898,5.874872,4.6802053,3.889231,2.8258464,2.0841026,1.657436,1.5360001,1.7033848,1.6738462,1.4900514,1.086359,0.5907693,0.3117949,0.21333335,0.16738462,0.15097436,0.13784617,0.101743594,0.101743594,0.12143591,0.13456412,0.128,0.128,0.13456412,0.128,0.128,0.12143591,0.06564103,0.016410258,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.029538464,0.13456412,0.4004103,0.82379496,1.3292309,1.782154,2.0151796,1.7263591,1.3095386,0.955077,0.6432821,0.45620516,0.36758977,0.35774362,0.38400003,0.3708718,0.27241027,0.21333335,0.17066668,0.13456412,0.13456412,0.13456412,0.14112821,0.08533334,0.0,0.0,0.013128206,0.016410258,0.04594872,0.072205134,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0032820515,0.013128206,0.016410258,0.01969231,0.013128206,0.006564103,0.006564103,0.009846155,0.01969231,0.029538464,0.02297436,0.026256412,0.029538464,0.036102567,0.052512825,0.07876924,0.11158975,0.14112821,0.16410258,0.19364104,0.18707694,0.17394873,0.15753847,0.15425642,0.18707694,0.27241027,0.35774362,0.35774362,0.26912823,0.16410258,0.23958977,0.35774362,0.50543594,0.6498462,0.76800007,1.0272821,1.3883078,1.7526156,1.972513,1.847795,1.8018463,1.8379488,2.3040001,3.0162053,3.245949,1.7001027,0.94523084,1.1060513,1.9823592,3.058872,4.201026,5.5696416,6.7249236,7.565129,8.310155,8.461129,7.8703594,7.131898,6.6494365,6.636308,6.38359,5.4482055,4.59159,4.164923,4.1091285,2.7044106,1.529436,0.9911796,1.0305642,1.1191796,1.2307693,2.3368206,4.2469745,6.5739493,8.726975,8.736821,7.8506675,6.2916927,4.6276927,3.761231,3.820308,2.6190772,1.2274873,0.34133336,0.29210258,0.7187693,0.84348726,0.6629744,0.36758977,0.3511795,0.40369233,0.45620516,0.47589746,0.44964105,0.38728207,0.39384618,0.44307697,0.5415385,0.6498462,0.69251287,0.8566154,1.1355898,1.214359,1.0732309,0.9878975,0.96492314,0.9485129,0.9682052,1.0075898,1.014154,0.90912825,0.7778462,0.63343596,0.5513847,0.6662565,1.0962052,1.014154,0.6465641,0.26256412,0.15753847,0.17066668,0.18051283,0.18379489,0.18707694,0.20020515,0.20020515,0.21989745,0.23630771,0.22646156,0.18707694,0.23630771,0.27241027,0.26256412,0.22646156,0.24615386,0.53825647,0.5940513,0.46276927,0.27241027,0.23630771,0.24615386,0.27897438,0.2986667,0.2986667,0.3052308,0.38728207,0.47589746,0.50543594,0.4660513,0.40697438,0.39056414,0.36758977,0.33476925,0.29538465,0.26912823,0.30194873,0.40369233,0.49887183,0.58420515,0.7187693,0.95835906,1.204513,1.4375386,1.6311796,1.7329233,1.7887181,1.8116925,1.7690258,1.6869745,1.6771283,1.6968206,1.7296412,1.8346668,1.9856411,2.0808206,2.1924105,2.3663592,2.5271797,2.6683078,2.8488207,3.1474874,3.2951798,3.1343591,2.7011285,2.2350771,1.8642052,1.4998976,1.214359,1.0305642,0.90584624,0.78769237,0.702359,0.67610264,0.7089231,0.75487185,0.6432821,0.5021539,0.36758977,0.25928208,0.190359,0.16082053,0.16410258,0.17066668,0.16410258,0.13128206,0.14769232,0.15753847,0.16082053,0.16738462,0.17394873,0.24943592,0.33476925,0.446359,0.6268718,0.9616411,1.2668719,1.2800001,1.1224617,0.9485129,0.93866676,1.1585642,1.4834872,1.8084104,2.0742567,2.2744617,2.5271797,2.8553848,3.0030773,2.8192823,2.2580514,1.5622566,1.4703591,1.785436,2.169436,2.1366155,1.9790771,1.8281027,1.657436,1.4900514,1.4145643,1.4506668,1.5031796,1.6968206,2.0250258,2.3729234,2.2022567,1.8084104,1.7165129,1.9954873,2.2678976,2.349949,2.2449234,1.9790771,1.6311796,1.3357949,1.3095386,1.4375386,1.5491283,1.5688206,1.529436,1.4342566,1.3193847,1.211077,1.1126155,1.024,0.97805136,1.0338463,1.2176411,1.4966155,1.7887181,2.1366155,2.5698464,3.0162053,3.508513,4.1813335,4.7261543,5.093744,4.9854364,4.2994876,3.1113849,2.7044106,2.8717952,2.9833848,2.789744,2.4057438,2.172718,2.1530259,2.3696413,2.7470772,3.117949,2.612513,1.6738462,0.8172308,0.3117949,0.18707694,0.128,0.07548718,0.036102567,0.009846155,0.006564103,0.0,0.0,0.0032820515,0.02297436,0.06564103,0.21989745,0.5349744,0.80738467,0.892718,0.69251287,0.3708718,0.18051283,0.07876924,0.029538464,0.02297436,0.049230773,0.101743594,0.20348719,0.37743592,0.6235898,1.0043077,1.4506668,1.8707694,2.1989746,2.3893335,2.4681027,2.537026,2.5665643,2.5337439,2.428718,2.2908719,2.2646155,2.349949,2.5238976,2.7503593,2.917744,3.058872,3.2000003,3.3936412,3.7087183,4.204308,4.8049235,5.481026,6.170257,6.770872,6.806975,6.363898,5.7042055,5.146257,5.0477953,4.2502565,3.9220517,3.757949,3.5905645,3.387077,3.2328207,2.8947694,2.681436,2.6880002,2.8356924,2.858667,2.612513,2.231795,1.7526156,1.2603078,0.88287187,0.69907695,0.6498462,0.88615394,1.3981539,2.0217438,2.6978464,3.1573336,3.4494362,3.6791797,3.9844105,4.529231,5.277539,5.796103,5.924103,5.799385,5.733744,5.799385,5.973334,6.3573337,7.177847,8.188719,8.946873,9.524513,10.003693,10.499283,10.555078,10.584617,10.706052,11.044104,11.733335,12.786873,14.204719,15.78995,17.073233,17.348925,17.004309,16.406975,16.200207,16.633438,17.562258,18.740515,19.817028,20.548925,20.929642,21.202053,21.382566,21.31036,21.69436,22.803694,24.474258,24.960001,25.606565,25.429335,24.359386,23.2599,22.79713,23.450258,24.20513,24.480822,24.136208,21.710772,18.389336,18.760206,23.043283,27.057232,28.931284,26.164515,19.30831,11.336206,7.637334,5.4153852,4.7950773,4.630975,4.417641,4.2962055,4.9427695,5.481026,6.121026,6.8365135,7.3550773,7.712821,7.384616,6.6034875,5.658257,4.923077,4.519385,4.3060517,4.056616,3.7415388,3.5347695,3.2689233,3.9680004,5.077334,6.340924,7.8112826,8.713847,8.78277,9.127385,10.246565,12.009027,13.226667,14.368821,14.943181,14.572309,13.013334,10.171078,8.323282,6.633026,4.9329233,3.7218463,3.4658465,3.620103,3.9745643,4.276513,4.2272825,3.5938463,2.8816411,2.0676925,1.401436,1.3981539,1.2406155,1.0338463,0.827077,0.6432821,0.47589746,0.5021539,0.48902568,0.40369233,0.27569234,0.20676924,0.15425642,0.101743594,0.06564103,0.052512825,0.04594872,0.049230773,0.049230773,0.052512825,0.06235898,0.072205134,0.08205129,0.06235898,0.036102567,0.016410258,0.009846155,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.072205134,0.18051283,0.32820517,0.4955898,0.6301539,0.7384616,0.69579494,0.61374366,0.54482055,0.47917953,0.40369233,0.36102566,0.3052308,0.24615386,0.24287182,0.23630771,0.2100513,0.15425642,0.098461546,0.098461546,0.07876924,0.06564103,0.036102567,0.0032820515,0.0,0.006564103,0.009846155,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.006564103,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.006564103,0.0,0.009846155,0.016410258,0.013128206,0.006564103,0.0,0.0,0.009846155,0.032820515,0.06235898,0.03938462,0.026256412,0.02297436,0.032820515,0.052512825,0.059076928,0.0951795,0.14441027,0.190359,0.23630771,0.22646156,0.18379489,0.16738462,0.20348719,0.27897438,0.33805132,0.37415388,0.35446155,0.28225642,0.18379489,0.24615386,0.380718,0.51856416,0.64000005,0.76800007,1.1093334,1.5556924,2.162872,2.6354873,2.3302567,1.6049232,1.5097437,2.1103592,2.9669745,3.131077,1.8182565,1.529436,2.044718,2.9965131,3.8695388,4.699898,5.8157954,6.8627696,7.6767187,8.297027,8.3823595,8.218257,7.837539,7.2861543,6.636308,6.0750775,5.0576415,4.2601027,3.9844105,4.164923,3.4198978,2.1070771,1.1224617,0.81394875,0.9682052,1.2537436,2.422154,4.7261543,7.6603084,9.961026,10.262975,9.278359,7.2270775,4.8082056,3.1770258,2.5238976,1.6180514,0.7844103,0.25271797,0.18379489,0.19692309,0.2231795,0.25271797,0.28225642,0.30851284,0.34789747,0.35446155,0.33476925,0.30194873,0.27897438,0.28882053,0.32820517,0.38728207,0.45620516,0.5152821,0.76800007,1.0568206,1.1093334,0.92553854,0.7811283,0.7811283,0.7975385,0.7778462,0.7220513,0.65969235,0.5874872,0.5021539,0.42338464,0.37415388,0.36758977,0.60061544,0.61374366,0.4201026,0.16410258,0.108307704,0.118153855,0.12471796,0.13784617,0.15097436,0.16410258,0.15753847,0.16082053,0.15425642,0.14769232,0.15425642,0.18379489,0.190359,0.18379489,0.17066668,0.16082053,0.16082053,0.14112821,0.12471796,0.128,0.18051283,0.21989745,0.26256412,0.2855385,0.29210258,0.32820517,0.3708718,0.41682056,0.45292312,0.45292312,0.380718,0.3117949,0.32820517,0.36430773,0.380718,0.34789747,0.3708718,0.46276927,0.5316923,0.56451285,0.6301539,0.8336411,1.0043077,1.1388719,1.276718,1.4966155,1.6902566,1.7657437,1.7690258,1.7723079,1.8609232,1.972513,2.1267693,2.3269746,2.5238976,2.5928206,2.5304618,2.5009232,2.4320002,2.3401027,2.3204105,2.3696413,2.3466668,2.3236926,2.2777438,2.0939488,1.8182565,1.467077,1.1093334,0.8205129,0.7122052,0.65312827,0.67938465,0.7384616,0.81394875,0.92553854,0.8598975,0.69579494,0.5021539,0.32164106,0.18379489,0.15097436,0.14441027,0.14769232,0.16410258,0.2100513,0.19692309,0.15753847,0.12471796,0.108307704,0.108307704,0.14769232,0.20348719,0.26584616,0.3117949,0.32164106,0.37743592,0.4266667,0.446359,0.4397949,0.4397949,0.6629744,0.9321026,1.2635899,1.5786668,1.723077,1.7591796,1.9528207,1.975795,1.7132308,1.2570257,1.014154,1.1454359,1.6410258,2.2350771,2.4057438,2.1924105,1.9692309,1.657436,1.270154,0.9321026,0.8598975,1.2570257,1.8773335,2.5206156,3.0391798,2.9505644,2.6847181,2.5665643,2.4943593,1.9265642,1.3292309,1.017436,0.8041026,0.6498462,0.6465641,0.8041026,0.9944616,1.086359,1.079795,1.1027694,1.1388719,1.0929232,1.020718,0.95835906,0.9288206,0.98133343,1.0896411,1.1979488,1.2931283,1.404718,1.9364104,2.6978464,3.4592824,4.0041027,4.1452312,3.9318976,3.9745643,3.9745643,3.6890259,2.9243078,2.6420515,2.5238976,2.412308,2.2153847,1.9298463,1.7362052,1.7329233,1.8215386,1.9396925,2.0512822,1.7099489,1.0666667,0.5481026,0.3117949,0.2297436,0.15097436,0.08861539,0.03938462,0.009846155,0.006564103,0.0,0.0,0.0,0.0032820515,0.01969231,0.055794876,0.2297436,0.49887183,0.73517954,0.7417436,0.51856416,0.36430773,0.24615386,0.14441027,0.059076928,0.04266667,0.06235898,0.13128206,0.26912823,0.47589746,0.85005134,1.270154,1.6771283,1.9889232,2.1136413,2.2088206,2.3368206,2.4615386,2.553436,2.5993848,2.5731285,2.6322052,2.8225644,3.117949,3.4133337,3.5478978,3.4625645,3.2722054,3.0949745,3.0785644,3.4297438,3.9548721,4.640821,5.431795,6.2030773,6.5969234,6.4295387,5.8486156,5.1659493,4.850872,3.511795,3.5905645,3.7448208,3.7218463,3.498667,3.2886157,2.8882053,2.678154,2.6256413,2.6518977,2.6453335,2.5632823,2.3696413,2.048,1.6213335,1.1520001,0.9419488,1.1618463,1.6114873,2.0808206,2.3630772,2.6978464,2.9604106,3.1540515,3.2984617,3.4166157,4.0992823,4.8836927,5.3136415,5.3727183,5.4875903,5.586052,5.681231,5.9930263,6.7183595,8.0377445,9.31118,10.427077,11.172104,11.556104,11.815386,11.483898,11.260718,11.191795,11.477334,12.501334,14.122667,16.009848,17.572104,18.602669,19.30831,19.426462,19.268925,19.042463,18.81272,18.514053,18.68472,19.272207,20.004105,20.70318,21.284103,21.861746,22.596926,23.890053,25.685335,27.480618,26.896412,26.177643,25.603285,24.986258,23.670156,22.882463,24.12636,25.38995,25.728003,25.281643,22.534565,20.030361,20.719591,24.106668,26.25313,25.75426,20.844309,14.145642,8.372514,6.304821,4.9887185,4.1780515,3.511795,2.9046156,2.546872,3.8728209,4.818052,5.3136415,5.428513,5.3924108,5.4416413,6.0356927,6.567385,6.7282057,6.518154,6.3376417,6.173539,5.868308,5.435077,5.0642056,5.100308,6.6822567,8.841846,10.535385,10.650257,10.246565,9.567181,8.887795,8.241231,7.4174366,6.3442054,5.5729237,4.8836927,4.6080003,5.661539,6.8463597,8.090257,8.260923,6.9120007,4.2994876,3.1015387,2.1891284,1.7033848,1.529436,1.3029745,0.9944616,0.8533334,0.761436,0.7122052,0.8041026,0.8336411,0.8336411,0.7581539,0.61374366,0.45620516,0.27241027,0.15753847,0.101743594,0.08205129,0.06235898,0.072205134,0.04594872,0.03938462,0.055794876,0.036102567,0.04266667,0.032820515,0.029538464,0.03938462,0.055794876,0.072205134,0.052512825,0.02297436,0.006564103,0.0032820515,0.0032820515,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.036102567,0.13784617,0.256,0.40369233,0.50543594,0.5415385,0.5152821,0.43651286,0.38728207,0.3314872,0.27241027,0.24615386,0.25271797,0.23630771,0.16410258,0.06564103,0.026256412,0.009846155,0.02297436,0.026256412,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.0032820515,0.0032820515,0.006564103,0.006564103,0.0032820515,0.016410258,0.01969231,0.013128206,0.0032820515,0.0,0.0,0.0,0.0,0.0032820515,0.013128206,0.0032820515,0.009846155,0.016410258,0.02297436,0.02297436,0.006564103,0.0032820515,0.016410258,0.049230773,0.08861539,0.06235898,0.04594872,0.052512825,0.08205129,0.108307704,0.08205129,0.098461546,0.13784617,0.17723078,0.21989745,0.21989745,0.17723078,0.19692309,0.30194873,0.4201026,0.4660513,0.43323082,0.3446154,0.23958977,0.18707694,0.2297436,0.38400003,0.53825647,0.61374366,0.574359,0.77456415,1.0962052,1.785436,2.5107694,2.3762052,1.3029745,1.086359,1.148718,1.1027694,0.74830776,1.0469744,1.8970258,2.9669745,4.017231,4.916513,5.402257,5.9930263,6.678975,7.3353853,7.7292314,8.123077,7.768616,6.738052,5.3136415,3.9975388,3.3247182,3.117949,3.367385,3.882667,4.269949,4.076308,2.92759,1.6114873,0.7811283,0.9419488,1.6869745,2.176,3.5905645,5.865026,7.6767187,6.432821,4.6867695,3.0129232,1.8248206,1.3850257,1.017436,0.67610264,0.47261542,0.380718,0.23958977,0.19364104,0.18379489,0.21661541,0.27569234,0.3249231,0.34133336,0.28225642,0.20348719,0.15097436,0.16082053,0.21989745,0.28225642,0.33476925,0.37743592,0.40369233,0.4004103,0.39712822,0.4004103,0.41025645,0.4201026,0.4955898,0.5481026,0.5973334,0.6465641,0.7122052,0.5677949,0.46276927,0.4004103,0.36102566,0.3117949,0.28882053,0.19364104,0.108307704,0.07548718,0.08205129,0.08205129,0.072205134,0.072205134,0.07876924,0.08205129,0.08533334,0.098461546,0.12471796,0.15753847,0.19692309,0.17723078,0.15425642,0.15097436,0.17394873,0.19364104,0.21333335,0.190359,0.13784617,0.08861539,0.0951795,0.18051283,0.318359,0.42338464,0.48246157,0.5284103,0.48574364,0.44964105,0.4397949,0.44307697,0.39712822,0.2986667,0.3511795,0.44964105,0.52512825,0.5349744,0.53825647,0.574359,0.571077,0.52512825,0.5218462,0.764718,0.9682052,1.079795,1.142154,1.2832822,1.4867693,1.719795,1.8609232,1.9068719,1.972513,2.1989746,2.5107694,2.8455386,3.0752823,3.0194874,2.7437952,2.5271797,2.3302567,2.1530259,2.028308,1.723077,1.4112822,1.4309745,1.7591796,2.038154,2.0118976,1.7952822,1.3915899,0.96492314,0.81394875,0.7220513,0.7187693,0.82379496,1.0043077,1.1848207,1.0732309,0.93866676,0.8008206,0.65312827,0.46276927,0.37415388,0.26912823,0.20020515,0.21333335,0.33476925,0.36102566,0.30851284,0.23958977,0.190359,0.18707694,0.22646156,0.27569234,0.33805132,0.380718,0.32820517,0.3249231,0.36102566,0.40369233,0.45620516,0.5513847,0.78769237,0.97805136,1.1749744,1.3292309,1.276718,0.95835906,0.81394875,0.73517954,0.636718,0.42994875,0.512,0.6859488,1.1913847,1.9035898,2.3433847,2.1300514,2.0217438,1.847795,1.5130258,0.9911796,0.9714873,1.4802053,2.0644104,2.481231,2.7306669,2.7175386,2.7963078,2.8914874,2.7700515,2.041436,1.2373334,0.97805136,0.8467693,0.69251287,0.6104616,0.6268718,0.6432821,0.6662565,0.69907695,0.7417436,0.8763078,0.9353847,0.9321026,0.892718,0.8467693,0.8566154,0.93866676,1.0043077,1.0404103,1.0929232,1.6410258,2.3860514,3.2328207,3.8859491,3.8498464,3.4100516,3.4166157,3.564308,3.5938463,3.3017437,2.8717952,2.4451284,2.172718,2.028308,1.8084104,1.3259488,1.214359,1.3226668,1.4605129,1.3718976,1.1257436,0.78769237,0.5218462,0.380718,0.28225642,0.20348719,0.13128206,0.072205134,0.036102567,0.01969231,0.006564103,0.0032820515,0.0032820515,0.0032820515,0.0,0.0,0.049230773,0.2231795,0.47589746,0.63343596,0.6268718,0.574359,0.48246157,0.3446154,0.15097436,0.06564103,0.03938462,0.059076928,0.128,0.24287182,0.53825647,0.86317956,1.2077949,1.5097437,1.6410258,1.7985642,2.0545642,2.3368206,2.5961027,2.8160002,2.9046156,3.0194874,3.2689233,3.626667,3.9548721,4.1780515,4.06318,3.7809234,3.4888208,3.3280003,3.4789746,3.8006158,4.2174363,4.6769233,5.1659493,5.7403083,5.901129,5.684513,5.2348723,4.7917953,3.7087183,3.8038976,3.629949,3.2853336,2.9965131,3.0818465,2.9833848,2.6683078,2.4648206,2.5009232,2.6715899,2.4516926,2.2678976,2.1530259,2.044718,1.8018463,1.4703591,2.4582565,3.5577438,4.010667,3.508513,3.387077,3.4034874,3.370667,3.308308,3.4166157,4.0402055,4.3060517,4.3290257,4.3290257,4.6080003,4.8147697,4.886975,5.464616,6.7577443,8.513641,10.331899,11.631591,11.9171295,11.388719,10.925949,10.486155,9.7903595,9.380103,9.826463,11.720206,14.795488,18.448412,20.900105,21.871592,22.567387,22.715078,22.449232,21.874874,20.74913,18.477951,16.78113,16.531694,17.092924,18.097233,19.43959,20.624413,21.78954,22.948105,24.247797,25.954464,28.068104,27.881027,26.689644,25.110977,23.072823,22.754463,23.397745,23.40431,22.386873,21.17908,19.751387,18.031591,16.059078,14.50995,14.680616,14.532925,12.757335,10.528821,8.4283085,6.439385,4.9362054,3.620103,2.7273848,2.3040001,2.1825643,2.4024618,2.7208207,3.117949,3.623385,4.31918,5.149539,6.0685134,7.0400004,8.008205,8.910769,9.472001,10.043077,10.610872,10.811078,9.931488,8.651488,6.8955903,5.287385,4.1583595,3.508513,3.1442053,2.9046156,3.0523078,3.4002054,3.3280003,2.6551797,3.495385,4.965744,6.3212314,6.941539,7.003898,6.6067696,5.5269747,3.895795,2.2121027,1.4933335,0.955077,0.6268718,0.47261542,0.4135385,0.43651286,0.44307697,0.42338464,0.37743592,0.3052308,0.20676924,0.14769232,0.108307704,0.08861539,0.07548718,0.08861539,0.08205129,0.068923086,0.06235898,0.06235898,0.072205134,0.10502565,0.19692309,0.28225642,0.18379489,0.15753847,0.13456412,0.1148718,0.10502565,0.09189744,0.07876924,0.06564103,0.049230773,0.026256412,0.016410258,0.016410258,0.006564103,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.016410258,0.07548718,0.08861539,0.118153855,0.17394873,0.27241027,0.44307697,0.42994875,0.46276927,0.48246157,0.4660513,0.44307697,0.4660513,0.41682056,0.28225642,0.12471796,0.07548718,0.03938462,0.03938462,0.03938462,0.02297436,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.0,0.01969231,0.029538464,0.026256412,0.016410258,0.026256412,0.029538464,0.02297436,0.013128206,0.0,0.0,0.0,0.0,0.0,0.0,0.013128206,0.016410258,0.026256412,0.04594872,0.04594872,0.02297436,0.016410258,0.016410258,0.016410258,0.016410258,0.026256412,0.059076928,0.118153855,0.20676924,0.3052308,0.17066668,0.072205134,0.036102567,0.06235898,0.12143591,0.21989745,0.24287182,0.24943592,0.27569234,0.33476925,0.3117949,0.26912823,0.190359,0.08861539,0.016410258,0.03938462,0.13784617,0.29538465,0.4135385,0.3052308,0.23302566,0.2231795,0.4135385,0.827077,1.3883078,1.7296412,1.8149745,1.4441026,0.7975385,0.44307697,0.27241027,0.9714873,1.9954873,3.0720003,4.197744,4.6244106,4.7294364,5.175795,6.045539,6.8496413,7.4010262,6.557539,4.673641,2.7044106,2.228513,2.1300514,2.5731285,3.170462,3.7448208,4.31918,3.501949,2.6190772,1.7329233,1.1388719,1.3587693,2.297436,2.1398976,1.913436,2.5107694,4.6834874,4.086154,2.0053334,0.5415385,0.24943592,0.15425642,0.16410258,0.2855385,0.48902568,0.6301539,0.47261542,0.3249231,0.23630771,0.20348719,0.2297436,0.28882053,0.26584616,0.23302566,0.18379489,0.13784617,0.13784617,0.18707694,0.20676924,0.21333335,0.21989745,0.24287182,0.28225642,0.318359,0.36102566,0.4201026,0.51856416,0.88615394,1.014154,0.90912825,0.73517954,0.80738467,0.86974365,0.8402052,0.7220513,0.5316923,0.27569234,0.16410258,0.08205129,0.052512825,0.059076928,0.04594872,0.04594872,0.036102567,0.029538464,0.032820515,0.04594872,0.059076928,0.08861539,0.14441027,0.20676924,0.24287182,0.15753847,0.108307704,0.098461546,0.118153855,0.16738462,0.21661541,0.2100513,0.19364104,0.19364104,0.2297436,0.55794877,0.92553854,1.1684103,1.2373334,1.1749744,0.9189744,0.79097444,0.7220513,0.64000005,0.45620516,0.36102566,0.3446154,0.40697438,0.5218462,0.65641034,0.58420515,0.5546667,0.58092314,0.62030774,0.5940513,0.58420515,0.827077,1.2176411,1.7001027,2.2744617,2.7995899,3.249231,3.242667,2.8488207,2.5928206,2.556718,2.4024618,2.1956925,2.0545642,2.1530259,2.1530259,2.0217438,1.8707694,1.7362052,1.6016412,1.332513,1.2012309,1.270154,1.4900514,1.7099489,1.9167181,2.0151796,2.03159,1.975795,1.8149745,1.4998976,1.1520001,1.1093334,1.3554872,1.5261539,1.5491283,1.6213335,1.7362052,1.7591796,1.404718,1.0502565,0.69579494,0.43323082,0.2855385,0.21333335,0.39712822,0.50543594,0.4955898,0.42994875,0.5021539,0.6629744,0.7122052,0.7056411,0.65969235,0.5481026,0.6235898,0.761436,0.7778462,0.6629744,0.56451285,0.47917953,0.48574364,0.54482055,0.60389745,0.58092314,0.5546667,0.5481026,0.5546667,0.56451285,0.56451285,0.6859488,0.7811283,0.81066674,0.80738467,0.8533334,0.9517949,1.7263591,2.422154,2.3827693,1.0535386,0.5513847,0.446359,0.4266667,0.36430773,0.28882053,0.21661541,0.20676924,0.24287182,0.3446154,0.56451285,0.73517954,0.7515898,0.761436,0.84348726,0.97805136,0.86646163,0.79425645,0.83035904,0.9124103,0.8402052,0.6301539,0.63343596,0.69579494,0.71548724,0.64000005,0.5907693,0.56123084,0.58092314,0.65312827,0.761436,0.9714873,1.2800001,1.657436,2.041436,2.3335385,2.4943593,2.3762052,2.3958976,2.740513,3.387077,3.0949745,2.7831798,2.740513,2.8488207,2.5796926,1.8707694,1.4375386,1.1388719,0.92225647,0.82379496,0.71548724,0.61374366,0.5152821,0.41682056,0.32164106,0.25928208,0.19692309,0.13128206,0.06564103,0.029538464,0.01969231,0.016410258,0.016410258,0.013128206,0.0,0.0,0.026256412,0.118153855,0.26912823,0.4266667,0.5874872,0.6268718,0.60061544,0.50543594,0.27569234,0.14112821,0.068923086,0.052512825,0.072205134,0.12143591,0.28225642,0.42994875,0.5940513,0.8008206,1.0666667,1.3620514,1.7920002,2.2482052,2.681436,3.0982566,3.2918978,3.442872,3.5840003,3.7218463,3.8465643,3.9811285,3.9680004,3.8990772,3.9253337,4.240411,4.6572313,5.1626673,5.3398976,5.106872,4.716308,4.7524104,4.768821,4.768821,4.6802053,4.3651285;
 } 
